module testbench();
    reg [29:0] src0;
    reg [29:0] src1;
    reg [29:0] src2;
    reg [29:0] src3;
    reg [29:0] src4;
    reg [29:0] src5;
    reg [29:0] src6;
    reg [29:0] src7;
    reg [29:0] src8;
    reg [29:0] src9;
    reg [29:0] src10;
    reg [29:0] src11;
    reg [29:0] src12;
    reg [29:0] src13;
    reg [29:0] src14;
    reg [29:0] src15;
    reg [29:0] src16;
    reg [29:0] src17;
    reg [29:0] src18;
    reg [29:0] src19;
    reg [29:0] src20;
    reg [29:0] src21;
    reg [29:0] src22;
    reg [29:0] src23;
    reg [29:0] src24;
    reg [29:0] src25;
    reg [29:0] src26;
    reg [29:0] src27;
    reg [29:0] src28;
    reg [29:0] src29;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [0:0] dst26;
    wire [0:0] dst27;
    wire [0:0] dst28;
    wire [0:0] dst29;
    wire [0:0] dst30;
    wire [0:0] dst31;
    wire [0:0] dst32;
    wire [0:0] dst33;
    wire [0:0] dst34;
    wire [0:0] dst35;
    wire [34:0] srcsum;
    wire [34:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25),
        .dst26(dst26),
        .dst27(dst27),
        .dst28(dst28),
        .dst29(dst29),
        .dst30(dst30),
        .dst31(dst31),
        .dst32(dst32),
        .dst33(dst33),
        .dst34(dst34),
        .dst35(dst35));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13] + src0[14] + src0[15] + src0[16] + src0[17] + src0[18] + src0[19] + src0[20] + src0[21] + src0[22] + src0[23] + src0[24] + src0[25] + src0[26] + src0[27] + src0[28] + src0[29])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13] + src1[14] + src1[15] + src1[16] + src1[17] + src1[18] + src1[19] + src1[20] + src1[21] + src1[22] + src1[23] + src1[24] + src1[25] + src1[26] + src1[27] + src1[28] + src1[29])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13] + src2[14] + src2[15] + src2[16] + src2[17] + src2[18] + src2[19] + src2[20] + src2[21] + src2[22] + src2[23] + src2[24] + src2[25] + src2[26] + src2[27] + src2[28] + src2[29])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13] + src3[14] + src3[15] + src3[16] + src3[17] + src3[18] + src3[19] + src3[20] + src3[21] + src3[22] + src3[23] + src3[24] + src3[25] + src3[26] + src3[27] + src3[28] + src3[29])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13] + src4[14] + src4[15] + src4[16] + src4[17] + src4[18] + src4[19] + src4[20] + src4[21] + src4[22] + src4[23] + src4[24] + src4[25] + src4[26] + src4[27] + src4[28] + src4[29])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13] + src5[14] + src5[15] + src5[16] + src5[17] + src5[18] + src5[19] + src5[20] + src5[21] + src5[22] + src5[23] + src5[24] + src5[25] + src5[26] + src5[27] + src5[28] + src5[29])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13] + src6[14] + src6[15] + src6[16] + src6[17] + src6[18] + src6[19] + src6[20] + src6[21] + src6[22] + src6[23] + src6[24] + src6[25] + src6[26] + src6[27] + src6[28] + src6[29])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13] + src7[14] + src7[15] + src7[16] + src7[17] + src7[18] + src7[19] + src7[20] + src7[21] + src7[22] + src7[23] + src7[24] + src7[25] + src7[26] + src7[27] + src7[28] + src7[29])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13] + src8[14] + src8[15] + src8[16] + src8[17] + src8[18] + src8[19] + src8[20] + src8[21] + src8[22] + src8[23] + src8[24] + src8[25] + src8[26] + src8[27] + src8[28] + src8[29])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13] + src9[14] + src9[15] + src9[16] + src9[17] + src9[18] + src9[19] + src9[20] + src9[21] + src9[22] + src9[23] + src9[24] + src9[25] + src9[26] + src9[27] + src9[28] + src9[29])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13] + src10[14] + src10[15] + src10[16] + src10[17] + src10[18] + src10[19] + src10[20] + src10[21] + src10[22] + src10[23] + src10[24] + src10[25] + src10[26] + src10[27] + src10[28] + src10[29])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13] + src11[14] + src11[15] + src11[16] + src11[17] + src11[18] + src11[19] + src11[20] + src11[21] + src11[22] + src11[23] + src11[24] + src11[25] + src11[26] + src11[27] + src11[28] + src11[29])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12] + src12[13] + src12[14] + src12[15] + src12[16] + src12[17] + src12[18] + src12[19] + src12[20] + src12[21] + src12[22] + src12[23] + src12[24] + src12[25] + src12[26] + src12[27] + src12[28] + src12[29])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13] + src13[14] + src13[15] + src13[16] + src13[17] + src13[18] + src13[19] + src13[20] + src13[21] + src13[22] + src13[23] + src13[24] + src13[25] + src13[26] + src13[27] + src13[28] + src13[29])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14] + src14[15] + src14[16] + src14[17] + src14[18] + src14[19] + src14[20] + src14[21] + src14[22] + src14[23] + src14[24] + src14[25] + src14[26] + src14[27] + src14[28] + src14[29])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15] + src15[16] + src15[17] + src15[18] + src15[19] + src15[20] + src15[21] + src15[22] + src15[23] + src15[24] + src15[25] + src15[26] + src15[27] + src15[28] + src15[29])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16] + src16[17] + src16[18] + src16[19] + src16[20] + src16[21] + src16[22] + src16[23] + src16[24] + src16[25] + src16[26] + src16[27] + src16[28] + src16[29])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17] + src17[18] + src17[19] + src17[20] + src17[21] + src17[22] + src17[23] + src17[24] + src17[25] + src17[26] + src17[27] + src17[28] + src17[29])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15] + src18[16] + src18[17] + src18[18] + src18[19] + src18[20] + src18[21] + src18[22] + src18[23] + src18[24] + src18[25] + src18[26] + src18[27] + src18[28] + src18[29])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13] + src19[14] + src19[15] + src19[16] + src19[17] + src19[18] + src19[19] + src19[20] + src19[21] + src19[22] + src19[23] + src19[24] + src19[25] + src19[26] + src19[27] + src19[28] + src19[29])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6] + src20[7] + src20[8] + src20[9] + src20[10] + src20[11] + src20[12] + src20[13] + src20[14] + src20[15] + src20[16] + src20[17] + src20[18] + src20[19] + src20[20] + src20[21] + src20[22] + src20[23] + src20[24] + src20[25] + src20[26] + src20[27] + src20[28] + src20[29])<<20) + ((src21[0] + src21[1] + src21[2] + src21[3] + src21[4] + src21[5] + src21[6] + src21[7] + src21[8] + src21[9] + src21[10] + src21[11] + src21[12] + src21[13] + src21[14] + src21[15] + src21[16] + src21[17] + src21[18] + src21[19] + src21[20] + src21[21] + src21[22] + src21[23] + src21[24] + src21[25] + src21[26] + src21[27] + src21[28] + src21[29])<<21) + ((src22[0] + src22[1] + src22[2] + src22[3] + src22[4] + src22[5] + src22[6] + src22[7] + src22[8] + src22[9] + src22[10] + src22[11] + src22[12] + src22[13] + src22[14] + src22[15] + src22[16] + src22[17] + src22[18] + src22[19] + src22[20] + src22[21] + src22[22] + src22[23] + src22[24] + src22[25] + src22[26] + src22[27] + src22[28] + src22[29])<<22) + ((src23[0] + src23[1] + src23[2] + src23[3] + src23[4] + src23[5] + src23[6] + src23[7] + src23[8] + src23[9] + src23[10] + src23[11] + src23[12] + src23[13] + src23[14] + src23[15] + src23[16] + src23[17] + src23[18] + src23[19] + src23[20] + src23[21] + src23[22] + src23[23] + src23[24] + src23[25] + src23[26] + src23[27] + src23[28] + src23[29])<<23) + ((src24[0] + src24[1] + src24[2] + src24[3] + src24[4] + src24[5] + src24[6] + src24[7] + src24[8] + src24[9] + src24[10] + src24[11] + src24[12] + src24[13] + src24[14] + src24[15] + src24[16] + src24[17] + src24[18] + src24[19] + src24[20] + src24[21] + src24[22] + src24[23] + src24[24] + src24[25] + src24[26] + src24[27] + src24[28] + src24[29])<<24) + ((src25[0] + src25[1] + src25[2] + src25[3] + src25[4] + src25[5] + src25[6] + src25[7] + src25[8] + src25[9] + src25[10] + src25[11] + src25[12] + src25[13] + src25[14] + src25[15] + src25[16] + src25[17] + src25[18] + src25[19] + src25[20] + src25[21] + src25[22] + src25[23] + src25[24] + src25[25] + src25[26] + src25[27] + src25[28] + src25[29])<<25) + ((src26[0] + src26[1] + src26[2] + src26[3] + src26[4] + src26[5] + src26[6] + src26[7] + src26[8] + src26[9] + src26[10] + src26[11] + src26[12] + src26[13] + src26[14] + src26[15] + src26[16] + src26[17] + src26[18] + src26[19] + src26[20] + src26[21] + src26[22] + src26[23] + src26[24] + src26[25] + src26[26] + src26[27] + src26[28] + src26[29])<<26) + ((src27[0] + src27[1] + src27[2] + src27[3] + src27[4] + src27[5] + src27[6] + src27[7] + src27[8] + src27[9] + src27[10] + src27[11] + src27[12] + src27[13] + src27[14] + src27[15] + src27[16] + src27[17] + src27[18] + src27[19] + src27[20] + src27[21] + src27[22] + src27[23] + src27[24] + src27[25] + src27[26] + src27[27] + src27[28] + src27[29])<<27) + ((src28[0] + src28[1] + src28[2] + src28[3] + src28[4] + src28[5] + src28[6] + src28[7] + src28[8] + src28[9] + src28[10] + src28[11] + src28[12] + src28[13] + src28[14] + src28[15] + src28[16] + src28[17] + src28[18] + src28[19] + src28[20] + src28[21] + src28[22] + src28[23] + src28[24] + src28[25] + src28[26] + src28[27] + src28[28] + src28[29])<<28) + ((src29[0] + src29[1] + src29[2] + src29[3] + src29[4] + src29[5] + src29[6] + src29[7] + src29[8] + src29[9] + src29[10] + src29[11] + src29[12] + src29[13] + src29[14] + src29[15] + src29[16] + src29[17] + src29[18] + src29[19] + src29[20] + src29[21] + src29[22] + src29[23] + src29[24] + src29[25] + src29[26] + src29[27] + src29[28] + src29[29])<<29);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25) + ((dst26[0])<<26) + ((dst27[0])<<27) + ((dst28[0])<<28) + ((dst29[0])<<29) + ((dst30[0])<<30) + ((dst31[0])<<31) + ((dst32[0])<<32) + ((dst33[0])<<33) + ((dst34[0])<<34) + ((dst35[0])<<35);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h0;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1484fdfc1bd5c3e75b68e6392c2124c74c641c9860679ae72543d5dafd639edb8f3d16fc354b788c977ce5d3a0291617d30fb66bda53144e5136b34f2d806de17848c28ee9b7d0eabaa361758b6934559b55933faaebcaf50980b873b79e233db8a8fc862439ba47b9abe327bfebdf3c0;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfd842b0d7486aae7e4d38d7c00f12239e12e77df6fbf51dbea5e116b28a38953e039570996b1988a62337a2136063bb4f2048ab528013cdf59142d00cedab05a931d2545a672b49d9728fc6e6221b64d3b8ad278ac75426fd4a3745c9cb99469c98431540932b8b5a8f1c096aae0cd1f8;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb4df62dce02d9d67b27469da798bdaef66cc474da52ceeabad3400a9e208d7c82d7c99baa74bfafca55f733a84767fa0892e0da430e740e187b2d0ad154d138b0c09e70f19fd50e375d87149203a74ee1b71d05c9866f29629ab919c169cc2ed6fbce1dd74043984e8c5a74db8f1ebcc7;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h12a86212b796c245e9399725a2c53c4f49e2e0191f82c3e2b8127e77446b3c21b79686db59fac7b5cae8fba920ef7088222f29ea404b6f9e4b719ee0cb2dbbe2cbdfc009509c0cc13fb1e424addf19f8dab3241ac7bfc3601481c23d514db6735a62a5844757ccd3daeac0606ad1d0397;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha068a94202277804c0f8f299a72f536ef22354437cc57997d7d2af8637d15bbd878eee3e83f010298bf2f33557db8a8bc483ad24ebc0bd8c5c41991f955b73d9e6eebdd6b573dcf094890cdeaeb0417e529fbd34949b45e447f646be6f4bcc3f2b5a6165224987924629c87662c80ec99;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7f5b2720528829ba7540f9c8b8f95e8bd72fd798590fd5e67a9e22f6d761e3127b81a4d8a37526d5daaaa953011972876e88ea035399141aa7570e780f77c464e4ff7a123b4aa1b4420f0c3934b4a492edaaba6429460240284e93d4e127797ab486f71e33420a16937620738388f9e5d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9e74773065547720ad8ba8587af1cff43d25d2d47df6191fb7e7fd93adfa5a9246f17aaff13746a930b405fd6ca57c9346afd8d27c170ba012903edee061fe2bb193d0b047b828a70640430cdd17c76687718dcac2b991c555ea02c4c737ba38a7dce7c4160e148a5e119dbf7f0306de9;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4584e41d59b581d489f39d785f137b4236f7044f038a467acda14b414c04e735eb9cb2a3d1bb707e6b32e649cbcdde8c5c74d20f1701fef9ad8231102616c3d8dca0e2ff2155c5f6eb14a5574f36dc282dbb63361876065b8b77896614af6ab2ccb49921dcb6530595f93033946202c13;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h526599e4108428c5eb21e3b8f2a2ae5c8b4dd621c90d6342dd4713a0558060e2a354a4fee0b9da9df7148acad0e13180937b76c450f965aa082680d577b1cd54afe626646e66757cd351a1dda3f4fbfa36266a43c4880b2d747fc1affb23fc0f513e9de2915f3407ce36cc7c288a7614e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf12fce69ac504af7babc307d553cde221e7c01d0da29ab3d3e97309dc4742350880491a72d7a55bc4f26e8f7abd6bcdd796e43ad8338ea9b1a4cc67b93d0f8bf3473c68be90573d9bd557af767ace20793ff3ec3359636a71ba21f777c730ec4ad6f73ae6a9a4a90ad68d9eb88c56bed3;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb5c6543018efa045a50f2cdee24316c68df7fecffbf4e9cd1540cbfa0bbbe01c14460626b1423e04a33bd9c67edddc1b7d727f1852b91bc10c9e3d6613d2bb226ac462d7c51fda152dd12ad1a13092b32fd6623ec13041c0ad9d4a3c90c3c7d2d793d29ee194db6e8123adf341314353e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he99df523f148277279b96badbe47b5ff25d03b1e063302d8d57e67e3566344968459c035c38d55fb8001594355b1d2fda1acff63a7921028668c11a04e27d476636b2f4ba7b3f93898dbfa46edf0a25aacde51a3b0009e7d41a12977c0e52aafdc8493a4a2f2704f2aa7bdeeb97748432;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5206a68aecc5b2cfebf56f55b13691e3d3ad3bfc8d1f673ab5e3bccace6f48a8e36fef71cde3100de28b068c309599e266528f94b5494cc9cc63bbe4f49a765274ed903d89d8f009d3ed6238e4ed9af5c5b644609ee9547b15e5dda706606e0ad5bffa9c141291564c8111948775c284d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hca925ab9f5068b5f241b07bd599598ab8fdfa8d6b088fe7b9e218f606fa87b195c12d397e358d8413ae2fb648aabff419190db18728f8924b65f83dc32b3f3ddabd8d73dcecfdcc194fdb4e1e924f1170b7be0703f07f5fed65f895bb22cdbd1184e34078a42a75404e44170ddb67e930;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h627620412a974d52c2818a9a038e16554b52a7c1300c9b2d94d9db524ddb18711edaa6e5b8a17308167c76243aa8dc77ccfb10d95acac848a3fee26059a7b86e6db81fb02603d859cdc49972521dc29c863551668b8df59e14b21b956ae9d72a85310ea3c2c3abba2084edf92e1078203;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7c78b081bafe113e858a06c36bd401a11d26b5d37339b90c6526e8b8694e4005d89dcfe335fda5d17b32503e59b5d298cab5c8f2642d0c3af8aa2a8fd9593ee6ccb4a113da16f0effdcce95ff20d97778f2dcebb690d10e6492bf6706daac28e8550de2f7da9227b604d4b82e6ac58f70;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc5a28e6aabc9b96962fddd6de609696be2bbd0bf3319cd796dddbf6bae9724b20c930c16446c702df07dbd3e1da88aff555b5e109c483cf8e2507f972d458d52910037a0470600192fe83e38d6c733326ad2422e50d886eee407626db38410ffe803f290cf0e1688f2cda030af8379b20;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha5eabd20a043a8acc145db02741c97eace1badf6c617712041d9191a639b68032ed37dcc927a867356fd2c807032ae2477f935547422e3a86ce20818669d42d7e81aa532955e5a3e4e91446a8c784ab952fcbd4a47a52ab893969800f203b5c37816e49eaac43bb9bb5c2356902d4e185;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9112e9e945ac4cd36a5593f8e752a842b9b4940499199c75e2fd33d911334cd588ade5c93709b9f24d9a78674d442373074f420f4ab3ee6464171322a07132f8de5c460d317347b847b7b87154767ffee543965b71dd1afcac576ad50f595852ff4ac8c5393341088c86017d0c0229771;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf02be6bf6c6000f710d7ebc2150c86f144d552e7ecabcc422d470a99a220ed2fd22aa96d6eab9f060a573087ad1d8257a50da338f37c6fd23fd83ca2bb12bf2eb7abe4c54927a090c8e55ea3d11b53f0fa8aa8328f48c3d6d8528a2613dca5758349a247c735580ebfc5a0e727b24638b;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3baa2f2506b24bc46247fc269b528b3faeac4fdf072d291b31431e8419efe2911d55d7ce4475e0cef7237e08c86bd225c3a692119970be07c5d91895ea3f5f627a21180c8eafc6ffbc781d3e193f0e9da3916ecfbdf37951052e8c3432faac9684f6d2feddc4f6f752553032e1e3e89a7;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb6e606a91335d7355a06bf53c96c71a99d1976006752396a34c7c0cb97b875b1bf920469c50458b37edbb487add96ea5d06ac0f445db2b536762fd169cd2ce7fc90ba728ec8ff894f55097af36cfb0e70d404fcec2162e0209a6aa1acdc824e5c86a9850486df70e8997320c3ec7b490f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6d8fddbe95fc81be6011b7c28235a8332f8cd0e2738eea7b3fdb518b693b1be7b43b5dfdc19ab0684363cef11c34069ed3036814f4aeaf536612a0f19997d4d771c9898d592f892665d91239f669591593f3a47e848fd1a8d8639d54ec2ee598abae03f138dcdb49d842378d48986bd57;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h749f2927c38494f0127d19dff62f1c9d46bcb5926b9bfeef8ba96a079cf3674dac3b7da8700d5a1e173ac551b5f377f0c85c491c5e1b8ca6ba4c23e244afe8f4855c21070993b4aaa293729f1dcfaa68cd239eeff704c94a34b49f2e11e72e280eecb9c6ca76a5bc8232a82901ab9405a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h38d313dc5fe42dafa852f64c016591327abac54ad41139386ac6bf6c2995cbc3998b549cdd9a6456409b8921ab7dc22e72d50e022adbbc52a6f930d5673eb43d7ceb6e6ef28a3c8b12d602250061f16185e46ddb7bd38b1aab9864b127b476f4151725178ce84d50fd1b1e0d7332e784e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5a3246854fd059403602af9895741fb89c20e96b4e803da63ee1c26bf61faa0a17c42a0bdeb059ebf9d054a8af5abf9bbb9a1bfb0ebc33c191a690a0e135c3ec2fdeefcdd70ff60488f148b804f8654060fce60962e9d1b2eac47f9d69ba3c891b0035ba923e6efda440cfe3b4920d86a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2191a7759a8f7442f6a26a6721f8cd7a5a3a26cf74877bcaab7a2ccec56d80d3cf00338fd9f0f0a31e90bba80b2d69cb659161add17a6272a322914321b4e6b631f553cc4099a4bee64868b0e6d61966eecf2f5252ecc99c547196d4e209f46c25f70742a21f4a430d93971e5f3e25a8e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hccd466cff4e0a504d0f62e382532b1e5f9e54772b97a75c9da439cbe39887a0029b96f1a0c125aff7ce8b73cf98b3f98c1a73301d95640c28e6caf7b1bb6666fe60247c94881bc2e3e562b1cd5c4122e1cc7d07e6a4dc859ef41b12e5c3bff700acfafa72110f32ade07fa8f45443966d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd8d10337f288cc012a92e18dced531f6ea8810abfe8d2fb9e30dcd7e92bf89ec174f1a5caee8ee54956cfa845115ed640ba7058c60a09c7c5337a364fe1d7e9abde9af7e4e8d55ab5bb01bc27f47b441b03f8aec30a6c6c4953157f97d50095c64d68cf71f6e578e6f92e92c11e16724b;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h37880ba0bd86f313106b6dcfb8894027c313ea3cf220fac65c238ff150fe7d0040190198818e936f453c5c11f0d073afaac28b45f23798b73bd6a2171c118a2c8249be0c3be6df144d3f845b610f9d6e3173a8a174dfc1d6a3b4308ff4039156103a88d68fa3aba630ac63368b9da3984;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5a8c616eb846cbf0fe8924832adb6ea1b65f60994352b5dafbc2d45019425d52d8a3a30cb1e31852eec174e0240d1ce93d7c919d6cd1d37828ec62e3a70c2fc1dea9ad274603936ba7ee42da0b026425920a48fa0ba964f71a5e5a1cdc0e8ae6dd52bf3acd5377e2f68a3d6f8711f8024;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8c222242f4b96cdcdc73bfc1556d5189ec9e9e6cd31193bca1975ee0e524a63cbb38884a5d8c6645c098423fb9524e2203e77283a37017fb69b5f7c93d9daf758786f7869ea463436909972f653462f75b2013b368ca1a2b33bfde28183eb35a256764c4c3e15cdc64dbe1dd6be4fd9ce;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3197f8121341f38100cfafc56bc511f167779c09246295d6609415d156b5ed90921d0c521553f3460d6a5dfb4791fddb4a171e3cb51e6c5e20682a5051af74010f418b4e4f5518d83768aefefe7bdc24b1e27fe497c29420a01cbe5f036e4c3b70d646eb8cccf8ca58f8f61888e6aa1be;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1c5b63afcd0ff6d1e883b0174c127c7365eed6f13d203bfb836be8313bfa836922263ca349abc1da7ddfe0002a2cc529bc1887a2231b28fdd1bd748fc5a35a20a6a61448bafc6785370dd4e81d374087ff9b688a55fc2adfa91f238b992c039cea00e1d78e2ed498139a3bece08424867;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h20ae50131bd5b032e2e2e744a142484b999c0201bf48c8bfeb7ad2c4a5d9e880d9b1bc4d961a73cca073d5241403e5e3023fea161787ad03ed75c9bb61ea674901822c04d926028c5292fd0e7ba77c16ca82a9e08bc8950788c89941380b17af8e30908273cc562216b6be5a4e9110a81;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd66f601aab6f401449cc13df9e5c624aa8c1c50e28f4203e59b738e6428141c1994f73b29aca04d427868219f30c8802b8ccc19e8e17f09a9991c252c64e70b92642c9c14f5d2c5408f04ed50d7aac10def65939509a62faefc00dc1db1fe964c35a9d2521c75502cbe674321923cc357;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5a83f8a77cf1a6e60ba053ab27d0a4868a5a9ea7db1ad7cd1d466db8957040634c437836276dd5cc08e256cb36e26d7c7652575ad2a75566bd0b8142a342720cadb8ae24d200f83343bf4ddac055a4b654a06bad050484fda0f892662835b1ba5e86fd25828ec71385974805c814f6319;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h24b721b52946d04426e41695c71220f14ab34999bc32b8c13fb35bd2e9395710ac61effecae333bb3335d89e4e4623605d21fb1c1251d745f6bbb30b32d9f4b2756dbab882aa8463f6a1cc89034bb805a64f978c415e519a4e9c3de597a3b51efba0c052fcc8cc2821a3237138d3c929d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha27752560903a1d96753b8dbc1db9a0e1ceb9dca54651effee79441207ad453654b6128e851ae8940e19cf5cfb9ae1e02c7418fdc3639232cf880ae7b5b79aee2a653509d48e980cf7c875a7659fc88a8c13eb34c744854ca05b29ae6aa04b072ed3152affa7b20d0b3557cb8735e09c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6cbdb6fe067c5561931c9914599e402ac6b6aa8d64116b8b6ee4ec92211cac6e118496558a9e74de4afece8dd455128ab74417820174229915f66ac35a3f2f4d8e6da85dfdbf7ebfd28d803838dff06a433f415cd0c8f3fbad12381e7b30930385697fdc94e55f7fb7d9bc37e32876768;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8e55e9618775134721eb2bb4b37dcd11ad180721a2aa626efbbbd988d4115b05978b9fd4ccfdd8ebcdd8e8b3551cbf23ab44c7e6413c74202fa048500ecb2ebbc700668a66976de17942088e38efa02a1b7e18ba540c59268cdda8a6622873d096ce03ab80dc36fbdd79786c51a25243;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4ebef98474c2462b38a410d66f0fdf3fdd332c57f870cff3c0401eab28250e4a0aed263172ebb654a5143908413ac9082d9552ba6739fd26776379e3986acb4d1e391504b02ad26ab8c82d40ae92c502beb35d7a17ac545892c0f2f06439f0a927c04be86d79cc9ad2d13406196ee61e3;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf85d14643aefae762302794a003b8cf123e84b236d97cab9df3e28eb29f7a94559f9e98421e50b5934bc9a318f8550d556a21a024c139edddb27165787be9d1b3917c09845da063ec65c4808741be1bb82a9592a99a260cb91a2fe448e97f17e90175c1c60c3a6a3a8969587a2e1e0565;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h806c354d42ec977a3090780e2de8660eb2318a4ff9206ed454e54d09d4058b6e8e7c18f64b563f9d3b19eea249c61baabb052a23b3142f241a3d054d861eeb1015112970c4e8a3f4c1026a3acdc485570ce4f19a889cc832dd9ea44dbea36973ffda5ef5c7a2c940aeb2bc0803cd2c827;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf8f40554e070928ccd8fe7136b6e3b22a1912902195ab17c25312e6c6a6783d7fca0766de70c3a158e8ae1553676a31f538c116ba25d9e68dad228c11d63cb561149e53e1a03b261425b021df47f6044763ead4c8a69e3170faec98e8bb99dc848184bd70ad01139a71cca5481602584f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7adb01772d90dab7323fce23cc032a615ec40dd100bb0e4879f928eefc9af583e0104e0a0f5e9a5ab5c30fbc268eada2077b2d2eb5964f09c39275f9a737dad5f5559c6451d977b679dbce69010c6e92be929950b576dceec8f9cb11864db74cf31e12670be84e6cb3c30b3f596f7644b;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hede51871143f2ffde07072973e01ed40476dac3ebb3ffb23b2f694184a92e39eb25f00501cd6660326ae3590a7bed3d02d30c3799acfafcf96157ba43472f9b482bbf4c2196dd9d3ece31330a9798be90aff825490b35a4cbd53e28a7b837cde3863c1c82a1ae1367e84e9c2727959a1d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbc3cbc60913939e3a06abe5930da26960a5d814d801ae1bd175b8cb77a99f2d1251aed35fb630c8b31d31a3d0f775750480710215254367570d197277ce4b45dfa24351cfd053325d2056aaaa972755ce6c62ad0793c83e8bef39e417aac3d2e0f2132e70a095ac47f7fd2b269b04c743;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h34a7a2cd23e68c2f850383d563cab3cfb112618084835501535c2ac2934bbdcb630dff24251645fd26cfa1e74530cdc78be32512b2c1a1ff9f94f7b00680acd78c05b99769e57188e5dcd2f23f866fe430de842e7cc38a79181b1a385bc722c4e807a4e4f8f208b24e908d00dbbf5491d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he8db065c877a4a9c3b5fa6795d7ff3008c116251802dda356e80695bbe0715feb754662457328706ab5908bdf74a569897bc23215a7961575c48211aa2822e41f84e0974d5d54a5481ab918551c23812f79f1bdc55e375acc593619ea97826e777cd3942ba0b2f476b99c732bae344795;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h665aaf2e9cbb1372a11005edcd97cda1902baa8bbd6a67f3500f1d862e9daba0c0b2fea06e2422e14fc906b220d63c57b511e0d14aa98f45f0e800ccf3210cbb68fe1ff3dd7b641c9dc40f2dae29467918922f75087ee52905b32c86fab21b3313ac8ffc3ec910290e97c15ce7aa947c1;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h30014678b51078cb442fbabce301e445e1e773bfd0500efdc95e5c96c8b6fe7fab1ccd31294f40a6a898f1d2e7041b1fed1c02e3a8ddf497eaff1380dc59c21a2620f40c7c9a8215c25fd424d21e63dc8f77a340eb382659243feb112a342b5e8915f772c3da53609affab3775b0377f6;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8933d9158cc9424e3a443613ba82d9c0376c6272b947bc55083b687c8241f1c4b36f5103c54773c6f0b22b6ebf854c4fb4051177a0afd5ea8676ad25e52509872a0f7cbcc938168c4f8c243dff71ca9e764aae83e41679ee64341995420b26175ace34da896ac24340e97dbc32a1f6254;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h97ba2fc5b8bf41feed13c7f49f98f7cb9894e6bb2cddea155a65767990c3ea60696afa873a72ccb93999d763fcb6114976e0cafdd09deee8387e40adb6ce9c9f6782575b7d228dd8a8fef9771bd4e0dcedd6d3283924a6e5f277df9e04cf1e19f863237243901e2577e55884fa7193c01;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7f6d11babdfc64371e17e771c7e833d6762e0bc0a9069e22f025eb70ace44fb555fa24232bc7e8324cb7661c6b5e937cf51b9092409a31f7835776a4c3666bcf9af21fbe83c5add77a8ecd63eb3ddfb80aa0a50753c7aafc6ad59f189ca103bc1e5b357ee8579aeca53b4cfc2b05f7468;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha333eeab2f803a696c5d25220d1f75dbc7c11adf595bac0ab5c2f5cefbeea4769b25c76748d33d3051b5a79ff98501927f8140fb0dc37b2d0321117e9b355e2d81c0d2f70ccc3e8b484d347d9910c88c525911a9506e3e82c1be4e3ed162e9780972fcb8ff453c1daf827a48703de7fe;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h85ae5b767b075b9c3d6cb6291b1471ba3c772774fe0a5b5f739ba613162378ef3f576b6f2c90e7be7325a6cc2060f713016dd60d9904266b3125d51922df77980ab96a3c7c655e1577f0bba1e5132617fd390e634f2641491b4cf37e823b5336d556275a0749a4e966e98ead46f777ee0;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h92e3bada74d042a37d2c2b70c8069a154c471f81e54f7c207eaa150a935ca3b042a3ca1fe3b8928778909873faba31eb6f6099f9413aefdcfaf136def534a3550a7198466db376f4389ef36729556919fae665f41117e259a2e2bdfc5a6ac283f2925b94c5a3481a8a27b8972a37bf0bf;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb3fe5f4585e8a55439325a474cde6ba39b52a8dd999913fd941bdf74942e453dc93d586b8b4c7e51c09270b6b73a65e4713795dc36148a5facbba9b2bab22502dca6b9fa587fd4330d1cfd26127e56434fa7f2cc583ccf747a3d1e4babf583a09c6ee7db30af9b44d0e793ce50d738c9b;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h322a707bd8627b01fcdf6a4321885dfee4f7c28115f03204d1a5c7ca91f60964ca6fdcbec7f127f3c7885b210a98a6d2a1ad6c71a530a6963192f15d310c05b607bea3b5e0acca720674e5202fe22d7be999dbc2cf0c25cbf61ea7e82589404177da6996bab9f9d495937ae60289385d6;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h957d4436163edc5961e1f52c5ac6c0e8a6c8b79ccdfeb992c04c7f550330daccea0a22fbd31ef7c04478ca716ae818b574a3cdc0857005fa60a51e9ff102035fef9291073e6904e203503421e197adcdca582f946a0a355c2f4fa321f101f8faa84b99605a5373680bf788c0def21faf;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h43423c460be3294160777500fe5fd8520d3e08de828616dd05278051775667246792ab98bb77f9127b19bdc6edfd2471ffb2cdcdf89b71ce563bb916278f44c9dd319bc9a70bb7255b09e8ec9905dd30c9cde3497fcf92c19c398cb97e069b35c4dd8ac533882fef752e88c9eadef80e4;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdb3d8830c965beed67f0372246bf9ae17d5f9c961dd19d02a557d9c7a6353147889db1b92792c2d5cc59ab05db90b6ea6204ae6637d8d72078c4eefb5bce18deb28fc99eee75446059ad231d407b69984f92be832e20f802e68018875350d0d8646924c8e872899f02e407f11e5f9c254;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6938dbe824700900edff684360511a087df6661c315dc3e2a4b541b4d33061661fb49a47d3992fc9206e908d77d16305e91c177c321db76f6acb09e93e7f94e9ffdc24e289a88bc787f05d01360d5f00b17f212ba1a7c6052122e94295dbbfa07f2c4750fca8b9ddd7a242ca96b6616d8;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5e9d27ba03d301ae0b6a00ba998b410759e8724215d308dcd3fad4aaa525a7db873dd36743ef819af9445a7235b6918ab21fbc8dcb661d3bf64b5865a3899092241e06ce7a1f4e48589b9526ec9bba5cbdd2ce8a26336911e80b31b66f398cdc77a2d164349558763d7835f804fa43c7d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h17c3b93afdbcc24733530013c81b5a11ca9c0d09f088d895bf2d2baa4a203b3cd1bd9ca22753fe4b364bce9af2d435fd654415af59644f7b020745b71230a2b63ebd6f99808d605cb802f3fa44a4f8308184386eff25923d8d717b28f646870c5121e81ef9800141999c94d812c89ddbe;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he0f7c177065fe6e66eb59d0a903d7ed3de61d8eb21b45686c54d12898a89d73e530226d3e1546dd96f5272c38169a5f48342dbeca6236fa4ac9816cf4734102e01aa7e9674a3ea562a5bb9f0e404430334fba85d3b80952485ddab300e782e000d9436600cadd4357f5f9146dcdf7ae76;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd4f12ccc4d9597699102b8e7adf29492e9272acf7630e14d96d656f650057d7b2cde26a14977506252eefa72796685b812bb7141a5036ca144dc6ac8933ec780fbe25af92b193ce9d6b6f24ff10adcd24ec69d8a3ef7aec8008b87f79cdc44e4fa37fa5cd0128ab20ae95ef8fe745e6dc;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he22185a138bebebb3a11c05e4fcb5b4e690d599cf8d67337a7df15bdeaf68e42405c24d2cfdeb6f588a7882863fe46e2df6a803c968a0d6345923d032307838e3eb2a2efbc51173ce59c968f65999f7c83280c5fe90dd936f604254c3f11bc76236ed358a9c5bb5b2b8ed27f2fab20e8a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h943eed68f93a1654edd01bd1c0a67ccc6191171c0f40a19e8ba1824bcace3e463ec55c3c17885986a2db8c88ff24b1bfde972e5a0b44346c05a477e352629f39f2265424e8e26b25abce0899ae4ee537dbd64588cf6ab12c79f005bf2418e90d7c39b9ab0e0e5e79fb352c0afc8de19e3;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5733890535374410570625880d1f8eb13222891e3aa19edd9d1780126049335c0ed6c0a6422a2a15ca4709da7d7741a562ff1f9ff556fa1925f8a4b6c57a429267fc3cc901756a0da575e68f6332545f8b8e9953e2c818a6b60ada83770c327fdf64c522eeb204951060c090afb906b48;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h119fb7a68685199b1a078c32e979d5df7d6941b56e773e0ba622b6a388d7d55e2ae0049261f79f42f6b847f96edcba9361ea3712571f2bef9b7fcf03c73ec5dab97ca7a21f35eb07b56b4d401622b0b54deb3a8e92cc7bf29276c9c5ff56f86843f7d7d1d3a30b19c2198924ed743966f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2d548c44d8981dc8ae65865c857e3d2d9d79c0fd6114d93573bd0d817100fa687acb8128d88161a18cae8ccef7f55d10101bde25a23cd0f0338d8153fa143bd8e5510f6185ceb9e927746f138cd5f5c8a609436104e2180b454c79793b7d930c43af5183124a31ece01cc233cad177e66;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5fa0ff231c004f030dc02203d34758193c04e69f4edd0ba2f50a146beb24d5b319eeb4ac3d89ee1c0648d181cab6d6210949d20f1740ffc9f96edb7b8073bb61577bd04396eaa1fae352ea939e17147086058f66deb5b1e78aebc44ef8fd39899d9230ed3c6f402bbbf88eb1e256fb9d6;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h72dfc1f507f76160bd898a6571aa28ab83499b229bd2a9ea3c7cf3e5498fbce0de589ca8d1e4a6b82ae5c5f0da29ced638630d3c0266514cda46942a4d0a00e569cd428acf166af2950c0b0816cfeb11c4a35a0b9973166f9c2c8fcddcf7009191a53e1c9a21ef4aa08f7f03e4b19b60e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8168689b7c60836848021cba61004cf834186900f539a1c840d7877c7f46bd675d33f6dec5733aa1d8a7748a71346f3b77ef28648f286eb12dbd12aa035b801e48a0c898a60f4b2d9eee4a79a2722cc8396f4a709e141fa4ed8bd3d855ca1d524429d344c5bce71b2ec497af647cff07d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'heeadba932634b5749d28479ef8c4b573747ff3205285d0297462e600bc3c09bc1f7b34f5589e396bda7d722e7386a7286a41d9a93f70ef769d52557ac0fc503901fca7c8659973ba2afae3b66e2d42d3abaf611d571028787916ed7ecaa87f6f3e403ffdf5b3ac1efe49ae621f9d322e7;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbc1e47cec3194585ccc0a6a62aa4534b413eee002d77b74101af7b2acf6e0adfa169354d45bcd826d4938734d9b3692a44d56dd3a78a13c078aa1039a5b7767beff90e1c257fb437b65f7a77f5b6a6e39e447796e9f561e9ddb4620d3c090aa2478325ab953351b706109519f89a6d771;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd749435855ffca53d8da6eff225928d5c1963435455e603ba94f40273705bba3efb5801984a4a4277c904b8c89c478eedc6f27018ddad1e5d6d8e17c29c97fae960193b566949b470fdf0a67bf5813c16df588da9a70e702825bbf8c8cf6a5e4cf6ac5587d56e2b82f0a4b319be785589;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he10b4322ac5c2e11ff693c10101b4ed2d86ca5e9c3b65b204d59dbebf8c1edd797f0a88cc824a5be02a6c41ee73bd41fbdf3cd2ecb66bca1ae2edf5695189ae70341dee15cee97b61e5890b3998f82cfae0e10d11c920764cd4b2de5b23533775fbb4708a3c7db437529e31e18445fe68;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h135fa721469e267a61af67c9da7a73628aee770b7c3a05fefb7e069233bfbd10c5b24f092a35996581efb1a3a1eb84fed023fe73b87beb9254d74b959f51c296cc5a22a907aae68f6239d46a5a3d323dcc95770346847d0db7c85c1c8d9e39c5d8d166f4169b85a09d37afeaba11be780;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h857d41f66a11a29e69ef66ce292c1a141c19f4e650e84ba33a9fc37bc02b726637f9f46c493183ff54869e28a31e953d0a1b0488d94663451d88b02c2a439049070d9399bce9e6a43ff49f0cf11524fac0356f0bc794c210e2f7725c4549e708766115963c65c7a5674fcd607e398d151;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6873aa3207d6dc8b0d57903011ec353b6b335a7ec1b3af6b7b5b45105b8535fe96036820149fa8d6ba522bcdb3c4fe1154b4efb04cb0c5494fecdfcd664c0c603dc25ea3381b52c7e7d4c36f4936bf96dda86560ca9d524b4df4a1b1ead42c087a5dd154d60796820d44d985c4621f7f9;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7a25057c6f5161e478c6455b744129e817ea6486fdaeca9f03205259b13230f4545c22313c2304905bb6e25929044cb1d0fc21901114b218c9f8e591e6ecb73105866ef2f41d35466860b5143d0da47a3fc9c8581371120c5b3ed69b070148e695e432f5ce9ab118ec9f0b0d3c09bb377;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h36444216a5a1ea5099d1bb0d0853895332bc8f8a25d52caca3c4d17bd818df23c4d3220fc061eb0193e23ff8c9e7800d09bacb71f2fdc182ec218f74ecf0f8685dfeb9cb46cb95ef44f12185c4c7f54661d976247718a8a1358e78cf517f8fea0db3c238cac72a874104a00df6b01adaa;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h778c51e08a216c08f575c12b35df4359f3aca2db2c22197e97ddafdcb603b89e3cadfc6a27087aa5011520f65f6dd04af3216cebd7ad625f103f081486386699bf695487529d39378820a0e616f81d37e854e25992126501ee59418f34537f31d1f175532894410007dff29b9090c81f3;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf8c5b7f44f774b1123a51a57450106853829eaacc0557f25773b2fb02a179c0905155a8fd3f796a65e0745381bf3c1cd53d55e4d50b2b5e61031a3f9d2d8fb3df4bf0c3b9026dca091b7c8feced644539bf4e0e585f9b677acbe0b51c599643f1a2932ce3a04470b84024ebbe8403f3a5;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8db45d3f1200449811187778380076edf51e7d15cf5c12807c3932d44c73b744b032bac2cacc2648af44fe7da791435b3df949826192a151e484cc8911ca39f4b5ba45f40abc80cf7e346f6262e5ee99e2e183a362dd30f14f229bd3c5205526bb28299e1701c3553b24be99d2d22d6eb;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h507cecfe949ba0ee00442c075c2cf5848d4ba2ad4b2301581300641a0bfea2449012f99fde7ed01ffd4f7f2a569b21443b7de1cffc5ecf64b05604f2347d42a2bf0cb6fae5a1cd758604a1491643d093c03984da0b2077ccec89a68b6b1486e77dab60e3e75aa3f7477c6c64ea8b87bf5;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hee5b22b0e23cf2b92a893983aecd18654ad1079a55799df46f5d35c2b439839c8ede8f710c080b45a6bb28bda837345d7f479ac34df66fd90fb922a052d250045994dba22a243c6dfe181ea05aa65a1a6dba030be69402e495be1c22b77be48fac723e105f542c60645ff507b40310aba;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h80f623de0cba4a61aa6600c91e914f002b2b0185df18b811b7e14619e0ad88a544fa667c57e9d425ca6cec44212a676d3eff7901002c6faacce9dba96e87b4aaa97cc7077af2a5feb5458fc079c4704e564149607f912003ac8fd445aec20dab73cc2e1d5a87dd21491a6945ea9d9d1f6;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2538950d46375df18219b9e52c03e8ce15cf8455dcf4a7fe09a5903e2028355383b5aee39f7e9e5f55a9cfdfcfc70b9364539837a3edbc1648a27cf67b3999fced16f3e586433915369a0b3a05c647dbdb708f632fed320f751e6a5662d25ad6c7002014bcb576078cb848fdc335e5e3d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h16d0d50d4172c4637738d2fb0239d515bb5e0efd3fc2e17bf8b2ffa3b06f972f08dc04fd3dc3adb309d4ec06fd191e57e9bbeee59bc6d159e6dde9a049f9b65abe553e370fb1b5bd5e3cd731e75a40bb361389e99ff245968a31a00b11a9b569967e8f702d68999a318bd200437de155f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdf6262d3d3cb0df8bdb71ee8848ac09c4679c74b482b172b23a08a0144c9fa4d1f888f16f97244ff2ce49d33b65803da867a898d5366a36e9cbbdb06c312b5ac2ed52a276368118381fe267a508881f4f9243f2744e3f1d84ea7ff08cac20043145f8b09c4342e3017232aa30349c29b9;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd49ec86e0474b39458d6af7e17bc6a98759abb334dcaa305c0e978409b2176405881110ffeb616e77c956d28f89dd1b4dfde867d65779cc6f89fb37f16aea9ac82b3bdde51f62873b13c619e8640a7bc61d025e449db4282a239691759f99afdf2dd9c81f2bb271b19fca0e375da9b74d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1cffa444d476ae6a46ebacd8f5fc82d598cf61a6989ac3fa0336f96c6ffa5e71adf93dd3d4c4b3a68f31af658961bb6d8df2e6b969f00496e49882cd713e25059a0c9dc1ee400a9373b3b302a1085d4274a5a84b7cf669626c11cc6e85056967f646c1f4c977eabbf053dccb6d0a4d0c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7f60646471a8d84386529f32165963dae8313f8ff39b2152751c2a9021568cc55e3839ebc42902cfc73ddd024a04a0d35db575727a275680c9282f62a92bc8557b2ebed7f3f3a710d67f711a2fd457697044fad0b5cb0fe1d6ec9d916073dc8e9a6906a286db87f202e755aa19a91ff12;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h98fb988c001cbc1d333c277c0dc0558ff05185a8216796ffe66fc933038cf9979e1faba9b7bfb76708e41b82948b39ed2a5075f10eab63df5a963d87812069b34f7fff273a3d29ff581116a4defe4862a694d81e5b8408e9fdce1af8308f99ec609af501fd15cab8d63794b3cf86965c6;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h50b859e56080bd032a3a9c77fd5fdce9dea23accfadcd74d7755ef7b3e2b5780a39c56e68e63211e7c328330aae505fa5bd1d59b5e3b1271d0b97af21c8e8c4dd50fe29ee060f12ae555f69e22ea7294da8e5514d17b2c312e043e75b908b4bad46fbaa040238456c445ae2165251a309;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h11d70a2a8d336f8df58b0b330adb71108492df47701827e65c64648fb154b0801b95069628ce290a069bde9fbc3aaf28bd089e6caf9c8900ded0676a3070462662d14b228b0cc15f1d99bbc6283abaf247dd417fd58132198e8a061c433199717ce542de523ffa46216ea21483b0004ac;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h872d1e3f14a8d0beed167362a79314c5a9f972364b2e130443e992ffadc57dae40cb1eae60b5e96e89157c66014bfdbffdad5d2e6bb5164b8daa5cb5acbcab61256fd12d7803d075ca3ff9250f67aef6abec7b134c0f035de289a5b6c1efcd5d1ed3c3d1e35d31d844996bb1c1382ba1c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6283c4a5866fa3ff147c4d656c130ee7935080cbb89e132aea6749923acd094ed9ff049d5c5fd96bf8aae6c35dacc3b69298d78074445131d6d1218e734ad2144b65fdaf2663a151169ee4e2d3135b42001cf7d873f5f7f8b9617104215811570f4ad553560d83a1a43294af2ace8cd01;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2b70e5a25b779bba91bf8f74145fc91ff10e07133cb044438382bce332d200413b9dfc87c01cfc83e2c18de2ed34f187b8d5b1f4f47d9f3b467a094ef89f786d79cd3d97fa3cf6a6ba494fd79a624cd328844084ea5ba163626b8d2113d87eeed514566b83fcce96a9332fcf365fa50f4;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7624159ec1a1d3f77363b0e29ada23969cc673c1b4961ec2d5ea88937ac132443bf7831c9ebd6aab8ac7d37f54ffdfb31aa43b67f1ff8ac19e68744aa74e12a6d7953795f114b5e831105c76b77bab98a199b1c85244566b2b2cba22dc44d8d3190f494cd4518566d5ecfac99b22fb77a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc592a8c97700ef54610edc9a9777a59ca8ad6d3c60331b2d45c18846469105256b39140503164c25cffd92371a7f64a207f6f5022588730c09141e85fc93390019bdba45210dc4522b8bf2331f253c4eeeedc295a1f915d6207961a79c340acd9e2a0e52b9397cd2322ff17db998fbe21;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hea1ac3f79c9a2c2b95016e587a92e8425e2fb695c8973288145146788e37342d5a5a0e3c44cc945777e380d63ebc075f11d2ae4d8c76d9c17139a2c37f938a23899ad771abf2c624a48bc3a12c807e3e447d1186ee8e680f579df1283627741bafbad9ade2962a19b1d34c3eadb20b756;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8bcb79a62c9254347fbce819ca56d88eaa919fed6d80f482269ce0e03185db3e374a9ec3b078010a2489287ac5e9f9d823af11fd7418001680bcfd278c16f3a63df4c3a05a817d129f9d3c5ab27f05b5deebb1f60ede8c54a6368eb9847eb469c0671890d3ca8b160396977a197bef9c0;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8248858a3cba944030effe9a5795e2d0871967da479140a3def2484cc9d8df8c4b48de849a36f1d6b4b8a0619856075efc82bd725d22f15eddcaa63f63470b019a8e7d7bef21255a2f623add5b62dde3d85076feea66d4219dba3e27caa1a7a6239e834946039a15477b40733309dfe37;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h49786b3f3fc48392983a77ddc2e796fc9c9a1877b445f15e00840aa534dcc435fd8b29c865c4796404c790ae7e434fcacc7de6486d24346677a859c09d536051b832a9e3219e91febda228423211521fbc868baffce684bf9c2791511c45a195af3be77a2d7e931ed1887403dbe59420b;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf99660857bd15ce02716047cfc40a8403861feca183ad39070846616fe690078857d5df4e0f70b1cac11b84e07a16df10e9e6adee0a6142a179bbfec7772661e32c75919d23f05bf9b71879e2c8c92f442e72fdc67a9ccd44393fad2ee9964f51809f3ae177fae9f5356cb52248cdcad0;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8f151ef47d383d09e71358b76902d419875b3733caece1eb46890896255806a71f7652a9b4083383484e3d7ccd6e535a3316d2f147e77b11959cedf4a11971502f73f9825df8ffdebee485abefea3607038e6466d226a6ab9e46fc555de4cd632edacc34dbd4afb2476efc87e99aad0ed;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5d64d1ed709d07a42553cf6ee4176459cc4ff5c4d4e304b4a5919a1f726bee08cc3c3953dbb13f547190ae884b5ea5659ced422a59ba980b562738d04f871915ee42eb72927aebc8308c1ecf4752f19020dde75f3f687021d5e4b98689f7e1b874c36704c88d45e19db99c93eb421ba;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h419e52b9c7572975ff65ded0eaec47c807a4f8d54245ee0e84ccad444fae5114741c3953787bb69a2681138a14bd9d242fc8a15ffb8b8ee18f8eb9d16f7e93df351c59d24bd76ce53d40012dae6740fcead7d567d8c8f63cb195f8b3268fda7cfa32afdc15f32d1de2f7534038a170b0;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h281be1ddaf3c84d5c13d2a3539ea9b31e29a3f616cb411fdf78ef69f7129e644fcc28f2380464dfbcb738f3be4159ac5b95642dbbed5fe60d6f6c25441b25262ac63c5389f5bd60f655c6b352bafdc1e55b73e05cf6f56b0338fc3995dc6cb0630bfb1fea91de8e864475170f717497d8;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4eff796b03ea52a6377fc157e137bb2ce74805545ec2b8e3e3a36b6075cbceaf49a836d3bec62e653cb1a4538b1f880826df83e596fd808dd240f0876756d6ef5a25140db1347370dabe9c67368192473b27e4a0c8745261dbb2df964653e4254087ee6c3fe24f7c21dac4e463a350c5c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h61115a97098f620aab2ffce8f91016e84831212a9790e0dd59855d1be751510f1f22e5fb7895d4724e147f63f2675e19e2a8232622686ecadddd797beaca67e8af9c589a75c947e5268f22dd4fdb5ce5f782bdcf8ded1d28951bf9e208bcb515a3ff8d073e0cd075d0dc2e9ee7ffe9dd1;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha7d58102d7e9be71e8fe61a6303807c6aab7a91ffa53b46e8e0d7f2ce8a900e16cf8c9478aeb2c6aa7c5b56181020122baac3353658f342e808bd72907dfe7846451f17886667082d9b9c4c8ad2c7a4a2f4f5ae24940bf26c8eeb6ac7844b8663b32f742ee020c564e4616a30da6df066;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd09c106a64bbf6653f2f561cc4552fc60665af3022353f2e7dafa704d0677bca10758fdd484a8ac2e514faee70b2eeddecc800a315d802782e3cafbba350d0a36552b9193c415d773f345b2272ed38c52c6e6359b3efa88922ec9d0c3584bd189eec38f977c08847b324e33def4c5a153;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h59af3ce8a92cf230a98f8a18aab7a77cb54534e988fb5f24bbb0c2451893bbe3b7de0c054d21de634fca0fb289942390f28439e6f35c130ee5427dd43c18c013cd6a98ae6ee344d9cbcaab0c3aae94afb11d3a437c72ec0edaf3800f202f1e146b4bf970e651251d597c5ee4695bfd6bb;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5f1fb202e766539ef2c4b8e21e0a9558d98ec35fb4c7c69337db2cf04a7c3895a8fed488d020adc3fd22f34b40626affbe838083e6ce178e4ba8ae0805d2d6ff467ade5aba54a3ba4b63eb00085c71c692d1f8d3c2a76f6e3a3d87b961f3166f81cfc9db698ac06048620e1b242e2ad84;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h542ddc2bcf160b96e65e54250ae2787428a7634033b81d05c612766b0c8cf9177e823bd60c276211b04a379d48ff283ad1e511358023f03d6a46451eb9275835972d4dbc600a9e420ec9ef91889893606eb90ac0a067576e3882b6733b9e273c3ddef6fcab196bb4bcc78b1818a50e041;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'heeb50826e051bc44616070abd9dc3f2c881fae00afabc141e9318b97a6ea747f1e2ec881c9d1c33ad74812de27c3bcc53445ec22968abcfb60755def65fc6441c4b9c08df92ff2acb05ae2e75b5df79149f8ff3e9b4ddf8a2ec60705e7b29bba6d5121d532e71bbc1ccfe686038789d60;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h60c488c77ef0779ff9b9f48b6dcefc37c79101c839b557afade8938ab1abd1ec588568be76e1e91df2452f634fc21f3ad6b8203136c6159ea9fc28d150477b7b248ff3a4c9597b51a5c4f20ccf56ce8635f3cb10ad460f6919da3ae1d2d8aa0cf0ca5a844af2418bc235247c5a59d7908;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h803c51e5497b1ba5d5016603da27e89258d7f80bf0efd4cf3d15fe37767b37f1c67d9a201af0e49c4bda295c1d41b3add0cfe9247b49646eabb3f1dc2b2929741772f607b04641b78ed42cceec4050a1ce8c0fb8d2948904eefffc2d375bcfc7e622debea96475d5d4fb1ee1aa16b57db;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h315a6a55262669873e29c1addc2f9ec4051fd61ebf94610e9811741cb82b1a2a736ef16eca316c8d4c58da13eaa2012885de50fc83b3cf395ddc976fe81950c1d69c5e1ebbccd09f0fb98a46ba2cfddc74855033ac2468c43405aee471ebb46318eeb7c585512f5f35fade87d6d8a3380;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb2430a1c94a9fb203c5eca50955763e047c120947280b999f564155c636d2a7f054912da695965aa8a229da63c760c547e712405f6148369466efae378a67885502204151c77f4f09f4d8b55e5ae596c56ef0ff97c4f747c3697811dd122c3489a69b010a0e00c302d70c8c2a1ba2d4f3;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h973001f134c7b66ec956803097553aa9b29252a7f0e9e8b01adfbbc19fb30e0cb594d8c4b2949149edc09129d55695ea9096984f404ad2e50723a3fb4e954b9d85bc5305eb033f0024c6bf416f28e289df0dad5c9fbd4b039e93706e95eaba6c2fc7cbb47c5c2886b761650917740f6fa;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h499ac7906385f0dbd2f4aa0ffeb821e09c148a0d7f5d7ce75be865451784d6c8d3aab9c42d670469fc5990f1765bf07fad138f469a73ccb115932d43c7dd059b5d225b95b5ccaaae3deef3f88228715a75c30ffd6586bab57c3a368d90a1ee663419385e77ebfd27bc8ce7ca6248325f9;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he02318a7761d3c4a0d7f2d5aacda27cbb0b71e3ac9f08620ae52ed83420c209663e2a32b3978ea573d5ecfedd045be5544f2003b41a911c16f3384e1742ec91daa5183a95c5f4c04cf7f28179c851187fe26bdd354deeb2e6a272205886a2c71d008cdff446d6cf35ce358ba1e29344f4;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd0494c60552e6e8c3f43005507147e789136eb81a916182d90c0ea339cc7fd28b7412c308d6ebd810450306d4289a4e5269c058ee70f3b470d5f3db91790ff219e72ba86be00eae3038eb32ad77f4100832934d77967775471d628ebd53d2684c3044716cf4245588ea99d00269269d8b;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'haaa71313869f857382aa4307fb5d7d3d71a15e4365ba67c532c9c57a4c8fcf8b1ddb6641bf74d579620818550bf562c5232740542a32b50d620531231dd8301eda43108b4b65413aa3d79ba8ede74918e551ac6485fd0cf8ccea42c419512f5573e5d8543c3f822f8b7aee7fdb561c5b8;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h73240f6b498080a4aff4cd21614da4a94e9643164292a1c3d839b59fbb40b95cfe09dd5393045f37e1a13f2ec05b4b91d399f703fae13ffee2baa015b79b3a06c1371385d9aca6991335fa22d822811adf28d3eec31de99d8dab9941163d40940874cad2760ff71cbf2f2a52f31be0592;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6f49b467f1c6dd9bfd5bed4bf1dd28b9baf6751cb79e60643ce9a8ab48da97a6b640e3cd7356f3233a0aa94e0e38b58314ad8d4d50610fe9943fc5e24ec072fa9a49084e422e474218f47848b0e1311f1aebcad3dde824810c3df6c0479c6f08879a625503d1cd302b3d6bcbbdbd51f0f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7bc1695d8b9211c8832a499839adabc4cacf304b364cff8bc37754ea9cd9c192567a1e9543b64df8df2f02f8e8e9cef2c6b889def6405c0c69c85d1e13a7157c8f83b8375ccb4646c3fc7fc93d76a0b65e67f39d166dad9e2ab42a22e71c75349d7820ee5f096422764c2079834749d33;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'heaa5fe132212556af06f8c25c35e509afb1a50de359f4de85a03a4f0c101df74633f0609498fd9ce0a2f5c1917a29a19d8c5de620ed5e8937daaee7b7ca7f925d089b64518659a032e55315f37331cabc1d546d0e972d454340647cc93678585664794ecfcdaa221570b586c2dd5e0f2d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he288cddeaa9c4edb8aab2af64811cf269b7122fbf4687f2f8dcf9ec6669af5b5981c835744c96bb4f3ea1f5e3b9cc5d81814682093f16c4f98f40930c47ed68ae6d77678a6d7f0f782b80c7c28634536b41feefd7d9979a6fd9cccbe12d22bb6f26a94b443f254823bb5376a15ab7058e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'haf47e457c7b1cc2147b616d9b4ca64532cbea22998b9f45c26a4a3dee3a53cd2203869815b75f7d55c6ef58f368ddcbeaa6635f4d5b4acbbc5b66b39ad777dfe11f5c8e515b59392ae479cc375dcec5e383c35891dd7ddb6784afc17c371d8ea08f6368ec0d6626b3806d00e885bde106;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h838606aaa68c991a5e4630c79be7dd0c84b64ef6f34fbcf5f4f524f4a8249757ff8cf44e2a33f795ab04922ff3c03d67d193a2c5339e181a53efdce2434c6e44f4f626586cef5ccb42908a3c8b204f7f3a165855aaf93b52c04a5acea068cee1d8a8dfd4367f506350c2be3f0ebecca7d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1beb05a6c3f083a752649e1a34c4554280dd03857bacb91b8b5da55e37d2f865fc00657ddd87c7c6000b642860452da3cdff4f2135f98564cc69eea7d8c85874bad9e42921c21a2d12d879eebd5538710bc8c609192975a0b7a819d51263b9c729509ceec8b2ffcf93348a7b59fb3320e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6559033f88a3e414550a4222a879aa9a4d4a96248ed27db9342cde0f10fe2d4e5cdba5479b9558b36945cde3ab2705dc92b3fd940b92649ac02447938a60d1495dca81a5e88f2064bdd27ce59eca5ced710ee4d14e8864ccbe62c8134a8cbf512d05405d21c3d1b0658f60caf919de3dc;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h58016030fd59506800f07a210042546a6a3888807bf51a3a79e71147cb96d377ea426e695bacaebdcc73d4421144e3f0255e08818321cffa936c43c7debc1c506e5169b0b71dc7b10ca4fbcb8c2e1b15c12f0bdd2e47782c7cd5035f1a481cd647d67c2101ee175db86221ce276289d59;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7c5a8394a090dd8cbc541500991c133f58efa3a6987ee7e02d66c391cdafe529a121da0759e0f8c4a55dc61f4bd3582be07b3bf7ad8f90aa256502c9b452485fdfbdc9c113094be050cfb56ad580301a0da374b40db9ffbea80c295a56da4c07718d8a882136f4f50bf8461bcda7a001e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h80a243d658ade9533bf47cb8ca033af904368a98c878427544e586ab5b16903d4254102c5313c01505ca6f2aeb8942655b249f5185c1ee38a8937f4dc094e622c22a2ebcccd2fb5209f9843aff041915b57b97c1c9e10661cf55cd695e569549699f1c0fca0d3a1f0ca76e523c1071683;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hac65ff4410be5ef91581cd06c8a0e411fbcdfe13743a4faff325299ad60af6f72235fcfe582de690fa07761fdc7761a559354284c1645e9b4b7df8d4a1ac0cc06addf2d016a1ae1e20598641b861aa5b682380445f00beabe815895af8c29ae212b9fae32531f1219e85bd9b69471cc8c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb4c404363ef505140847713ece91ad46d0acd85fd51cc93631c1d514c4bb66562763486bd0fd833c08c77015d223e27dce5da285a3dc94c197f9ebb2ef5284f703040d0fbbd361c3461b74b56e3de78b314648fa2b514dbdcbffe6f3eb1a28004b9e658abe5e54d304727171307c1e832;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hab90537f3fa341cda0ca6ed5f2cfda926faf900a3e6fa23011e6499ff800ee139f62086bb9787d7aa47b432d60e62e5d756b2839422d13898a10b8d5fd9178b2a5b97a80d327763aa18d3651f0d3583cbee11afad4de07cde434a6e3271d6fb45353edd5bdab82586eeae520fadc6c515;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc9c6fc6b46635993b3df8c0584be42e4212a7cf2136942583ec432af69d5fee66eff75ef366af568959a22bc9486df113a1d573d13f48e7866a0013dda06d17898a196166db10f22e9c3ba3b9541ee9ced5761fe76b7b7f7c06a237cb83ba89688641b32567adfd42a7715e8c6fac6d1;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc7aca094610a9ee24757a0474b984c521496fd4b5d73b547d6cb4a2d80e5da001c295da9ff36c4e1ad250d41118fab0335b12920fdda6cf9c5684f942034c7b18460f6903a1edbb89d1555c9cf0834eaf5061f64777af29f5bfb05b4e918ee97ebe70e20767dafba35119c8dc7269562d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h62c76287d5627964d21321bb348cd1df8e60c3a380a403be1cd933f7b8d9200998af59dfe5f2c8493f4a73538f791f2298588edd6791a6273e40d20795951d06bb09113b232d82ecf9f9ffca9fd2ac0da60b425c93c87a9d57deb2bbc49c80e68fb262dc5e4165608c7eb51fa1812ee72;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4f662360b83631504b2564304a435de258b024412f5049ef78d813ea6ad1b32e4e998327efd05c107202b98a589a752c96c70fafe1b1564a79354353826de383e472e3322ee9664c18338673f84ec5a485de9dd3a2c44e0de47f4d323b9c373298860247ac28650d10ece751600c78fd0;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hea975d8283cbce4193dc496df98c2f7e34f9f40e3dd33e71d31bf61c0fd56adf4c594d8422ef4cd0a8bb20e50b5f54d662add3abeca283d73597b6d08dae76fb880d93afeff3b636dc394fdfdc88a2946e1ef5c827d220eecad00b3c1ef9668890fc739af30b5f4e33123e9ebf22194bc;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb96d6ddf437fd0a3e7e29248a34dad34c9a99005a4f51c0a5ba4b2dc0f3770af801f2fe0ff1352a42b5a6f7bc51321f82bf95324c634151b85787248e51ce0d7001a57a5278bca5651032d1ab47c2cf774cdb2dbf11786ae6693b28ff431239a763633e9efd58fbcb12193f22c4681232;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h54660a897640cf514e2dd7adee6c55cfdc37099d505588039084c22b6e01e3a7da8a2fa5b8f822337585c42a9f6a1f0ccd67c684f462aee2ae0cc536476f4ae4018268807cc72107d1c06c3f57c20839bfcdc8e75e7923af18c291d573005ee45e9adc92d5041c6b6284b82717442fdb0;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfcab158e8efacbba1ed7c51fdfe7bdd946ad865c6418cceef5c0377f33e9d47099ae32004b33333cc516de140fe75b1da946b450004d4b2bf9ffd64155d346fdf4a3e6dcd689ab32a9a8b6b27ccb649c217728be1879d83a50ef4f85d504808ae4c0f5525b6f23f26c1fe7e09f1ecd772;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc638cb68f0996d006727102ca11adda9afa03e96d8e58366fa21891ad3f5e9bee5eb6d2a59b36d830f7a4ab8bb7d6c4ef4d5f22c42b788edd3898b9ca48ca78a0b5df074d4872beb1078b18a9c5442469f15b254ab63317c4497a2e452f08eb4ea2cbcbbd87bdaf415157cdc5206de0fb;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7f4c4d94a1ba5f8151ee86b8dec5c1364017b6d2b2950192330d99067752628c4d5d22f65e8c4aac66b972b17f8884613f8e87414933e168f56a7a2d4bd6266ae8c239eec6ddc3e79cf434e793bc64637989f6412aa730ff68e6067ae27f575bc42fe3b2150e831b27807aabe5df22f69;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc067de6d0e89e4755deec18482ea9209594db221c9fb8a6b7b4060e4e2f7f03f46ab91b55f1977dce09c30161b6d220b0aaa0be564e708c13548fbc007de3678e599c2db93f5835b1a2ef88f01a1337f316eeb51db779655a2478d4163ff867c3c156473bbd0ad374bd827d0f5206e6a4;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8d5cc7834989058c5d9654bb2b43ebae265d614970bef5047d24efd8ebd1e39b5e8b649704f77f368e5b37b4c3266a022f25762741622a2cb62cc959b7d97f4dcd4cdbb3ae6462671838cb1942b93ffaed739c957b5d4e5c205127d135f5e3df5a7efdf58d84cb7e44973fa3288629878;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4a5402d529532024b458c29a0b77c766390174a853843b51de029ef74ba869a34141bc46448c589db3cbcaec0dd40520d5ff810542faf6ed89562a834225fb5e2814cb6e31de0b92e32f833aae8bc77c8d80890426f071f3cfecb4f5463d21bb90ade80f0598a75b4a818cfe3c93dad7f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h21b9616f8546996772175eb163cd615ebd5f5b52243e7cdb78ebdd1fbfa1296aaac497693bf905653d2289d04a175dfbc2f4f14bd121cf1fe11150c017909ffa02c65405daf6b1bb168bbf6719a65221d3a61a4cb62e7295723b0dbe7fd28a61e2980b05d3e56d5c1365cccbcb107437e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he5db6bc407495ceaf3ebf885f2b9763679582dc1fb8f08be8b8fc75569cc25fe30c3fae06f66d62ebeaa788c21116edb1e01d2a39954e3d35ffbf75884163c1f37858978590dbd1eadd7cf0534f53cbae0af84bd71f72ec8bdb2f3fd81f254b3998727276ad86c140a8a34da5229d0b8d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdde908acbbba9dcb7dcdb32deed5740b34073197ae179a920149abc4418c722f98f0aa0d6da668405c6b5dc2ba35ab023c247f2cacc22fe5199b3b73f2ed66b292bb65665b09b5421eadfc41df32956fc6637e2bafbb95e3f6a71033b150e0620ee779f5a9f4835509d13cb919c103a51;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hcc758a8bee45f75572fd767bdfab37ce57b11b492e674cc5d77c5a7ffa87fc87b5919463398be280322897813610e953413dcd8c8c6f5ea7b811692945d734890721b60a0551cc50cc7ba60f62d9f242c86589b45b10f5bdaa94ee45230e5b850626df088b0ac86d1900fb037e4efce54;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h669f2c69954d305eda62a15e06300c942581894805cd468608b530429fa625664eb6508356c1ad51b02d6c90a6260f5a2eff38b49323076cd89887afc23cbe1fd27120c076f1f30f70a122c97308e66c95f90cb6cccc589b8b468951cbb7f157e4d24d4eb85787302b310dce12633e956;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hcb29c1265bb067958056bc9450040ccd40c44b96039e79e4bf4fcef18a6fd355b8acb2de11ae7679c5ca462dc90fedf791ccf54fd7ef2416ee3438965639825f0f1553ca370844fb4e0ab8a3c1000c4712afe027b25523c2b6e84e949bf676ae529065a0a60cd1e3b024b6780bb08157e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8f4533605e18ede3785da3d4a17be60d4eb38a8abbb62ccd917d24543390818bec3db2468b72aa2b96f04eab712805f4e0a99a1384af525da77a909d18555b9ea0b67dc65aeb26ee7ef11d6ede6036adca6a64f124583a11defdff601b398fc4ef4b307ccfe138288cbfb2f9c42c95112;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc8e62422031f757066d84ee27b806df3ba67861ceb4c5002ab54a829c2284f56a6ee71a828e945734eb0aef04d1de3f47144a5755462ee3eaf2fa68e959cb7cb77f84256a477a55ae9c8defa76db9067a6c62f1dd4f650dc67c4a47252898cfb19b2bfa8f16129cca2d9779a7f007f1bb;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha504765b1a1964688875b3eb0004158b698bce1162185319c5716764e73c3393885b7a1bf568df3ec902a0292b158729c6c5d8979cdfe35f3b41c3da32bc511ed9f71da11f2f7e010bc0e836183182316600284fcfcb4080348e8255abdde959b69574043fce106f8309ca858f23bc423;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7aeb42aabaa16385e556006a72d5138707d5daba41b5a6ba0313b65e2fe6c09d365639f3cd79f1875fafcb7c12c1625f2e60e25f9ff7ae55fb5b56e2cc972ca77cee38df9d3684c06a1e1cba7454baeb80c9a5e0ab2bf8c6c5d7e57364ef48dda2c01b4cb77f698f30442eb542ba93488;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfcc385bf8932333ddbd914526bd98927a8f4faafe9d9daff2f364c998f50ce8f3a373891a8d0532c8a85b5af0ec154b3007a0e5409e166c870140dbae9d25575d1a3f1dd8333d66fb490a21203c5b298c45c96ff9365f3c1e4def957cc34b1762ea87a9673900add3d35532b4b86f75b7;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h76b31d93fcd15dcb8e8252f93eb90bdf5e5a883c812e9a5d14fa2b69ceefcb8bdfe32db442748eb5121f49a9fe56de8ce091d3f09b9fc6c30070c8a58174a94b035cb9d353dc3346d4051e45c3fda41412ed80d42f58a6d4e4d11f67900f36f405c0d12f1c239911e0c88a7574d507bf7;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdf07b621a453d6bc630bad971ac604762c1d7b0a44669d36045267e92bc063b30a021053e8d5ca7e46e3a46cb26dede539dcad2eccfa3e88c5fe98486d37536d3cd099f78dc79bcb19620427eb25bef81c1c6333b76ed910f47bc0a956a706a299e165aad8675c26f46c0484132ce3fd1;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h878a5c4a63307bc38cc554c61b2bad2d5ef176254125a46c827502d5104dfa7eae0e46cc9d3af7e84178d80303a435c66f552b6157c512373438ff78acfa881fe8aab5ab1a06d3509b7354fe33ef5e03dc0f46de542d11f0eb0e4eb273dfdcf01c817a556b6a9ff2a91e3f70dadd12ff;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha36bbdb45fa30aecc923bc08e6a2fb92a0148fd52cc132f76286af4ac7eb3a4e2141298b1c5745a5cede8146d98c26c7a444a02b9a2a8d392a1d275e4914a3e1c53cd16353201f45fb4d7fff8883233d715a0399e529a69d66d68ef5e95a33fced030c464ab36828dd4b80bfabca39cd7;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc3f88d10c538dbcdf0b14667e3416db052eda52e6dba1d08b6e7c40ed2353e4a781cb815ff1176ac2189d6ed13e330fdd77c6eca3b5f5296e58ac2a4f35c7a378dc7800cea1dbcef807a5ca52ee47a5e3be3497d099db494fdbbbec5602c9e7e7a4edea9fc383fa8f2e95fa5c36b9982a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h91a7f914d8781593569f7ee0f430027b01bf16fae0e590583eb807b45bd3e06cae1c8f02a0f2148329664dada7b58fec1e78623557a7d55691d1a21561e23aada4f8fa01dd55de7f0d716c879f328b148ba97d0ceaf54d88a4a25bac9937dba394172f6853a36de742462b903961304c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hebba51312e2615528b31fc8cdefb1640444ac032781826aa2e84635c70d5171b1e64d2abf64119971623d7448175bf6effd9a9e24df89a3f41671cad4ac93c3d67a63ac80fa7de58634e052183d3bb843bd3f23dda0d0bca397fca2711f2ae8d522cccdc70b3b9fb23e591e8046c7161e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha1429b3189c108bb54628ff34e9873b65ec0c51faca26085055bf73d4ece61c04fd584c9d653154c1f595c7cb1a9e13726dab07ff9a4077d1fce2ab5b350ea32194768f5b020038e6924e843e78b58d2b5f5ad386b094fc6d0e7053b818c28e30e820759dbad2e6dd6c805b47b2bbeba3;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2e7af2c6d28f5d7101879f5d32ed7ded05d3ee13e691f6eaf3b7c9864e70cae83b27ab51382765af145a3ab09a194b95abb4dc53d670a73006c986ac691f84672652063449c5875a346b52adba06264f620cc3d21f523038f6affbb046248b872715be93399e079b75f9584421eaa31e3;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfb901dd7f8bf2647d8aec53850b25f2f1206f4401c9986a489a8c319076f863d746923f65d753c4e3e417f2da7c349dc6cf3f08e901d2963f888227c913fb1fd6ae1f89b21bc34878b150d8f60ff3b5b53a410b41e619199711da16300ade8131954cb783687a8bd230943288a24e42f4;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4098844b5322c9221a5ad0466b41e1abf1cb180ba1cae2c8e5e501441917d1bf1bf2f47c07a1b2b7e5064e3ad51693a4b650c0579940f0fbb99c1bf789d3fc4e7baa88be88980cc6114507a8570c793818ba66230c8a1f8cc6c7abc3ede037044b34baf33859bb06bfd829b38455461bc;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h591b76fcab209d0b7e00c8f90236cedbfb6b39f255380ab44c75e19c27860a8367c649c3b2eee66a7138b0ac0806e3ea6f5c2f61c72033bd71080e51644d475e174e740b2dd678ef0e7a7a8c1d6c3ecf6f8e926ee60760871f8eeadb107135981f7e632bd976c60a770475a95e9f9860;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h57d02cc67af16efc722e139c12c39ed7e06fdf35a1a6f97564e414ad11b8fcb3d1ad057a58ca4350b6111cf71c90229827b5af92e62421565a7b4e04bdc6f3043189ee8efc5b4e187ce61abdb011604742df4c10462546d23e6d1bf4906b3adf7d709dde43d664bba8e1f6583f5a586bc;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1bfc63185dc0cf2c663c83b08ca2858aad9ce8fd22c4e9d6a236a569b37be35fd1d21c975a8dea8402533120fb7b1a3b6745d59d311faf58baf3d57e8075c60822b607c66b29502d28b980e5a53e4641ea7e5eb9d81250143362c02224eb15d7f4af8c401ee98dd531a37ea43b0393a2;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h80a6db5ccd18dfb61593ddefbd5f9c769ee70bf0b47537e76b8ba7b3c3e1aa04740484f2079b22a3618e53f2f5f6afc1e81e2fc396b3c9988e3934199743fd1f7941b30f1c8581e9b422ccd17537efb6a899dbf59620072fe5f1fdae1c33db63d6f4e1006a3466d754cf57f3c3be8934;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8b2a099c5defcc7265eb9fca3e7a1b7231af2582ab0de9f34f10de2eea2f4f1512b6d05d11e2a8648b24fbbbbf75f13a1d2d89368721c323e1f050b95e5b5663aff3e8604fcf9f988cfbfa80a98960ab6b3153578642bef400ef32948096bad9bed43824ddaba182166bc750c64dc6053;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc8bac58c31abb30ed63e21ba041fa4f015164970f606425fd257dfc46870c5b6ea36d0dab449362b1084ac44417741bbb2683650efc1288e2e25a545e7ace2e48606bc859f9450cb4de80bc7bbe8236a0ed886ebdcda70f3126e8a86b6de242cfd041be03a47f4522f2b9e8b774d2e4f5;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9f123aa28256f48dcebc2ff412b1d4f0b521a797d246d888e5ae4155290966bff64860fb30c1040019ca9a19f2f11d63ac98b31db94aa90c79810c7048b0f1874802ae7367b5ab8bb8eaa9700fe656ef95bf7e2a0a7e80a0d7a282d9d4b19ad861ef7c85f0b9a47887b06b9f403fc8b1d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h928c84a76edbec842c56efe6c87539320242aa320fea8e5225714b5c568051d3c8ec6e1a67f8a5e502b27fd678c9d802c096fef72204cc0c1106787d03a47ad0f823431c73d917209d8b02090d996549b4fca2f20c2daed4f28e74d941c1824cb09ede6bf111e226f0c967cefa2befec1;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hff004665a32e0ac996d1a553c2772736d9a5cf29affe18f6e4f06aec2740f45b1e4de2f1ce458d230be60918e13fe8fc1dd87cddfd337ef906ee0e83c877b14e0cadd6857a471c74975f3f94d2c9f5b012348390976f6ce6e4597a8c6e0a9a62141e1de1e556d05cdb0b900a16a10b6f4;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h17d3884e93922ba85278498bca69391da0cefadae2a82ced353910fda341548e4877d0bda001e333bc20a50afbc83acf30283bffd853b38e4ee237d8bdaab39853c7e8ad729928e83ea760cf58de8f20b6185723144b2d0d3307cf4feab483e63b208c6526f5669c02180a50718872ac5;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8a6fd4ace0b42c350aa9fd4a5ccca4cfbd402ec621d6ed280d74d21bd324b5d41114ed0bf294cf773bb7090ebdba5136912880da96b58de70b07f9d3b4aa3f2005731e3d1ccf0387c7e4dc409c1b9dff377f809804aa94bdd0c2e94200de88eefafb3b7978a80d1335a37d11698ed7402;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd4b546ad050b007e4a005bc847c5ff0827dab8c630b8ca3a993a308fce75520f4278878245bfb201e778985aef4da6fcd6091e294d49c7eefc1d2229133691f5557bf0b0398c7ade4a472db6fabc7bf926a3e181dcf96ae3e11ffe89317e747dd577df481d136dd2e7a1c3e4400539661;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha0950b5fefc56b3c6cd8cacc72a3eea27fae343196aeb2253bf5375c31519a313997b119490391dad48baa361be011d00d1fa2cb0c9895b1f80a3e307b4680860739819394a1c4e6c44159fd87491a748e04234defd32539a26986f09512906af8ed66068afee2c087f7e83d7b5880f7e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfb6ab62fc49943002e6ea26c09bf921bcc4d7d987b3bfd34e067e9a6b8ab698f9d3c1e9b12dcae02b1ebf126a8e779dc452fc561158b65520767df491192d893e5762859ec82f7ac2c4098bb6588729f09746a2aa6e4f80e6213ae76da3c380c5ed974359bdbda9516ce1ac80cdab3159;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h31bb278211e9d50928183961d5e364f3027b73e038a48641a6614176b61917f14611cce8c2e33880752408b73eb59558fdce28d78067d3d4b7746fd8e9f2b79a0a8b77105e262b1765dfd54ef9d3f5709a4357b1eafa343397ad2f4abe268f8f1cf4520c645bfa6f39d506890558c1d9f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf42c7e05852af110ff7fafd0a28a63c320ac61147beb2a64f1a0b338113e166dc3b111c126b5a96979604ed7d8736453795c2f34263640d61c1b7509ac3a276d844eed5f8cf105c6ad569718b0bc10d8665adfeff687a78fe5790c13c5635d36f89bcf709ef0fe590caa08cec6809664e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4fa827ad0a5239278b1b26f45254999d42264a74fbb2dde1ec4adf2b65f9e8a5e320af59f9bc3c37e3f8f6d61a5f988aa799c3aba90e32390b2498ad32e6e5c96b1ccbc0592994976eeb557cd254db5bda8d9b76e4d5d8c04f700ba9f7aaeb05c8880e943f34360574e7ef7c4f54ccfa7;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4ed9706de588fe9449c7ba9f569c486828875c5308b0bf26e9cb6227c5000ae0b1e37a85d41001d882bdd1e1463358a61669db89dd192f5ef7fd31ba4d7bac9b7025eec3f7b104a124600106d3d0d2292275b03a7766a6030e21b61e783917a43adf3f993e2e1de5e81ec674d3119174b;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h686342a588558949c9c8328ddbe04305e4ffab709b735c30801c3bb735edae0acfb6f78c130f90b499834271fafbd1dd0321ef41d1d70456c4194199c51a45f154c9f773d43cee82f678e54e59e5054cbe2f1e40d54b503b25e0a19cf1c537c494f251a81bb7766f76d6f714f5809c4b2;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he8088373799d77cf078eecac604d5029b969de49f90fbda62b6acacdb6a8c7e2a6fc34cebef85ccd0a8e056d244d0ab4574f69eb447280f1c1b0ed05873049acf28191d0f4a2e463f0e720e50fa49958be886998025ce6c1a588b1f1539426e1542685ccf2662010011bb64a01bde3c37;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4bca9f7297932b2f3c46dcd4c4263b0693879471bf110ef7e58b41c1a26f025034dd3e52781643c78f5420f8d0f3b695fa50050d19ccbce0604e67e1808c7b1e92ee9e148bcfce345bbd23daa38b97a655d54cbe844dc941727a39e8809870f0a49cffa03eeca6af5a9d8200c96fe080e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h57d93e5411b729987b7bef2da0f3bef0286366762d7430f0c21199f981e7783a47877bd473b7114995b7dd0526f4fe4ccdbc5095c12918e2a409d98fc10e257cbd58970efcfa2d95c8bd0d878467e85d77293dd6d096f52f2ce123175f3d6a13b80f0bfa686d0e7267335fbc6493c0569;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h434f29b0876aff6508dce6f422e634535e68b9aa35b7de83180a89b208cdfbbf561e981140f59add5960cf20284f87aef3f006815416e381e52d7d2166d5fa3ab0bb1aaff787335f6c9755890366802459aa80f517e75320ca8127f8fe2e8886e38d73ea6034617fb8916b3c8963f2861;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hcf91bef8f739d2fef208865315516496f99706ee686bf25223bb4c9eea08d89dcf66c8d8054586d12844de7d97271dc37e84481e236ceabc668bac35fdba7eff2561487e911b78f9fc3459efe16b7e0851d4e106e092ea81da25e55219026769283993ba71f03aa23d81f6c24490d2f67;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf94bfac01e4282cdc25d7dfcd3d3aa524a28935de6e27a22d1b2c4381f811fe9dd9ef339b3d0fd6ef42618e3b9bba919cf0bccb9425f3b91c92496a8565c65a90de8e66c5c828821f08da7b2f8c25fad11ef9f2fef0407b47112dac3297f6a91e66c4ab181b9c50d655befbf4fd8e46d1;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h68929fb025efa4ab86d13cd383054c4258de139c242712240e33c06a44bc1fb96009d24512a7f95b374376b4b4edd01c777e7ca232bbbc7944084597823f802b38fea8b940a9888470bee5bcd1482021df1a0ae409a85cc239595bf4d924742471e84714eb38eb3a0c53ac1350fd40f6;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hcaa8e3ee735e26ee72eb01116dd125927ca31958ff501f42c16abad506bba1e3af164184bbe30d814e3bef36b9d024bec3d04192013186266c867044d894a272fa3dc561aa0e5116071e857fae3ecb96a6355411e2b6cb88957238a96663aac1c0ed43ae43e12cd272631fd2c5bea74f9;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h27e1cf0e68b40165cdbdb028b2d57a2005fa1b412447866d85d8bb0fa060c746a57fd5c0d4c6422e5a7aa42a1dc1c320c9b131f82f559e570d79dc99e928b8728afef2b99fa77d0fe1f8a2d19983c8b26818dea5cc63b046ef5c87ee53439a409481212c14f8b74cbc084d158ce886bca;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h51dc5c25250a827e5fdd3518178bac1a0138f33dc24c0b2e91ec954b14fcca349d88bd066dda5b743147099304169efc74245258578200d68496c2f0743ff50353b6753d6a49e636607f7037e9743a37f9598dd0087f7f5ea248e55df7861efa0386235a905ffbb7b2fedb8ed12f26c3;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h22a12128b124b9f0a6a693e805f8f8988e4179bb58074b7bd0108a0d81ae5e33a0256ee6f3e8d25382dd2ea63b56a408bbc4366daaf34dd3d0d12e07db248587058d20f9f1f0d8ee1181f5204b86fbdd69c07be5fe304ee4454e982a8961ab3bfec3142e900c3a588915de15d20f7182b;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha6d62f5b5adc5773a622b4108e8c8385aa63297f5f022fbd55be91f8ac422d5eee9b0fdbb203ae2480315142be6c1e3eebc7b574a1f9bb8cdde9e989e25de854ac88d82cbe614a1668cf7011ea89c0dcdbb72f957c2dfff37eed18174f2d8a1d90776ad03f32e352871ac04c1f10f8cc4;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9ab29d64dee558f65c94ff358ae23a06f23acfda6993aec16bfd98e96e0dc135f4d6b4028ce89397998475c991cef26a0d32a269f6892e761d1bdd505428a7ea8d0024e16b68af78e3028970762347133c31a7d3d71b00c45a25926d7bf5908526f90f08d4530e41b4c8b7b8142f5e67;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5cb8537c00799c6bfcd7931a160de1805c508ff5beb8ea1ca2133db7742207f6fe2b74bf6269e448aabb81d86438fffd094df67eff6b35bad0d6e9119e8803d6583c3c28aa7c2213388325ddd8dc705ae82be00cf4fd945c03bfa2c3817ed8192cdd341fca2c6a81d9bd8f0e5920a161d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8eff9bb1f60702d110cbbd6a4860f4c137bad73d5a596820c840cb56189af1a5b0f9a2d74fea402b9255a574bf6d490d109761f0898a605aad6c595384c89e2bd7c4dedeb0631784b04f3353da77f0538702ff6d3aa165ec65f019432bc2706f2000cc02c4bdcc5f24e473df75018841;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3e8157d388d64b2d61bf3333f44a33902f331efdba68733dc20a71e610ec1f3d72072cbe13251928dad545928de1010e822f6ce30af6c4ec897b7161edc54c131c5f2d408517687de4c5ffc63f1ae3a47a721a29d8b2536c5dddca8c3c8028fcb81bd1328d324a6fd96bad3da9b7c8a42;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h46b3d9dc0c7b004cd99bde060f83906b9d385a2bd7439fb17eac7e24179b8f1c636bacbb58293032d9f7bcd32adb1e8ba818db34828a0cd78eac0385e500e91d59f36380dce1a9c002aaccf19c2051d35cf22e2624819201815060f49dfa63bb1cb86afbf767fea3b68381f966e4ec219;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3c7875de3db878da866088699ca7e2ea823740a278b9f81f93e6992d6331dd20481a4ad31f94c3a38dff2dcaa98ff6cbcde8b6d69e14b220425165281a21a679d577c38bc2da781cecdf0eb3ab58f8828ee502506beea00f4c8cb13bc51f1a77b8a0f5d3a5925ea8c435973ea6e3e316a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8a584352cb53d9360051485f2297343166e89999f7e0791768cdf9f3f923d9a83a2ac0c233fb618018cfe29be2b4633245dd783fcba28cf0ef391867f44c860b37f7ec2d5483cc15593a4fb54d0329be4ee71abf8fa9a9bd11e5ce14784c66ba38acbdca5ac15457aadb159425e9f8ac7;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h88c755b8ebaa88adcc12a65a47057b084d1b23cc70dd0e58865746a84ccbd4a9dd2374ded1bdb56db622ca29961ca63aa599866cc2ebc72f56cd75f03b3312a638229bcce52f579e8f536280ac3f73448bb9df5facb1be9fdd84b857f579bb62b01268bc62e6d57bb40ebdedadc1e69f3;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hcb16e7379fa75ad35dc987f462f00c8f26661c14620d6c72be52ec8e122997276f820c3c0f8844b891bb241d42d37c874dd8d8a8e46ae7bbd0e3040659c4e8aa419333a576d8b74710c7bccfc514619103b12ac835688dd69e78f7dc9cd76ebe5b70a71a5c6a55152e08491c0f5230157;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbefd160e7c21eec0db7b9df737a86365fdecace8cfb587425174d88b1039fdd41534e1b43780528594d1ea8432ef581d48d6bdb2a700aa61417d3b196d45fd00b6328e05afdf50b28f62b8e79cad3486e425bdf2336f870fbeb24f7fb45abd9e8460259caaa35be427ad09ba601db1214;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h58f79155ce359545821323e774becd6c3f85d12f949ae338642f4e792d49bc03f4656a2eb135ab439a223bb6d179c26776754b05a7e8dca397a8b9858fb42e52f524a83c60f9304d1981894acab79a12aaa1b3503d839dabc7e244722b280759dbb2d7e489b0bca3139f8e7c508df7051;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5e2193702d33762157093d1e647863af6512c6430f234374bed12956390d40239a7f66cc2c7a656eaf6faf1b7c438cdb788baae353fc81f37a8605de98bda7e834cd10400e0d29e24e69e2fd6a704d208bb61a2e3b0889eb92bdf1ec7c6278b8545b34bfbefe002d01cd360da306e3c7;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hde07660509eb0762b09caa40be0957195f1694c000d0d07148868928a026f8f7438cb8c98f16eefcc98d96e11c45d7f6d281ccb391d2c5fd4473ea5bb860ef5a746f521c9096fbeb0bd479a76fd78181420b5382c14d341c80cb2f0c3afb308807e86aafe9cf99a9db00c0f9785e93b3d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he0620f2d9cda01e65619d4b637b1a26979577e80dbc51364ec9d13854424542d0de38d63ac52c303f1b93dba2f636f3041a9418238257723e4456167358b39e5e0df8fca072daaa51288996648de1fc80679672640c910f540892c4e24f2b48971cf0b2cd7eb404561038a20a8551ceb0;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hae77a90fb7f45f871364e7d5610cd7956f15a0b2f6087c2f7b89a948b1c85ba33751c6452e38c67a5804237153e005454144fbf03b65508034e3aba0eb74a17596bf65393557d0ec89998a212ecf589d7010727c38f2dc998ef741d259af8d5fa1e4d6a8edcb69515d50a99f486c5b10a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7ffd04f4f1decf3841d4cb95c02e569baadb23b017ad8885df056407e21b8a5286fbe753972b3cb202d2cfb4e9a1758b81ae216500648a337d45ec79af525830415cc18f757f220a31fcf53dbb4aa49237fb90ea6a2e4aeb74a35ee7a3689aa9f93bc75f715e1ead579ef03883dc99f7c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha3a59e8d07507507f6955b1103e4139bb9fb63ed09dab4398195857d18137c6e2a7cb6a4e0dc067c8b84108e9506d4e8720f6d8f8f84dbf03c70293b99166db681725aa0bb0f6eb6f9cb35c842fe4ba4ad17bc550225e84490269d38840cd6e20bab7131a5ea119177f91d60b9c12fe;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h823e7925df29777f2cb6aa45758d33434cd86decaaf902c03e89d7d60aba102c9d2da10b34c12a2a981a925b872b4a1e37eb306700d280f25eb5b3c3ce8a02b1230d5524b66f851543066e9b97940fef0a0efc49f204d08634611fe2aaf4b478367ad5748a6aa1d6fc90b8fe99183b0f1;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h73ad8af082721f4cfb048bbfc327549a27f51fe003db3fc1a51ac7b052725f8510b51df472d16bc9aeb48314aa9be36d29bed91d093bc4f80811c080dd039df7fef425386e0af35483d3b3b093cb547c8ebe6fa36f9e7ab626d33b55d1b16c9a4a9f72f6a81238a6c7de69b0a882c82be;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hec4c3f98d5ec4292c2ca5577b03dc1156f5c2bfed5de4d7ce5396392c0abda93086aef79c4c9eed3d523dfbe5406c379e98ee92d44fa07bfad38e72fe6cce0f37046f3043838767d1184fbebdd549578e06d2609edf49c79953e0f151b9830f089f13e0df3463b6ef6ab1d9f5e0a5556;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb320e3de14008ab732abcc06b2be498eed9ed1dcd119325030ede12f9b4d170527a3ee9e9419ff84df80f7c78e92565755710fc72b1b1f16968c9092885d38c5455f496ebf419e815234d7e6c6abf9a42b8744c503f45654dc22da62980cf708d0c751d08fa12aab1b43b1f7429041730;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfec7abda140d7355f689b2e5a4940427e195598d9848dad9b73c7eb87211b1073e4d0f5c46f88116f1882ccabb70c29ea7c71112ab06b8c34b67dac0f09322cabd4ae4f934508a9f0262234ff6a311225900b6d2f21cdedfc18fb24ad70956d6c68e3d1a038c010f40f334fd02adc2f39;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5efc360bbe3f85c5338437e565d77933c99c5792b09bb35bcc2f4a0b32784017115fd60778f010aa2dc9a3e76f492c45b38895e396e61afa1feef73611a5fe1e661118d6b07f84b32b76be833844c23b4dfaa27b8d7c400030dd14529d0ae70a08d87f67ea4eae1624ea94278f18220dd;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb6b2ac57bd15b1473618a0fd6e181fbdc9c01e2f3699be85690ffadde0d4384017e9f7b92dbc454468a42d50931a7b44cd8ee31d8eebe1453c39523cc5abd2b79f16a8e6d8d4aaf6ed217d843f4b278d9a49edc1808f2f4194d069b899ea28dbc590684f610a627c69dea5bd58497b697;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h67c7d978e7fd331daa2f75cb4dad75902cf45809e335e39731565c6fce9bdc47e1834f6c7a6801e36762df97f80a34fd9b5471ce60829dae222d3bb31a2fd12328cfe819fc7abd9799165af0b4d72a78e192be7e1660f7c15ce358165910cfa91ddf9101839f3e3f74aad990e7b2afbab;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb3321a6e85e113876efeba0563db5772268a1f28156888c2d009e1dbec29e853d7c2fb54e12226814dfec9ef5971390a95f31acb887663240bc23b67e991e5c6591a567e84bbcbed46dba0b5c3f1798ee5ae9e132e7645ca32a4ce09dbebd87ba103af4adc4824ac20ce3bca4de475bc1;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h405ae793bd94b106cdee3dce1aba6593b4e0dccab1330457ed203c94e1317a777109a62fa17b3f0f73f47efe543245929310ac64e95c2f54e9a2a073eb0d6cb0108af36f2ff28751895de713ea21daa31f28417b74f69bed5979a1f29d8381ea1fa18c2a0ef77125498ab3a7206223834;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd16677d5a86e682d9d4549e6c88030f694ada63cb0a9d7528fd49ee6b906e2da3b7283aa5f6ebe8ad28c9d92b6b5148563f97a935b4a2baa491fc6d6b8299c82254a65ea091c3dfe57dc6aa405f38bf2bd2ec5536a2676e0acad8aa10805be71420035528ea8aa6fbc54096fc0918746f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h35aeaf3d34231821f0b8e7f50f703a99fffba7b3c7bae398b8698a611eaf5bcc0c7bafb5af20ddea33f1f242e747bf1e8dc9fefb2110632290cf9eebadddbf263fe825d46c4c92103e11d342b18630fdb13af25776b7e5524eb5f6131944bc6add59ae5235e44e74988b950f59c24f2b;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9d97ff13c76d06c3668f07ccbfb5452aba9669c0cbc94356956b400f930b546701747ed3a7fc17415fa98d33575da80bed2057f78b72476c5095a2f2135963a9d617de742d8494af5ce3d84f5739c0d07ad6405e1f41c91b0ab7c4c580a968dd47b632bde9ddac49b3fd6d5c69fa42501;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3e8d03bb876f104cda55087f03601365faf05a99f7c01dace526970dacdb06c3814ad6936420bc686533f1d2b27ca992e92327a278c0e921dc52f6a21839ba601a645643763498a56debce8e2f712b2a2ca85d130d1c21d8558a4591f89d17a52a4200896f8ff44eef3a0a41c1aebb103;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6855ffff79f67eb2c73e5d9caba82b6d4de92bc3b90b1d8b9bea1c11bf00bc44ccb2736867baf116b5e3aad62f2adc647d95fe533f70177682c3e9b839f176efc48f4c7bf3f72080adc496e1c34a4ace88c821c93a7aee5033ef6001f53a607790e2d8a1d7950ce26dc676d8e3216d2dd;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h33a598c5252269ae3f7d25257720badec664717bc0f93bb3d66e5aa2de4280daf4445090bd30f07d5c3da6e216c064662a0bb55e4d847acea13dc0b058ec5924a0c08d7f3fb903251f508b9cc79fea8172ab98eb94741bc7bc20400cba7a36baef12fb43bc4435020cd3693e919aca392;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h841b61c6323b0d8b2eb649cbd0f4398535cc4824604c69b187ad140f25719028a20d022ce3ea3689217d28703729e4d64288d83ecddab2b3d124b9af2ccb3cd714c56c96d355832c062e624b9e0498e593cf99c2edeb487177e356cd34b1e717141a7f9c5d363ced979d9a00e61c7baad;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd62cc3b7fdd21ae9004297fe16550d5bac22ccf47d35e9cd921a0d21691467df06fb4d28c1e556c1ff917a02c0d1f8d5bfbd893fe86f9545b9f3fa7d6a9e1eceee14368139899415525560e2d5a9b7c715e3197c784bc2cce86c0785ea57fec74ed8dd2d56972bf4e149b4baf5a9c3159;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha2b416f3c943dbf06de4a4ee63443c07436f1d394f1c46101c36d46e818714a47a076d79b881fb0bdcf9b6fb206965f0238a6937fc9049cf896b7c822a6163faeb5d0cc66c2a52654459506280e36645d71a64be78c9049d147beafc283c986bd63cf77f53c9a9ba02ad176d053244389;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he433a74a0c221be324f675a94ce5c3727301776ba415f568c72bf74954fb5a41e662a316442d8ed610ab5cde50152948bfdb2fdf4ea3cf8dd452b0e2230e44bb4ff528eee6a179d443da9dde2c695d3f4c874e234033e5a2af1ba53a8eb3eb0e63c0ee5c6e4032ee02c169b1dca578c78;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha0d2e22cc3cebb17f89066daea2346b9037ae02975a38b376fce2f9bd857bc38fcf3d7d9a9d4b6e0fca2664d42c85eea402bf5c499e8210ffaf1fb02a1660af382de7f0bff0d34bb3885f92aa5da220957d7213c9aa9dc6eb3cb013da1e4131b82cebc5841623263555ac2a4adb70adb6;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h28e0bee2f176e0466b094519f9dd505adb5f4096b10bc68d2c15af1f40e15cffe93ce1ec5b58f6e41cc20e94ac5ced685a2b5a4884bfd12745ee3e7fef0fd1cf2fd1a47de1140cf8845bb0339670faa865e298c5b8f32abcb1a8dbf0eeb1bdeed79cbbd732776e84ae07fa7b289ed4aa6;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h639d91d9777396f36d098f30fbf5fc6a2cddc883d17589e36c4e6b53e1246483f6f07b8c7e4d9cbbb161d7b628c7e98e48004da5c488e3f419f1dd59fe51438ec6c24f11763cd38bf5f943467f1c291fd8857e73a9c2cc23ab4fbe73b3f6108855c827d81bf106cc29a21d7a70a6b4c54;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf31eb588d32eba9efcd18ecd9f108251ce75f1dac7f739b605302c17414425f79b4b40556b248b9c0e9f30c285e88766e6192405e78cd103f731d14b43bdb2d49c966b5009d61db0d6337bda5fadc9651c43a4408f2fca9e7ac5793d20f60e1b40e1202221f2b5ef5aecefe3eb0bbfb2a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha193c8501c373206552c6bd15c0b631d5703dc519ae24d25846b82676f5764c4c711772ee7493b6ef3f7ef321d3275b7af0650f1f788f02bcc8d45a854fe247c18052ec8a672820a012c9ed5f8025510b1b3a882c3d0de1d3e94a2dfd65d8274bca463c7226f93ed7abde9bbfcf1170f7;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9826a298087a7c75043eccd4138c32d1fdad6d0991210a27a5204b56a1d9b08233c8f14fe3c3ff1642dcf1d53d70546f028ab191741d489d2bd13cb199f0470db14bc4fec0961e0984d9a67379f39cae902b10508b2c9d30444f35789706f67ed5191234da7d3341ba3febbc9ceed7a47;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha7b58540ba614b03085ffca4a3fd6a979c0f974e024f60feadd38837bbdda1b767b47835b744f9c964746dd2a6b93726e68d2a73589a85a89e6e51b83a8a06995d58eace75bcf5dc8175ea09c22f8b50036f92a5147f7910e4820e1b11856430371120260bf4122993ef0f93933a0ff59;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8a756a99502513a386d16f647f0a05953fcb7d68d568b06e3f001c8a84ac58becbc497c7f2f240802241133af48ad37dc688afe075525182a6de18212c74c2ef0b28fb2e92728588c9d761759c6f2174b08ca45b5fd97a2128295af0a0ccdb3ff8076679219733e81445c894887871938;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfa4252f25e56ee27f1d970cb28a7a715233a5054c31bddecb2006fa84f3c3b96a554172c2b5d1b21be8b4674ff40c571eaac8dfb358f90ec5e2cc799402e370381b02b8a9af7dcc2e61a3cc1fa0a3ab261ab3d335360232ad73662ea567fa20d25cb0dbe9c8cf3db6eac656d6d3f0c36b;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hba90d5629d205cf54f0f32bf9ccd756bafabf8349d84aada9a70a50753a042e4850af4152484b16d94d2443b4220f17e2cde89b0d6a057afc6d550f137a986860858beabf12526555d7a026f13906e4fa694818cf248ce616f570bb0cc06a58bbd3e6d9d23388fe328f7ecb2e073d51fe;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he8f0b6bee41d8bb608ac8c5d68992bcf079a6367f13035a19535b912aa2805f0a9e283e4d1d074e42457886365ee2fde99e3070f1d13feed2f4669c1eed29a5adae4695bc1afcd7524e313d72dda1e2b80635a182b2ac8cb0cd1213e01551de7228510c72575de44a4d5c944b9538f228;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h70faff3c48c0f78e95aed62905bc925c069e4e385c1d54953190cc65c3f7c92a2bbca19c7eb9dacfd056386c8a62c72e4afcf186ea01abc0932aa6527869e7156693a03ef1c35c6001e41e16f68a3e85bc95530e50076858687f435175c54991929e67b1e78ba1451879abd0767f04bc6;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h70e5403923722b78c988c6b149e4d23cd1790ece1344f1cb943ac4098123ac4c8293b4889d700ca8b6ed121494bd780737925dfcdb008083ed31a5ffc31bd2bd2e789cb2819e4a1255027a99e5dec949eb315a232cf6f85e3b5111048b48be9ce4bbc78f09d4e5a22e328099ca007f52f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha3674893bc0609e84990f0c7f1466130d8f33573b3aa80ea642f97e295ac84d2a425f55b717db73a01ca9e63f6487d0e78ee5d558dfcefa4b69d9c067817f745b262046dcea1b4c6c2d9237aa7ed906d564b98f513201a49eb60d96dc0dc2806a68ecddcf1aea775cc77ddfd7245dc729;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8ea8af1d5b320db09612509d3fa7978849e1156dcb383ab91c915959ac7e9a6aba23f235534ab3f96466e9e4b062f9887877df04b06cd3abbfae40f77ce17f35d69ef6f80222e229cb0bd35125f203add69be6b11e38bcf5f71a05eedd84d3815a6be8470e07db09906a13cdd18e6ec7e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h11a15244e28231be7f97c22cb14b1c416c7a47f6c0c1b153fcc8d77b78a455f4a54cd139d388d459dc6409bed8421c2ba448a2314480e10ae125c6be97098dbbb2963ae2b41e0f4f1c3a25cb0efeffd29e45cd250b2783d0afd6308b7c13edb57255e3cd176a549402a6f8f9108a32755;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4d1ddb823ebf99de573d3565a59305921e648b816649250f10647c7367b36a5ceeb62e56f643b9ac56363b2a9467cff982c3b37c8040956c460304c347b749c7ba819fe4a2267bf30aa36625d1135c7c8f227f4f3f33630228fb58570fee295626aff53c4f7b2eed1f3b1f63866f3bb67;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3b22a57e635178606faa2de458fa5b37da8a619b3759fd2f34872a629514072836d430a6ba6677969c494b1311c621c1835b57b9716ccb6e0fab7ca12aedb43ecfaf77d2c14874dc65ebc5c60a9e53e7a38958f9b9673e9d101184d9987cbf4cf02b29074ddfbd65fd2d203942d38dbd8;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1e79ac854c6b47557c1730c6e2e3b86df735d3b487a2c269c0353f398c927a3896945e645f3eafa2223f380bf4d283d66a2515cdb23afdfd01566b1e8243f79b703d713c9fc542e3780d3fe77e97293ed15a32138f1d977d71562ea809af8134f6976fe8c98fbbd6d202f0ac90aa2666f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h52935727564fac9f943b67926eb0b7ce614b05e68ba893cb903feed71feb67420e078abf642a2240315bb7c9d8b35f12ed1b237eaa13a57181c21d4227ecd03815549a4ab158bbe19081533bc4b7e1e86ebc97bb72813f6e89b4f8906b3062fc19b4bca2069113b7c069351ec6c481fb7;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5909cdc0c92cd1d8c1beed15a4ebcd91506cc06b6af1a1c22023eedda3c66990951ba0b1029d8e5d0b45268809644c4d072c0660800e1a2d5d37744970ee2d1969fffd9f333f1cfc1d15709d9acb3bbd644d4fdf6ee21503ae0d8098326dec90deb7c3d1b912c2acc65768193c5371467;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdc3e097cbbebaa2cd8242835d2139f00cd7c9f38a5991165689b0f5e9661d0983a524141616a35455a46718c85d55d287cdb7ae6531913f307265a121826b88b025d1e0979602333e62c06951ea58151f1ec12cef29ef4b83602e9f9e6075e215d6851995eecb8f5a3ef174dbb09bd940;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9b7e0b0c73342ace25b7d5758fe0de262de9cab6fcc836974b0a184dd575af1fdb3d4140ee73cda117eecced5f3eec9bd7dcc8ea4781ae5a2b6d085a1d6e7946e7acf9cd84bbc2f4e3b30ff79c854d36816048d8ebcfaad1fc363099c40d0eb58f00f276509d203f43049289c261410d1;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h42e9655c530da5403eb30b1ce8d6317370bdf6af693c47bb22fdaec143f9516c41f24cd81cbfeeb9aedfad153bd521dce169ec3e7f4536316704b8e3fafdb8d4087048794c3b251b41a98c42f42bebc82a156f0d2cfa01f320910a31c162b1eb0ae7f9870b095aa26730e89812037dad9;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9c048b587ba090e9ff80f5d3fb580190ef0f28fb7271d8bbfc2be116ad923bce492d289e74930b350e62bd7fb0ba1c12e69606862db4a5b6cc99d1a3f48b189e5a93623218d9dea942d0973936bedf2c26311cefd76054cd49705f5937cef2e885568858eb713fd9a620d4bb9b1014ef0;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbec2d68e6728575087b619a942adc5ca7a0d19b74105e63cd2a72aa582c4915d4e0c6048e2e182f1a60d970ba6fa434325974ff7ce36f110d4b091c99db11574cb4b5d56e2bcb307027cd0461a63d1609352f7bc8078636374c4b178160fcd8ebf20151cedaf791593038a82debf418e2;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdcb037811e2ae3a92696efd15aec1dd012ee3841d154001a79a05c395368fa19c5aad5a01fd9d51fccc7f0312c86c6dcc08aecb9cfd023dd4fc4e83e2d71a1ab25e043a1b43d0ab4101db78c7fcafb042c8bda0f7f58e0ceba6bfe12e6921132464cdfac72d004b49c28199f1e713c68d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hce29849d45644a75d6fc232215ca6345b83d091f42adb406185a2d05005d88d2e94374a8c851612331e24b8b190f1e862331cca7fd3905feefd7ae2803ce8f205667a29802e6dac89b8157253558f93307a7ca25de9ce3291641b0d3be3f283ff530afff86265a29f762837d3986d1806;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb0d810913219d184e716aaebefe859077d0381cd925770bb29ca88a33e9a2adc8a7743be6f9805344e0a99cb541720aa20673cf5d8d99ee8828583eac5fac2778aa852a6d94f6b6a7090f78831b0bdc51e343d9e8a0454bc41bcb02ad1726b9205cf273d6bcfec5c5fb6d22a8ef881baf;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha10c83e56f49a141bf492bd03ca9222e46f1b21f8055caf4858fcd652d620e06bbce59bf713eeb766455a2be8f34022fd61d173c48ef185acf37f9974ccf84eb99afc9acfdce26d9d2e741bbe8ad7a4a067d708987f838fc5834ca61dd3cb2ac7797b47d2830317f4618483ae8528c337;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h47e7ffd6fbbca9f478f8c45a89ab9e043b7c29ce1134c07d62c47016fa27505e4251c49c9f2a6a60fc1eff2b61897e18c48f6d136bfd25294703fa8e596e218e30329744138fd259bcdd9003ed8a83fb0afd814dc475b2760dafcc20d6f6f4111a6385092f989d46a65cfcbac10e37b89;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4f28abbe3464788316c17eb78d90ed059ff5b67ec16b99582eeac2e266cebdd47c794018a6047e390cf31d058b978f2f1217663effb404fbb811599903095f971a62e8b8f74abeed4628b408baf0363e5177fa30350f80c6e9bc46e2be4bad5021bd558ce367f612bb865293616f64597;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb6484058431de16dc82783a0626425f7708d2a6077e0784dea25a97c2f6815d14a6d5fb9588d9584911bbdf42c751310bfa8704cbe93a2a25f245bff7a944fa0a5d7a1cfbd011cabad2977d8b109d2d4ae25dbdccfebbd9736e0c5d293fbb7c88a133dabf9ef5e66273fbb6dc355fda34;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h30b1642370f65c6820de18de0d0e7c7472effb8095276c9dcef77c30220184f57a7babb0457186e7821a0b9c701781cafcaf15f7b30776688f125c6f7e4ccc29d26e1dc211ea6fe80705a08ee982380e5bbb16aa08273e103b97e195356e1fe916eaecad2914b1497eb8b619855251860;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha77c4190181967fb3238b243b2836f96291923072857eb6233bc0d0dcb1465d1490fb80803dd3a5331d9a8b660ecaa5b9b420c45a5ce72f4dc5c7b613c6f1069ec90aa8ddf3fc44d8f41a4db8538a0538466d1626cfd532a8e4ca9bf908e68ef6fb565a3114d52db70e7a55215ae14fc3;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbf36e05756fa8abcbddd79c6bf4958e995941aacf2571bc2878629a8b25dfb3c01f23c7af88ca6e274a965ff39cbacf2422d934f5cba8d157a45dfc8d96cbb3aad239f7314c0626d31bc2324d8440f7384d4999b232997bc7c9fd839af35c88e94f98d16647546935ad511d02c325006e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h337906f5dc93e03e8cc8d74211102d8b53c7b775fb0075da3ef8c5db7ac72b6a409a7c2d127b2f93624c6a464b24ce09b715996dca54f8a7bf8f831b2d6b5e9600bd7e02b7f49a18f4431598f1b52957458196fcb80e7a8bf42ac6a57114637170be7bf621e7fb8a28516af7c202a1b1d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1fda0f83ea7e248f165c58b7108f9ebade5e53e6fdf35abe427a402f720e6fb0f0104d510e921cd272cd2b22afc374b99740d6db6a5480ac0ef1e9fec0a2a1293fa6b98db735fac443a8e698e5480ce89ac45ea0d439698d7743039506e6a1d34119f1a15afd48db14931eb208d8ca52a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5e3d08edca93283e631e2b0efe751fc846c65b8e9a08b39797baf618748b561e5f070a759c889b2a7d25caeb20603de14e1d4eb06234f5610fdc5dd96d12c0568982da182254312b5c79e5c74b9f67aeb84ca48c91c0a9aaef21b2463bb9e97db971ca07bc0447518fbcab95bdc460337;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hcd684e2a82aea27b5464a8bccf8690fe994bd657fe07386ad5c0a69d8c14805e80cb9a390c784d73d25bae641a19d7a4a4aebfa73881d84221cb9e79b9b1e45abebf6460bc86ba3436ffe72dddc0301f2796638cbb01fb83c64a40c56345aeece1796b6865f0a98f6117580e87c05c8d9;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h431398cf6b1c9cb61fd257b528dc2034d8bd2d5596029a30e414b67a11f63868cc76cf3fdf596218c00151b83c6df3a963730dc6111d82f2c00f3c6fa81b55cdb6625965fee26d4b4f40aff375d18cccdfe324fc318a2fdd5123c17020b9661c42724fa1452bd531d71f68b4458cd7d61;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he076949d481118de71db9b046d95dfe5d3ed37ce5221ec808fab813c1d0bf340584fbd1572bc66738a47a97d7cd381252ee0984460103300bd96d73c69a360fba51e604660e08c8af784bdffed4af6e232a91564e64066d3458bed82277fea7978d6793b577e72e5f28d0077e51e259cf;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2f7adb8a675079861f56367f5949d25ba21626f5aa346a944ec599beca0f9c391c05a9e38ce7b37019eb9b8cc4d58be21370b808a01987b98797a6d17af29bef7a4a34f2dce3883fed4e33d87e3973db26494c1bee2ab493bcf343f8ea8d2e141b28dc78f8f1cadbf039c8462e5d2941;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6deef0db523ff007273ff2d93ad0b736e88cb62bb1067c23664841ce3405858d6ca6ac9eee80ef4312020d5450abbddc39abb4ccdf5635a748542b2a9dc204acae4a811bdff884ffee52c73cfe29098f33e170253a4fbbd69f9dca9b027048d204baff63e9db840288db5a2c2cb8e4eb;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h743657c7f758c59402c9621e702075dc6ff8bd0c4e937a47409a4d5c820279e485d2d50725e43b06c5f7ba35b45ce1798d7fab43c9ca8aacc04e8178f811d6fea5fd0a8b62ae54a68115e4c129b0adf2fac06163d1cc027fa1519f252c18b0cb0048538c2a2b81cf87870d1e37ee52381;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf404ba1066d035c6cda9fdb31aa31c792731e7b4eb27e0d0996f672136f4c908364792f539749e147046290cf90d3200387898d1ae52e602830a283d28bfcd305462bfe6538bb75848e39f32ee339951f2f7139b5089ec3ee652e0db9e60a05530731a3da675bdc4c9e2a4b5aa4df2886;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h191e9f8169fc93e4adc85b4910d5fac4d72f25b83ba491c108b1b3aef8c420b990fb7a9554d13e840b2805cf85137ea49f92600f5cbeb95e97cf1884a63d65d824f510dc679bce2574f81beca5c72945e6fb4dcff9c98779801ec77b7762aad0877a407517bb919a19f3c2b80e608325c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h77779c85a53ee0f58816378dd13f2a4464e83413c04078fef096ad2ad577fe26eddbb0d74c5039093beb3effae9d796833605e4ab58255b5ce506628d389b461da076bdcdba27616b85451da4e4708c35930354642a080bbcffd2d10a67b7494400990a5844aab4e68e2a660fe871ef58;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7d68c65f668d277d89139c09b3e8b6e820c56646263680ab3d176b5c579a2c215939a5a65ed282695aef818d4397316971247b9b5dcf21b543b60c49d26a2f1bf707033284b384da4be667101b109c738660be1b59d2a7bd827393fc11f6b4218970ada3dd78b7ee1bb468c859797242a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h917a101f11fe996b4c6667de241e7f8f3daf160f72ee293bb50acd41c43b18fe05023a47a5df70512e930652308695b1001838fbb59d1c6380173d0d3f4f62e200f711e116bfddb0d889ef13618fe7830feb3a868a9aa50086fdc7ea6d367840a78cfd8b620297c2a61016d4f1bbfa841;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9af1ce39c710488d55271aab8ecb42a2d3e9219db446fde85b2a65372466ce419fda73fa88d3e9899f86ddc1bf6aeb29b983cc10329ab668ea15a2b25f082bc99466bf53d4fecfb5380bf7c6ef71a2f5756a55dc5d27184cd84566704f4c0825e0ab4919fd1f251b3d5beb7051732113a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbe6850118a56ef5ccb20444cb9f5efe454ee30b7cf0b3d88dc2ebbff7cb947346f2a3d5f41ea705a2b863fdec5919fe3c646067b496b9e40dbb6d1a01039f49aae5b75020ef6f56e3949fbf6afa164e2c40761ca1e59f1505723fa054d3d92406c58c715c99c50d2035f2655b3f655983;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1e2183567c9b826030956f4c068cbfdffefcaf3fb2801ff2e8e07f166c148445e03f25554dd7d4eaa90ffb3823c2ea350fcfabf2b1c7eceaaf687c570d56b621261de8c02a73dfe9d09fa643e6b5f4974c56d74a3eb12a5706ffa2de2b08f4a6c90f773d88eea40aaf90270c9619a8ebf;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hcaeda6a94bf8219e1f5e182135fdfb52a9284689d7215a021dbfa353e1680e6253b27b781c3b49908a81fe102bc12273425e7064065a9a90f16a2cbd72427d3eed40bd01770590b2cf6dadcca1200be9735481a5293b2e271ef88e4f70a616cb70439eaa878bd10d6ecd30185dad2ec9a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2d50cf50ee69c9c7d278592f921d8e13b770cd77ca4eda8a1171dfe7ad8f9b9bf8c3bf741bbe8fac051d553e31e7c245a56af54dd02cb603f93e769bbb133d89f9abac16fd216c1fd8cd230c86c54e62002c19ed47ac7d0311c8341d4f4456f43127fd6c3f53a1ea0b5ff911c162d35a8;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf0851f095831733db0dd85dce67b16416dfb14bebf6a8f6b286786823cd36fced4ca72b3447decef857ceaa6a5047a83c6443fce148d59d994f6c9fbf6806b86364d75b5076f3e308a5f3e72f6c0957711a385969a8b25ff465d112c9f9bd13eabb94e481e88031eed71c83f101528f59;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h56e7d0f08d2c408dacfecf6fb3ae53f351c6701295e21e8534c40bf8b088cfc7f2283f01e97d1a6726dcd37d64b2e1a8ea3eabbd42f5fbc3f0793498c4f88431ee02a090fa5f5c2b57c92270d2a5ed528bf8d6d8dc14c90b75c95b872a906b1ccb8c0db8bcb8f20ae7b4dad661658ce06;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfdda8f893a5b661c70c7c0582963adf1109461d7d2d183473b2077cf77b17a54ffd7a4725d8a15e351c95bffda5540d1da4ec3eb5e36c039855a135cd92304407696b83945d33efc827375375aa3b9c00043fef8622c1389129b6c93b17b79af188fa18560d316a98a7a59d168cd62777;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'heea355000f2036bb2e9e45a527b8366b295f60f3d811a24ad56e4ad2d41c83689d2605c48de6c7ab7ecced6ba5a62a4d4a26aa4bc47b9b9a8a07ed80743dd1227f28dbac6272287fd3a7e780dd7e046ca2656da3445024e8e274083505e4d338158ca837443a37c17af953949a7f6f4b2;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd6c8a2d345a0b2c080bf404833f208406d9421ad7931c2ec65950ef2193950f67e561289ddabde91bf3b084ff976dcc3667f47d123f0ba131ea01b6b6ad12dc41e78d0017da200fbfbd6c31f6a64aa0684c6d6e7d55d1ac45a4866fe46d58c89316038c80024c176e34efdae9e3937800;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf16b98d6c224256c1ba36b3e212334601a9cabea2e17f0f6a6cba5237599e69d237652c63766c21f6e34f7190fda58e8bee2f2dd6d7445e773cf5ec547e97197a49568a9b58387dbe015dd4ded9bb4962ec55f7c80733cc49f9f1a17201a083bc86845158a4b2b3a7117662dd05ce568e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he0975688b91a2fb76ae82f61208fe9ae6180bb3e37ee3c71a23bc6cd2ed9bc968dd9406c8188fb2468c19b4b568e7358f136cec40fb1236f8f01576930e6efe16613c578c9223c2ea6092fe6707f44973a4f1b3a7c832c86ddf89a77756463bce5b2fd4c9628362d3a6a4247cf93a3e07;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf43ce5d6b5900a226b8243ff3292ce29f95852eaa944a275cc699d5d00de227dca9cf6afaad5b507fd8411bea8c267abd1539dc81ca207c61a78b89e080614912a95337b92993496e7e9629333f14c03d893fdabf954173d13d33f45f8c2f1fa5cf8eab5bfc8bd763d8211c06fae53008;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h348918ad9c2d46b3c8a9b6df08ecd31aedafcf945d347d89fa34e0a28eeb92cb9d01cc0131f9e6119b49195f49430a905beb9204e87396b318c60da322575979f83e7fda43429741cfb2afabf02630cef3dd436cb17156d45df8c5874d5c20ee8b40ba9e835b90a9d02e1b363d7556d4e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc6d634041868543bb6b0c34eba0714faa1f63040cafe787bc0de10a54b9fce1c47085cfcb91e2f97907f6f038d647ec921b01c776e3456ce467825d0a41333aa70329c17567798379eeef22e092d79074eb7f3000667127bff572ebbca03c97a1aeb2bbd9c6552fccad2a0c7a0273ae9c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf1e0b36c0c15d0f40d2a67ebc8353ae20666bd01650fd142a664c3e41dbb8191e63886f31cf240e911c3c077dd604d556e9a3003dc29e3dcc2ea3c291749904a4130521330c174a2ecc0093208b427260635310e225266daeb1cfa967a5bb7eed57f2fd99af0afdae73f080c5a459c2b5;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7684aebd76cf5334b3a328809238a56fe1f3d063bfcd2bac7d0c78b830abae57d5073a6ccbe8d9d811bf32522debf5efb82460bd5a48cfa9f8623260682db5544956a1a6654e34905f611979cd3c29abcf4ffc695b3bcba13c9f9495020a9d764925d9b4b2329c5e5e67c1dca1719bba7;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9941708aad96b84c108019ee0c173029d265bdff8cb7bdd002baf0e77d489a7ee19d8be8ff9153dd8eaaf583dcac05ef402992e10fad79d96b013fce8e08818e46fef568512f3dc7d9f2c40c0124ab5e26e6dabfbea21d8ee8fd723aeaec3e24d4572f27608ba5f8afbb981fef91dd1ff;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h31dbcbe226521d1adc139d36233fec5f42d4c34461ac26a737cd8af41b04149519c0b1a2fcd4e7f2ca4a90647790e57a6ae81741974a3bfc33fe440a65378b6d2ebb38c7f3c917b79107347cd4c23cb6d314b1fa6c8b6e28ef23745232bcf19bbeac4d19ed18a228aa91e388c3f47ef34;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hcd9a6bc5c0d8a80a02c43c8eb96848934a3b8a1ddfb9a075b9d4cf638cb4d074199bb4515135c10457855a445d0e55282bfb67e12a178a2106e99d35a4c32570b75f29a5c3aeb55aaa3e662663509a91ea31f007d157f4b0b03f7aff80f68e8e7f28fb8bee0054e287d9928364c67fb0d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc2ed4ec4f2be5167611b72f2d77ce09698fbfce48a8d5fb9f977af2d5060cb8f611dfe2ef546435e00acf5ce38a1352ac6228ed03623f65be31437c84cff5e4c2fc879854b6a6319a282c79b19c5a5ef00bf181d417b97a1e2a04f16f45d7473085707d2f1505ffc346a1f26c4ee403b0;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hed81b8763d909601b848da0c7e7d23ce970059db352bf8a1044f8d3b1f27333576be7c303d83a8788d805558ffd1e915921c60b773ed9778c8ac88911d11f3e66d7a5ff5daa0ed3b7df78f2b6265c80ab3c646e20bdc12490a928aea9ebde41e147e3df4c09d0d4dc7b87e41d0171d0c9;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hcb402a7163f5f7486827ec34bb9ab5a425a41374a493fe9d21d1903ea0989001c892cddaf0e9c8bcfad8cb221acfe8bbd7913fd7cad9868782c18751d23375321f4325896a1aef4fac8a056e1035faec131903b1d8ea3e6f1b6aa0156214a63041fa8123d6588f429648b34aa47c202fb;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8f09e3b4583572abceb962ef6a0db87b3fe35da1388adab6364e7a1a0d2178b850ee0b060b77f6cfd5197ea7377ca15c05caff63aef0b75d77be8c6599c1fea599be44afa188f1d3fc864221980b645979cbc9b6eb4432fbc1862ffbf0298f393a864a87d9866bba1a6b9eb020757cb31;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc601c5e6f46e62b50f9eeffb7b4b031ec9641801a7321810bf61684909ce8b5fe5b79151a253b59a2ac1e7f0b94d39103380d80d6b1d40ce9f3bb6967d954df92f893c5ac2c576009b429fee49d9a23047f3a1ad1388a50b659b6119f9fbb98dd5f5a9e037a59d323e9fde41eaa9552f1;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfb76a4b52405c5ad8ac639bcbf7866dc1dba552a71a4ec1b3d6512016037bd3d9ec5d0e7f881c18b8c6b2b6211996c4d73889ff365404241ae262a5e9f3c0975f5d7096409a1225c8c8786517b1e1d7546c7cb47485ff8ca2b4e4bff5ccc09971de57214c3d3e72cf959e4b2cdc661b90;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5d3df162ed0091f3092b15bba15a34074ad39d76b9612172427b542aeefc0e70772fd38cec2dce3d583b2348b9071867347f668a853d2f1b00ef44d980aa84bad14c9bfa556aef80fccc842e7dcf80363b4d546f162d51b79045f0065afa23d495e959873ba0dadfa8ee60272763039e7;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8037b8685c4cc5821fe99063511b432a960b93c4141169fb4b7b38fca35912df4046c6bb9fa886f2cf75647936e122d32ef33f088bde34c22c05f2b514a3440f1ce29aa6da5aa29617ac024fe8a7e0144196fb968e1b074381d8658ef587305d07241f319bdb5aef6be01fcb4806ef30f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h655781badf65b756c00e001d05f4f35a0f772acfa1e279a0ca4d9b2494b701226ff305edecc9407466ff5ae6b03ac145b835846933660669ad610df9e34919bcfc2a259ce944a8d0a2813c2c8c603e86084990d1d438325121213c5d21a312e4f1560319b4f315088376403e7b048d302;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8a71ce6603179a7542750b946e285fda0a5470cbd3fbd8ea94c9f91137bc66d17736763924545794cb04c83d7a48bd62a00285d6677f5ef33122d0f3a47f36816d7c7a9bde1a00e2b3156fdc56195e26f05cfce15568a8bd1d47f9ce354b73115ca6df84f4d7df8b69629d3e5965714b2;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'haaa82452348c98cefba1f150165dbb611b26f034d0df373eeab399a778293fcd369e19f6fd9d7790f836c936c6c5714b4d91207a3c022dd6b932b37fa5c7fca2587af52a2bdf0be0d80c53294a99b3f63cb58d14a4ee014ef8564f85a4f76ac3a4760351b967fe86e81c8664fa074751b;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4673b244c836264dbcf5f693b1a9afe782878ba436d8cb0452f5db18cbde03eef4ce4e4f36db1c90ce3418bd5fcfa4e8f1a3f9202a86a7b6f4c8b150edbd6f7d84eb34d3986902b5a7214104961d98b7cb69eac9a8d18ffee01997f5bdcb1bad428583ffcfa6d17ae0e7cb1ab89ae7677;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc16ab3230e79ffacb1076ecf6163f4a0eddf090eeaa93db20f9499310475fa71ea528f2c5b2c23347886960b1a5c276085da955325a4769057e5741029d52bf3d1f81e7c77ab6ab9ff78ea8aa717d0d2ecd7437fad09f9ce0e7034005cd4b9da6ba55299164d23bd1cc2f35b6b0119d50;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc9c03cc4c49935fb6ebae4afd8d74ffa660399e3e095d7bae94671e30d70d179cab6d554f288df165250236d8497492271489a4d3025d48c7e7d336422bfa05a76a86770542870065db4a3149f620fd91fb1df6398eecf8efa2d388de403e425d939756933aecb758f80678b024e1db0f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc3448e7fd015e809fc92cfc947dc48bcee629ede1483ac2d40f5b6d17a87f7d1847f44aa1b25388c7dfb51ad5680d42c3d5277ea638da365b9184ab0bcd0d4ff688d0634fdef350021d8967d4a95b34f8a045b3489b6c3e8d16b4618be09ce284118e156d3d26c577c8b518c87adedff6;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h45848c449edc60e536d7679ae2d260ff30c3fd0954d8d8e27deff2397bbc16b3a77047e64d432bafa82daab5c831b060461c2239f4cfa1bdbce081a5a1b800e69b888c8990afb2a1a105b518890f0e149822b8317b3db8a363b18cbe8295e112c04789cc53a63cf44d16b0037b3248562;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9e7ba8caef448b67ef10e5a003e00d828ab077fddae48d6a33fad40805617c3e17d0d22c8ca9835c42c8c7c55e50935cc55385c8d809081ab9bd129b6635cb89603af45fd725591f8823151e9b10089cb8dd61c8143e3a42c63c49a4c08ad191a02275655e04ebba8fe887b9ae7e0fb4f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5a3f322f3d20031dfed790c3afe2a737a0b5ada032bca1206b741ff574d250b44154343a11a89a2203f8e4c0cf0e4f9ce9e53043167ff3dcc474a33cb246e213169ede2a59eb53f18477c2f2cc0c7df234230529fa9677edf76a27e55af829b1ec47094636147097e283b02fc3d231f58;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he0194eb52ca08e2e2542f4f08d5f4cdff8d6cc7966083f133a143095081495167833f53549f22d596ca69135c428787f9d2d442ffecd60c86250be7bf5eb6ddbc4fc02b92f3245ec02eecbb58135b43dbebb3900d4c0141821c9a224bf9316f6a6117e541d2e578342d8b4adaff3e6d9a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hcf739d8945eb9ca71ec6017a4f7b3465e0ab212dcddfa6399076f6024b1ecf3881b1278adb3e20bd53bdb58bbeefb3b8ef82d0e5d843a291f1886705e7adc6176f17b5b2d574584cc0e9ebe54b0a31531936dc07b8437023912649db44a30ddd2827fb2febb0b0b52929a0fb569406e8;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h841d7917fd3e7e419e12bd301fb3369cf4338f1fb4602ffc4000efe0356a863d11dd09d9ec78ef167e5e20ad32b0aeb6063f37cce0964c0b8083728fd9b5996b049b8d07d89e00f9b67bcaa5bc0c1572882c5ff55a2f92b99aed951dd3490204f4e0a3f6f34426aa0839d719e7ec043da;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hcebb8d28fc5fa90ee53e1b2444eb345ab75a4e370779b0860f44d16c4218e8f2db4f6e30c13d048f97e853157788709e858de5039b9a2b7bdb1f665788f985356a1cd9bb4fe3e78a9b60772ed7a12dcaa6b378367d9621cf982f1486b70bd539dc7cab0804289409463bbd4e3ff805831;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h916befd83d11910bd4827c77cab68f7c8f8ad7f441f10a3f578567fe22d7345503dc48fed18c113c89bde505365be26404c3d65f165503896f05d7b6a32d587c3a3e493b07afa82c5a70a53e04ef5025104202907d5b27a41c60baa6d4b721d303a6d0007298bea645ce5ee8798d60801;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1adce8d88bf0841a45fec39c121ff6cea24b4dda8d25279b18310a543f960c7c3d1c47d64aef1d5e8899f3e0d30f21aba44026dbc1c72098656399ceb5ebfadbd07ec38db30ebab90edbb869bb05af7b23dc2c3073ebd4c011ba3d51b0a821bd5605e8bb8c2b07219f6a2dd30773fd287;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3cc4032676150fa8119d3261ec34d38d74d5ce69b346f618d7027100b02e4562b4f0d4a766a0826178eac9ba7f0dbb2ef85708825d34a4ebbfa4f4f0574b319defbf181a3873f0b74ee9890ba315a721acac70e8a6a0b2f64e38e61a8fa5798b7089c9232c0ecd54da11d715af139e1b5;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h249eb4e6f5bd8ee84c681b67f8f9cafa60b9abb5b037feed607e022bda46d3b2630330acabaf47dcd1de7de8ed07cd68e3c65c17a67857587bd113cd6a2ca8925b76fe0024f94104aa343eff29ab2ec95a9e7e1c315b608b03827fa11b0aec59b0ea4143eadc24c6470fab613a7a76ee6;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf1d3efdb37edd78324507f7d026cc8412eab75295559c8526e9ddc53589ecf0376930b3bc09e0eb14ee743fe606e77129d9a2ad593508e3956fd83810ea5a28a417210c45c3f898ec3e5b5c1c6ea5116577c29a6ee5f8ab20a194c0c53c0f362bd8df17d8b396e4c95ca55180b576356c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf16fad34f837f3b4dd79b728b39607e0a9e8850968305242d666fbf3d11ec43cc1b26f5e97862e9f8d3e2956338af392a2a0705c708ed4f709789908aba60f183deba695460c93d8a0173ace400d66c8f1ac5f2b463afa08381e0c2d08af76b47a9b735d08906d22d8dc42599cb05eece;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hcb764de9aa5cdba8b21b29769016ea708b48aae3a76ebfa6c6981aa15975a13c3479de7e2ab4bcf89f36282c4dee2c3a1d657d8ef658b50a292c247bf2cdb6b9ffeecd904b8576fe33486ea8d88483b6a2fc3bbc2f1f771f64dc8828679aec45925b6e3f5733561a45e8f569ddf81360d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1da8b77ab6bca1db4eaa57f54cfc1e82287a64dc3480ea6fde5c3e0a57a88dff2ee87c66344f42460217b0e5cab64770ad538e2c94cfee3f8f9f0ef56eedf7a30854eb08d1dda833aa48adc2c0c75d27caecddb4a40847e5c146b70d5fd08fa25639cf938aeea0ff1175730d30fa9942e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha72a5b9f00f11fa27f8337bb752db9d1efc767c95e28ba05263ce39780bd749a1b7d33082578e996457304f414cd1fc59aed368ec4f83f0002610ee2bc3c3c3df08563dd877ca333f2162c9855f75a1c0eb1830bdc8ef0e2d13d2d3cbfb95bea7c63a2d219c78381917005cb07293086d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2202120e8d437135182508e08fca2bc2a358b2c1de66cfa2af99cc4cb83245c2b960e9338859535ba44c0176dc866991d4d125c43558085f6240cc1e6b111e5c6c8111efb3f5ab15427f169ed247501a15276f45c0c9781b066b69e500212c1e99cd97ef279f15a70d5b3eaf8bc997bb6;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h902dbae1c6697e5fa2d0249511c86547f909e0ead9a9df1966d69740b8bb6266e311c3d0d8219cfffee16a00f28c6321df5d442dac90c6e7a1177d1aa64e52a61cc95d01ba0b675f003cee4707a56d030cecb6fee5bf753bf75375329ba6d522b8af63fc87b3510e194ea8cec6ffee79d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3d88fc7761532a0c3080c2f05255ca513b8c85e5f4d2bbfcbe540011723e878fc6a8009e2cc788e3e14fefe402c948e6a9e8f512c897355262e8849bafb564d8b9d19de2efb4ce57ed2392370c76d970a87322686e93a860ac5477407df7b333e39db2f92eb9b84124d50bb5c442d05cb;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4a57358089f95c2bf1c676f75416fed8cbd5308ec5d9c8cb3e18c0fcec6a1b3bd576113202eba43ef91750afb1c9012cab02cdd581a619735393867dbd9f6dd2dee991fcf54287d15504d43db37eca667e4feeafd5cce5bc57cd08c76c8ab753ad699b8d54e4d27fd72259c1a4a72e8b8;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h95d9232b23522e36e925a42bc8e7f06b6c6796881f832eeab727a9c8671cc6ad4311e07a05e8dfb5c0698fa5d72f064b49cce9a47d62dd55327929ec1c5857b13250d605831d525acc7f19eb15a0c9ce55b7469505f074634e3f4ae9640c87b2d3f010cae05f05b7e4667a440404a9213;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h256798a5923b371606c858d2323bd0a1c314ef8cfdcdab97d10b98fa29826df526ce6e8e94fb53610c8edbfb499387472463214469689d6156f9eef06aedafc4979c5ab6bbb0fad37f7bef67f31803fa72db0a28e56d75e1359f78fe226ef28e5c2421a9acf67c3827a3bfa13d273a1a2;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha38c3da3555dae338829efd0b308c1b531454c28dd40039e49b9caf1b9e10e07c0c20d91c9d5a7eecf60bbb196eb8a590e2bbf5209bbf5be8a057a18886bcccc55c0dd5a25be677d2f6a0ab1174adf2a83d244ae2c1a9f26076c9d84ed8de608521a4d6572ccb05dfc5ceeea32915a9a0;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbca1ebd612ae5d6007b31dd30ea84a64c21d599314dbe33a138a3251589ac1273465908eb56161412e552408bc4252554eda2ca6b103275a31a857d233a85558193742f2fbfa61bd5fbb9639d50085a24027dd8d02e504a8e296e77f00ac6700164394923917c31473036c61e19a31088;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8696beb68970bc205cd79d72e3b456ac63fb7daff8636d2268d9ad5d1f14d0e1501747c972cbb6dd1f23d776ef4c1a548237227f763614e571f6669eddb7d1235f76ebfe50e68c1ab39c48a961706fac6a798aab366eb21c8daf2ecc5c2839789381ce274818ea48c4ef9ff3db196eaf3;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h72e3ae7d092545716e11ce468470dd09548843d4b945987241bfe822424b107d9a97afa35c702313c30955bfc5cc9e3b32a52de086f9de154055b388b81897010405dacb03cc5aaf7ca5c2a8666e1c92cc698738dcefdee119a47c2e330e35303203f4108d99ce201ee4d1a911557ad76;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8deba4badbe3fa07592374f7cd5eb23daa30319b4be6703f279e385dd81abf350307ea2d319414880cf0b205915c3057f3ff2a349224cf09121dbf5e42cf0dec12e4a19767c8c408d19276d0f87e5e2330088a488bb2b869ee35374c3b8758ae84a01df79c5632b663387426ab76f6304;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3fe4cf6eca26f1512ccd0ae4abb23ccc8a3835e48d56d7bb0015b839a29dc5c3185a45e3205716054c9378bec85aa61dedaede5c039f43af32bd26bd0b2119f84662f38de2e6e19b5ec917b1c898666cf41088f22cedd50e1fb16ce869d23924a8eee31f3776a4a49a4b926038ac67a3d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7502b83b09dda8909aa899b37cc0517a5cf8a31275cbee3386fda76bcff9a363b9e7965e79b68d014682775a87adf3c7cf29d491eaf4b7d8d06e2495c1748169007918a9bf7a0908963e40954c0035f4218f5219eac0a5196ad5a05ade6c4e477ce10da13369f5bc4e647e7cddd4c57ad;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdab7d4657a92e89a2044e617811e8c22343a76d5d48eff7d66f817ac4619db710c2f2374f973f695917e0102736f47c5cb2505ebd7d4aedce6ab6ca02fa7f3c36f181c3057f402e1ed9982f1ebcea4f4f5acce3eeecc51db7a2e8a8c64f9668a269b674af39ff0eba72b5defe8d716587;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h30a4e37ddbefcd522e4c17808da756d25aca0fb2e3feb880701231816a57635da63990bdc66474924ffc80f63488a7e02e3d0db0b1c643bf5c3d2c253a73099d6d944be8ce5eb5172b3bbc41baa638fc47c438d624db022f32984ad12de4b7e34e4884d0e3da6d5b9ce71b28bd2358616;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha9fc546ad1098ddcec1c25565ea0c3363658c3bb7c4939559b7de7205c203f5b54e395bd715a93a66a9ba9dd938a9461c5439ecf5093180715d1103b3afd4ad0bace9d1bd5e9a57c241051343630ea8ec488238344515ab66eba3a0e765c04482b4e696aa95bad3168ecbcee9936314c5;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4af9b5427de2e7dc7b334b5cb6dbfdf30efc825e1eacfbffdb17def88db100a7b2240646b82d373ca49ba1ec978f8704eadc41fe943df28cf9a9aa9f635f35cae3cb3cffb5c972b2bbd95fb4553be10e0d9f1d190775f6e76f97a8f33c248058858ed3c725eab5926789a0e95dbfcd50c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1b9bd8de08abe799701fbdc3984c59942b523edef6f2f9eace46ce4261aa60395402523b3b7a5840ab438400145dd59dc2802b57257eea059816214724284be0a5e7342f9a34ff3c2cae8a91ebd2857c307cf52a96889dd4863068494224221e3ce7df3b2f30af6e01c640b0eb77dc2a1;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h90dd624ae90c41da12d654372d585d7bebcb1fc8a0eac26cdab1f8c1fd76226411558859484320b39cdb9b3a065edd2f85539e67497a7f056f0a79d169414f13fd4bf813b303066d43a9c6a072a9fb3b34466df228821a8539ebf5b295b06f765226adccbc39fe9d168f80f6f254b43f4;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h580154cc1c38ff931ed4a8d0671dd9a7f245dfc5b4ccd4107ccb633cc7a2239aa6d1489faef5744d7fef0ddf5cad5ddf0cceb5df376c329b590b1f3bab612802a0a8d9f92b132b869986045b91dcdb630f9dd26fcfd37e43bf4495d59c141aaa585c4b39513a83d54cec3eb5ea9d71270;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb6d85605b47999ffcb4ee7051e986e632abf91ccc32d506e484a8d9f558a6fcaced058153578432b0b95d1d5e5da0d32f36a92ef21fe1c8efd2b49075e7e7bbb827e61c9232517ab9023eb8e0f500fe47481c7bb15c48f6075ad7c2c53ffcdd0c4b8ac8e7aa39b56192f18edab84c2f72;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb06601c679b074b4e069dc3651e78ee5b407a802adac85877862da62f6f51958df28dbf207503cbf34df35358d3db9a786c571b612ae3109acdf66cd5710f942c1d63cedef53a9cead10fec6aff339ae9a14b06638fb213b3c3d99a933c8a1e18b27b9c21e48ee7658917c0252a40b5e6;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3fa0085126939d9fcdb121a50a495412357608407562d054f4a3980cf312a6d2b46b3aac15990b2685efa889b2d2decb5adad0fe015ab8d838d962bec94142dc4fd50df3eb428ff6f1774bae7596dbfefdb3fa0be8ca8c94d32515fbfde64a44850555ccc9e3ee49a4b408f465b3416d8;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h24125d98ad0dd822319aadad40c527c2b8995ff63a06888bdec2e043be800a678cad1a90689de5951ea48493d5c02f5be712e30b884daf24618457e9a0d567351b9b7e39eb44e06be9e31bff7d9c04172899eded96a37f67420e8d46c31343e52ba706e50141ee6d70c9d57cbcef7f699;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha2cb5ab9ec9a5f3679e8d30cd0bb67b0a402bfeb1d91b495748dccb0c786e094a203a449e7ce13e5e8f7d5b12acbc65b50ce0dc9ca18805623ad6f69761845556b6f5275e0fea31888dfb8eec42aaca7b2daf077434beecd4ddefd9057646ed69157835d296d3ef459a876d8375054d9e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8d469e5b4c87776c7007cfe4e83e4e4d1b52a7b53fae1e36f6c50a3cc9329469ed4b150f2579bcf989dd1a7fa0ad41c83f106e8c72e69341670795535e5b02931271b7d83d504ed3352454ef0960820f7af8adce5b9026671e29e671f41902e5c2eb24343cb7284be3d71eed17be99f7;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbe89cde62ac1508d818a99a3e09919efdbb36d554445a94164d973be553c439a20feee307b5083cdf7bf9e031c3897b802260ea083300cee85fa8625f4cdff09f965473fe46a737f06a59fc56400d811ba9a7345750310f689d9843557ac0a6dfcec71dcba9c9818b1dab4706ed903142;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h72309b425dcbd61219c4e37751503e3fd4a3ed695f629d40121250f5433be7357c92192d65da52c52385e5c1eeeb67b9181155ed47fee0eac2c1f91dda9fe984073433249f766b823270da3a4d28cf97cc438aad4c78748ff1a391a283092e8a52c8617e1d2b5c809bf4cc5dfe0037477;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h30c9b716ca9ed291b6b932c734994c68b8122ce9feb52b3f0d52d152a2307a6647a820d65fbcf6a0038931e3ccdf246f795decb64afccf7a22231a6ab96ae885b5d6e7e7750f1f2040b2fe541d1afd18df688f828dacc1f4395ae2517a4574ed43c58799737586fb389981a8c48a13e68;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5bb1e33912d142c24a7a86d299431f5feddf9b6e9225cf11eadc75d194ea08d1be371dd51f0c6f9f06ce9932df2f2a2c7638453c012663beab5310a123d6035d6de10a4667e72a53601e5ea7fe573ded478a8295f41a6f50f6dc8372d4bd802359a82a70c6e6d00051d35232ead9de38;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7019c8a07e0bd41a0cc347283b3c9f662c12e43fe528f6da25b5cf85b12a891ccdfe1e0eb3013b65d968746b4b05299b63983048e7a1985d6221aff579c2e9ab7a656dc6e51089382e2c3eb4f90685672b0609e1a993095ea55fe8aead67beb03c343f0fbc180f7689bb8612dfe991a76;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h208a510811d2e7788d1c478814a0db4fa8fe774cdd8cfe8183ae5ae16d3182e6ce4940774a885808a68d7aa5783d2f9ade209ae7fc8759c772b78880c66fbceeafb2061be421e161c8a4a92775141050d72501594254dd050db972f9493d15436260cf3aeb4972249ee62462459305287;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h395588b23b48d4303b7943be5292e80f352ebe1df0fe91bc120d502856f2dd0214c55d814f9f6fc664a906c152c06161975f083be02007f77ccfcff11ebce47e3bc07cc8c6c11a1585fdea6065d03c8613d54ef47cd82c95401b728b6be668b41520a20b0e98c146557839f3eff66c0e8;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he76f0bff75c602f020de22dc1be5cfd29bb508be70b0b4129b3330d2105bb8332951b6c61d35913fb016460a75a592fed3a5672f97e1242155b1e0bac1bdd59bcfc6698897d47b021e4599c38fed2727039d9ad5d1e778329e8bf3c2753cf0fd43e6ee2ed58fa1048d0dd4cd80ff31c03;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd98647ab64fea64f0ef699b8f08b2a2d8e49664b2e5317f792fbb7cff9ff90327574151ccbe8748bc4fdb8ae5bd1e5828a139315f92eb61cf0acff76d82c2ac8e016f4b26bc8dc86a24111ca3df6318370c9f737ee99c04beb4e2a4f88d22cbb0b3c6b970947234552cac371682add5d0;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc86530edc38e9b0e927a8fd9a5c9820f04ab5d54e8bca2f3e07541e1e00e60ab5df8e5063b51bb56446b6bbdbdccc45c0ff154cf93249d9dee83bc453df2fa42d48e839c975cdc7da6c1255f15ace7d7bf2e5fe9406787134f8778b0128d237da33c21e7c58672d787b1b6702d8ef7023;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha931bc7edb1e080f1efd2ee19971ec11705844adebd3cc116817f8ecbb48f8f880d27611e9331b097782a8de8908fab895ebccdf031da32eb43cd8482fdebadce80627086ab90abb224ca157d05dc3ee98bb4ecaaf3cc0f2ed4918981d38f3172b2dbc66bf88f2f3e354be15c2d081368;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he2e7be427539e57f23e3249ae57d89d99193b9a6bd76c7b0542f9a2edb90cc73b33024149cc237df80e2f8db2b46559740468fe087feccebd9a7a3e2aa856e3c6f456a6600d27c71c3d9004dc3c830f0b54d7896c83b3986af96c1b990221f620b187e281cac7b9acf97862d36544a141;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4fbefdae06b2d589babe2aecff9b21ab68e5757b1f79b8a82f32effb8c808f0b2d99edafd63f808bf779d8e3130f4787bc452ea1b5fae240a6dd7904deac662e8b923d8e47703f9d6f3c143016b881d44fb932146132efa345578409d2bca860e9b5c3f5fd558e46bb38dad750ba336e5;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h14b6b7565d0a9b7d64031799e87e496b4a0397263055c158d3e4d99ab8bb9be10f3d7d223e6e1ffa9b934a7bc8acbbc76c1567366f964a9825f7e4d36442bbf9a6cff136eb0c2646f6142cdd60ce21e634590162c67ba4c1cc9267a3c51f665abf436ae2fd3b46a6ea13046fe2a10deb0;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1860e8aef527dfea62102bb2e24d94bf863f2b9ceb1d7ce5d93cfb62367281a65f08bda61d56d8554d289e1f9cd4caa428d73f7ce045ca3a7143feb450334ae3b37132e1e30d0c47b9c4645bfeb139375d499565128046321301d7fb24835ed31da0d9b036beb93aea231c3402603a6fc;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2986259b6147a5ca11d3f55735c6876e49a5e57e323c84173319e3cb4d2c4003b983a0eeadf2d6818082c1da3a8df6eb91d4b7d61fd01e6d888b97ed6fd22a690517acf646775e3a753357aeb1455dbba7ad7b92a0d9b6e22bce82f645ec8af4519465b20574a6bd3590ecc6d6bdfbb68;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc4adb9252fafda069fa541a09a34b5af534014565153410d77fcabe209b5e0910df09438efaa8975803916511a1929422467d739da34c64da37cf41e7c94675680869ce4f25617c43d5f4f5b7574767bdcfb65f31c5fb5049716ae062f9e461d238040225438bbcc1d39db77ab0289889;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hffb1ef4173ee212b809e1d586a18d5ffc4e01ef690b7006f4764e8aa9393e88eba6112973e28d843b4aff23bc06dfa24efad0b9506e12e8bb0a1ed710662ec48b5f6b8cf5df33e6db140959deba36d4a23c37073277209ef7886defd65c666c8f70900326ff5901a98cd5cf1132ecbfa1;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h21c7b4a561acd051cfc718767bb444c451a9dcbf62e521261e3073e1127b1d4d3fee7eb9b51dfe8b2bfbeccddb871e6907f015be73c76d12285d686e3bbc94ad1ded427f7172e403c35492c3f6b4f2650ab04ecc80c6f2cd6b8677ae41bf8e315f57916956f22127bd7958341ec1a0bd8;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2bd08ed55b492def894ab7e602abbb8b5127899ca02a30c47bfc8187bad98db5636850d9b8e185fa1d629f8264034e1dc9ce0c6bdff62c415461fac7e35ef34daeec8211891448da11ddeff1bc0277e42a737b4c762244b0ba970802982cd5be8d45c8b3fa1b16ae085cb4358b730e707;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7df131cc08d71577148a9ffcc65da3351fb9630063e53265373e94f966fa447dd160ec449465981becc17fa169fe07edad83d9017d9950219f165fb2b75857709b587de29d5b9eafcc75dfa3b5feb7a422e01d0e2d9d069bfee0c6eb924d93b111104e83d40789538e51ecfa27f20c6d5;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7c2d394103aa44c850632ba9ffaeb58c918c5ffbcb244287650be500a549e1cbca8f1bc0a8c1e97924b8cc90283efcf25267fbc6569b449ae49d4e84d5aa345bdc0eadb7edcbe77cdc44e3f3591ca6ea7fb1b4be0ef6b3202b5e69e25a686c73aefc21c2bba26310425886c6426488f26;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h27be988d500dcda0553b024a7aaa0c21c0710e8adba446d2e85946a9b4ed060e94c6b424dab0c97a48a0597a878b4058bacb49b18c7aaf257126ae8a1b037faf025dd436c3439d40e6c21584f5535f58729286420e4b48298ef4e121a6462dabcef8f12536577c1e15c56f12288646138;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2a88e62739fd98120d41f5ae28c95fcc5c16c7fab2d1181e9bf09d00eafaad00a6afb92e67629010df4be3b3554aabddf992c6598fe08c76b3421722d795783b38ec4504196f3490e04cd915d95ecf00c06b5618b0ffb6a39da88a817798ad6b5666caccc500e43fb8445a57856056ae7;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha943714b3dae26f99baac4e563f9e2d229f82d78d43d37b9f89e9bab64bf0c96217396da339de25e8f41a9a0fae3d72db711b1d75b2ffca218c851420d33fd8f8b46632652be6b6f53a855172e6858ccb249e7c3c08faf60f365e254eef69b022145e35a60e501d7c7535ac1734624ce1;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9c01b3a363e0b47c34ec8ce6063d46066fa600fca06eb0a3ab16c3dd3679c21c486f75eb441d3a4926dbf1e99c5818f8d896830186bccebdfb5a471af51e2541b6c30f6a2284bb4535ff865d17717f73507df6019fe97e842d2f27335c4de506d512dfe1c07031c8a7b40dd500ab53283;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6a3272baf6b7b358ca7ec7645c009794a6208f74b3c574601d612efbdbdf3334a32b8c638e131d1ea610ec3b13f25aa664cdfe3b8534ab723bd7b2d9b50dd0ed2acef74e5b4e9edae9950aad52665be106e25e1c179566ac0c10362f24796604bdca1e9b4bdc8ddb33f733e34260e5248;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6811ea7fcc1c30d7356afa1e63c91f0ec03d85122cd79e8a0224acb92c337a95f1f931bcaa6aaa714ed58ce2949c6c8253fc3f84bc5523ff4a6e66e8526be94d9015f35dcd1c456355c4fde88346f5cc510730772758dbffc40914c58565a1d7fc782cbd5b0da11d908b5967f02545cca;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd2b245f03ae875443746fc785b8b29e52fe73b13476b470bd8ef995df572ddbc62c82a202f3a37a6f3e986a76d1ef1653536a36dd312186b3982c70255aaf462aad490843db1d4def855034193f003e5efe0ddab31fe5ac854f1d2e78d6587008a04206df097b1f471ef1b9d26a372e78;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he2457707e90093e8e3fd343b939f90b64f9afc6a3297aa56125dfc65b5f30b197478751535db9187f1b05a88f310109dc03b4fc68c856a2de1df7142d851bd72706c616654ea684e588443a805108103e3b183dacc532fc641877050a71e0de108cdd6c113c318256d38e9827e5272b62;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h289dbec552064e271e07eadd7cbfedf32244f57d2be41102b1f8de1690e255560e6892df549f6ab93814edb5d0b09b5762b987f60836c73ca708b27983a8de05270ac58a5c276f25a7080cc4458e3b62c1759aa5fad23948ed114c396bff4194a97ba9471b4bf0317f3c63a3e434ebed3;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3f10df8d3fcf4c79672f87be5673767c28b7e35195f8797158c3c3b9cbaafc9e84c859ab1b6729ce0126e9ba68254fd49cd04cd6517d76163f41681ce4f36b0fbe621f0a2d0d04a963b32f200f3bdc74b7d2e46f965853bd9c57e5e4ccc678cf81158fcdd3096c46ec6344a33b138f85b;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6e0d040d7441d8a335b73c1ef23412fb363fe9cb7ac769577e330ce514652502433a484c08920252706eb383bc090cd47c1cbe047d69572e9eab3f5c8cacc811b49bd4ac9c4f4684748399a37393a27fdfe98c1653afd236b6b89605b8ddda37bbfb3551534d28b43815751b2c138c1e0;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hda70917f81f729305d040bc76b80ff1906ffe5f8227de2667743e0b3df778d83f8548e14ee83178bd11a3a4b9abcefa1562ea42f4c4fa460f6dd522dc8d581c0220e06f091a3e6bfdadce1444a20de91a1ff736bd5f2e9fd708ee9eb57afb3726963fadc3f543086dd664a9bf0eb4306c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h128147d1aa61817f32b0b25f86481b4fc23f8a9fc1d9edce81a351619d2bc64b49ff38e9524f75f2ef738faadc02ec296a9eb2248c5bb6ce9a48f12ddbb193b4b8b0955a00f5c75f360a5b89dde22a2b7d719b9cc176aada16937255dd8e393fc44e4f75a93b0df7cf23cf574307266e1;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8e81c10b51391248447fe4c2b32a86b20d7b7c99d9063004fcc1f765e00a9b270591f36dbb2dead12ef321131a271ac9bfb19c392eaf1130af9eadd34fb15c5a436cd646ebc7a640ff1a5c1e3756e282a98fd3e87bb8138feb036c9b149f88462e0cef9b2c146866a72aedef6bf84003f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he6bd4e38eb2d51f18b9e1d02443df6d3910cbf64dc2806a5db7d002595376f88edc9699c2957b36546dd44a8f9348f26883fbbd95c2e32dc105ec430b8c9a3ab136f46147daa0cba35af351d28e4c78c87378b74a3fc57f786fdc9f8b13a601a648326bb051ba0c20e9633b6f0b474178;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5aa67899135fd62dda13bee93fe0b90351c7d4812dd54517172753493da86594d4e5e19a8d0539a8c0e569c13ce0946ff22226cd9c85330aba7a42d137c7167b92dae6de31a83fa2bed4165787f44b0e8eead5e3e46cc54fd90cfd52e25891cdd0ebe4e8a9e7a3537c9dbe8c6c9fbfc9e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1d68de7030188d5a23f37f2a976836a8c0f3f726ec54a7fb707175a4c34e1d8f05a9c0c50f94d325e7cb9769d22abc9da57fe196d371f84ec27e6a1daed8f9be197ac94c5b3c40fe99501104ef1f894a99c871ffd0b4e4a5fcc5698d4fe1d5095403ecaef8b373fd265d8f0098c17731d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he3be018546a479c5f5ba0f8e19bd467267f3554fd30768ea953ab8a12792bcb2012d665694dfea84044a133d804a37bf49bba52033fa1a84e8ad273103dfd1a8bd725e4a190b91256c7f52d511761621180211dca15b57a78b2460887b264ca59278c5e3e983028733c7cd2a383456df2;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h805d27029bb0820b583b55f3046b548a28c637dd3cbff79b1b96632c08e5ffb13b48667c2ba061df452cf4954159fda78556214cd9336e8967793a68e361b3440dd77f211c9ccefb93438e5cbeb3cddc484014b5976fc6179ffb56bd090d8c2d79d2e345368451eabbddfdfbf82085ec6;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hedb1b18a178b22877423216f6e9b3513891789763a39fd1dfd77b91f718a35617ce0161677ecb2e1f72905b56589e77dfdce31c85279bf00116862fa264a259ee4b7f68232a06d5c5d1cc3a4ef8b1b0389c47d190c5a0f3044cdb5c9982433e6e458ea9f0050eb939aeef69b51a8a2895;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hed9e8e0b3140c0bb1f22e9f67c6663de18e94835f8fe6f3be721b97bd87afcca7e07a215d4c463f3f88faa9f96dd5123e8eaf49a12a7ff9c2d2e19bb564b7ecce74e26d526277c6589e3751a02cd7830b9954499e24404608c247b5aac5f8b264ba0d871473667d739a7dd4efe806af4c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha735b801d3d22f1bff22ee100f60adc490586d6e69fef31c61b0de2dfd5a1f8f7de8dda85e69670cf60ee739f1f1daae30670e0f1a57ad43d801b1fbc9e864b25d141748a98091712b97c67a886f565930cd8be84e75101e9bd52841db24d11450fa138aab2156e1c01b92afcb9ae6793;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2845a30dfdc385da07b58b594a24890cf1d14077c6898450f00a1691187a929c288918ff7df5b0192eb2b60dcc45db1209e3f3fab59d0167f0010fd9eb9306aea7088180cd7f5aa30401e8c3bff68967a1cc80dec1307d9b841de85c64f4ebd6cf1ea1ce000ef5dd4cb8f5f1b7893a6f1;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h488decc51361cb3390bb4c8e806161d0842da09ac2f22dee631a60b8bf52e1a14d223a3787dc0cd9c7bd7f353414beeff78fe237ee54426f049e8103ee27676d5cb30218f717a217a7c5127a1edc285049ba21db71da0768fbbc13f0ea4d73243781e72e8391f063cc9c34c51b917ec1b;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc4f6bd28fd98ef3f97cc226867cf4cd605a076a2d9c165154ecd3c7fb5d4dfd3bdc9b8a712a8d0cb8b9f0389fdbdf9d74bf82c5da2bdc507f0e16174c0cf4323e10855b5055942d6c7a3bb578109f8dfe9b1b89bc8517376bf890e6ca3ed0266e3f8f357d8fca7c58daf780fb7625079d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd13b1deaf5f0ced98a5d1efb80fa188d840955a896fd85257b9e78adfdc3f30d17c598f56b43a73afd39775a22986c8c69bb75d95d9d8fac59ba230a49181d2642ba6bd10ad7c603a7cda2abd2e86190c04e225a5f25ef8194049fe4edb46c37e6835f781fe768bfcff6f761ae990fd13;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2002261403324a6dc5c2dca47b1cb139b0f8f3230f34c96f5ce482304c4f3367d0e7b209749b4868a661c71145b42c833400f0b0b07faf7c00b9c7484323f73324d4671dc93c7b767a7aa261fa83ce52525985bd00be77aee7d71b4a876c291b553df22d6a765b93b88b0a6a9acc477f8;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h63c16005a0fe598f99470c66da30ad93d4b7fb4d3dbc6b6c8a69530912620385f09bfd6aaef9d286721d1daf10a377e3ed44295d2e005c480acec22fc0fd68439e294f69642681a8c452cc557ecf6b50fdc96d6b2c95c9f8e5e340b7a9e8bc085753b4dbb648e75f36c3d3a573ed281ff;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h87278beda5f1c64252a5c6eeb391495ac016a442414f94d916c612f737bcd830b532c2965abb43a2e5c0e200eed2c07fd79b244b48fd66e00f8206e975cede5326873736228d7fc28ed2873441c8852bb084c12c6b430ddb96bcd9fba7468cb85cad583fc4152346503d0e7bc4856d3dc;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h864cd526462eb84d0edf2e1fa72a6cbbe747789f122ee8ea2b5e7022d1822a4b819c8178d49b940b3e4fa9b0198e3ee883dba59f62706240e0e14f75c924b818072b223413d267c1b006a4806b1b36d67a2e2537215c9a14a14e4c733168d978d7b9c9f5c8a6927d45262da3e014a456d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5d628bd75f18f19242e07044fc65f97858a9ee5604bc744e832513f3c504901fddbf766cfdb88b6c717160e13e7464876a3ca6981c58f6a5a8e7cf37501d4b66186a7257aefb3a5edcc9d5ee3c46ab3393fff4741f00759428caffdd7db6fb1baec69fd6708cd41efec27c9d31accca8a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h22bcf8c7f52eb20abb83665d4f4ad8e043ef9f4fdfb9536992b0566950580845b8b7ad77f78ad0a7b07a98252a78107668fcbf08a9570e244de0e13c34634ff6a38c676bdaf83dc506a7475ee24aceab0d4a30a09f9566d309ce42b9059a08e892c3e36b76f58862431c3faaca34cbb60;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8799c89b1c51888ae7ef03f9e44b1e835a6349c7b4dcccfe90ab9965cb97c2e342d98602244a46b754ef4437af75facb0626f34aaa05d4d457c73fdf1027f0837959214cd5a382437cd10085d09cb95ed2f40f736b7ea7c8c792e697801d19fd543b7fb240015bc2625cb1e31d85d4462;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfd25faa3cd70b6f75873c3a52e7ed0adbe59b30319d7eea45e073432fe84db74a7654ee708d1751a68bf7cc2b39c9afc6904c2e165a7d1bee2cc2435896e539523e184d965510a8875d6de58b92dc168fe46784a642bb44576924fa8725229321f44d9d5240c7e057fea0908f9202bcc4;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1e5258f9ce0aecab954b09f64a3209649ed83bbb791f3878a6c34df446eaaa3342e11c6d7eecddeb92bd80e5293ae706a459ceba0636966b9c7d60e674c69af53570d4724ee5e21b9aaeea8821c2a56aa77df5db26d2b7edaa53d6d816b9425c6d5fa021f6e5396c54e362e95d8678926;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h63959218de391e4b8ca1d3f053cf88d777fae496360a3fd593f20c365ec5584f6183534a43f8036b9d966c24395283394a54f05d48639932adbe6ccfbd11b6a1f5f6170b384222016c911a98d7967b64f84eaa34dabeca9a4c7fee569b2ef4ea187943027fe360486ae4c10651c3e3f53;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h44858e7746fbdd96fdb8cd21da271b053880032022f835b0f6e21dece993585d8ae874b5d35406bd61e89d8eca8da744c3f1da1a6372f027d99e3d7eb882d912cbce9db56001108034071783c619eff0647e48489f84def15d3bd27a26ee73abd1344c63d44e573edc9124f87b0aaa24a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7430f62134b10d3ca511d50f128ed5d64019e418baded09e2a789a8bc4d6c4336aca4d544e36b3711677cf841d633e4e96322bd8ce6c090f5c8a74587e2b8333c8111e30be58286baa2d02c5ed437477efb24b5bf5c26bb37265ec7190232dfaaab5241cd809b6f677c92edbc3ddb0d8;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h32faf7ca59693fd0c084daf38ae4cd1835409cdc50c5ddb4e95321fbdc0b5cf7fecf637583a75358c46a11aba5001ee11f4e5734a48353ab3764b63f5d89efea188d25839f30a24cf404b48587dd570861977dbb8b170f76def72006f3b72e7ac33b43339ee6346149f20e1dc8868fad1;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc89dc1c06ce61c918db7724ae3172ac9a73f3bbf1fa0ddffe5dad65286740e5279f9ee5c8f2d4765ea059799db4ad8ae8a1b756fabe0ad9f68a1a47ad3092ae61ceefb6824d63379d564fb5350651eac7fd2a43c2b509a0e2a45f80252fe06a2419fab5645962f7bf65c97f1f29cdbd47;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h96e4406cde78084123efef69cee7426cfd12d4fe286f21d6eb5859b7373757ed9e918c0f79b9001b5a9e54beee9cc5467cd3ec475c2e9fb4fe37447d3805d83aa005587deb2983de78e0c2716574d8ee81ac0d806e78bc4a99b45e55ddbde017cdd76647d07464ab1f023dd0c8501764a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6e044f191da9c64d6cc0366dddbe15d4fd6edced61108d097470db89aa6b0989468ed856213a28ffcf47a2ff5a642d555b2a5d40127b3b219cb9abed22deace6c1919b23ff4ccc81829c81db45a96b03578913922d56aee9ace1643df6c03250a59ceeb18e0a5f2f39d8558ac4d59a43a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb3f57468bd12582af2ea59eb163a03ef578f70970a0ddc69c71790d676af003571eeeff5eeaa792fdb4c1a991fc44e31f77fc323ea19b9b2ba820eff44c59d07ce967f7730ab9d2dc0a9e5473e5ee0cf358762eb43f4dc320e621ef727736cc0a7f40d49868a0c3b292225228d787b805;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd9f3b1a3ab5b5eb1b22770686cfb2a9b6ac130aa24a32ccac3772fa1cf43b91b7dbdee996cf5c46b0d17fb8aa8e1554a04dba280660bf9f9907bada82198a1e79c358e3f0c7792648b8ae2e003264ea1dec837cd0ec9e5d20216003c966c4869c23511fcf66f4f43a2f4689d6292a4f90;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7e5e419adcacb11e6254a8deb2cb0ed2952ea00633210208ceaef70a905f20c2511807c60b5eb722df68395145d4adb72aa802e9305d5896aa17ad36b15dfec23e7e07da1b9d7c4e3628d550376ca3bfd12cc8042f1d83018ea29d99345f9aeedca87c37a5320b1b83bcb63003bb455ab;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc2f4472342ec26fd5bc5c0b315264eca96398c3ae1ec723b21ef9af5339648fa8f56b2fa59e8a213e6a55e1fc4442f6edc864279d2819e9753a751624f92477a6cd779b1256fd4211adccaaf5b08f3e957a39fc35ba46bf1cda9013cc71e748097d8ba2dd12c25d2e3cc29b8b6b2861ff;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb96f6bb78ecba4218d689997b81b14d77710fdaec4044696c5b3347f44f8d2543d7dae50226a1a6e6f1847f4329bc05128bb0969b4b81076abec3293e38b631a0ff8a7fa0a86b1158e3842a595587a187472ff37b0b8ac878a6f4b9e8bf4f1d4dd1f2466bbf91f1759e01d5e29e145fb5;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2d6fe846e2fdc5698b98f5fe28458745e92bb48516111997d977b784fd3b068d511af54c5f5e789969d8535923512c94e5e91079cf461f4bf5c5d08690e49680b4a22f0cfb9f4cc0f4099e95de4921c1cafb59908c4fccf396fbf764876b7c11989146ce6cc1c1c325aa6f161366d7901;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h97016619015c4ea16a8cf5af1e2d651418cde1caef8025143e156250ac3d24f2344b81026cfba6136dbd9983010a976682ff50330360d1e50c0374332aa834d8c781ef2548b2f0f2563ff1c413d2f2cda42aeffff6710f73873f792138f070882dca529db44fb38b23bc5031a1259b736;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he2490338381bf5dab3abdd68fe9076812d9edcdca039db96559cf8d5715e362086bd83dd82bf7f95581af8e2b56e41b2a0b1c5d26d9cf892b2c85e723fa89d6ef341ee0eb757eb7965d9b3683821fac33e013ff0c8eac73d4e772a4158b3ccdbe73fdbb5e35ba58be1dd253009293d897;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdbb0cd7c7e4d1016a5a2429f3cc1d9f01364ba30acc4edf75d39c4e53c7b48cad5de88182fe31e59c745a4a924be6fba4e01e2a32a03a3ec03338124704d5c2f8d649bc3863870d3c4fa3d97d2dbba334da95108b70c24ff9bddf2ac0fe82dbac474aaba21b96d5ee03faf8fa62df7383;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h81783244d9515be176e7420f027025cb63881049dc1eee4507387d91f773330d9b00ab8df6610a78fc0908609d64e189853aee47899ae3a7d335f83c97c838ead1f25f5599e187f4d7dc8403260397fe9767edcb6aba8ee7c8ed77ff9d876d3faba23a228d51ac024bf793fef833f507b;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1db34b7135525b5851e1172d6c1d97b1ce7da5be5b5fe27d6efaf902ea26433edb93b4047785eb34b9dcf981bf7ca24e7cfae13547a2906fbbe07064cd68a9ca72677c2b48873fd77d6995924e70b17a68f211160d822a23bc6d87494b1f3d4ff4e348bea79aee89b3eac1c79aa5ff472;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf8b4ee36c6a7b80808f6d6acf6aea384b049d627cf35fe4ad1714259d9ca52f7ef6a1bbf8a8a93c9cf0e1180349c254877819ae0468d48c77425c0f8854d0d3400efb0f7c3e3e562317e9df271a780cf7403a45d051ed9ba6d93e29ffb9a6532f086723dfe8c960cf24952a4d9be5dd7c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb47f4009807119b00a9bf8c70bbb0a64fe6e09ad2a590dc7b05dd764ad37a13620156345189c009d6f904103b1483940f8fc87f151e8aa804035805c216677165e74a5eea449de71628af36a72fd3e3fa8123202feae7314335335a652287e912dc6fd2349e439d163a29936e3a76253;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc927b8544c5bfc3eced42289606fa386cfba754c56c19eb4ae36d658a1f24ae548b9923386a221bea89636ea7ecb60cee055689f5f1a002bb3d62dd0e6c008102d8bd3ed92418b2eccec7accbe649db3a391f640f53d67e550a837a6e3fdc8a3ce8ae1b6d69ffd18db73dd7ec695ba4e4;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4cdc5e8a9f862775789455e22820a2abec104b3df8a03a3cba5d8fb0e2c3a1f7808aa1f4acb2798b94a9622d94f35f1a35a37f0a686fe89bbe6a0ba2fd3787557582a5b8f85e95fa2cfd8d5ac3535fabf826b542f0184c195f517ad189e2ebca0fa1fc7e92aa50fca3cce7b19de3d43fd;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he836cc76db9b28a48a120b42af7ba428afe5666b161c09501e1cc86cf9554b217ded4902bdd1ec8c24fe1957d3a1e80b132ecf6b1941746acb55eb64430a97d05af095d22a725a63adc5a8664cc2f3b856e37a24a7f9d1f964cf774f7f9890099693c33cb1da1da116511ff1b3ad741ff;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h33cfec3dc9cef93f037b293fa4631462f01b7ac79b70f5f5e3d0bead421f18f49a4e92f9bf411e62c87b815aaaf7ef2a0697215baf5f899863e303ec42bf0f6a5745f46528b5e0f84be289b36774ea4f6a10e53ef8c227d05fe333416b1765c59b9bfbaea6fb814f2fb7ba139a4ecaf3c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h29eff8b6aa43735ff20563f9c2f98f727abbe3b87d51cad22ecf282cab502aadb8a72f1c69f43ec7dc245e890d91b8aab820c6da313dc72d1c8f94cd3ae651052b794421716c36310a458dcfa2c811b261f36a7014ba8d901e8ef245a5b92a36b6ed66d16c59f14d261268e356a6b73b8;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h73e7e97e69d5aec98583353829d56474102f0f790fdc8522dce83f7a2fb2ea75327d7da5c138923daafca58b3ad5a71f9456d3d64871c753b994b4193a9427759ada8c28f8033eaea2498ceb7a718c51addb36f073ea01b843f16260d0b56230bacb26467503401504538ccd61b1ed556;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd469ee50bc85f9e24192f9836178a852cce864ea6289b2cf6c3708cc358bc1abb4ec1fb3524c25b5e3d8c93ae617edff8aa5909fbd64c732169473a261c92dbab0d595386ddb9aefc270aaff0531c038a8d24b0a351be5f707439ebb459c0d5b027f78c996b822b8ef0e1b692353ef7c6;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8f591d95730ee7d18dec9bc21833cfe82294f7ace55cf6537e8357be519c2d150857f2293166748df9c0aab3e26d07d88cb6462f554367a266eca60fd069292c3e94654d13e31cd9acba29b21a26a5a92361f5d9ad26b8c94ef06a19d668749746e90f4d6a0f6f7e24845babec22404de;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3f23b5e929e6c8f0b76476abdec40efd5f54113e80311b8faedb709d7bc5f5b6f5c488a4be6deef4656b9110e4c2231334c33b2837b720afcf2f9bf9564f2fa50fc1da3762e74a0440005eb1dfa8011591a09ee81d23492d0922fe25676bacce8ba191329af08bac895e4630d18e0a413;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6c24b76022b034dd7fa6c2fcfe27a29bc63d11a6f12a18258e54069a242e85da60af81ef4f897ef0a05f0b7f1b4a619f675d84cbe11d7617c3a55f17793861a8d76829c030fe6431d3c40eb42f16071d4077ed16d43ccc0affe2365faed32ec686e92488d6111dcd942745433261cf9f6;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdf81d9be23c4e4f62d35db71120000889dc4cb565f2d88ab593f1378cc99171444f95e58f05a254a025a409532ca065f8f3e20c04bb358bb8ee116cb0b4eb056b8dd7aec897340d828e2af18172150e95a5af532a4869733bf43b3bdf0d848a8ef9bb1457ae59c034d3d0c7dbd1a0172d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h18debb1d8c29aee494efc61d151f38640f1832641a53d1f569d8fbc5dc7f261c27191e0269133c46a1a07560906cede022cb05778e17fc19f109d3429787e899de2f9206c158fabf4d94af703258e826998db42de276c0bd884ee257d48f1c28a6f3cbe23f65437f486db492ceb9e6536;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha14f0bb94e186596882820aaafaf24a2397fa64eb76bdf5a9df51df5c5589459297b15258b234314f798a17e04d599319d56ea81a874d35a81b37e60a3d93c58fd8bb328af63828429b20b22c752430a606f4eded1d39141af52d5c0d3a8dca2054f9e1a00b6734f15b93ef057583355b;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8209fe6c06e86afdae85cb7a12dca0f3a20bd46c0670bec2de7924f118f75ab707b0a73076a76264396111b7b731b26fd198eb52eb754d4ec0d45c596f4c98fc33bc9a466d7c8956d7ce121973c37f86575e6b3a4cd2c71b3722e076de3d981c7ec96c22b4bbe9e5c81cf1b8e4e283108;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h64f961c2ff13f58e2729be83797a8b6bf064a0ab870657190a443da0cbeca5259ffd1cac438fac51e5e3d2b9d8e9d05a44a28f2c477c61e1bf0764d5e7ab32ddd8c979745134b229e12a5a748f5a278b6be239d19d034261a4a5457e6cf4a425e1be118d1010b1df0450a68224f9e5827;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb472d21e960611d552432d072cac7480f35ce4370c4a4ba4ceb73c73631d1c7a55465e6612185b358b2e2fe36e7302907b0519fc2e3176ed550bfe6c16255c6e997594ffe240289aff8976366fa3abc4d583b1ca5264fa1d7177888cfff7dba47a42ee6c20ab0c526af1fc04f4596cb1;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha6b53e80befd962198e7bdd9dea78ff301633e52f7d09c5e6801cca1464cf16a35ec9002db733312affde1c4622d7d38ca31956e3e41d31234e42437ac077a46450113b96c82af7ee8411428abf55f6bc508e0628bc9324d7937dbdc22b9fe658e93137e8e8017977f91dbfd12c5240f0;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h19ad8449721cd41cbc6f1a60ee131b40878f3d613a0605ee527f5a51131ab952074f591227691f718393102f2cd66ad860044b2f28f609c50a3ccd9aa8444f9e8f09bfe968349f0ea6e2cde6d8f1c77afee7233acff52ac8590fb3939066903a92335685b4c9ac62b8f3b02e76e84f654;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he20e78e6d3d3f2e70ae291d731536d6baecfc199086a523035d93fb185d8a47532d7982719a4bd5579fa22c774e3e5f55641c4c3d61da8f117681002d8a78dab3880cd8fee1377d8b2ee3265e03d5289ac73b916807295ba0b5753ec77040c73373f090696a0cf25cf0c7efa3268c1c11;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h116992789e5fb0067e2f28d679e2438f7f9a46c7ca9d1f84f58b3f2e6e03677b550566451d1b3ee2155719cde427af7015dbd7329625770b69b8d136a30b7f6009f2a466a203fef1e46d6885f6e9c54c2d8befeebcb42bedc023139401f60c0a9ecceab9b8d3821d4c56584763506ad83;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb3ad712a098155f71b959001c7633c5b86f306ad83400da39c8a568da6e4c8c6aa27fb42398499c44e179c442ac4a6ed003214cfda8ef99b3ac1c8656b67db7d48deccab9d96e88679ccfdd8438863ab2d96fe8b8417573adbb478b6611d55567e4d2ca8604c237f26d6578300c56867c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2a00ff6aed8d30d94bd46f4d2bad622752bee9fd768d4ea9b37b6008c13b53b383b69e66efed3d5091836e46d14684ef882f8b22348480f3c96fefd4b53e5f8064e695870243ca0b309871738edf93219e6a81ac45d1eff3f9d20a3b63eb462e6e9870ff0b1aac817ef288d145559001c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h369db6c44f84449aa660927337fc79ad49cab84239ce12c64bf628387e21dd6ae778f593cefe2d12934e6b6cf4d6ab73e590b56245b272a4d042f98942a2b865dd3e56b219cb8faf7dcb835117e9252ed21abda76e0c0d634645c3f5f33dd3fb4f1e04009705d33fecd9766a0f6b976d0;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h524d56300192d1bc82df005b560c99a99cba7d80e192bf429b8369d60261c9d9dfd0de6d70b999528d4c119b447141d36412a1a7675b0c3c9bc02e6dc5c76152d93d9df111b4ad2f7277f61f8d051886f11a38584964144c136ef033a316c7604fd72ff948e28e7d35a3499e9bc7d33ad;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h76b77808aeebfd1a1be02a80dccd51a18fb4c8afec56d42a72411b6e412bfd45cbacd8020bf75fa9dc7b6b5e3d8fd4fec707eb3bbc9028f0a85a5ed22a128c86d0ad6bb9cd23c444cfa5d321112e857c578727d788faa5409d49fb4373f37df7c6a21a230f73b5a3a791e7922dd99b1db;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h10cd7b5d10e95edf26472029a36e717cbb11ab044013b88b06b0bbf8c94f552322ceda21936141970db0b071e17da692acaa367c0d2d3dbcbb72411e6fb0b4b74a760f834c5177243d7a0979709b97c5fbea88ec987d386fcae4a6fa0bf864b50197e58b5b5caf7baf99e9caa846bf319;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4accfc5b3e157daf621c8e77d671e5b0e554602caa610ba745fed80655cfbc7177db357ff90d464ce14a32870d6de65e19d261b886dbf1943275f70e60ae4db2989d211a8723573a0c4f2541aa527466b09cad9f4675b15d522e767deebbf6cf05b200d5533249f0ba8898c6af2d4cd37;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h42e1b3f96950f3a1bce74a468560a0993ea71bacbcfac6f60db46d079ee9619a4b2b87e17f1eaf0908fa1a15b46cdfe8b3c3581217604a0d50340a93028ceda2d4f3b9a3e0ca5a1a760e77946c15ba3a190c4ca5b474fd2594dc3d40c81ece5bc0c751eda3cf719cd5e783b5eb2361f7f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hcec7606238cf7a9a7e977b4dc0c84ba496f08f6b96360c332b8bf38ada33aa33348cb47985fcb8d0986c6bd9f12c3b26265fbb98f2dd02c5cae5e46bd58d116f19312991bd100e142c0cce57d9aa9e86d0518c753f86a2a0141bc0418598152cdfecca78d8aa291198b8ef04bd4366c36;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdeebc69a9acf681c9bdc895aefe6cdccd80f9e9c93b71388b58ac2985ca17ee32f1ca7e81d780ecbf43f8d5d96c2d47a0719cb1911b28c5863218588b54fa7ef46c3d177d3906078ce559d4b7ac72215308ea838cecdf16bbf33717ad011896eef95b779471e36d0ccc49b429889f70a2;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc6cd41a6782ac3376970736fe9539d2e6c3b39f9ce4f1f7664f46d11c432b6bb00821f53756c759abffccf407a5cd38db5d52ed12f44827209c2c44d15a6f3e17ca8543e88b87d0d011f7e9697329387b42919665cd16d896cfbf3985043295f53efea9d0b647272d68a7e78e15b7d5a7;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h87d93d8273d0fcde5c3d291ad65126837d6263b38638aa890c383872114caad3b143daa2076d215d752efe71fb29a4bbc023063f24c77ee26c797af9c21e226431c037f40db168d380cf9352923dfbc182559ac5a8d332ee772eba28698aa3b12e60c2b4a0a6b4c5acdaa2d84a4bd2055;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8dcb31cc94b0d86e6aecc15d4ca000d7d9c6019f7cd2b90293f3f3f069fa032aa1d81115e46a3417c32545e78b0754c0c420d5035a22f4832f7f3f244efd337b646dbd99d1afdb553677aa41e96f87c6f6e85132d2e9e5bb7882c4862cda46b5530d5aa0f4c57db6c7f4cef6618ce1632;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha179127b84ee2f2bb096ef7c0f8b6d739fe7b9a079f8c5ddfbee3cd7bbe66283017364c2daee9a428761ef5582943afc990494303dcb17ab3ff56e9ef3b45f3851658cb85246ff267f210094644bdf94ff5b450d5e12e62577f1ea8bb2f71ba10a4b98f6904fabc742c91abd509af8c54;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h683af7e9460915f17df8fb31c3b40295d6571dd997d52efa3b4d8832f6ef67e0cfcc7c942f348efc584b3c13a272c3d2f696479ab74eac58523bffba4d449a466ce53f6da928d018c042557e0dcedcdcfd595cbf0abd2e412b33a48677fcb9e4a43b8c529a76279e6c5b0a2bc02bf0720;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he0976d2a091afe18f418e9ed18b6983729dd9bded0d209591e8c6803fd4d40189605749055fe6f3e36fd8614bb5c4b76ffbbca8bc43162e5d3f1c01eff28366a38568ed63ba9324c3a10d27edc59bde8cf4d212def1b1a66c1daccebac5867d4dc92032c1028ba75fa804f654dd1b38dd;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h57e3425170fe50420066d98ce7d46ac1af9181f0d5fc07fa9ed1cc52b116fc78385ab0699860080b8aa33b01d4ed8dc687c207b5285b7cb8aae9e110bfce43ac1f899ad4737a8c60915854eb618a13b03c1c4b533e6c0085a57d0f881a0922f6051ee8b887b0360e7f2825e7cd30ba571;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7e61ca86aa3a8e28155f5f43e4b94e2e76812b6b578d95d2022e8cd6166804f07db0a8a2d03e181a4beecc7f5bd0ef771ccb2d46c04c0dfffdeef9167f6143d85141f9adc95358d0fc0842bdf80ed9bcea849860170bc3917b50817229cd2f1a39b6da5c5a7df532da64b97b7bd8c5c9b;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h32107ab970b11620f49c5de6e8fbe73067744918f4a651324c4b47c02b42c60e4432f340c41e575102a0334242762d53908ccd4559bab2895689450d4b5ae9df42550abaeed50c2e8a79ad8e614035170b199d9db10b74f213ec6661a4d66328852d75a5e0e2a33a18b4ba4e510ed9ce6;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbdb2b38dbf06194c3856c274ec6b6673302800d3d9c91f258c01507638da463a1bf860e26fefb9d0e9ea5980088171604facc77dbdbbc2b31f00ac1b875cddd6ee776d32b9d91c88bb8eeace6532289a5084f3c0a62258bed15114f93848529f0a898faa40c5fb76807861420dcf7c05f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3e393ec7e448025af17e5e427507db1888c1a0418dd3552f96cd785e85c83e6e0481975f6e68f6b8091a87c3a8fe65b6e597048bb135d9c64176c3547df9bfc50c5c2006dd11497a9f398200a6fe1329ae2d78925e7ab8e6d6598069f20e11d85a75794879828b61889f622de6f1e7421;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hcc632ef43123954aae69ea23db01db4cbdcf183bc81a42f9cdae02ff36b3f0fec9f1e9f39358ff7ee335f253642eba876009f34dae18e892049808c6b9cebe7f7517d715eead660d2a41c06aa25cc16943bf1a0170732e840087e9c8fdc0ac40c9742874a69dcbd377b474835ff912eff;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h80641f378d144a0989807ed96f92387aa45069650ccbe8607980b0006c729e689ea64b86ea10033cba54b31cba4b4262b08027918c0a0199ba4ade7749db298a8181986491b0de1b3c4a079ca1274109d49a8515864f51ea80284cd692678bb88fcb6c9d00ae73ab76069b3c2139401ed;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h28861bf8f9b7d92c2bb73e6832953b126ce10c99c4b1c19452e2eb7bf15d2cd95bd74d4e80fd7ca0d523cb695850b002e5c87961a815e82acf242d9c1bda084e36d898cae98f5e3942051055ead0d11df287a49384ef37c14e91ca063799b7586afa37661c212e38a317c2597d6f9fb03;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha92bb31a8fd9a3568ee7a8bb2a269f6949d2cabea7c424b186a77a73d26306071d4ead5a0a5d51890cf6b8af0379300a58517a317ab10f64067959c913b38be17cdf55c38d9aac7278327511f46ee02ba0b058580be549c737f4cc4e05ff4ad3f58d93c924a11f6f04d33f45cb0232e03;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb0a6ab099796f4a2fb26deb0436515966df5d45e75f598e9843a48fe335809dd21cefb1fdcdaf39464f7fea1c6c8340f2f64b3dbe85824a3a54fe9ab84a5d3c76c1501b73ba7c4bc2a1fd776d89667c0f88468c833da74559cebaae67ae70e097b3d70f6e67bd5ba144d195b26a6cd6f7;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd9482356ed44139fa8b92e280cc1182a15f904efd65047d29562ba5a0391b02d47911ebed9b03fcf264f3f5a25fd2335363626f3a5be8579754b4c730817d50d555cfedf7bf95b0dae9e5227f7b305e2d5b35a37b7ad56dcb2981f31b11cdb9f6ba175677740d3db85c9f6e86bed17132;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf8c24eb587d8b5911211b345b61c89121e0060e96474c7d972118e1abed32c8eb545fddada7bbd1f6bbf94a755995394bd74baff27ec243330393ff23947c941dc44e1cf3031534277afea2143c30687998075a53638e3aa4efa6803841b8e1fb78e93a4a9e9719e91d6d0af3bc7469a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h278f48abe741760310f63178488e1b82976d610ab5eff13840cbee0c5713aea1e12c02c57e0dddbe6e9c01c8bb1f656eb66d067dddf9e580fb2b5e5850678e9ebe53d3f68f9d1be397b300d17c3ee302d6cfb049d17e7cdba0d4d449d202cc5e7092c1cfad043ff250941fdb0dc53897d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5645326d451589bf912691a33bd0b91d5cb141059760de33b0a8d59fb9d6d975898d1174c55146cddfbb0ea07be41429d6bd827d20cc6e5d2266a3bc5fd32a2f0df2ab3c8ba704ff8568f64faf471bcae3efd67e240d6a7e6766728d89b9bbd43bdcaa567138f0707f4f63873dc016981;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hcfd53ee903fd1568beb0af62cb38cdc122c2ce97007d38075407da4f718f08007bf9278a8cfa69166db79c0cfe6729e7df0364a10681dfaa47f6909a27e3f75af18b5f285f7acc8b46fb6051de43bd8fcbf6b2f4b14cf122c3591887bee9062dcf86ccba59336b618b7ad1a1fa02536f3;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2e74d95c9132a9a6088354b65a9cb19670224229d4f20ddd43788ae23d31ed54a9d173bae6e3beacdec3c415cdbdc6a8294d93fbb9812d38ace2198426717a4e6c1cfe773f15baec9ce569ff94a50bc76e6bfc05d4b1981745fa9b71c8ee8b0bb5bcec1d7c1a89b151c0e2c96d01d3ff9;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7c6355df2ebb6f1e361eb4597f36c4468d705eff4fc20f89b8901fe633c81f7740c296f734aaf32d877471f63a81b11c1393feed5d5e5d781ab84622f6a5f7241e6e07d46fea2427d745a4bdcf5c9e7e4484aa917d1d406242b474721d1ea39e961c3fa838086671d2307d9ff444708f8;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9af9e5a937b30f196caf71f9ddf64480a63f9268de0b8abe88605ac7a2495d60166357a08dcb0a67d76bffddef30ec7a41c227bca617b2f2d4198f85d17e81f353c52f3a24566761503f839d35e9c5d1a0f1423b840957f09c3ccf76f9ae63f48263aa7fdac430614c3ff0e4a1daa0180;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfb2f37446aac507b7891403a5e6bbc8973ffd14749c596cdc229f188aa4a32eb7a0a1a4dd8110a498a2314a89d60e4bee9b8fa4163f0265a351d7f7803e9d82b2aaf3f13826495eb61a8b942c56d526dd80124782cc889c29d1018315a5685b7e2e25221051fec76c489ee24b99afe69b;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'haf6aed3f823c8e433d2bd83b2a5be1cf500ae03b0812491a32f81b29c2ba990d6b15c2746bf5565cee031be1ecf0858a32b11167121a4e13e507c0b498d43d2084857b12eb918306d7b556a628f80246ff0ebe45824e0586b6420f7a72afb96488eaac0fd07cdad8c281d50036b89c300;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha34aaf807c06b316762a0bdc2ef0c58afd25ace92748a73310789cdbc99f52ea09c4d161d49fd35ab037b7e2b1a49a72f85eb9b3a9d803449125da7627337e51be9cbaaa9c3523524fb7a983f9e568762b77a1d251ca72b0a0c15c6809660ae21ba7c50f2593530b6df029636429d944a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc5c18e15ae84c436b0ec464d5da7b2532037b3cb4edffddc3d2e14ef41b468f7187382f29c59e83dcd65fbd3454abe557c61c497b9c4d756499d28cba950bf7738f312dca9e6dde84f6dd4296d6d90a5af62750b7024e10d6208f36c19558a2d49543655c5f1ef02567aa5c89147726b;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7f836f7f68662dd8d98401bd80d7224092ab4c0da1587f5446a657185aafbcfe1d32a2d50820f7b00fc064a98511542b17bd71fd8add2cf86590381f89468731d0f18ecdaa2eb948cc0fada6651d0a9ffb33f320b6840947d3704e3559b9300963d306187b8710d421c02b5beead34fc9;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hcf5b8a0c268441bde4998656e7f5977b7fc8c0718c7b38fe1101a687af1c5020c6f72dd20e934e3b22035131219dde0b561f0c21f5c7f33447ae2a1023821e9241d4f05d2a2741ceff03b4dbc039d6efc780f1495b62cffa51ee67db7d32953bd0b28240fdce8352826b480c1080b6c3;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h686722e81e5abb27d872bb568deadd7625f96f33f017dd144f01d331afbed4777c1bbbc0e7ba7b923ed3d539d1d743f4195860b10f62d50796b18d8c8783e3047471f488a70de046ab8a1c5b0fbb7a82ea2cd6d661fec421474702d234d6fd1c4ad69e80e805a9c7e5a2738d64e872541;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h73e9c5d2595332069767ffee8872b19dc3d4f56f178b68500507bf5f8f43cd1d129b44438d95ecf588458c05acd07b7e6fc6ed5ee866fa31cfad07177e260e03ad76853b7e648aa78916c2fa96bbc53959321f166bfa6aa6100e2fcccdaaa4f180c4c5b6d368322a5e04c6b23c5542f2d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h49573432918e3b01f28bfbd64a66ba586badf3eb61ae4aaa461ed4847de1a7ca328261b63a19b779730f97572d797a591c989090c5721973bcd27fee3ec7f7f4312aeab01cafd0feba65d357cd37d762d053f2bc5ad04977f9094d9143a81b9b499fade45c3fa72b011132ae886f2b3ab;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h12194a9784cd7cd89e1520f74903ca0bd72a6b74c59241394b91541abdfa32d8edeb1aa249773b7daba1e3737ff8d0c388d83de39cf0a4f534471a48fc94d633bce7a98af452795316116855af7709fc474aeddc19ed5d92170ea84762b35b799d67feee68cfaa2a51f0a243f78013ee9;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he71ed82af277040eb458002200a728ec4609413c2986f8243858d80f49d6fb543b0678d2e72d3813e96d106a4a5d7e52c486acce20976ca86fe8ce3af4f8fd50f22e88bd87e9c57445680cc3dd98fa872241a6f66651ea48974077cb19e0a2d6666ed2120dfe3b69c1e9179188662e9a4;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9d3cbaf7b87c5813e2556a198323a8d811eb818d15fe92c476d396e1904e2ba2a85465f0184eb311e7a4c4d7e09381021ca70cbf10a565ed6df429d1b3d0a5a099c64544fbb533991c50d610bb3739b796f985ab98ade1bfedbb74c19dcd2a25d860b67bde1555a428ea65f604e0114d5;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb988ef408a3773a71938b042a3685b361ef9cfa189b56c5c530e9930d8c49bc979dea49f0f4309bec653ae5a830d756be77d5c5018eab7793e0281182b1e082c1a2cc4b491f1f129f4df78221ac8716cd11248ddb018004cb703629780004506cf65cefd91a8a0ce14ab3b653a5eeeb7f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbf4624bea520eca08df8b672cb8163e6c9424ea46a011500aff2993bdb482bc8d98c1272a957f27488672816597c050057e5eb4181c270f804b4e93201b1865d61a1892bacbb5a2dd408cb0f5e35c89f1f4463e13237e16d763eb05b605ac7a54d0670adcb5de1d4346b8c52cc7ee1a4;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h693f8026fadf5fef2953e6d37f4967d034eaca834e7ba3a95630b69f965df0f6b552137c5f5862b827b4bf65091c7de9b61295b6a7809bb64e3bc7c41a733e9d28476b9d2ed1c21bca554aa0cc31a7b67851a3aa360307ad4c58494a945bcd989c46d3cec88b54d0eab8a9e742c5ddc65;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5714b4359847f93eb2c76ebda0158ca59ce1bd8bc8cd36f8f47bda6894097f055dfb11238861635eaa4b2f585db5bc8744c5228119c6fcea58f7e9aeb08bd106e20aef781df232547ffe0d21f115923b528ec149a8921cad68da242a7a51123d1b0e67e6d5aa677f15b7248323b6fa87d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h41f1f60f46845cf2cf0d6d06840001641319f31e2195dd699b7eccaf084e01a4a2ee46f6001b74d5f6e1f75e4b975daaef18c839695e077501f3e2d5738bb0a9d26d95110db7a914042ffd9f86919225e46f6dbcf7971b4a9aa6013e07b287131d7c1ab9fb0fb5f1dae6dd63e4de05215;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf847f5bc9d658cb2d0537bfadf421db0f68bbe44ece8be093b79058946c0ad19cfb9c136f19d5293825b0e2c1ad7ab213fb03abc1eca1732e231e0c9383ab6d1cdeb9f4e0d9362a519a65f3d4a939255b973c44ea662387501a8265c55af00e94da7d18e83fabc327c4818d02fd32d2b3;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'haf1b7e06c5a9b1599abf74b46e81657096b8923d06522a22030986c6c3244c23f02f25242fbc11be5d93eb0a077b08939b7e585b382a56eef183c7a0c5bf222f68750e5a5f9f3f1270ec4ea15b56e78edfedbdb7edc8a269e92457d85af81bad338c98d9d9e90c8ae957a8c15a924e7bb;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2aa2b607bebc60e2cc7050689fbcd1f71d9e5fdb8579f4d2c67f0ec957b65d2f6a503474ed353992e7a0041c2be557e6091ddf97b8fbf1e814925910f34a421b627736c0574f6da6ec62d32583d2a1d2f6c3cd5487ec7930a0703471ad6fe33b83ae150244cf3cda085a0db332e90cec9;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hecc11173d64627702ae1db7fa1f932edd78b27e2870e6198d38ba752b1544bd9dbcb0025b8176855c465a489b9d40a1e7be8eb56394c6b6adaaaccfead1eefa7ea951f18e2e17f6b70486c251d687f53613c19278ecada66f3d2dd3a4e5589133246bd94132574c8e1522ee59b74b964c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc1610aa7b361a4cb5de198f407e2aa3b62db58de8d9035e6113814440fb659752e4c64ceb234b21c46baf03575adaf0e711a0166c469816c2eaa29977e514c3f2b419830b60e537bedeae9d7ea2a819783bdea7b46aa02125fc1d29472e69b3fb6fffcf6aff15aeac6b86ed61b287c331;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1f8aae5e02d21f747fb9d7a206ed0a03ba7013f3629a49d285d63b79fbc950c0c994b075135cd711af2715436b83495038d4f2f786268ab9162ceda206c6315114e0579dbf4bd51e89f01ed315d4a6745bc1abcf1a307ca042fdfabe23a6587bdc6035556589862e2a1cee63c79707bbd;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb7c28c4cda59e3b1ef52eaf1c5106ccc701037a2ee14b7df79063c814a720e2c9bd737d5efa879f603ea5b856c09f405eb51a86b380daee002e5af89e2370eb3b4041f00de6a4c37ad19b9240bc3577ea3f68dbf7989764a160e5a6ae40c2f25fc37a5c9dff7e505208234d4311ecedbc;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hddc9342f20475a906ce4d434a10b9aa33f604a24a56472e66205f2b61385f6539cd0fecfc491def4aace23dbe7207492a02d001a5e92bddffda74aa0a49d47df14794a699f7adc98bdd0d9d3353a15f024da888df5ba11b8172089a22b9a85b3bddc0599dd5c23011db16c17733e353a8;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he21cf5485c1c7f73495661aec352663493ac35047863387062884d652c2afe4a75d213e0803328ff9ee680d9f3ef66c8007799469e225dfda143d0fe87c5fd51520f69517c77c5b7f727a03ec46969914e546a0c3dc53b3c28658766879525331ba9c8fa98de01a8068d66a22320547c4;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h314ce76b405d15b045f133749e7e1c425d3ae8c82b03dce54d720dbe959aab53aeadbb140d9c60004254b0fa9c23172cd397b26818e8ebacaca0e28b83140bcd25dd53e99dce2fbf31109ea25a73b5c22e52e243cdbb6050a7f077a4b85e368acc83e12c4d0a9ece7bc4b68f036761dc8;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbc85280c97f1295c641db029a84930c1722c8990d460a7291ae9856523236986f029d4c854d94586025f54507a37b57484d1a9aed9c866452bc30bb043d346985468d37d313e5a7d280540203a0ea9023be79c81e7331d5d851c1cb167c42e1b5cc6e7eb80dfdd1f065dcfe398001219e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he5fdb49f911c35693efbca64816894e9d95d0a4872e7bce2133c219993bf14d643226b5283a3321a14a32be4a8ba4aa492ce50386e91592944d26248bc5ea44c41eab099d9e846121a948cdf7ccd40d7b85e66aaab29fcdaefc519e8022223ea8df1e7c91e790ec41fb296cf220695f1d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1dd05c76389a1ecde06470f2e67e78c973f793af752344bc5a3d9d69ccade86d12aba09728d20eb54a7c46b44c3c665d5c9d0ffa5412ecc219f53c84ae2fad412ee3cd8dc1cf3104ac3b69d61e3cae3485edc10fce2249814aefca155130fb9f2c364699ff6fcc4067453cdd3e444fff4;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6da1727029a1070d042db07ce72163a9fcc2bc30536dfc5a8eeebe97b36065f1345b3b348e44d0ddc24ee70fc2efe5fa5bca98a35d9ea655f4158b0a26009998d557dba624931d66611f8e068cfcc89f31fae8ac1e73a8d8a36d10191382804e653559408567721904533807e3fe7e820;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h494647f9067c7100531f15b159782fa39bbe40b862145991c8dd1f59ff494e6c4a6b649cb6ad4a6c8b5cbb09b7cf1d3724817b28d8e0a5602d3bc3e5f2b9f060cd43ef0903c28b1f2dc01484090f534cda5af400e684320b9e9dcb785aed836b46da151d446eb833ceacf3aa4c951802d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4b4a4745af3631a4b0ad206bc8e1231b9f5186132308fd44d3f77c9be4bc9b54ada6efd06debfbd545b02f212335977570ee79f5fe4169cbd74dd9408fba3236940929091b1b681d446055e12548af23904212492f514b1c212febaf86a0757a67849257f8253056a3a80951346fadf4;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd15c08ed7783128fee2cb6052ac615c684d6ba66c741696b06c8e572ad05ab30f0b54d384639f337d806921acb9f5761e79727f5fc647bc280dfb5b8c204b6a94bfab9e5cff7d1e349e1a2d982f33395ea94e8f1015bf2bfdaa7af78033dcffad4f21da4c31b01d08554aab7132c16981;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hec3f097287ed06f2b6591bf374cad80baaf56d1fd683e334fcda827bf5255f6209ddbbb538e82ca22176304f3c1782db278b8267216f7bc26e5f649c868c6ee9a2bec4bcf618a6ee5c81639252bb9bb4d88f6aea340f9e615776d6813bf14fe9a5d55bc934b22ac0bb28a43aa1c5beee7;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5e9ab9c1b9b95491901c2d52984ca2fab94b84234f2e14dc5468d04a1b1a66e1a4a2bee1baba392102a3f1138aaef8efc4edd9640bb16a9c2329e5e81f07958bc660d925e4a16043980c16f127632deca217c6779819a9bb1c3fcd848e7852db6ecb7d2104263d42eaad457bfdf3b4077;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8e6e309d8f84550d236d1a6b3690d8b06888a56cf8bc99ee528415e67530ea94e670f25cdb6f3ae1ba2975b624c26ea07c1d2126c40c2fd8af964b00ddc1b438558353a76c7e238d2e44a0151397175121514377550bc26b6de9a8c9ebeff2c379c3eb75f0cb0ec76221763193e415f91;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1fcc8d2465ac45e131d3d8134c622dcfd4977ee2bc3c564c521bcca10ce3d27464f9a9415147a96752b9ac531bab28966e8b4dfe68a5ba010b986dbef7f2ae200204ca5525afe83bd44cb8ec8a100416a13dc2cb59b1dca0e9d91b58210e4633dbf4dabfa38bb963748be6e929bc89ae3;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2ab42341d2bd8bb6965d4a6cbaac95d9f0ea48a4d603772c9bc1001bcbabd4aacddd5bd9b10e0e95849bf80d820109bfebc84f6b0ced2270638aea16b972eb4b3174e4189bf5d1c999c9aae1ef9d3fc027a601a1823bfd34bdb4c21e22b5356fef9d4b03d17d8b5d4b1aafbf45d34ece;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha25eaf5b018372c81fda52041571e0024691a6f814d5ba23da4982ac2bda3c90825519dc92c9ff5ac9ac10f55d7700966309035e05b7db790c4b07cb54b75d09254650149ef7ee6d71726bc576bb3f68d4c2623971c3df45e996d58dae3667719b010596961bead7d436d5b9b4077a64c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc73ca328a93a89cef6a95dbe2ceb4b5a5bb60b69ad8829ef667980733dcb2a7f854f7ae6e4d296740db2ee2d4d55c03c71d2ee0247a5e28450cf08f23b504af912a133e0b61812de19481587efc20bd781527e1eb9066ec3e704aad166b4a2e28e4f3beb8fed0ea2f155fb182eb2c0b20;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4b967c40beaa73f36b0a9308d172dbf6ff194466319e8506182d0c13ebbb2c37f7a94311872bae7cd8719d407001aff206908c41c8cce23722d451e42abb96122dfffd76e7316e0a071bacc56de67b28bd3d9186e78f37b5cd7ce5fe0bb29eb51c0d787f6feb88e097d8674633eb41185;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hec66ea8eba616913e1538618e243a0a2c14fd556db66f3d7b9fce8f64ddab70f59bae1ed872d17b9b34791a853e89a4cb0aecfbef14eabfee44fd83f9aed87674ad94192ded206ebb5c653481a2d217591cc5b64809b0983ebae6a0259053fa449d14019c15c75e9fdc3b29111177eb09;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbd70b40cf38267237dd092552d8c8713dab065dd3b517e1043ff3320b00166253a338bb99603721c6fab08bef983a41215170d95418a739d7445e797dada8be8ee91fde1b3ecf1dacf20ca9b420eb3db27743fc455cd402dda8fd0ea72afb5db0e774d136a0a8b11eca1d79154736ca11;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1ea93377a2b93a221b6ce84cdabcbfbdc23a1e88994fababa3338ceb8ab19da3ba4416d4041db9dd170bfecba98ae79f00d89b7469e09c389130bd9c65afd7e8c6df9536e088bb024a7a6a06e038b38506fe18b5cf457697b5cb64201d4110247e2457cdcb0057711133ebd46b8939c34;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdb4ba2396483d287cbd3afa7c30494f50b7c933927017582999c19613e8bc98d37f9a2b1e575617c1691dff76c9b97fa33a5ea611120c6d776420b1eefe45953ba649cd8415dbfb1c096d9b202b292bd0557c9b516fcb8cac5f0de72f0de15127f545e94a3c9d8a4538e75ce6fd8ecd65;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2aad8a0f52f5a5ea30bbd48cf9a9b4bfe34b256dbc245c0ac45fe1ef30069c3dd196c7fc5baff40e099b0fa21fb71ea3566a7a61cce243d49d645729ac5126c0aa39ddc3feb12d07223242462a3cfa7adfc175627ad1be0d8a1998b16b69f55b165a4f3dbea52ed674229a6f85b88f7da;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdeb5316033af5e55481c5cbd230135a1cc62f7bf6e69b4ae28b5d4b7f571d3ee44577ca0a44891f221a8acd1de3ec658c2a2ad88b0ed951f23767038669e4c1569931a00f73f4826d8cbfccdef14f02ec06951bc519ddc7d133bd24cd3aa79817b6462456e9644d9fe6419bd288b45524;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h28fb44033154e50d6754604ef2b83d6626771068d8403b045a6e339b6b2f5951a317c858679d5e7ffba64b147841e313371885ed71a2b2024b2608ecba06024249562acebfcb3314361ba5c950a57e6f0f3a6557725509596abff2e159d35075743d58aea151a1e45e1171d2bf1207554;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1db8956e43b1e8fb1fa9f4dbda4582c05c5d4590da4ca3de4ba7726676d8ebd0badd9d655913c28a1b66db3c1cbb69b6424db3a212bd0a11dcc6e5ef595b55bf09c19de8d1f19bd9dc26b0b5fb054efd06f10111bb6a364051db21236e457ba29ca2b395c3b3f4d73f0924ceeb47eb011;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he8042deccb0c5179c9717201b352b9ae393ba6ae1fc9c8d67132d4b837d8d81e23e12ba3be79e96047a19b1e2abdbbed525bf7404fc0769a4617f958b664a83e18b3757681ee0f3e7432f58f7e794717d1b5942d39767f5995b66d95288b32f96bf906ba378fee9d1f087597507aa123;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hba08ed63dff81a2c53a8da37a88473140a918445aa4caf8969442bce2e0cc46bae51e3ae8d7e54f47611b8db7a043250cc921dc65c1d8f1f8876792b08741dbb743571550d361d95cd6302cf1a6ccb390ccc61dcbdadc1d1bc07da65701412c87b8ce62d9bb39972e1f9cfa7298f26dc;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h865a3feae2d55c7f8016241a78e6ae12802c6596ef1819a78e2cf71ff76a2dd622c712948d764466dde18a50acb51a3b8842ae0ace7d8c952c2fef80317186e1cd46d625c9a1d1c7a527ce218da5b069311d315007cdf9e3574eed56cc97785f82e48bd1cdc045bccf649cd719f9cba2c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hce8b21f37acb426952e3abeec36ca7dad1d0b3c642aa3fe07972e4ad70313da1de8c89b0e78806be628566238ccb3b021942226f2d8115ef52d5fb64fd0a4ef075abb288bb69690d90af5415d03c3e4a12fa46a054cccfef762cc4c029559680e413fa0780cc4d76a15016fe65b7c6d7;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h99f8f05a33d302eb99ae40888ddaa343550ece29911582ff1bffcf49832e573e02b3f9dae4408313c6761ba9f5fa9b785285b65328ac049837591fe468621ed7d4d2b4277148c6dbf3cf148ed29f82495959dc85924b5ac7e603a14b7622d04f971e64970fbd84d90126d62f1c6d0bb6e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h32b1d0537c05104683d6ce82c0bc1c0e9ed0991513962b1865029c727f0b4ca605116151cebc47cf689176f13925171e81ade299047e3c9ddb881dc7f21be9d4e54bcd685c9e483b48d7387036cfed52a30097c906755e8caa9d4c54e432ebb58777ca25e6bfc83f67591bbe3de989c28;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdd4e22cacfc5bd7afe9623573908f0e56780516a3f860788ff15e984937d8117c62fba61ebf0b0b4a97db14056d54528a3e5fb342bbe74c53fc19c9b3ef32bfb557e6426d7ad3706a44ed3616ea48ad46f44d6ed424adb94a96302e62b14c2df207174020340a526a323df29519346831;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h59237f6ff2513b8d154579150928f6898ce0b56b1275fff9a44ed764968737f4b4eba04cedb515c99ab9ecf8d48da5360ccfc25804c01fce202d3b60549c526a56066e432221583eb878390b6e5edda41b7d548b9e5aec20878389d110364526b3f8e257bef6ac3c8167e517abc2450d0;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2f21e0fcc948216d0c0d672da00e62aef3960492e5940747792c34782450e0945b9caffa681bf4caf636e575220429d9767bec68ee5c975be5450a7a081f44677b619d90334bf0411cb00ce8db86f4b748f241dfe4c24305291382cb4d995610f2a4715c7053c3a4cd72de63b84bf6e9e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf948d778d2f6ee515a1056c5a9ab050c9ea24ac7ab631a9d5ca44ee52853f14c54cb8c678bc3abbd6d2316f251ba2580d37d13d7b30183c74f4e04c259aa4a365f8c37716674fdb47371acd1dd1e2de3a05c8ae7dc8bd6c9b71af3da6571e1e2dbb029142725efc8d34ceb7ad58a00605;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf7d17afeed58ec3df39cdb1aec3ac0816edfee878efd1aee2b9fbfac1c6e501981377900ecfa53040fb5771b759a1cbcf48db848bee046ff0bf64b06243d4a5b66307cd3bfc23d15e30cb725b7b1dd3b438609ad8c9f5d5786b69664bf4e434b38100cc4c5b611b18697401e4f6990b53;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb9d58b62945070744e2bdbc23aea43c6723323d05dcc0511daf712c9e5274894e31605e4af2d8b75bf82dbd9bd4d5adcea565fd45ddc2bb30c2ad0f4b41905a7255077bfac7cc4b367289b862cfdbe3df52a7cfa24eb539c63c7ffdff31caa663cec9b867331eb87b497fb5ea897c6f9f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hcc812c22a35c941ba32c390771bbc414955aabc6119d472baa6e1194f35e96bcaef9022501e2d31885c7046f779df9ad10baf7f9fda9dd949319753fd1b4b7c0b1c1d7dd00bc6ddedddc1f953abfe8f240c7f4e4a08dc456982d7fe82a66905fd059ed14af98c073db447ed04b1e714e9;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8afe9c90a4a367c87f7856ff1fdb28b341df8e2d6d3f21fabecb45b812b1d1d3602184e67ae4435b3ce5031a8196f61c710d837df54653ab008fbee097c238ade0b6c20acd77b4480bbd0e64d926f6935231d1be5b5abb6166725edd071b047dc15d31ba45effc9067dabad0bb24bd084;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5070c84abbc467b550be4b845094da40fac9905ed8d9b14fff26348eb5722a952f19a2e7036123160bbbd28c945486fb7694da2a8e16e203cecfe64ee34b679614d5beccb6f3fb966da0217a3b2e2b4a8dfe26f871a49a67717241bb4b2338d7618d2ac02bd27a523a224d6f0c2c19fb5;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hca3eca4ecc1b78eb73ee76365a9b427f4cb85800f536e9d6d43e603c9709d83e1710ac995359a58fa8abceb11bf42495cb848617d790785c151f396589a122f9b6ad7cc449c6482f828c2f93639ef9316347b26408ddd332b03a3d088d1be11d9119b30db3f4758253883d8b5ec479eb7;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb82ae376998fcd3ee0a087f542fca1345363c4e4a88a32bc15d75e1120ad5e8200fabbfb5da5ba24a71acf3ba68553cc5d50e309a9f647866765748054a436442edbc51e81387353b4c4106bba0246c829c09410545574ce9c22fc129e395ae11bdcd445c1e82e1465c4627751ada55d6;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h31ae2753d917a9c10bf4040b4aeb9305c4c0e2e377f55bac83730ea0fad4b22f968d8119d7b97f006e0be0a0a3783980934397241647dc8505de14aa394a2f192d56c42b626b675c7c83bf3977a395841b27cb185cbfba9e34bcaed9b4c23e6ab9f4ca3209625438daca345bca43c07f5;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc1163a3996a67ea53942487ff352ae0127c24a9e65884e9bafae71c277d72f0bb8390b817d265da6203a73ee243c3957d861039c8fc31821cbe711645cf360a079e4c19981739f2918a1be6a8b9235e89224be027b3323723ccf735b7f8f98bd4c4a20b14335fde439b3fe18917a3e400;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6c35d6ec819bdf941ffc4bef947b234a2b1be387a0d57511f109fc1bdf5f59514b28a1d1015469b310d0886485b44ebbed97f3b59600ef91106089a7a3fed7ac65bf9886e00b4f55e77df2e0d7b8330154ec8e96f700a4835396d50362cbada310345fab1a5ed1355440870711e031cca;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf4a5c40f701031c6ba6d70deb5e6d546e84257b82b37ee34a6f03dde51019a38156d409ebaefa98881efdc968c2a46abe976b2c468623079e1396c8ec36945c6445bd6c986261420a46a06a0ae11f146545f296f5598f38bd6bc01d0501431b85b5dc63896f198e662b9fde51420dca99;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf135563805502e51587ba2b341ff88772a9463de25fbf1f1ddf8be0ccd645438d0a81d1e8c3c90804f1d33a63c6afb446658ab69d186b8867b5d2470ea1eb9dd4e5fe2473523655cda87e8db4cd05cff6a36449f2412e14941c3832cf5960dd5d3d72637c9645362071d91e3780c83cdc;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'heb3ed863c9821517931f4102c6e5635ad750d86c400df2fc0419e2ddd132050db6b5630f13c210c30b32f4fd11508d88d63416a875ffc651ffd270f06b2a8f0fe5178fa08a13d902e670d4640ae840ade08b780f0dcdf5970ed2a73b56539b244d1d8824a0dc611ea59cbda29d44da24c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb1429189aecedf4d7dde238df69d62d1d076e8a9103c70202214c79d786dd141db0e91f4a8c9ac967305b29b3b6ff9c82531f3d9e613b441654e3a4db1369b2b23ba5dcd38a7d68d1eae72313df5ee1549f8f849ccd1ec87772888ee38fa76b3356d41821a665800aca7b75e2a949e21e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hac1a824d3fa51ce41da4b28c47a9ad03e672d8f7ac8f9bf450d9afaeb69603836bea91d76c9465cfea7aeefbe7589449eac73463f9c507ba794dd228bfed18fc104c1835484a71a2037b243d0e031e9501a8c69c8ca96aa5d01c8ef28d5a4fe532eec39f8f955b409152681c3d1755077;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6d853f54857a03392cc4195a66ee1ead0099805a8278781a332fb3c455e671d5f9e1e4ca72545b1e54de53590b2898ea2d61db5efb63ca352fcf672eb8c39f696240d3f21d5021130429ff582322b097b835f0091f99840e1a1202e4ab55d4dffed7380a46ea6902b9ad75ab427d2ca35;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1f86af6740a571b5db3361fb8e963ad8ede70142fa24487a6c2bdf54eb0375e2d1006e1d44da72a32fdb2b66fb74fee555f2bb02a718104ed126763b9366b8617b70a671eb5744f6ff731600f20c4c9701305bb54137e1c02d1008e04afcdd9b6b9e60794f9d06bea7e0043d864a3ddc5;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h216281e5774c9aa6043c5288b4eda839f056111635b89aa7b74eb14f585aebe431c116a59bc091bc65eb85f82c3b805295b06868c286f657a83cf6881eaf951206ddf0f2c50c017a17272b156a4caa85d3f4e08683f01ae8532e8fba623b40bc4e5b7d2c99fd5ad856cd711796f973ad8;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha04958958b028aa7f990cc92ff76c549a7483e01a0126b35ac11a13f5fabb8517e39f11e355a4946ec7d3a5b3edecfde89752dec4a520da642dc724743c068dea8e154d1b1f2d4b04a7b7d9d545ae7a078aea3bcd8c561a9c5e9d627ebd9477a8573265aadc9d462606b279a05faae6f5;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf12618e9cdd5d6b0b0ea241a86e730b6df43bdeb983e6d4edd7632e225ff42b456ec2102921b6ccfc8b1ec21df645997c4f19c84bd9cd4ea38ddf78275bc7e18ed665da6df8138ab4bcf3eb6ee0a61d7dee3d9a6d0e01c8582962537b7d8ac7ad16c3202f7e30ba7b9df3764e126536f2;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h24e861c9ee96abebefdbe1d6ac540b54f228df30e6957bb0368d9f444bb762fa906408d38109ecef7d5009cf3bfee6a0311697086f8e74ce7f6ff6a8308c912741f8e70a0e35612b9320d0fad7ef55a5dfec9522c589ce8f981eac46584ea57bcf8cb9968efa1412723131efeca841f00;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h84c79af010be6c5c0ed109a86d6950960c97799ab9b4c1179e1592b7f347f3f638ae1116455080aa145c8cc8734e6c6edff28b4fe72bf78eabf3745037634179f07afeeb9860bb41c6739f7e3b1826215e95785da7feaa9ccd10d72a66e1ccf2435416d64e0269730adcb55742173b193;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha56a75c02f58c00648aabc3899e2dc613db1d9bf86ee51d3e01e118191659995ce4d9ca9ee48da20241654af633e50c5a9a659a42f494a884bbf707840ab00e52354675211ba4fe74dbba568804cf09660858039ae980fd2e98bbabbc9c0edb4c61342b817f1e5e5359d83d6d2f9d5f89;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbfc870c411ef076cc4cd61e845c6d3dadc890253c2a0976a8de1d7207b431948ce1051d8ff3fddfdfa9a1a91c01db6c2b174e57f1e6f0ef3937b992b2b3bbbf02e551712cd874b9c224ee3ced7adccfd542aee34ed11b31c44dea96e2b165c15a4986d091deb660e00a7f56679081524a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha321e346b31975722d944c8f49d449317b4f12e89ed3feac8c193e06a7296d56a159082fa240b6afb43efc5182b50c1e7c2007afd93ae4caa80e90c46fb703b1c5650c9cff3dd62f770e3b67c8647286f0fedbc8129adacdc3f9bdcdde4f77a047306cfb14eae1d8ac0fcee423b52f609;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7297544b05d983cd97ee971d28802731f476b8d185ba776eed529c903d44d989209341dea50cd489d6f4762b17751449aed56fac28948a95f48e9d368acbfab07025ba58ecf718bb5886a3f54d2266784f54e1df00444acc469876fbaa05bf06faa87d88850589562134081c99d9f6b2a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h343c3d9a2065ab910e98ff63ef145ac90e515aa63f63c7a1613e882e6537e5a09367480344901d4fcc38ffb8f975dafd4f4cd495952b3dc520e2f79dacd4d792a21dc34963045c663e597423995e18c3be541bf4222b4a9d64f07fd1074b01796f53133937f31b89503204af5773c7bd6;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he095f5b1f49b0833843f0c62682ce2d65651312233f259396836d679805fc356744264d9121acc633bbde336fc00edb471784fe4f9c0173ce6b32b08bef17c66c6aa1416a583236bc148b4438ceae9b69e5b11596b0e0f6100cb156d1e72fe661af5e95cacc7b0e97483482ad5104bece;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4df7f1d0701a88834a55ea899e750e218b51c3da56b516e1e222104c0a1d0b4295781ae4e4011aff2f412436851405eeba28ba07278679a22ae743b1cd03977f5a4bf4a60c28b7a1878b32220b6f80825508a2821b133d06201664864b2e7c7aceacaaa6c55086c5307e6027ae39ec19e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf6e9d83c8a548bff8e60ba8276d8ef0de8a8de111355bcb3f28db8dd8dfd652fe9245ea473c9119eafcf7ed2da70166d55a66af850e411a17e4701cc0dda633162186a15b8877e4391481ec45795375e6df07b89611c8cf6bbf2adaa96303dcacb27c3189d9abd54f22b51f68a164d466;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he26bb1ee84e280afe67fa996465e6d6787fafef2ffd758188799000f44f711e032a39246d6419dcbb4c7861a6f2869e4a22fd927469ed865c222c7c8dbd4258973c229f3e9c5539b0edd40874eff0f06456c6b87a99b39617069ba9e5ef2ec1cc4e67ea3348e0f39251b390b81728df59;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4fb73972931e64995770fc5b58bf34f2ecf7fdf53461c6c90278ebffb42e1b6152ee7c6c8c4c2b18a668357f8c39638a44245e3e60f5d6eb4993dd5b61d45e533395134970d84dc435401894edd83318707586b451ca11ad50916411df9de95ce1e19e26a5cff3ded5332d5c73fb2c429;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8aa7bab9178795711c9082e2875883fb651c34b0b3898e87388c8514ab2538a577662b1d4d57bc5b202a0d188f2bb12bcbd038f18bdd5e19d69fe6d7702c1c65baa68afb214159cec31a6845925d5c4888b2c5cbef1ab228464b9650785cd0c79f97d1fe1b29cdabb3bc247471d4f2172;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5c7602e8327cf9f6677f0127216fd38d6c3b09af77f4374c50796f330dfaf9d63050bdd182348982b8ac2ed37604f351de65057c2e8ec62e8d61e3e18fb691114f6b06313ef1a326985aed5784672e93cfa82a6717afec492be11e9f73bc8aedeefc9b3d439ec5f1b482c1366f9f4ce8;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc0babfeb317547a0bee71904b8a2096e13bd16b601922d3c464cddbc2f8ae0c8fc3c40c61f8835d9f72658b6356ea3d12f58f6dc86577db04daefe14eb25c27fa94e3f19a4987f9a0a37e49911f37274747220ca582702e2a53a2c22358c443c8d9529ed2d68143be7d9e484ceb768c76;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc4af2d591d3d22e18bebf369fa183bfded11b31a49bf56315c149116b492439403fef68e3d49e81467d280cbd1c85631ac463a98e712c706f40d7b6fdd63462fcbf1d35a4e33712e8863c42b1e0c69f3a5d0ad32657e3dc129f9fc5eac284d7d4dfb754078c3281f29efb28a48b912948;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdfd4828b2ac51501489cc4ce981c17e6f61b26fdbc3673fb0cbe54135dc9d938d3c99c4cffda3f513a5e26546a76dc8b7f56275d70afa8c14eb9ebbdd2ab0e2537451c1757aa69573934f12bbf1b88fef79b4a6e66194d7fb1b0b060a8522eb614b09c4e815e18d6e721d966fd934dc7;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7f93e58965b0cbe61a9fc6e4c758a1bde8f93f3346b052caa215140983cc947444c6d5248f6a535c4c46ef15635eb648cbc019dffc1de41a4cc8c1d478738fb1586884b81a8447c39c6402e94c9a0eefaf50b4594a69d1704f726427c26bb981795768549b4b821ff3c2caf1cb7d5e437;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h10124daf124001c3b684429fcdb0420425655576affddd83656ac25c65f8b9bbfe69bed9e028885f3415cf16f6103c61afb9394b8e0a7793327ee75c75499f962b7c525507e2d9f4edcbfb3f9e97b070af0214177bc42c44d58878294445a18a27d7fb920913c44be70a26e6b99bf7887;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb32e5fab370441697f71546ae73cfccdb7a5a2b3781353b40035dc97520c2f1d86abca77d4f4c7eff4ea32acc3410fcea28fb2340c61963e4a27e61e4a55cef4dbd2bc1d3f35e29e37c8a88bc3b151dab26b2595176e1447a98f929eb3253d3bc19bbb6e7d0628b8623a3954a85f8a0d6;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6383a32d0761319fdbceb4235b1b4ac962e4831d5a88a3ed4cb8463c720bbc4f9dd2c20a1dbf431eb3c761356f9ae210f6fd08a521adc0ae760ea139b3b7e6724bd3e4e679a4ea5e1c4a234d31239c770655c1fbd1e2b8dd5344e752251acc5bab222330972604ac53f3f08b448ce6e27;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha885d10244dbb45d839cdb1208ded8895f3d3084a6173e0f78c54170b1cde0b6bec6585a1f954e3419aa03c799d3901fd891ed425fa5b58b4dffa27fce546571b3ebba8ef0333dd94f0b687e15ff958caf342766b1251d311e087a6bda017cbe7e59508ca01f5e503ad886de22e0fbc31;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbb0863418a197bfc0f44c8dd16a232c60c8411173e7ac0e62101d7a5c2efc16855416b62a5b1301b87c1ed838b7bdca61af25c5e6274fea383660b7f3d2fcd4afdbda548c744bbdb025891c482171a9067fe434930712569649417dcbd323c9785e95b5064198cb42f6db3c06d1540f0;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h306448a8206f1dc2220a59e220687586a4f37b0d8bf09f8c0271e8567d6ade1b2367195a95d8bee6e5d8917eca32c41f2ca8226683eea08a61847e71c53ac79e208f7ae661f7432e447d809ca30e1e93051eb445a3b57a8890c52bf528203b9d96262d23b27e72409f1a3144938742ba6;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h554daa47a96cf5d12a1bcf0c9c5590cbf7a9d236459105bf0e1dd308b553bd8d2df99719a87fec25b17fee3adc02e87a78cdcb3c47d8b19e070804da403010ccbf0590f5dbfa02a4230b9cc079eeede9a8a678eef8cf2aeb7d919936dfc71cc4c55bc71bc10dcba3f0166111baa0d3201;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6b9c033efeb303a175d467bf57db3eaa5af3aee961a94fd502b921ee031540042be4dab29f12b08fba9676843a418401ee4ea1d3ab811284f63e838f23b4d6d9cc6137c7d6e987430c688634ce52a2847d7186c87c6ec512f128479185e888da3b575d29cac119417bf0ed61a1c01517;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h306992861cd6e9c1a207f95cf837cb9367fef46d1f3934222782d3c43a0e8aa0a795b2c37267cc01a8dd6f031cc525547795c2c8922b29a48fcc21d8110ba0231cb2153960a8dd86adccb663124a3f54468a006a66e58a9c01a3d699e911b5a15d7a3f3e27490f0efed21fb2098a38844;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd8d1e7ca0728dc85949b4e65a172a3fb0bf80555e0da571d40e99f98f42559274c95a910660dad9a025c373c887bc83d9a204a4f3ff19363383ce79d03f07d00b97d26f4a1e391b244da2cf0a47f790ec69f29813f2109259b141eafff917d8913c16896da0eb7e4bb94321ae440b6cd1;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5e98e86795ff5e03b31b5e44c33f0f229116f7858bd7ce2977944c43cbb06d398e673f51f592caa40711c98a8ef2dd7d96e542cd4603963cafb012f372ba9f215f5abd5dcd9725ce21f473884e974d03c49baf15e13c9bb5d9d3bb359947d96d0d11ead2919f8fa36744af7be864db1ce;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4237085370f06e759e6083aec4062ffc2bf6341ce129c84614d79db0f8ee784cf95d22028f3dd230b14b3cb9bf322a55886f2bdcf21452b0b4bd4a4c874e6291d09e583446682fa6742a5569b6353b82dd3fd2b0f029355715f3ee5c0a995c6da9f7d0224d5a29dbf40a32e61139f48c1;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha7ca90b0ac44a15074d24033afd6def9f2616051f500bac7bb66004a98a3107b1f7f5a5dd0ee858154aed9c2ae29e6370b20a7d5e21227a686322ca0b204fc1e41105d2526022679b9848f671f438a3b10b4c20d3827040e3b12b1d7f5d1bf1262b2a3fcaf343e5ecffbd67ad00fb3a9d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'haa2bf08c3af5c836cfeb800e5209824101032d1d2ee6eee6e79ae2dd9e7b739db1b3de81e525b2f871b62d959edf4d89fc4336b1260463b8a6c20722d9ca45886bbe11cafcee6ba07d4b9caa58039d07a1b17b26b2baedb6f26bfbd498f761bed986dda647d2af64d2301888dcd146b9d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'haef3dca6a1d76239b846c2e73c7821d504e7dcd573c7b8851d85b4c09c83f3b79ac766b875be534d1105c3dd2fd7f74197215881a51c27c8c471a190a73fbd6a91fd6170ac1ccd5f1e043097fe1f75fa9276890b09bce800916acd9362133f4a57d86685dc45fd8fa1a934a669fb46e22;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb87025408ca6c79c15d72ccef2bed3afc042b41a6cea3bb2aa0d96b0459bf3c5f549a9a7c3c4f9c6d745d63c2f19f9721bc6c6115ca6973f2eafbe8eb70a3506382db6478335c272d7da8a13f24605fce93846ff6f3167f568bee858c598a370654a34c6947b7b36c5a74f0a5705405b;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6548221de33aa88c19aa72e10d0163fd73c35bfcd4fa302b5a8a99c0e8948dd96a53e96ebb406c9e0472335fbbc17f197990d3a5fbfc887c3b7c27ab6fffe90ffe727beee647d2c5064a73e5047e1f9a51d8e1d2ea538a0ebbe6f63c7753e8426cd544a76f2c4342d7b0222948e8296e4;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2ee88d36a8432df95bccf01d8034b559428c11804eb9b5d976659d493a3a6544ca5be2cfbb6371fa3983777dc976997fda494585ac19e572b75335e4eb861c2dc9f869b2eac08a077a9fd1433f25d5f2f436bd1a603312408b23277db0b1e85dcfe26b5b766736b15e52385bb8cbe285d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb008ac816729172af529ac3638083dca8790d7fd779742c010573aa772de57dd95621752654896ff2fe61a60c192fec013cdc03f4a6a9676b007c23de5b97db20f0d729755ea0bdbb83ec616b71a375271c0f665598cb589d4629ef0d52db11ca0d160c5e2042e5f43556f37312c23700;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h11de3d1e53635cfc41a36ba6b7e6b6706e13c3ae1ce0392f31b42e68b8f9658a353da3d9efd73584cebeb6d83573fae9a552f84de3b65733879045facaa7a0ebc50d17b02037576739505ce4930b4d832fbad774b75d6acc037ecc0d232a1f2559b7f87e19602f55f3264936a2a29569c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6e18f071f58d74f0781429d50f2b37e5ddfbb6108439a21efa102aa5ab9c59897e33ed1edbdb0d4c14895a1aae6173d3819d493177a9aa9087b60f55b66dfc1f05a13d39e5160b463c52622c9eaa932384e8d060aa190a75ea30cb946ec8a844c7c549ce50f49bb6684488315a5e5485d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h35e4c42798116e9cb868f98dbe7873ad060b5a25b5c74a6b28a9d8e3407aed624ac4dc244b89962a4f1c5c28bd482db9333cd83b98fb23f080a49f052cda8b3fff65dabe2b71dac942bd7df2e3ea75ab4236cdda596ddebe6eb78471e7826a1b0fd888c6c1ed09496bdbc72b984f178e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h876293e1cb5ec51b3b84515b4813c7733152f05a9f271103cbea24376b7442a7d03c6d79568786225903f33bf8d680d3c49d7edf45bcd514d09dd96440235a8839ee6d91394c2f6f7fb404fe15aa2633fa121ca62d02f73b95a65f050e4ebf9e68c0a6b3ebee2864018085047dc09eb33;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6be6fceb5e58cb32ae287523e76de880104e11ef6134afaadde14fb1074b2f9be44e19b253454314b34d42dfc3fbbaca404e02783044591ac7f166e0cfaf4a4812a32db781e48969660bfff9762c38926609fe82cd81463b75a35375fa96ef4e61f7a9e18c4858c759eeb6f4bd77d7a14;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'haef758babb57f6ae84c774afa2668655eac06041b670662b8ef32292cd34e58ff482d2f0954aa7184f477ecac5efbac5211a784b32e56f1532fe82c6742fe995ae3f251a80287b33af8da6c28149c3c64fb4a77f19dcbd3c0cdffa5810d782ae6a2e51cb4c1e4940144b6f228597e0266;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hcf6e683ef8f601f48104a193903e12324705f5b6d66d1e022f10971454e71c161c465cdaf712779d2c3c47766f6b6120139662e5e7b00578cce9d1feb9d431de97ef7439d42daeab19f065ebd602339add2ea0e0e65af7c61e77e147f3631286d068d25b0b0ae1602e022be432b5de694;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9f4dc5c2cdf54bcf8593781bca5194986461d685371ed5960d7cbfa85014946a5924276d535169ecb75b23520bd5590b14b1dac0ad804361924fe08875393ea9936022c88c800b940228c3735000fb5028d1e11296318b0279f3efba8826a490aae872aadee3bab7b0d013f86c3f060af;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h98cf9a9ee61d80c8efb1009a8e92ed3f3080042fc000e932af2d9a72f95db8c8f5a11d04af18e700a93f4aedeb605e64bc555b108f2bff0cf85a68b286382d6074d0aef55f6e3539c72a1df2cfee03e12a9de9f46f9baae12f3ad239e34789adfbbdcb0b57bf918889ff12e3fab2b1206;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdc52692a9f3a863cdcbf33ed3dfcfe8327a0282c4dac8d8f7bdd4a6c206ccda9b67051f78d8d6d34e8bb73092be44006e2e1b6e95253dfc98d03494488fe01a3e924c67da8421a083d43f88086d6a08c082617cd7b18f447f3e071a9f63c097e418bb466cf7021d07009ca364d08eac11;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6694a813544b1a2d4ee43a78f5f11e89ade962e7d252ffc42a6d09f9bbf879da5207e2e8791cc0f49e73d46a85ede2f25f62b077b650198ffc39785880ffdf4c974c19c49217d3eb1774e0838f80319d9c2a360f51e6f9561b3d38b9c4a5ff25a64a87b7e63fbd486eeb4f8b557612069;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf9281cc21434422866aac970679fd4bfc578c09372c7f66b5c1e01f386749361ec2be0400f3e2e1e6676dff747d2c61e60c8e78ff1a2bb7f83b55afd3b75c0ed078411a60f7c5e07efcabb48598753ca9722dbdc9b98f95258db74b5d50d670f94d0f4030ee981915c3060fba7ce9d783;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6c5b6655c6c07894406f2a809ffe69089da7c6c343038a31fc235ca1161c006298c07ea496c805c3813d2af188d60ea32a41541e8e48a191a5a2a63318518a8d63a7ddc5d2231140e4132089e15d777c10cd9656e3f013efc44bb995cdc1882cd6e8f3e16b1fd40e62fb1ae490d8d2521;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc770e882611fcf661f07d0f3063d6396fd589fe66faf4458cb0baf59582d48b0957391dd898206b8547848b3aa834bdb1d8219266e3b8b18046d60a399799f8c575418528cb6e23a685d31371cd1bd8ada354acb5afe261a917d6b5ad678dc15c1a24087cea1c1048775c8b55fd63554b;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1e5e385d6bdfa3e370b548f599589f7d9edd9051941530fe06d0574d75572045b10be863bc5abc7916ac5639bd341289f9f3c06944a13a51382ba45b1a594d4ac3a1a5c8aa1ee102453798531ece8ede32ec438cd99c765516b031f7f6ef0ba118ad7e5554585bc3a36d564e9dc684424;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7dfbc1d2addf2da178239e5eea13a7220fe1adbe2dfe23619dd45487945b24da0df521317bf4e017c68eaa7656404d2818cfb824318aa5e70f7bfa01824f2514fbffb17cc4496e22494356dcf2f0e5fa84f66a71cc441efecca6e3993c1591c69da05d4dfd7f4e1ce7db08406261a3261;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4ae6d3b2fb0ee4808b5442ef93c49558d113d066932ab44e25222e44b60954bdc5d724b5d7dbdd0c57f414f8235cc0620fb1c61c885ca3906ca4a5faf4296cd4d40816aa05146087e052efc3e252555d10e3e59b832044c1cb84a4af7a5c4ee6a72c724c4ea5c4c2974a70e85d4a5d093;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5d11a5f846d3e43677c1a5b2915776d55f508dc81936bbe5ef4e678f262146e82334f08a15f39a8d6abd2172016247936e557e5a8531cff828c558976fe728445dd7f7bce28287af69b3bd91e6b2e6cff5b04a0fb6cf780aa76fd66145716c03b0bfe2c802068beebbc1d6be549a71db1;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'had3ec9bbf6bd0f7b137d6a41a5dfab88b1597c5dee9ee39967bf4124da068cb3a2c6389a874094f6de547ff6642359cea8503c975c7e53f88d9f68059f89c77b00a43ae5c76cad00e85e3e05ef94b55691f09cdea373546dbd3336d3bdfdb88c8baf91b1ed0c6ff9f5dc1748d722f4dd0;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf816644f083b411eee193c8075e1fe36fc16c35ef71cb1a6eeb74f55088c35a8a36d000cffe7608755493ccc1eda67c5c26adceccf556dad1929ee1f7e5b538f4b5497e69d19efe2a24e468819545ef1aa40a680e4f7d2c60fd7ade903dae1a5dfc24e6b5715566237b087fbded52c14e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h14759d0d212d56bf6a34630e319bfc0ef2690ef86e4ddf011aebbaa8ebd4bdeff1ddbf6703c0dc795c6261a4185efe4eca3ebddafb02963a3251a91f9271cbe04ebda11990e4a37a2bbcf349ee72e95baf40d65b1c0b7f84f1bbc93b682c0f35613c329fa8d46268d272677d810943734;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h98997697aa4e5343241770f747d4dae995bc8559913be849635a911b36a0a5ba2a6855c22666200838ea55a18b5ccd650981e7dffb039400a4958852bd21499e20c4d4f53bc37b8a40e67443592e79917246479d24fb0f50333b69c2512bb2ad5b1b417b55163d70d067394559804833f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6c9099d53cbf51e672c59f7c6061d5f4effbb3c653597f16916cd752b618905c512d41822632f4ff80cdb8f2ff7c88dd69626c87b66c983cd14ddea8c149e0483e67fcc4d65cb124103817ddac7800c128285481228803af07830e570e69348073aa5f6058ca65fd49082398776d58118;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h418ca98400d3085aea493f84f79db2ccddf7365c17ded34e8cc698588b0334532bfe96caa864f60565f9e023f3a79c257c0195b8d87b0d336e51c1b24055b09edb8e312b4e19348c42ee97f85598eccdc67ae378db711b54c61b6ef65c1ff87ecd8e6b3d03e6ab4cb0f79ac6dd1167d21;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc9e0176deb4bc4493b0a5b57f9cbc0408d8148b136fb0779944a80a02241e70c95afa3ea6bff477ede33eb4880505e2fa9c10bb6a175d65a56f336e2c6d7b987972f604ef05d87463f3b30ab0fa872f3c6678034d2572d934ca5f0e84361d252dc2c3bed5687da302f18ebe798f864a97;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfeffbbdd8bccc759c16841e103d33123340c81028b9ae62c30d669abd74cf17bd3e5151d1c3935a1d8ce754f16f1ce79462eae1a228164376883e9a9f29410bc404ae4fdfa20caa1be71814605fe62525803fe83e4f27600bc524c4255c2b1bcc2aecf2cdcb29961536a4139576bd3cee;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdb9661655269f4bd96c9c259d314942dcbe7ea835aa82e90866b7745d5c1840b6635b0f75da428d5f131adecd9ea46d2457a2a5df799752234135f1d4022d94d3a407e63048f21cfbdf750d32cf2ee625c2e2582e6368e8de7ef29894eaf1ebad1ec56bb1e54cce0c34dfb0ede42ae9ec;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd9ab6bd115213691ac3f6fa9a00e1697ce8488ccaa5f58a78eadc2e70ff0bf6503aec7400acb9baba46d31f68f7fa947844c33560af903e57947d92f687bce897a8526b6d877512b1a1e006030c01cc9a222f30241a6b54247517d9fc7b75281778ad6d1c0c4cd503127ad298d50c3d01;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hec4648fff80a5ccc2a1615bbe9a24c8e3f5ff772594f9c420e6a09151ad119b1e436c6a97d15db193af4aacdafea6b15402c763034c0b72a2b45a86df72880189da495a8dee5f962e1209daedc07f090e43094f166ee3875d4e5110ad06d66868b69d8e55d212657629ca71834afc550a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd16fb1d6c7abcd4227e7e032aa071c5b3e4e1f29ad6249074847a6a658bb8b205e9c31bf361e6369a5d5762b252af473436f26a80b3f6e54e37a9e7d7a81884c64d1b4be354cfa59d8c57795a0c05990994301c4797fa625fd3515ecc47f647585567017c904b29602edd89f14daa1ba8;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he3a9946994b0c41987c45b1c4e372802dec789e89fa37cb8844d49075ad84d89248e9076f8c35d4de18c85bb0ca0ba396b391288ab5d8a86e62ba8220bf201896461aeb797b0aa289a54eeaa46c1b4bf78ab5f345e2c15a3b69502c291f37ab940b320d7410730fab4e3f5f8cc7686016;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h911c04387636bca39ddf2d4db6e86b94fd520fd85d49f84508da7209ae137d5659ee88700fd3306f78504cef8a865c35b4c6b194d0d701a27d4046093a022ae8993d86db1c7e190cefdf43b11d11259fc70781b212750f67620c7200b0b9f729c3810b0b32e495ace571729c00af6af1c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h254697ae68ea5649bc2d2c86f98fababcf01ceda71e28d25ccc923bba4808111a7ad13b4117e5a92ac5b792e5fad21402d72605fd3c54be47be0ce37ca77cab73224fe1460abd97682d106c63cb74769e901d6011ea6cdcb59a84f4d828afecc0f5329e7e7737803a5eae844124c49517;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h72adac10af0ad1f51cef59e62ded4fc7b5041f06ea7971ce7457e48689dfebbd836719b88b67a9a4799af453bb601f1ce87c3a5209dff87258b7aa6c820cecfc7bd62086c6e0817e96c6d0a2da8b5b01a584b7b946fab52701014ab74cc876497d23b051f82aefe0e2c29bf9a4b49573;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb989492ae757b28fa7b1b95850c25c0e58d0efc4068e433445b493707e1295b95b90547e1d310d1c75e5addbf7e379b8318f05bb4e30044ab5f7461ea55565383c798bbd6d995d21f6a3b905aa90fcf9a9a3eac16a6522719b97d9b15323a51baa8b5a3ddd30b01d1e3e0a7661ae148e5;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3a69b11d1ea65b99635051384636b076c6e25a0f2c16446dcef0b0577dbf5c46b5ba38c892450b79ba909d712649ceedb4af1a452452cac9072105776a019dde9727509ceaf87bf7df991371ed3085947db79f4f5ab69f41205ebc032fc7a81264563008e95577069231ae6b65aca64c9;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h940760401248e023bc0368a214ba13b13f48a4a795e4c207ba171dfae161c4332c2d3b374d1a797997dc964cb729201b877c647af0a92db142cdcaf2d5466d5f17c16b9a81b984709916e954a28799909429e7acd8f7acb869ede244e32420fa0f2a3ef47108838b98b6b5a4e4e8abd99;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9c1b172aa7ceeb3d55cb15c521b844580554399bfcc1fabf7916eee3821877ae531be96abb012013c069906c6eb791a281eab0a464d8846f73fdce471e7a57b81946feefa40d8865bc100cf9ece37bbba7eb1412458802e5a9667be9f8573ffb434592e1e53866ed7b9e1a8c10c40fe60;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hea5091287c2013d21eed713604c6b4c194c9356d1e78fe1f9217b761d4fbbdb50044d636c2dcc41b0241ffc47248bbf50d4dc716c18d50a1c723d6919f40df0336624dd276d1cad05d69087198e9cf0827ad3f5e8ab6f558bbeb892679773917084a1532dcc6b9a22890e1f0d9b08621c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h69f59152ce4e1a50e3b4de9870479f87c3aced85ff80452751c1c0e8e2074ccde280e24de890368a2279a7fa95ae8287cfd744e8ffe631d4e15ee387369e97cf87e685442fcd92bc012a5c7a6a1f24a88b9a124b6bde281c4b32bd031a5bbe14feed2654faf14894f6be6faf8207ddc43;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h95e04be1d8c199ef698195af10441895f4eb706c51934877214756d9c71215de98b9aff182807d760c59cd300fe0aa9b791c169ab6ec0a2ac102a74245fbe32d93d01ac3a49eb9a64db2497a44b782d3d3ca11e08b8efc613946439348c6257067d0d0dbfc9562a89ac1de3f560736c24;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h366a41ee3f17b0fa02c41a40b846e00ace2765d523c52294524b135a6b3281bf267af235837b4f707fa3e33d8271cfbef38ee5c4b512302db65297537b3c3fc3ba768103ed9718158159f616974c01945a14b988883295b5eee2611bb154ec89f529182e7179d8158fb3272b55ba370b3;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8ea67e66a9fcce69d6cbe87cb231fd73a98a8dfa6a9437a7765b512081f61e378327dcfcb01c4672b5a6a93732aa586b88a9fb41f33b7d1bae93656a370c075e9e6e44d3887a3329cd9ae3da717966241b55adb378532cbe0b9bdc0097d7ef184c938c59b208aa5dd20df820994d73f10;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h50d1c732f6a4f3b5738c0b09befca8af590dd5da1db21265509d574b8beb9843e7f0b2d33cdbb38e6b3a0473e0831b9734b6afb80e9efc6e21561a143c693db5352854dcae56b15acafe59c58d3a494e6efcb3ce0129ae1c76c14e8cbf142941e832831465a0f9952e56eab991aa6ae7a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h36dc7fa7fd5cc8e673aa218c76869ee82f382222b56b7b44b177da2647bc3b7ed92275a52306bdf06541e8bae197f11d59810ee3a1e4f7a07ff18adcf7e7d2f6287df170b77ee1ac06524dc4543f62d22994027cb9e9dabc61e27efbc7e87ef9a908f60501743ff868199259225ccb419;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6747746455201bdc2d32b47bcb8ac781aad4658b9342208acc4ca413707f034d5f22af26efd1d159e554d439188b338baeafa9f47ebaf057524cc906dc860ed74fea1406b98e805e3213b98a69b5b45794f3ac6a015fa611c164af2c9af0efcdff8e19e94244a676efec0169bf9704bb7;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4ecb0f95393c34eb2a2b70627a6a1a8e50de3675cdbfdf2a8d6beff89aad81b60b22a9c851cff95c40625f41957a1e2cc87af5eb9fdd46166e4b27fded909af151c876e92fb0554fbc3140f73eb27662360304929b4af5e8f90ab22b7b59b2a30bbe60ad2a0d27f67ea0890f0e51a86db;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbbc6b616b61ec9dfcce55a8ffd622c343b835d6f670041bd4688fbf3f707e36d5c742389d16b5e9732bca362536c1080d5a168109aa65561cddacb4688574550752d5a424208edf1d959c3606a7e76fe40daef1e0999cdd83ebcd141e872d1b0cbf9400413ed67509dace6bdf06b0af0d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2fe637a6383a5e9cbbd3b7e53288df3d73d45c97fe066b6c880a521345108b83b5980e2674b3bcb22766b737894a8934c312770d0d24a4a72842c41714d2e9409b1ca202129dc4363e72f5e5731ec61c8e0db350f283f665bd2fcfa5ba54760a24f621ba6beff8484883469d5fc0dc1db;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb68e4dfab180e1fa34373590bbec179d279e2961f9c86829aee8e856e4a30e6f3d5d5ff21d1ecee882058e80df07b60b5618909028604d4f7789995ac5bb55ee63a6389198411470672e48f84ec8e699532cc53b76755a177207c76f49112bd57fb81f7f2fae41be03fe26745b17a2278;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hcbbbe16d78122d82ff1238e68bb618eeee58a3abebee99d9a952446ffc166488543b815336f030d8c25f060a034e3bdd76050fc186e740a4c68573bae2e0f3a8f36bfe85272a9c83cfb5cdc62f9dc9adc1f282a358a388a2aaa1f41f42a1dbd30ed9b99c2c5b4770f98b0f8a99ef86cd4;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h256c7f8e77b8f15236c4538d5534698ccd383b071462f1c866ce4321ef8a973f7432d65bd81e76d3ea943de5640d4ecfda2f5f3ae4c2413119148d4c70bfb58e735cc0437c85c33c4715abd2536062d46769aa7a4e9d9f3fe593198bd8cc30c392ab4026914f28708a3b0be5756ac2c3e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h17110f2f49515b88d34b6e7244cd3bf40474e36202227cf78226a832005dfff4185a91127c188ca8c5ac3ce121c16f5cc70c4b080df899fb8bfcb9e4b35f30f2d2848c2518f4030ff8eb7c8aa649c37671c9cf74d6a0350e9c8fb5d48bb323339bf1b04b3b5747d8fd255667ebbfc61eb;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h351e0429515a41eef12dc7fd76650bc111e95898e5205b4a540054d6a6ad7b8df1521e1340170aaeed3d494b976d736d038794862f80a1cb12673dad900f858d4ef0620504d42f66c0dd04a5e2527870d5ef72d68e51348dbe93740674c4fa8713c32fb85115964cf895955ad1a8ec825;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6ff11806e3c1d9c5bb1b84bad126b215bbce59babaec095c60b25832b1feeb1290bac2ceb4ce8490c5b10da36ab778c7c83922f8ee17db7db4911331631c86142f00327ac86f83397d4101253f269f952c8c6434a8a39ccafbd2d856ddac68f5fe8dd22250048576a1a25007504fa65bd;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc598aa660853c3679ac365651198af17d9422e6650052e04e56a948820bb09fb5f6c6ad591f7cf341ce854094ca2a0ff6df42a47d23243b956f4f0f1867f073c9307ceaf20c63cdced2c0722ada59b6520d51128d578574a053e670696ff1c15e4670a28cd447798cf474ad6598a11731;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8a3ea6d3d58b3ae48e5fdde24f7f131c4bbdd49e9fcc38a6a05e28caef1bd79811d0ad7af174639eaef167463ce084edb769fea0b09e8a3e1691a0d4e305daac2f784cf87a26126644373f9e5665b40d5f50f5a128b8d9aaf95923005fc370af53a91889999c7614ec43b4c0e9ab03e3b;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha4b66e84d7b5908625df6e585b9a5c90e750e10348d94acdecd127f0af64463173e2a698795cbb243b35cdc487d995fd51b48e4fd977ae52d5894261cb5e13f7ff3b6e31a07dff3e7fc32d96dc535d09254c1d0ed74145f239e0c5ffa81ea81f5abfa27b23861098fe0c0bfc43a1a01cd;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h966b81bd8ed1f16858b481803c74ee2dcff2217d29004e24d08b048e1d84b1b7fcf03d757fb95a7db1aaac52a5a93defb7212fbbf6ec6195c7e4490b4c9fb72093a9b174d219503b66636902bf0fb4e1b3bd451c96bb7cc36e8f817727d15a5c85dadd70a42caae9381946e45966267c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7087e061c92c5189322b0b415d2bd12ff8260a3e13d21ff4a1be6ce46e055b12159aad860638bdd48355eccd5fc80df524c7138e456365e19c68e621f76a93d778d5b5cc1c700f3ac4c40000e9d795e76bc3b4076b3f772ee217591e16628c5132bcfce6c38f4e2aa55444cc2b21f8477;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5a936e328cf9b4ee9a87a493cea7e1480080786b3be0971cd92a32be4133d2c76c8bbaa56cf664d65359bba31d1f71fc8db815dd99851ffba333aefa5715919beef7e6b17c5ce9fc4e5c384eb1b16d0cb14b0e3bec62f2d3e08db872469c3166eb6fd0726bcd903c0a6318eea3f7fd18f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3837f0e1cb69b41af0261c3712c83399b5164dd33cacd53748227312a0f9354a3e59070a517e41d8a1bdd64c09310cb79ed153467124731f2b08987c1b4866aebc9b2ee71a5e4a8778270f786cbb2fc1c31e65cc5b3eb9e358ffcbe060d792776221ec9c3340f922754b859518b98d0e3;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd131a87e42462ab730c6373aa46ae438f74e3d1e9968b96e0ba7f41d2e2c73674f0f8a119726645a4212bafbf9e2e4bfac09f7ae5b3a76633546ae2115849b85692c148b61bfc8d8838160eadd2fdc8870254567f981101d720cba926e07065934f8d01fece0dd449188f1206454d9b10;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h26a1f91f4fc9c1ea3a7f4cf11917e8b0dc330f8b36f7aeabb0573137628549bd3b460c463062acaddde135ca8c3f10a305eaf7e3a7ed24d06b4db1c555fe830496b1c4449bce9537e3e5e1a2c6cac198ca5471449ab7bce470b3cc1ec2652d642b78d75f7d60b1a74793977037c1395fc;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h92d120c5d2ef2c455a24d619c71524729927e42526f2640fa2e6f17bc8a5a4796068593494efcd3121d2cc6362aa403808a78cae03b7f328fb909f382a400383d429a2b684d1bff12b7af7e59781ede2a80437e9cbcc799db2beeaa72e0dff49a35f43ce745d8b9b7d72d6392e782fb6d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf443ba5f3133bdf1c16aff7f9269daf5c344be5442a28dc377f41e5adfddac8a1ccc8054a26e0be2a35f3dbbfc2d75133095cde39b79490c58d4ec82f30092a77e2cb49ca0734f0526a9cd2dca907ace51e15908b476d6d2a7ec0eea7ad7c3313ec301838cd484a221fdd8fb9c8e348ee;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha8cbe0718f6ed9409e382d7296f58bc13519bfced7b20eb4b3c36fe6e49b0a7cacb2956431eec675df24679e4f73baec486140a9f7f4a5e621967c3c591e7a49e50c1fbb1870a3c4fc87462727dbf39081f37a24d9feee8a2a704b1482f4c49a6ff48d54c7606a2871aca9f1ad8943b0;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h14055b5b19e9fb0cf0194fc9b663ef54521061f92f5145fb8db3407baf8b7e6981ade4d2460526419098697b8a73783357045c21e4f14823b71b1d6ec3102ade8a4e2ecc4c8f0541e899bc1ad2fe7ee3aa85159784759a31fce3b271655631379e75785a4dc8d30fab4afd66d340f3743;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb3af7ea9752f19af79733099305bb7cfdd4396499240238451a5a04737d540d76f13f7542c37691c3a3a20925bb3863251f7fb2c69965a83e02dde88c0b521e2e6a4936de177b9dd7a7bcdfd3d8aeebbc64c2732847c04f01b8344a45d87e6e0136d9e7c622312e101048a98edf1c9643;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb29586818c7c38d50c55d01687a269ec81f5a0c74811fd74eaf9b63e8f89ef79cc3141d3a08594f4f84a561d92295070665a10bd5c6b264fafe81b8144ae0281674c9c8759223ce60f6eee83a62c71938ae9101ab8ff97c2fa81b7df090c746e763be3ecb1b3a145efe32026402bdc896;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2bef94c515b9e9623f1d6a4ae2b89e98ad9196dcf0b44ec96e17262824c205d9af11f9a27980ac52642927e6013ad6907c7c51436aa0a676f1ae020075c8319270562e1b551e5680a02d42040f283bca3004d8157428873abefc44d7a9c76deef02e69c9d4cc4ce00faf0adee8b8d9fa7;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3df6f994180091365466173e045a28c931855aa664c19bcf1487b40a83db4305a49a6abefcad1dabf0fe41e7abb26ecf034f706218c6731304cd23111a3a44c1e9708ec8498427818cb23b598f58af618b54d53a81ad20356a5fef482f6bd9ce2d4aa27c747c7551de988ad91eddc54a5;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h231bd6c224d19ee6bdbb0d5ce9c2f47d05f7bcd17f3b99c2af5e54562171f59681cebfa06973714ca45e2bb2c104f39b711eabd133db34a0c5b2ebfaa2c88fc0f4932eb0ce42e67f03d833a3d50d8b628b8c8aecb507720814fe035374e29f4273cfaaf57ddfeca654547f55775abf741;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hce5408b58ea0d9a33e03ededd8710540ed641ef14ac02d5dc94c1b706273fe8df4cc6ed47042559875faa44b59d0f45efc8a4f163bda4e9f10e10c2c267b691c6b8315bb3323f7ed89d635120def1c6acb24d13dc3fafc9f8a4df0240dff7d143a96c088faafe22f1030d6a905bfddbbb;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3f18c91f1cb6e3855b1070c594227efd06d18dd04a628570a41d081a27f49ccdbcd07fe38d945f4d2cbcaf4b310b885de6a672fec8414b309c828caa92194c5d5eb96bbac331e58a9ed406ef8928eee4e9496501935549e6ec222b03d7d7674b3505e56970bf6b0ccff99058f7d6b3d0d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hab698f16706133c60719960e152945438741fc29e195b8a784bdf36efa6de5280f8e75458d7108778dbe8d20e1ef5f2d6a949ecfb0aab6f72eebbe8181d63d0e5684dd37442367f3cd6537b50671f6687c99f3d926884ae10ae9e6eb7821ddd46087192746f48b349dbd42cd356ba46e4;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha58e2aa0ca574918496b323981650feb3973363e3a38cd4b16504bf63810b20957dc7fae7fe8f0a7c813ffcc6d00b0839dc12218eeebba694c33733e75b1fe95df7d2dadaf932b18f6031fc1f358a71af991e3a840299a886551ca7486b88482c64a339eb0b2fc3c72ef47faa84411425;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8e15fc8082d56b108f56a92a98dc4e6e2ea64b99566b7ae539bda99417c0b8f10857232c03f9f3845f6f69e5d67d85031381cc2dd6011e5499c825d8f08d68d49c7d0fc5454b69cbc727eba871ff4f6abb0f6ec4fbde7e1e12d6f29dd193fcfc07a39f5c95d64112186381c909b31c658;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'haac80b11f81e0aa300529433ac8e151d39fabd240accd85edb1139accc6ea6c9a49f6a14294b2d613a067ac9198ad7679da6b269d2abb023ed300977e8209febf6805c1d6cbd5edae9cd976bc01233f2b4f712a9729ad5fbde3c71d0d0f1cc4302d14f61f70a4d03c109b46423e6c1e0d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5b3dbe6fe684136f85cf162b93bfc600493607d091b3d04ac1d0726d9d93cee3ba5c4065b4b9b424451d20fc877d37657c4b03204526b14850472e671f3d1e31c85c7ba547d6626a5335f6a60396d6088d5468329ca09853811fd87760308c2e016e9a0246aa81c3d359070bada940e36;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h677f7cc76c0e049bbf02db8ecb785261096898ed4dc89b130065dac1c93a078db6ed172363972cd59e275cae37f43150d1b5df4564c2c84f38175d03047c858a78917c72556d1218d74465ca9bb1564e305f8719d038144558b4498384a875e2d9548beb2482f6073c17160fec08faef8;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb313e3b78962525411b27d389e773ea69d7cd4f11b937e4c6cb7cf1ff25775600e1909a2c85f94f89b588ddf03aaddaeb2bb8c08b92cdabc448b538abb6f2cfc19bd7517e4c66349291341b39109e99d29674560f0e7d69a0b042060c4d35859192d5241caa080d4dbc9ca5f7db230343;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h56efdb20a012342524340b79b4a63dee01d5bda1662c3de60bc2becb3b2219cd7dedf18de28b07036dd92b6ea65a0f5f999faced577b694c23e80f0543444882a94fe8fe3f7ec4a6625ccb20f3313440d3ad67ee6c16462d515a221eef8d91422a3092e52fff1100e7c086dde939a8e56;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h11e5c19fcbed0d347f691d33b5be4c8028792b26115dd6c6549814948dc175dd5f18fe87333761dc69c3a54b1802af30e2aee40fa7c027697c22ce71204e2d4c1af73666fbdd6b4a3fb21340efbba10ffe4b14ce22c9cb6efa108351c44ffe9ed134604f1e2654f09b3b8bc9f4ade02b9;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5afa3dcfeab2125bb0fe6129165925fc5f2b5f5685501d4af10aae9a19340584d48bad7f039921af83607913fc1852d5d7b49085efa8e367440b440fe820099bc12ff59a3de9c9220b2a4b0ad7a3b63a51d0eee1678e692f474aac3bdb2f1dd2e7c5961a133760fe57c14cbf3a7332da4;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb0e3e192b1fbc97d09f6212386cab8a63089d2fbe15d7c82d3cdfc41769d6c66cfb1340ff11f7b3315b8e5cc978527cb2fb407e4699a573fb84d685f19fe997a7e14335a3bf5c6f5f3409fffd55aa87aade07345bd0fb8350518b8bfd303dc7d646a793a0f49702c95ea2782ba7583672;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7dc6836c12c36f5dba3603088609b5f7dc873b21024848f9de950c81cf167e4baf68c16bbbbbad4125ea6b8d8d65eca19ca6ab1b7c8207f79c82f3a3ac871eec5d4bd60bff7b652f403bb4dce496c6a9acfbe633f3cf830cdfd2d91acd7383420761e8c52d030df36eb6c4964c9e740fc;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hab63cb265fa17ac61dcd4c9b289ccfe877a0c3eabeed7e6c2e33e066b0a29d6613257872c8889f2c28bc489cf00a35cee5e5076067dd369d2fc23aec60f815bc52de97979b6d9ad963ba00c72a01f5f434c3ff0b5faea5aca84c9232b96ff46e8aad6133e03088fc771c978c169e36ba;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9e7da5f59c63bbe0c52361e0c6128eb897154430e7b17e7dfd1adf1b437b5e9504eba22ab6f49b66c0cbe955967fc019dccc3e1d28dcc9a2875e64be0ea7084cc79a9704937954c9d732b861d3da00d3efbfb98318b597d7e053f5610dc255101a112204dfc5a63282403c1eb344042a3;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2745df1da0a152960c354b9c4c9ffebb46cf47b0622213cce65f2f11456f3f53bd156a9c28412cfa13c8fa5ca3ea86a09f833b5da37fce630311d7ecb831f019010085e5e03ed4b5a7c89639958efd1fe58bcbaa06930c09a8364e22775315e4db43bfb5aad3fc8cd01b12576cd0dc72a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7d55e3ac635a8bc35c5059a442ad9647544215410dbc7d7f6c247d7b9c6ed81d653060e7412bbcd4c88947fee28cf33ffe2b61140e6e50fbb7d227688ab7654f1d5503b1054c7039624d07b2c5d9f6611becab8e79458d199769e29b3703e31f0159143bc0093af502a823bac35a0aff2;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h61762a2ec4e17a11c4edbbfcbd27c65e8c373b64d39a89ed7fbab3644b48a6de138adcceb682af23931301f91767054076eb846506b61270bf28fea5513cf2db2cb9def1d170dd08d5f4bc85c514e116225e2c302a0ccf0bc55cc5fc3ba45b9f4752e62ca5069cefb27d0fb7588697712;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7edb8c975da4fd599270e1683c5ec15adc2ccec953e0225befc4b49be71bad8e9cb51fb11ecec702757f47ce6c7979baa50ab85c54327575b4996c4ac1c25865de880bc60a360ebf02d53e3dc674fa0d9cbb248ccceffdb096dfdff6d28cc296ad87b6fad55cd059602daebdeb491f93c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4cd614e23fe3fcb33d2a7730fb33dd2002aa547e6e2a7d6e5d89ce035ad84edc297461578319a65cba25048a1c61666ac65f5cb5add81d55ab5ac0cecb4e11c869512beac0693e376b869fadc0851c7bb9b545ecb343b4425eeb8d12be3c837758e6fdcaeed0908cb82c03ebf05ef6901;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h35c75aa3fe04f591d81bfdaf3f691546f376d4f5b9a1ff853c433a3f433b38404bc823999271c9fef193796c8201a7023bd768540e35c33f9d086901629108156f097beb65708d972c4543d5fddff2eec2593aea9471de1e741e893412adeba7cd0a21dc882140fb58604e41e4846bb85;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hef155594fc07de42d6c3a1be82096cf3e80d865795d9c3a5855c3d4f9694e6fabce7241fcaea58037cc8fa739426a8a99403e65a375775e977919a9684d0266d8995320aad3edcb7d899bb8af0312f09767b0cf7cbfd2902aa088debb5c25c959b0ac5648a7dc76613adde9691b196800;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8bee9a544814e1becd79e7c8b3ef44d9a2e98ec8a562776a3527ce67460d59bde57142cc095bba95e37626ee37b39db6098664aec5514b0aea26578d38d8d926bf517ee2d1472043375e6155a6489fb099f41e1e7498782a36f7f59b1a542c3b54a45624836eb92477ade38ad5607b0c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h768e64d541127cdecb52d28c5c1b20bdad0ca20bee28b70abb48b0e8188e586ef202eb5aecaec61480360011eaef2f6052e7ab9fc8c72c6d04daa28d8e75e8c5301cf8ef43ec2c8bb7c43a9d8987a0e3ce21c74f2bfa7de989f4f2b9b7e19cb8a7ef4792a4e2aa5b68989c82c7ea90361;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7f3245dfbedfcb60301c5a366d43fddab51228a2e91c92efa2fba2a8fc616cb8943be4f39c82a6a56b942d099040766225970a51acc0baa2c35169e171b97e7b454ca08f0a94be05d6e97fbbb3ea33a60082988a3581d3182e2f22edf90be742c950ba09310b957c8d848b4373a34ccde;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7e89c5fa23024d6b2a9c60e75f10f9f550de621d233371b72fb19c19f6796cfa513a5aa106bde47af41540b968346b3d7bc9a8b3bcf35490c262ed96f6b917573f76515cb68895a613b3021c48750bb1f2ef5ae765c03957661d23ef82223b466805f2601e3789f73e38ba4fa192aa42c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hba9a4a4998d93924ae88035afd827b64804e361bf05d2ad7e9b6e2416122864c1562c5fefd63f12ff66b6f60a098baf9489feab46d2c76270bf5ef7b959e85b800aee1aafa34f33be7346eade7d37490943b58bd2d52e4b1c01760d94cc1408da369565920e9f9c0fd4b162bf4333113;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb8c1e1e2c55af291e68f5615c939edb1b52f4c11ba13634e54c8027a2661fb3c922cbdf74c171f7f70c04b130daef54926fff886172aac7f6f87b4be6c686e633415c72728e8fe2cd7769f9b1e81d6ba58d00c79bec575336a2aa365ac8287d90238564c3761f607b74999a5798ef485d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdb4e1481d8bc0a56581015873cd5e94bba3e85bc8d0d5e242d21bbe804c4caa0271b8a85d06f2153c4dd0e78f4201269e316ae82dfec27bed91dbe60d804191f363e3ac5692056935fac1873f7f01c7d79b79a09db1d4ad8fb5e8fce80f517a67dd5fafd6e0280d3e676b9633729d5a8d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf2ba40734f3961d3fbb6cc325836b530390eb699e6d12b058a902ddb6355472ed88a73d659b8ae2a318b6d87dd2aa092a4a194c400b2d0d85ea2719e3f54eacfe83433761427be07866ef07e54b2f7654c80e8c551e4c2c069c0933fd0edca80918cb9c6e71927a5de5799862549c3c27;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h63cbd15c858985ddffe30a96563faca7003dc93688aea0890295b5ce1e9e2aea73697f93ee224c825a3499f1c99934653954eb6ff830b0bfbaaa985d8fd9d1620a25c1bf8e98441a0e6a07ddee5b93131aacafa72bfa7ab3a26617b6721dd79e3f2bd0c15acc55d6a52dd673ff693c25e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfbb789449ed019f5755c628e71dc8aecdb1342f8be4fe29f51f15bc8727f3c2b1bc2d34c82bb721fc928822600ecd747f59cae0af1779fdc289a56e9e82acecb5c92b2162e7731e54001c5a1c967bd72d6703fd5e54ff649761737604108b4345bf98cf24ab475b762224aab8269c9b7a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6c0a1f9c4f1f61667c851eb054e31dc0176c78850f4dfc5dd5e0de8c8a9af0e01b89f49e3e4344ae96996ecbcf6eea1ec44f5a28d9a16082f85d014c8fbb8c921dd817d4ea8ae231ee1ce0e07b85c0dba17cf636562bacdc42fa12d1810d79763ea107f0d5845f69a7183e9e091afa4e9;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf00b7777507a197380d9ab227820f234a63042ab86a1631f3568a6352d958eeed36b078307a6647ed10e1b5ce81dee5b90f368c41fa34e5ffd5ebd9aa764309e52202a1c788e979bd201299d271d99d671953bc210828f1826e79278126c20b193dd1d7108062a5ada6e423f90dab7a27;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h73ce0c6ba112dc42095789f438d8f75e9193fbc0b45f8520b555210aec22287bc55464be6847bb2bb303157374724fccf4bbb432ee3ea4781abef8fba6718e4ea2f8169419e4acb721ae5bb0a3030821b9df8e7da56f4b62e8191a590b9e6dad8921d95b71ea8de1a5123126a311049c0;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1d33b3d25c4d967c194b63fb4afd48abc87d50568704e684a2052d6ff75dcc73562464276c7dd938c414d1511899af40cf10d0d0c36a37e4a4d891006bfbd1120db34ec9d6af7ba6ea31efe3a42c654ba7052013f46791ff921704105f03f8770be0b72e04a2ebde3484e837034c176e3;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3114c06c480bc1560ea401f3f30c498432a3ad5a76349df106349a70ab650ab6ba3827f4bf86d36284305c31cff32bb62122e36116ccf2b47acbcac8d83a6f402d92e2ff9c91803d4bf8104d7fd48e6f9ed7bc2bd3e35cc26d7c0584b3f10a85fe57b8b7d62a403d2a06730e5c93aee34;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hae0b9727e623ebd688da344d04a1eca0289e087c7b4acffc5bfd0e6ab028666583072f3cfece4354a1501439afac8e6d448b5a1fdc6bc21b795fc183d2b0c3811a1e35dbe5dfaab2c2e73dac9c9c718b5fbf5209bd736ad40c4f2f832232cc5d5be6e61a81443c1d422892813a5cd7e34;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h90d3ec3264096f257970fe562cb997427062e318791404f99a8a8a7809b72c62c562a80678d39fa31748ed5973c322fe2b170c509ab1914b6cbf627deded5d3d48f80d3337bcf5eb4eb115d27686cec3b272c3e274a6813ca022f27dad11ba911b0b6619d04a14dcd5e1d38a2ae4b352a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h985add8f8bf51317864b7ef9bc8714ca8dbc7a10aeb85a77e1636ccae6928e5857cff2d5bc25fe85833c01972e46c394b1f28e9c3d6f3d15b50956dcdf36f3f0fcdff20fd437ad3e3cb40e9e3d6437373c3f0a33e46de9807876873f893a80132fddfc60c5005f9a95b8dc3dc27d9f2b9;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4877a17c6068c3d9a019b88135da18eba803f22281ad152fa497413c6f652fbb6528c87ac821fe3ed5b3b3155427001a87828db0d6a3a08dae0f8358d9c47295515f9bd90fbba3b4e6228052d9b28cbcb7197908cfc0791c9d03b88474104b9418e9cdbd36467502e9f7ea62c4bb1220e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h793ffc69948ec4cb65351e0083b66da017026ac3c45b33fc967a9e55c91963d4e8a64c7e8bb7b2dc886459a1ba43986c05dac98ca76e5afc2e24cc5964db57e0045e20217cdc7a8dd2ce438233bccedfcde1abe347e1cda1e5457320c360b9504c4061477d92cbdd05837d22fd4f4d1f3;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h99c8736c4b7460c6054574e1a4363055ac50a3d2140cc785682b17a9b2a12e4f766ee56bd9b33094a18d608c3eeaf252fe8897a30e3c7b8ff54ca9f1f95061a71b4ca31abcee67e7c2502173a27613a7fc7af2c822c08dc0157f402c79d2a96d0ff59db119944229bfedcfea73eba378;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd0639a78afcfa936af809df86a7d6a1fee5ba32e77f2657b5b2b46a61e4a8193532ab03e8340c4732b438d105c41077cab86e0810a178994747adf0aa27aa9a8f51cca5070b4632ee5e65cb9b53d4778655d6d366852ce1fb5c6152b09a07f65dbbb9ef24298a37c19239d3fe6f0fd702;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbd503f8b589053045b1f5f30820ae34533367dae62e0c1d4b80571eaad54c6df22f86311f8a2c2f963dcace941fb9222f90e34a0b1fcfc8d27033c26b25916f05ba9593645a3080bf8e0e79107dc4cb84c5f822af2f3ec0f3b819a140b1bfcf451cac6e35c16a16d41294e2ffbc0db39c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hce11bae97828ed3c0f17c6b786ec723ae9d8ac449f2f6165ad6d40e584d219652892b07ade785bf6d668ee0d398228051ae60ab2fc3a17995f0b6e344c1e357b070cbf80a23dfaaf4b71d3688e3099705a8f6a721b8e9ae9d9d0276d6d953fd41268722eaa4dcc0da503427b5d39858f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h825c5b3167aa8d0f404681ebd59b76ed262b1a55fc6af067e91891f2b7fecaa0b62746b7657a43a76f02e6a15c2793de5dcf0be4ab050426f23516ed1914a83119fb1f025a66a7c32759bb4c2f84d5a84920be6034a326574c01c18468abab9ce31d246f412576c3898eeb02c23776b68;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5674d1636728e389c112c749965ec206e9c520b7d6044129bf94b92c035a9808297a39f911e496f33edfd807fb9ea5e6a030974def942e874075039da0cf25100e5b1b8e87c2f872f4c1fdc009065ed57313f4b855f6024ab2508ec7b0d2476c2da96799d2e8039348eea81ff291f490a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha2281758e48976340e5094bdcb605719f57de3b2a6f23de737db90b0fb55502ec3bb704fb1588d7883a80b55c0d71412a3d2a0063b373e49e123094397bc0292e0f849efd03bc8037d2fdb1d55a5b69cf7247db9c190014c93ad82633c558fc7717adacd3e13661faf236179ab86b1a8;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2a6180eb9fd0fe16df4841018c516e773958be854d8fee110194b3cb5fa8e4768a1548559ffc4c23e584080fc20149dab6bc0a6f74d04c660c9fa7bbfc7641c101a80fe40dcb09f79d8e904d3a01ace932c4e0b17bce1e0e967b4a224ea548582c7232f2b1c417dad53f36ad2f5159069;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h92cd06d4895c058cc6966dee94ab025b9cb15c631ceda8011a4962d1b676bef28fcb513abac43e725bc387d9ce464f468cb90e4b8f20ac35a58954280ae1f8e005f67392b010164e600cc7759e7192df70f11e01b75856486dfcf8efca7e958406d7f211afe836ed51d29b9c557c0e217;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hca5f101ad7a15bc581f72fd62d551c70213d1bcaccb881dd627184d4f28b84ebdd8f0571c2eaa26f3a3d224825a91176143cfd6700596cd2eea9e57054ef4fcbdd75024423e78cf558c294ed2f5123f96363c41692335e696866f76793175802f59772f5ea7099ae1c48b4712aa9e5bfa;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h249b122332aa8f73581f9f471dee8a5d050853f3228036b1db9263317aa42a7d31a97cb685a2d894701da5fc87e432dd61695da5b5ebbf4f91fe8581d909ba4df39b63721bb09e07071fedbfc6bda0721bbc3fb52348b3874e0f71196925b70a57548c3b34f453efc57a416fafe7fb9dc;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h94eede375ab5ab4550209ce7aae2fadf384444673959f121fe5d4cf02af962050d5a114921f5d27221f309fd8fe04d1228165b303df6fd930516b8a256a697363b84003cbb8f3b66399c00d16c172fafc3d54354e813df460f10121929f231b020a3a7bad0b438e35d6fe2efc56a0a344;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'haba3c975569ea94db06c09a203be8afde7b56ad4e55ed9bd38908bd52bba6409b663919f2803113e4f9f7323073bb9e6b5a721d6997b60d51117c1513ea271ad0b61965cd389f1a5d55463e62b41eee2c98cd49815bebc46685260e3c607006efebcc1f49d7ad20de14f3a17bfb314e36;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2c5d03f73b1bafc988103ef96beeead257b28905f811f5d6107afbbbd3ef442a303f058422f9c28d324002d312896942397620f235915f8e1512db55c1491533d61424b6d85ccb1b3ef9e68ee40c5e94ec81e46490198124e0f7e2a4f8d2ca639ec63e554c76c0670f56c29dc51cc68b5;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4b62715b42cdeef556ca5cbe5791a7ee74f0e91f708fccf498380d477fcbd1e2841a39bb13a2a6cc14874fa5c5d329efbfe1aa31b63607ec138d5b8ab62f1d180536633825138760bb3e9a2df15ab59bb10704067833062c1398f477f691ab94c97241787ecab91c1f29ccb1f9ab9ee84;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6d700b98da1f0eb9f749741a0dc2b75d587f4f44004afbe0979df731cddcbfd1ade3f9d93923b90eba1b37fbe65a76e826fec97ed70a28ce83148f6870bf057cc12cc63260723d577b0cf5c4b2a94f74f7901ce7670ebd069d4bfb35eb8ee9a4ab139879e5b3e9bef09807145a0a08187;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6da2e6b3b5602ba3ada93c1fd8a84d6f1be4a12634271e422ca2a5d35ce09c1f9b8a5ed0c98c8f48b7703f9ffd7b8c81d24c132797dbb62b76ace767f642f7e4b5132d6ea0edee7ab6918e31bd40532a86f64447d249028239bee9cf166234e167d574d1d736e3796d3060b0212f5d666;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7928f2dab05d82f78b6da8e8401755bff97477a31ac25481f81f7464ed42d2aece68b851686ef2556e9428016a1a6f6618aacb3ace1644061231fb06515f721df077e62385f30182def8bd5ee41d1545706c74fdf46234e6fe08ea5d05afdb0033375d9a67bdf8ad6f621eb79a75e28fd;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9228c93749af4d1f2969ac41938ddf238530b5453f73d5e21ec5828a1500036b74b3a8ba33563a8c1981da8ce8120ab89a9a9fc43ccaee8ad893f32296f5cca057a521638ea8fd031994e15c0c0be3886b361fea0b57dcb2abd5b1e2b3b87e831635d4c406b755d1e6a8228817a542664;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h44975da667e639d5eb2ef1840c3d0aa2c759d0d03532dc043ed436e9affe73934d66d1badf55577121a52e426b93ca48902208f51fd7baae3d6054fdf202e82e8539ae54cc5f66a1f67e8d4a063292d0af41829dc537dd9619bf864e2b489fc3b9ce37edacc0cf8c9b0a7d43186693b8;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfbecb29dd8345391b3c61df91ab983a7146ae776dbb3bd125a7327afc31b5c28e499a99f1c6b5d5e639f34bb00a9dba5895ff601c47fdc536ac7269008c642eba4ad2d035e915a09a78cc1e4d1fd2790908b0b28bf63e22af8996603eb440b74e0475bfb1165f50c98a8d38a67f61bec;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hcf52e1bea3f91e24e67ae0b8c6d8e2585cd12f8294c081dddfd1d6b8351dc8b6fb4437376d4e86d87670cd8989de25b3a1e37176c580b2d3ce8b175aad68cab96f1c8041820ee5f51a91165b82ead4f0661bb8ae2634339be1ad84fda51f45d31988883bb89296e3fbf24494216f6cba8;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h95a395be8178b61a1b3f087c0e1710bbaea6e7bec6f6b2d8eff38dba70244cfd427b0ba7bc7d8610f9a335d914401b7d1fbd60bc506ff48b76b39ddcc9943ea02a6cf9b507c28d8c2e6f988bcc13e94c7355c500a0c0f1f64794404bd510970211fb234f8349b30ad8fccc2f61f78e56e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h35829229f4eae0e6d7da6699671a25cf9c4de36d7ef1d66f9b50628e8b1168e63d0e3ca1b7abd5f7610a7991932beecc01565c47464997f3820122455725fab8d25a8379e7120206540f279467a8a8b3525ac6af1dab36687da4eabe2093b4dae5c31b2f3a24c9c4f50cfe72bd14fb829;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he79a435e79a785f1da028bbb49e26f81db46a49f731cacec8064cc9c21aac0ef52dc0e35fdb45225c108b473ccf80918fb58d37f2d92eb91b760a1ade2e7aa8c113cab64fc80b97dae494a7b163b31ee4b9e1d415f50dd811e82e8afb93e06617951d949eca38f813333b44b505349955;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4ba554c16c76bb284a5632c00a8d6a4c803b40d0f227a4bc2eac5707ae4ba97bca2d9f930edbb1d3d23396579df984936e502a4c1a08580676e39082f0666da46992708e5f0aa38d50c6941cb2f84098301006d8cccd346602fe4cb0d8081f96823e70c84b33b2d7d51757aa52543b3dc;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h861737e575821f1ad25609d1c967da5ffb23b8f78e586d97ba77ec3c7e0a60f9d8a3ba09f180979e93b66a00e72f765437f528de20279c0550eb77af2b8d8bb81f08513258de3af4ce8afcfbbd0ebe1b870fd8534da3a99f5ffcfc2ed89c48cb7bbc5006b3b79c46fc37e6bf0fe352222;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdf39c0dc7d53e7dc1c4219e85094679d7d1427a04140febba2ef3b7b4b5ce12c506f10fd1f3062fff4d222b1c7855ca763e8ea7b9429e75772f802d56ea4f20cc7995023c19b270cc2122058d2b370dec06271e29ba6aa636266c96a11ff1ccb5bfc5d14b5c8b516aad43cbb85e2c4751;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h61aa51168e9ec58da4e4dc1ec68a348ccaaba67b88c2de088ef1abf8f77c0013afade1e0776751feea3995914e152a630d418c6d2a600fbdd5d7ea5fcec1201338495f05612eec30fbb7ed098549e4745f638744f804f18e6c5487763468271adb1a9a2af81dac35d63d3e5d7464bdc8d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf572f00a14786a074fc0daaf6ee54c106f87bc4f2d1ffe582a8c1843d3cf7ef6d24bd4c3a05239d0b64488dee402747a9801cbcbad66a25fdef649c7df476c147e9029d3006f351989928bf832a090b84c700672e767743abf9eeab8a09d2a0a02c678c9d1140ebde6aaf1f713642b5e0;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdcd0fa1d75bc53651ee9e24da49ca4ea2371bf05ea1ebe97cd3175dc7adb408dadd735603b060d05642d2ac247f46fe85c861146e1b8bd9abca1f1f45140e4d4746525d5e4b1d9ce2b40c0332969e63225a803eb053d6e0db22c665876d469dfcb392bb6d7530b47dd8174c78271b852f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6ec52e7c621df047baea0e93a2eaf6c27421a4f77423bdeeb2f43c83bc086431b55b9aa072de384459df6161ab9a7938ba0921326fa1bb800dc5a3317d45f843dc3825285b75c86d3ab3634147cb70df98adc2bc7da8248bba0403121cf7ea221de368c7b90ae821169725277d108507a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5b6a9675eee3c3b1e5993d18dde674ab444ec78c9642757b210e6003a4401b0e32a0ba5c364c445a7a979423eeb073774619c54ce89c1007d657b36a13b1ba99867f1b2fc86a0af0dbcf36ee4245754539209088b15b653a00ad82c85fe2630d4fa55cd1896456de08d4337428aff3453;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h25bbb0cfd9324086f8f9e19c332a20c355a82c339eeaa85f6c25bc4dafb7b3405d2eb7125d9fa8657a0b1d0c17d12af0581e45c4f5684aa1f45fefda890e1a411e18f2b37db942a2e93480823767a8a5d429a96238a6d11c6a9aba1483bfd364ee629d706ae251843807f8da2546e91a8;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd4681192589cba8f78466ab51fea22791907f86f6e62ec94893ed7ce1ff589c50798554d340ed1544a346aa3e99147e433fd71ecaa5ef81f489d23a72a1e1c8c3b46106b9dfc25a5bbdf635d0de7f6e447f5fae50d89d1476f87daaddff342e9a3b1d518ebe909d45a859c99e4f99da56;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf25dc37fe24a68523d5fdf84bce94988ffde1c5326b13a7dce3e0fb569ff7fbfc696674e5d7ef0d40e9d17ab2581799fdf4d984814a78426f259a9322cc516d767c9258476c46b48152397ace732154450d5c4fd804adc16d4c204ea513feb573b6ca7217b5f8e42759b8d2af358a032c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha44820d54a168c65d2d4d0ba04ec6e57cfd6e42a36becd8faab78f4bce6eaa12f41d4e1d5930eb7b3a7f22025450712441b16ec1edd1c1490623cb7c6cc9b971890200449445d6ec46ad58957787d7f6819b45e52383713d6c46ee8e16d494d09205534a9fa1b6985c51d328e1fc55c3c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2bdb627ac9848348decd4bc5228ee9a83b48b0dcfc339336cb38f47a3b7fd2d38385553f2de678beda3cc29d1e92a021fb8787af034466181823617139dfa1432d3b820fa9c252d6ea914cf9257f4427857c380e46311742c4fa75298c71a450cb7bf3022f6d1cd5d2b364c422247bcfc;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1f6cf29c7cb19e943323daa4edc7c9e27f07c0c9af8cb9b36ba74a66220b0706ce3d5de3187c3a981f561c558b49be931733b2e83ce0d5c060d2ebf159e3f36a5df15d551c9d1ad20c96e97add88557150dd69743ae607135aebbe59606c82b1eca965902242bfa26ec960d42ebae3ffb;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h583e094cfa1978c9ae86c44b68b6cea8ca472f6f427f193692b7b792a3d913bfcf53139d13a02adaa9da2f8a293feac37757ca448f954f8dbbeca74094ad58a5743d64b487d5f0f3c5fd6ff87d62f8ea028416cc7bcf29cfe6489d02c9753f4dacb64ef3a6b24a12697280282f0791795;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1d0b4f0a225982d2fb85b85d4bf28ef5c83d49b9ab322cd79eee358138108ec211f9cf9e89ff8d4a76eb86938fa907c9b1e4b9aa2dc9dc0255ff57d07898c070eb92e8a7d3e031eb1b48469e68b426e5bd700457b5892a3ebc663010166295a9ba4058cc4e88ada696b8210929516cc;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he2f142cdacd14a9017f1356f31f30c7fa9c8b102a33c7d186f11e15fe14a9a742a52a1c76fb1a2754d84656d2610c052f91d69fc40d5bb2ceba8694399588f71bd25edbcb745d23331f736130f8212703e9dd3f48928aa3ce8f50b7ab5806b9bbda1bea0852835dafd53d7ea6f2f83ce7;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb3d1d3570174feeedaffccccd1fc0b767e1825d32bbe77b830718f21c7b28ce001d51cdc7b161b3f25078c3eb8c7f9536c5cbacb1045dcc9db04476a7ee4deba564169d769e35acb4bd1b250bc2d099916a460c970d3dfe8266ecad48012409d86c62f221bb63ddac8e1987620519dde;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h699dd82f5ef7e1492c593bee946de819702ffe3dde63d196a322ba646cec86ce7f015a62a3ccfad4941b314461d590db249e39d5efaed0cae78c795da10107e483e3c461800515ce93ec9ffb3b2807ae9b665431b28c8a2cc441d634e7810601f5a3e606362f1c4bb0afa850a6fa2e837;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1fc1525fc760a1e3b11a6cdb6cbf105700e515f9928b270c095e1d7de1c9bbba3df17725d8d5370f727a4dbce661bd889b839b99cf67332f26a3c1014bc4f0fa3658bfa3b76ab700362be2251ce2f7a15393128c886bbaf564ba0dba645f04cd80e56e1a3d5bca4450cb2d421b78407f1;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h50db5a78adbc9fd4ce9279da8312aa5792dae4a447fd5c0c7a1edfe75e8de0321ae56114234d3921e534316433e56671c7f852c4d21e8b59e6ba11c20395a1bc96b4def4642643d67dfe2b6ca417e268af76461cb467c77c5e75fa858e139fa08d7f491cb0241cbf8c608efe9cf7f9d32;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7273e1d0d6c389dc31295f444cf449ee86bea8ef24e7a5628c8e611f099bd86da567212190a1f6ff33ca1a628b48d7918ff30f436344a91abaa9eb3a9facba4c951e950d42095026366f20938e386a4ef595c989150f0602c5a2d4d311c5a68a5da348082be25db0a614e6073f5456f05;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8064dc4a48ba7d5d03a28457c70f43dea798ab82a45bd11ed1c8324ab3a5c80eb05ee84aa4cd1f78fd3b0476b8e9f59d1ec777106220fc8495ae2c7471613e2d5c18cd9fa86d9c9a47598f2a3e82a407a6185286e87ac5f1e8b8cc467764de7ca6d86640c03c94223222a404763d5bb70;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h19d565ab07503878f87758e6d601ab05f78df6a2e9e4182a2d3d96d8c220c4f282f3135f112a38709b0515c178506e69a4df98d7cda8d904d5b12f61c74f50969835362515b64c8bb7d1eaf469bbabbc04e9172543f459b39865905357b5434fbae0477a7406e66337b3ea5bcbf6a5270;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3cf92c2bfcd2aedbeb04481a8397693208783c0de819a67a5a2ce066416edc21f6a6daa62d4a0a10df33b6359baeb6e547bc5fcc83a407ce68f70b615a0626bfdf44249b2babc05b288bdd3c0fcf5284ce3e6b7132d4ac823eb7e86e94e0ebd5cc88e866c25de4ec18dfbbcaeac15a53d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1317437bffdff9e96b651fb9caf1079451e914bfb04dea3c54d2f2a07cfb42a3830bd0bfa5f5457bd47edddf3e1be32ec722267ef69041277d1358be734aac31c4f34a81a5995d3d4fae9671e24321b441705d9a7c708e8f84ce57e0f8814703ea8cbe77577b1d524fb21e8bf321a1704;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h95861ee298d877d1ac069460eac01152912a8ef969546c48ff1ac17cb9d37de4d16c0eaf593d5dba42eb4c3944a26115e6e577103dffe1913573cce046a0e7a9c92bc7ab8d31c1a6fe02c8db2e656dcc6802c30a5cc9c19524434312373b275fb4d836d3d5a21f2461cb1d19ab7f31811;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h94d564058867d8991bfcd5e02dafcb80836fef062b623653fbda74048eb2183a2f0e045bbbef0cfb8809151d2ced1123401fe812211c5e8b84826778f1d900da889ac42b45d3f3890ebe7dc18fbd7974a0e81b21e29131e5445a00c459f54264dd69a8280d8fb6ea9afec9dbcc5468561;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h143be83a50c020d5eae7b574a5eee9cb637ef4249b75cd3ded2fde82baa5341adf6b68a5b68ee79610a30a1c9d5bd2931a3af478c99355ebdbe13733685791f766709d7f2b09a32b17554004658a20ea84b0d3c78c4038c0cb13e0ad4febbcc1e9d8a6705a16009399fe7bab259baa6cf;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5d14ad08d44666314d01cfe49efa611434573482a716775b144ef7eb30fa193c3f243068ab40ccf6ed8b74d7c29cd48d009df14f1a607d8908343b0f2589706e63abb47f7f11321010eac334f4f73b5ca66b7df8182e5e2efc3abb59c3589aef688e895dae668d5fee22c4a0c0a1b36ee;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2cd2e5740380bcf6adbd3182a1fdbdfc4547d9fa7c1cb6ee667aefdb681fc0e443af738088a1e1fc717da8fc053259aa822f36690bb7a13290072540508ff327ed7faae43e81227a6f5dbd91015b5f960e1ba92a85351750644946f98b4121df4839c44333a6dd95200192acdd558f70b;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h84d2bcad50a89553338fa05fac49a86ca030faeaedcf7b66ebf869e5eec7fb89a2f27caa61017e54fcbe5889429978319b240b483ab20d057fb81c6aab0604b87087bdccd35ed1434c60bd1975b22d279a5ee9e4246b417f245dc33d52e2282e37738debf5825ed072bb2f59ec61d7792;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hab7477645320bc4c403b64a978d9401a7cd5ff5c0ad946a529adbbf83977b40de23f4fe3001e118eac91db3b235a131bd60cb8ac94134ec7ff64e23f93a75d47b5249cfba47f6024e397192ea19a947c83a023c47b5a69ff508de74c2d5f59e048c54926b9fdbb38486e5982a04b34b41;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'haa3d14f430202fd0f4319d937c22b4a33d2594fb8e77ef44cd5935f3ffb44cdebe61c148da9ca9f2cad281144239a4a432273a15a20df112582fe0033633becf31ae166b94cfee48bb0c15b4240bbc7b639c38c57f2d2aa54069bae8b05049b4a0476d7fe50e9eea11e7415bf2e7b1a05;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2b223f1e897e8a0b99c7329fa3892409711f2886587daf22b59ea72b7eca53e3cfc6d07c6ef07f40f3ffdf0ed9ab604305701874c2978f1529c2195950dab820ede0798dc2d72cf553ead4cfd53bd8ce8fb8292f9aea73c6d5d47626791b81427cd403e4d0e63a5373c586ada28c7e3e4;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h23b4a711b6ae1d341ea5f885c0573419433dad35464c30801a7789bb56bb2a280e4d3d0f328d59257b27a2ebed1d39e8e968908ec09fe6004727d0e24315ea946d8a5b452ae837f542396beefe10c55b5508cf7fe9f6384374b6866159745fa6e4d404b71b1a01087a7178f30cd9640cd;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6016e7f40f4c4fa6f7d02241fdec7941de1062c5e6ad658051f65ed656ad3a59ac7b9e83721861e62ac85283c2d0946138e1145360b0b994e3bf78c47847434ee7057452cf5b5e6747b38f7d4ebe44c4ce109d9d71d804268eba6dc64c6cbd6e009f5f8a2f798f4ccb5040c9ea9882b3e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1926c4ce333b6102dcf295ca109e4ffd4691d2ce4f3f2036d59bb766cb21f3cafa7a309a6bae23299692ae41a7a24d085e9f7a6044975d3b3b23828bc98d0b30e932633990c70822d8fe443f784a0c698ec2025d7cb1c5452fc6a99dcd7d639c03a5411883801911e532f3264de987dbf;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2f8fa76b9cbd7bdf1f9d58f7e0df204c837b8a07f72105f241729d822210c25062c118c125c15c836f9cd64a48d91f55ba0fd6de01ca1601d4745ab908a8a5fee926891a54fa25479e874dd0b49641ab0b76ce8d84525c04e57af4ebd7ce77ad8edfa38bd48bf70c3ea7d322f779a5d0b;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf3ab1c08f0afc5d1b616654858d2dbc6ebf70402ecf6cf19b8dae81346093bb0abd373b4b9f1b03ffefc47ebf4bca5f992b85475cdd144f21611c75abed0a498a3bcf99d1763e85b88fee7072aa1e21a50742893f3ab8b17f2393ae2cb7c32683ed65488a25799b4b798a78423ad99475;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h891822ea5cfaa345572fceafc4d82a69b993e6f4286a55d70912e09038d9a39db95ff19e8fd484acec8ba536eed62bed656b49200053c5aa27f33a1278acb564be0a4063dc68c3310573c6b91deacb7362fa2ef4259b1c9f95c0471e740c39d4a94f89c645815ecdd0788a2d608227a8b;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h89f76ed8d5da448f7ebd85b5c802ce0aa48a4399f839d97d914b87d0d14edae39da062c7b5f37d05f898ecfd1c20a3e6d1eee477f40226428b4ce291c6acd5605129ed2eda0151592615ce46cbb5edbdee95eb6d0306419c43047b8bcaa03d303f010468b74fdca08341d174a79741258;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd351f1ecf0e43aaef8ee0c8d95f6a291c60045e5372c8e710f87b41544fc5ce2f9b7ed4f8f224f5ca943d0bf2f62a59f8a319511314b5e53cec6be4619414964982d764821c7275167675da9ec5cd457bc00b2a6bb77eff890a793ce9508bd4cb1cc8a3be3b7c289eaa8ded3b0c42f8ed;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd1310d3a0ffa172c7166616899d34cc7dddf94741449d8c1768ad5a2497aac2a1968a689434db5ac297b580ce854794e60ea115a79556b096eb9adf48096b3f589c7ac69fe4d61993d2f33d7247e99e4d01b5943d2f004b1cacc2c397d79532a0cd52bdb38bc89e7cd6f0ad15a7953941;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2bc48652db8a31f7b6661841123e3ba15d9c34a5c9a161874a859d3378d47f77a2402362ca7c76458c4c28da48a075fd865500f7fcd2797f40f73a273b5ea7f91f26528f11323625c6a4d8ba8d5888789a5aa66c2293069cf85539853be81a8b974803878b3e4ce583aeb28f416ce576c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'haf47fe5db507d3216702d23f1c4fb2249de7caee0e89ae91dc5146642ddbfd2b4e66055ce1e2314cf81bc3259a03089a38baf19cce1edb00b2de2020955112c4c68b2b8cfe6d4d5a3f25fb34c65209ad23c8dc982dec9b58fd91ffbbb980b39b516e5aebe8d149a95f94bcd74515a0f1e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he429caf065d67a9c053881c0b7c6719672ae28802c8517b19045340b83f1197d5309c8c3761f433ea93b479b7ce59b5512f2002ce5538fe2d6277bf4ca9afbe8bee1fc5b5af3e04ba76ba78c2acc295ef1d194f3be43dabe8e1ae8918971fd611238c56f4d930e5cada44c86ced039936;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha39dd1b19d985c75725f983745df01ec4cc396c13abd340808de3d54801b1cbda2dde1d56ea296baaab5011a9aca6963faaf9a06f47ed18337d5cdf580bfae5e500a4bfb3eac7455066af00ce8e52b80ca022d8b247d6973c99ff295302886881e76524c61fd45e1fe745753a6bfb122;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h31528fe99e80fb51b63f2c36eb22175f3cbb0cfdcaea92aee30f819c3708edcd42db1476f6536c77e0723ee205e7d3c40cb4128c150f6af8ca196d803dafee9d2ff8b70da5e056a102a0f50eeafa33d42b30597cdf3bedee8f8f36a2b935c3cc2cfc0177cd422c1a9bec6583c475d95df;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha46ff64f3605080c5d45dd8d8eda56a23612845c25bf3fc944b8bfea78e252cab3a5cad7da492e473ccbb9314b2e1ea0027185bed839e77688d242c7b9cc95e209cb1b0454ae709540042cfa853170ea3f539b3461fcd5bbac84380a2557034c5c48ddebbc6f03f3d34159382a96755c1;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8c44dbd03f44414f921f54e9596e05eae1b27c88a0c6184bfbb9e73d1a04e702a96346f9de536c5a645657c19758973d2246f6a64196104b8b2b1420cb90b744a4a5bab761d94ec8b3ec48aa8341c31929b75701bcb3363ec7a88d6db17ecb8d051929d67880532007d0cebde1733805b;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he0bd318d328478ba2eae4042f1957ff03fcec4cbacdc614889005c72f8745f7d906a931f9b64a831871086d2f80d28dd21b44a5d0e4b2649dfa5ed79ec385dd8f7b583766d47133d5e8dbcf6bb3db1380595411e749be4396b4ae46b365393f34869a28f26905518d794f9b28c1543aa7;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd03a98f23d4853e94df2f450ed19bc8555d96e90da0c4f55c07af59079cdc14e83f4aca95652eb31f495e3308c7f7d1878ff61eb82f1d6af61eb05141e08fdc459308f888ef2c5941d4db7f78a39476d592ae0eb3acbfc5702504eaa8df384ddb926b5e36af2e92ae17c5eea187fddfda;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd8cb6e7c53709f220ad698b3aca61cdef6af2d956ccdb112662f21c6699835577ffab657f5446d4389896fd83c479a20f4f97dbfc371c386372c932c14e8096379603b9fd35bf1eabc42922e93482bc701e2b9b57a1c45ee882b688a869aa6341746eafe0852fc29827f1964a1d491525;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6c4fcea0ecb766defea7947b42b0ecba12dc0abd98f3825f3e9041438b78aa201f9e9ceeac69444e04659bf167ec169994e7bc1ad9c55d06bb5d32b660b2a127f555cf6a76cfa7eafbaaedb2a5804b966311bbaa132a240cd3a4f5d2ecfa952e975dc8d6dac34cd05b206942ae1dc6430;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h516b0b5fdf47e5711ceff967feafd5d3315a3687aeccb08a4dea9d155fe4b781e844be728656266a45718eb25e4ba2d028250b8b29a3422dcdf9b4666080bbf6bf66195beecdadeb1e7adc3d9d548ce254d7e0d7734301ed3023bbce4684e48137b2032f75656151ee200a6463ae0e86c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb93f1577896d47ae5b8ce97ab6dd530bef2ab51e19fb5df4e7ef18aef092462e79cc6b2f8a23f79314f2a5231d06970196c91fe4460272cfee2752f566ab16ce6c7dad0ca2054c66f1346ebb613a381ea5788ffe79408ed7e3c9c17d81e9e124b85310fdc0e7bf640cd88baeab83319c4;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h735a1936e842dcfa569f4dc8a7fc88089d10a99436d3effa200d3e14a349a4de5171b65e03210a9f9b9a49c050c06e7eed75c4b8dac6cf03d72e595e034751055c9da9f0b52fd9ff1abc8096e048158f1bfce5dcba92eb4f37f2d20dfaaa727d7b652bde01e02cdd9ad0a7ffb20278ca9;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hff949205bb3e8c7c24969277039892c3a815829bd0bda2b81b1e72a9aa1565f3d0ebddd93057b761c36c11a67878da554f25af0154877a4f22428075da0f10d105bd0175be5332b88b008b1bf5b8323e5ab9ac611aded0eab9123984ea5c6ccd66b2bf029d3b52c6a970daca113f157e6;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb1f0b8e0c75bf46877a9d05b40269a2afb6e72bc577b0ece99811fc50c62840beeb9d37c9824299f2af5b89b7ab780dbad1512c9978081a1413641398d651899ac44838ed6c7e2b1bab1ffc4f1e75c460cbdd4d217e1d22d7fe4e4372d6e1dce95def796f5d046c06ada00143c9cc34b2;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h51ed030c0e3b93c469b9b52b0ce9c335bd9ae34577a1e2a56e24ac8fa52b59bad645a940a3e2743485bf84a5b80f71829f11f16d67bf074130b0110f72e99f23595f108e72a17d4e02b045aa85e278c1217d0142c6257e31511e82d43a341066c639edaa0cfeb37d862f3a37d488bb39e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h933511436d815d136c3fc38d860e6b54a927ae0b0a801a57a583f4eea1298ec9a6718a52a87cb3c6cf590b77ac176d8b0a09efd4a35952d91eba594cc3f4878f68d71526657c4b930d104e7032706b7fd8a251ec76a438f0e9037ba374c04b3231f546aa03265570aeed956260c1190e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2ca9593507491e1c188a674c3cc40047ea6b263718f42bda96bfda6fd206a61da86a1d0b223a39dc599a45b3a3a9353fc3aacce18a6d14fa9becb56678bba830571059fae434a3322c08cf16e2989940a6da3d902d3b9a6af36ebbd4912f67044f8eea772b1c690e49c8f0a3e0d59d459;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6cf531036fb0d6cf93e38fd0f7a691a0207871eb3e8a099fabccdbb6cf250a7be83bec40d45ad175e0dfb589bc81ee6c9142b8d5cd8254341443ea567f6c36d1c388b0b4cb6a8e7f28b2f54a75d18fecead37c79fa2410b1569de8a8ea6bd67d219b35cd82ebd1651b1729b97132cb62d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h250444f4983b19211ae8a30dfa3a6987de8edfb8f5c2191e5ba78431fe0c4a9f2accfe2f8efa68af944f8100d5c80530bfa86b724c25e5cbf80b22f38dc367b5dee1f9a2d516f44a109cf4e82ba57746185db598b17bd6c98fcf221d5a5872d8846338220ef593dd193ee9548c70c80ec;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9f9103763919f6fbad8218364feffdf1740146bf8e5e6bc1f9eba72214cd4e2638f81f4973cf85d1773d47d047f5260a9cc1035227d64a68c402137257d264cc90607e7c71253d0e98303d2208ec4fb748fe7a0413cf81f788ce0ac5a7c1d161093e9cb172324541dab3a7ff0d64d6e7e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he9524b5ce5ad3178c3b59b8efbcd52d4810597a713aeb6be2400774c6838922f849f5689733b7d946b74dab7e437fbf5246cb383bed979e25030a7a3b8d3ce62af827a057b94a155f649c7d6e812189ca80ee1f9e507ec11d8b1eeee7f91ef3fa4eddd6e00dcd5690329f7727d051a314;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h220e0796cb6d423c3a3b01b1139a299b91bfd2b550553126f184e6d90c5a3518c7924eee251cbe85ea92cbdc31fe5f97af5a074faa65a3806ac7b502aa337a0f9039a5bebaa79f61a178f573de876a577148f07a720650efe368f19be49f49e5c30f3090c8171138d54377dd97639f16e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'heffc74e17ae2879d77118fb31882151aba36f289747a4b77a3735ce133e8d4a71e2550d5813c01608d9436abfa6609f2eff973d887604f54297652985810f8bb82aab38097f090ead99111b025759b9a8104f683c3567605638b4abd4a68de32e0a5838c05d226f8a32d833ff89abc13d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hba0417f2d080ab90895294f1265074ded014e555effc14b3741a4eb982bdb0033f52019daed928df07a85bb07fea156668e3134af09dcb50780fbbab58b082ccb87916126988d28daabd502652c2105599d7a9dd1d4ffc27b954b58f7b4989ed85c6129a8bbe4eb48e90d4cf42e5fc10e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9ba805e37860e2b44d3c32b0245de16385cc0a7e971948467fc57a7c3c7b4317d5851e25a381c02db8464a8e1af5bfd3c9fe43c19a10435edad64da617808fcc6bdf2cf35d4c41f87537ab3508ba6b1c1ae538773948acef3fe243717306940a2279177db3b7e50f513952476399ddb0d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8cacad15acfc20f28ce514be4b3aba9248d76f4ace89bd7a8edf7961bb1dd2d311b6e410c63de83fe71477412a3b28f31bc51e7c1bd1a326a7f285b5fac704da38392fb63448f78cb38bec225048fb264479e6b2e062c2aaced158aaea195c0b0579d5da3146e3b705f58468e0c0cea0c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbef18f0fd6bcde4b5045092434905fefcdbe325df50219f2ea57836c1f68d24b88749058c8f7dfe9d7848283cee42e1705802c3921eb7ee7783bec8175bd1eb5340d029dbce0b5989bf6fe83a4446149d88968417b223cb03436cda821cc58abc93460ff05c53a8e381b4ae14a516615b;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h89ad7311c18c1da1b5cfca27bb91295f5f89602c7253198bdf0ff6acdb9a04b815a17d4dc7b611ce6954f34239e4eeff9ec68fa34ec07ff60f1de6dc4fc173c5aeecceb5bb409ff1dffe227cd5a62ad274ce87c7ac8bca1109416c95258735d2dc606dbed3f6ecf808b17f312797d67dd;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1513b1191ce35b2209fd65e59acb4320c31b4bf3c6df925b4611cbc6f32b67914cc9a41ba738f1c4f59a9d0a79d6d90c973512bc4e471dbe7a501765c2cacd4804d63430aef522bab501c265be83dfcb187ad93d02a1d04bd1621bd8c83233f0ff4db0d0f94e094d5007c38c03fb414c9;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h66a0c40301ed6d502652a453ea8b6b44175cb09c12a88b50e2d1e4b733b673e203bd626aeaa76927bbc22472ca45ddba9a32ea42dfe2110c8fa6c9e21bbc00be60aa5be07c07e2e7e68f69a865026300d9a51e296342e3888f8feb6bd4c0e107c2dd5e0a1943c6eea2894111c0123ead0;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h34efbbddb208e99cb06286049a5f95788d7e0c12d3ac77bf219a26f85e3891810d77c2153994ccbbc92ac1f2646576896a6fdfb88bcfb13369b3b98b27bb2bb313439a8f3031a7aff9d5326b9e9ecde9df17acfd188daaea479e426bb3de5cb166d707db932598db6aedf55361dda896e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6cd8c7dcb088e3128de66a59e57b3d3efbe304578bb020b4841ba017f737711a6d1fbb23f973b75b45e112a089626f2a058166402dae26b8e1fd31320c36f98dcd4fe3d351595018d3180224303b2e6826424839494097e60817137d1cc7ef31df7ad99db58ad66869756526c83c2a101;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5a9928d9e1af25030f53c688c8be7ad20b0ac32137e3156e43858644620822bb28e33930aed5a3c872a1f2075a35866ba5c7ed7d002ac9ddc518102dc8c2554135bc9287bb0fa5994cc6698dc93403fff2e0ec3cbcd47c800c3f7261771098686529b101378749b7a29c51f33364a7818;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb96793a3f1114811b63f70c22df8274f7e13a62cb7bdea749b9d9007dd03be760d414cd42f3570fa4e772f821c48dd84469dd23610f4220f02a9cedf391e02f22e81694dfb79e09489ecf0de811020c4446bfe34a148a6d3b3d740596f93f9c8b4971a947f127abf735e357e5ef8c6e5c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h956d283cb1dfa9a0d5b9924a167728dcf4cfbfba267dd5471fdbf98d384ee32b54ff3f7973d9ca0cdb8e28a45f715651013d3b56741c8f6593ed8693521f929d9462ffae0e7b6425778568d2b4f94e0e5fdb6299eef5724d844f68ad1a7f1f9fbed2dbd5afb61e5857a12bd81b131704a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he6eeb955af2b831ab8be845fdfad8d71de0d39e99704f990437fd746ad389a4ebffe5f74610f25f87ad61067ba8c937c2a09e9ff15b54c1b64c5687021b0014f33379c6d6cb3224d0ce04b82ce3f63949d882454da85dd8d9552339285397aa61fd1c57e72285ce7fa092d9996a413de2;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9542215adb7e22f95a6cbd0c063e3d643a55d9129f7da8d584d0587a87c8d2928cf72d034f6b86646981acb5afd25dc5e05b24fda795f151b7b65d2ac4051647f79d2627af51f451a5d09f406ce7ff8cfa988e5bc0edc96fbd5b32c42b686acec6b00625de73694f4ceaf41f8cf639d2f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha9482c0407ce60f75f69468836ac882aaff5e2c48f10f3514e1438423b228864cee15c09f64f189b113d69547d2f10deb09c4267759589ea7066171e31d62d02d48ae7fea9c53e8f4f2fa1d429cd5562ad20ed6a3e7d13714800ab3b21f82b77fc26c2f4ce313f3b4d86bfd1474de6899;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf9bbffe108668ec302025bd1742deafb70f78de3acf24d726a29452e548246e4494c5592f29cab96caa707fa1e7a5076705caa93d4c07fc0e997c31ad6290d00431100b809788209f9c402a67b7b42aeaa40c7b03d8cdd2e66f8ed701f6b945137ac6a894df4d02e880bec80fcb2ee300;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9e131e84af0204fffd561995d59012920df906be046d8cbc1a71d40d883e7d4e37626d19dbebf0f36e7d4f0f92811650b266b933de66a83dc569fe655b9e869ca45dbc4adac689eb0c83cd642d8a4cc3ece61113b312279e96f079d85eb949abf8a686b958390001a9d49b5824bef100a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8eff8c4cfa15cc36c9afc4a147e550d9b966c80bb1dff0ef89615c6671d437c63e83d44819a6fcaa5bc8989b99a86289088a4ba7a0e4d8b1c51afcdbf86a6673487e29139011ba4df6f18f7e78518a99c5573b885b4081ad72fbcb293218de0988f342ecdb5cb3d744633a0257f3986bf;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1bbed2063f22cc90ddec1114e7654286cf09c61570de5adcf227e82e6393c800e6d41e09d0a456262ee974bfc912219afda801c71036f3a0cce2c09f84038d6567a19dd859aa9d4cea7cc853d0ca8f8a2e74ed9ee7d0d7319d692af3abe7938b38eed6d115f5acab33006af3de652725a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2af4ffa9d2fec0782dee7e08a74a3aa5f671e64356ac9f96167e774348ed1684077c93a146911af099dfa86bee5c49e5a05acbd84757ca810419cf93b04f57ae91bf31271dbeda69aa447c885f6da1f45ebfad580ab7bedcbc528e33cfcd178027fdd28ad1b6cb823ec1635b8c6a5af47;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6fc83f5ec129d96c84f2b4441babc9e48cda3f003d0dc86d321cf555af6ee3c961d5fce6a3f9197bf11940685b7db762af80062992f16589f6259e269378524ece46b80ed1920961a922e0746969c2287ca00f188666c281659b1f39f4317fa5c9619612ed8c8a5e5c99fa95904766137;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9b5e247745fbfa019f65d09a14e0685ce250f9854d7944d16d27bca3cda5f339063a906b9efef6b29643c62a769f01a7d8483529cfa03ddd74197e7588fa9dd2c42335adc683a5f8be449d88d61b692992accfcffb576061c671ccf0cea2422164efb1fd19aafadcf92fb4c58017d4caa;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3043d7ff11aaaff5863271498f2ddc10ea4e8453b1c65286301920b6d0c3f7fe8698d1dc843f580f6bba64b6ae2cca8471705d6fc3b8e1772617ee795ceb8bdbf3908297c591e1059152ec86e07316254d03053af1a4249603d5f75a46247f3b8ea21ca9613d9fc11d7a15855a53ab0e1;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3a87f3b163b04c2e6973e80fac4ca5c1848a1380df72052de274ec81d2b97e6c1fe9d101ca0896c93e544e56e3a90417f39df991117fd6a86d3894fad46df5954f84d2e266aac180124a1468a36a3a525d92a7529ff2ca8ee613bbd9d623994a3ad2ae65c4d486217c2a370923899a370;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6f1d76595a0b33e9df0ae8c2a88956118bb3a64ee65dfaa9585de93a296d41755d900b01f2de9c1908d693b7f5c181ce4c8b5c74ebc872a76458f4d8462e34a7c59422a3e354cea75f52ad66c85663486f5190bf878406a1f5983566e2d13b0181d413088a660e9b82d510a4a8cfa8995;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4566dd5ce3cd48a1835ed25accf421943cdb0e36209680e5b1f5b72bf18a2bb227ea5584fb1120c39a198919e954f246fc41fdef4b747596089ec3c12e542918221a49734773f0119905b7ac4865d0974b0c12633e171fee5d364ca34b476c57d27ac7eece9df23ee941ba311061ed92a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8718dc7f29ad8b014d5ce719f707d8a1b0197e6a2efc6b876feae4d68741bb20bce5acfd8ae0f6abd9926b72fd5746ad7bca96cb44c9e1769c99816eca7afaa8116ef380afb3f526ba25e64ad2277a327a7e393188a2f20134a76d2dffec2092248477711738d28a607846292035263d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7ae2b108df856154f88e577e43a24e3a21ead66ae4e99d23403976e957f4f2b537e129959db240993857d5b18bfb57321bfa90aa5b7902b87a00e19a97775a33d2c1057b34a596783dc472fd45730a3290cfc14071bec967d6787fa72eba2237b8e5b365ca6c9e6cb3b66b39553e03f8a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfaa77d8e75550b9a34de2ffdb52e3c97adcf1e92d864e9138f381602136d4d5f429c227548b383d168a80c2ea2c8c4e43bdf803fe1bae5347fe540ef0722819d60d635ddb9dcc25991f1829959ca19fea0579ec0d7b63d55369e321e2b129a9db474489f7e4d536def07e99005b439a88;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8e3ec6ac9464fb858459d27b77e6a7fd9cf016496b95556ea658f4f6f657df3a6b56834464365f52cac85b5f0b5535a4f762e035b9ad6d3c34f6113fbb8967df8700ab301f00a972e428f86e5f7e054c0903916a7b4a3c6cd6f65306cfd15319f46de7f91a8f363a2023f97ab41bd1004;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h62ddb0f383fcf6884108a79d01889bba147480fefe2f645134bb3bed94d9292e1fca842a4326b988dfc036eecd718d9134d165b9030000714913c864c327900d6a0cd496d6ee4cd016a81c0a5c942ecaddf107e37fdca08a18d181ef2d003b945bc7fb5a7365d80fb20e800e124da90a8;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hae010f3e657faf154f4faf4e39bbcc4a853905c38065508e286e00c56965c34bf2a07fba8a2f67cbba2ab0057f29b8d884f840e84c6678184b15da2ec4bc27064dcaa08b773ebfd995ab503b376f7e084cdaddb66e58a087ce814b0647d2e342be16e7cfe0990ffe937e8f0c8c8d524e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4bcae6d2186b74d0ec7bfcaefb301a6171c9482f9c909b04263b9a2a0352a133d69dd4efbee0d9fef24d244036e5cf9a520b44087d9ed184120e9adf7c6059a4f4b75484c1ec768fd7b6246683d2a7e899a16abccf9f3bd07d16f0555c7873f98a857596fda487f84fe18d8eea488db79;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h51b59a4979366d1f6ab0c18bd1a04fa76ccc5a4599332d6f93b922e2b6fda00ce16ba5e4529de3b30dfbb71073124196a4659654aaa7651db7ffd3fd98df141c94417541c42f58e551bd6e1c59db5d501cd5cfd36ed380009e3bf48ffdbb6d3ab2b235acfb55ab2044710af35ead350b9;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h79b650caeef71b9a4ae93ba99ede5f1ff4c396f5a267964021daea539d49aec701987bb556d8f9ea0e9da560c7070896b109ea1610a181ae765749ab7b8253a7df48db53fb113317b91ea657c5d9a62a7dae2f98015597802779ccb55f42dfd20f8e59a14bd7b991bdc5cf0a0868df29b;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdce8676adc3cde9b6869648a98fc1aeda99c231b2e6f7609f5ae25541d8697c647307fdb4a769ead34a90c30db54e752c28649c1cdb615d5fc579a50e9c316ce9177289185a69f6e724217380bebc8ec3ed8dde43e5ef4876ef12529ebf0755aad4ecbedf2c00e57ce8e599ff74c71be7;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2dac2c3afd12331d962bfc7a07d1ab7aac8c74ed2e4666434ad64e8593adaf7d71ba25b7eefd648b76ca3fb2afc4d58a99d526c458b85cf5d9ce0f19d33c7b79178be32b58d25f0e79424b7d990c53aa3e3433e1309f4458e7e688c3c1424da7f912fe67dbe8e8bc1077c185e3c9c0dad;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hca2d6602c1e9fd5c0baf752409d1e1e817543630eababf57c66ef2d727c0c6c1a0ce7d82ff85270592277ec28c730941ed4132913dd6c574f104bd8372eca909e31e113219c7e6d53bb81c813e7ab90c38dc85c958128028c677e47b851be2e87294b16d8d3f4056bb068d85231d9d6a7;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2e729668ebd3ba4676ae4214eb6bd26562457f373231d11b91a2a6f5a3e446071219d4a0779d54a7451a68ec89907780abbc3905b37d016b2706a31a1aa719ee4cfe98e84628b5738b209582e9c7dd351e6c3643ecd22c0384e1bd8598745b2318aa7eb46c51480b3d7e93842ce7d8666;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3cdd6a4aecd617cfddd9e96e8ee927e60f7e3d549f6d5f5772fb6ba74fdb15b9b2606fca55a205405059736dc57e3d4f9b88aebb7df51d59e1cc4b82fae754c65c3e3448f83c15770e804b7d5f85e3f788a27c9eb7734d7f46364dc43a06090bc251c961fd29b568102865f344f387756;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h43d043a37cd25f4c2c99e16da83abaeb09358e7f94c1ede785e53800c503a2780133939f175e335405800eac1948bdc8757a3eda0557a5c771c51d02c7e87b33c5c1f7819bc7d2006937f312bd8221ddd33094f5399c72d9f95480c9e1a5d9891ff57eb9f2dd71a5b59d05eaad31c4b70;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'haf93cedcdf2c137c4ac9e673799cf60d6de7f53a5341c3836223b3a41e9bff91c92a1725b7f1b0307aa4bdff5ffc3aabc45ec4b03ee2cdbaafbbf378d59b92b5ab4dcda23fd592aae385038afe60d89e3952c75e0a5effd85e0f5306989de00250e5e6380f35cc83591f916a307bae338;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4929323bbc5ba53f476d38bd88c4bcdeeb68a5774708162c26bb29ee15a2c675ecdea5dc4d9df406c1e35df9ba9eefdf8ee73aead4000100869e6bacace8ac5b013486958257d4c77a518c1fd00375bb681da06ce2b5bf13fec3e52d5fd8e313f164035ae031aa4d2a29ff84cb717176b;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h63e4b8aa7e6004968c62cc74543e614a63f43df0eb2a15773bd7ac582a3bf272c8ea6eed4fbed6a017f415e4890428b208a886172524ef5f27d05dc799cc1fb981579014662c86f81546db98c74d2d186341c38437705092c2e0a4460bee44eafab9f073e63023c3db4959807e37fb0f0;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc1f2357206135d59f2a6d1d7fbf76f9af79aa394f427b2c5e46db6cadd3e0c983386b35249911609e30e428fda2fb00518511b2a9a6a7a27dfb1cd285fb72bfaf8080d1f01dc08faf49544af697c58caa2f0ba1d893240e7e5758f6adcb8c61c4d5258cbd413a79629b821a753eee2554;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3aec6218f6905d97cf2d11d74fd419de2972f1e82185429a7badf33fde2929434aab9ef56e2fa05b6a9cee27a8a329bdc06a2dbd028d2b06086645ae44be1096ce09744f84282513c9120a4f54eb70c7c41347a7fb5a23ea31e507832a3b1f859fd62f1bfc94ae1283f49319b8bb1aaeb;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3d3aa232b1fae024add0d023c2666d24b2941c0ec1c6cefbdbf5edd3da2f255c5967e75d4c9037b1d60a88ab73028d0107887d8f1af7e3c7e67330467c09fba757b90c33be0924505a18371d4a86ae5493ab61682bb0890598c9b757b442fb1e1c4923fe0921a4094c491bbd34394ddd;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h24b61885a4a43b3ddd134b3a2fb33e3fd8bb27f15e410409bc66415eb31ca306e952eebe47c7882ba2fe39981b515e3f9b9b013393b4b94e0f060e973af5192da96bdf05587d1748baa988a32da2c26449ddfd56f45268fb45f18f7304cae8d6788255f5a7bcca33503cb2316c5635712;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7ef46d630b6dc8be7552e99aec70e053d6bc041b4612421a8d79f233caa5629f1c405f6e4c026c5a35861164ffdfda8e8842491a78d5c1702b2e535847fc54126ca775b258e3cee18385882014d9c76eeb5e6634e9c6cd7cae6989f2c7c53f8c89e7657479ebde26ab347e7617db2c40f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3caea91b747cec29c8e90bf65b71ae41f63762be7e43a017f72b28d4f00c47b93ead5bb06ca6878cf9ff3eaf437982332e6511761adb1ad51e349507344f41e125cdc920cd204e757b840a931e9c43280392c8b4eec3b8a368a5f30f10082e1b32c2728122dcd31308465944bc6730572;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7d0e62e2a8ba16b62b4a41285f1d2743904976e0e924d46186468a5be1839605057c21bf1a81dbd2e68329302fb8a7f31c4fbfe85764d71ddbf0ddb0f62ba6fe3268976f15786788bff805c31801cd1c561b6fd6078ee1b6ac4ac954274a20f2166a7855aabc4b8ef20e10b112011beeb;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6f22b060b13e3d1aed54a8f5a753046ab97d9f3a1a271cbd66d02af722b91a10bae03d549865fea5fc8fbac92cfa53c6a5857d607531b4a95ee23c9b45c31c807525e7138b9cec1e579f9a841f7bc94dc8c04218e616e9b4671c4ce8594e1861f432b82717a569d064d599d92d09ff479;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1cdf5317200eec3b9de08db742c0de6e5722311baee4034f1b7fb693b08bbacffed3b56d052f787c7efdc6d845ad9269a79d2e6ceaa40436d058e6adbb4a813f61bb3af2d393110c5a900c9eda2d7ef12b44e7e45ece243d26378fc14156e6c5184d2e1e86b1e97aff37d25a8e16d3b61;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h995933fe18c9e3c775c19e19c25c1538f0e2bc89e35e07a81490b612c0539385d0f6da20ed1450721f61bbcaa6f68021cdce4ea339f312cafd5d4a5af61ae5f073b3f3a5d7a4eb123bef01d0d9e2836e0a2256d2144cad746214f68ca9d9b582eafebd66fe46bcc44432d80c1656c86bc;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h95681632ac79d9959badcf8f4a8c001039bef975ecd941d2284f057ead793affc222b00aa0d40ab1c38b7ac702d48e0fc43ae8600d5ba8fb82f737191f8536b142c1a55696f5d873211cc92a3116898d3ef4d2bc617c170d26c94c8d127c24ef7540e777029de4a5388ca11c008dd0041;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he3a8040dda526e06e99fe6fd4a5c3e7387c2345d8cff644d6a112ef0235622c7ca0cdc8a89e33bfa476c5b32a5162f842a64a490037a76cc00b31590d0169cd766d03b82f8ce824c54ee0d97811c153712860d07804deea0c27afa9ebf6c69f8242bcfb437d8f0e46bd5e4255325170c2;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4fb65de9480d39ff00e8645f429cb9ea192a74fb0b0f138584ecde033fd2890f56915c3a01dee2975908a2d687ac58dabb0186f384bc656e76d459ad44eb5d7bcf1bcb7c022eb2742f1e995e9bb0f11827fbe23aa0c0b38948b475a55de0ad52ce35b6b18bf664913d5547e969ec6d79e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h35c455ec9a7c583e3801d0d75829721c9547cfce3d78e650d976246354bb1d2dfd8e2dc9a89e116654ae9dfb82db7a5f70fea32a333ec2a90a4c9ed008f612c36f24cb78b393487dcde0a50ed50f90b38696337de8ccd00ebee456c363d3d9f344f72f3b521012a538c17244e219aa3f6;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd9d69b3203b5d50ee93783499ae14acfd6d39ec4804fb12666d70d8df8eab8dc498eee53ffa96fcb4f69f624f0dbc7546b61f4fe7de4adfb858c9fb1b6c7de8520c5fa2a83c92f0c385de52f849c4f806a05679a79303163fee65db042ac30796c187ba3098f07d353b0c49b7316f3b3e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf8f9a0974a05458fbb478ec203f862f3bf6ed6df503b5132a159954b695a910e63bd64ff54c07beaa0e0921f85afe562b91908d490f8e6402af0a42bb6bf04289e8586442361f2565346c4ef8bf22ead572e1f63b73253c479a78508e9151ec78e61214ee4602cb203adf7f3ad2caf859;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha06dc0aeea715552df2e3a9a87bedbaec6ba207bdc1637dfb7e00509ccbcb56121f3c36444a2b02f7295ff1a2d63964db3d29eec0eab80e8753d77496188b8a41271433c42051d43eaad1bb4719a6f0dd18616dff8df4bce2834ec60ac107cdb55de9931152dba14ef57f31d3ba4cea13;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3138fa03555b6027476155e7b84e00ca4f28dce91342291431cedffb645498b9a74bb0e5fcde2a6ab3dc768ee89a156d774c4c3e007195f0436b84e51213293829a1cb57eef8e0e1ea39cc5bdfb181bdb5b44b65e3239499d11a2d62f2126db479e03cf4fa9e57cfd45dfbabdc8b07b4c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h60bcded2d54d8c8e2094667cf641e200ada47d2e3024456d4201e37ab024fdda4c1babbdc96be4b768dae74441d31b8a238ab746ec60d72ef15b48e8e9d31752a3db06a1a1810d1c326d4218449f852824d5cb69afc8f56c13567de762d205ccfbed4b5bc75ef5f513ef807af88b0e62f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb19b780fe7d6299276979f98068cca95bc3d3baedc7104bc6a371db24b208b709ac02c7929e4e323b67c93cc139fedb8e5205cb8582a0a73bf1f6f7320e463a1db3cbaf9f12c5cce6c64a906198ad27fabd3ecb26b425b697e47c96ff9b58d6156da3e10ad4fdaffe82f039403948fcec;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hcc73a5220366a1c898cecff98048149e2ae9b7b368eb7dae7da06210dfbb409192bf3c0c406dfabf3248a641e7d980ff7f1bb9c2ec3eb4009afd9db9ff0ad9f43a80e986f957e31e954bf3d2a65482b2e01b497ec8fe7205d21d3513c813aa1c841658cb30e338270823a6658bace6533;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9010574875029268ae6e08d3d08868a4e661433f28832c69a221fcd9f6351939e5d3d05f18cabce7b6e60c40d94cd80a27601b7aaa05d9d4ab9b0d868ba350d3d0109e90ce5b5c2cc504ac8f1b738997c9234a106fa1b8201048e09d0febf4ef3f3c34baae5cd9fd59b9fec5ddec43d4c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha51d95b578aa4e132b795066daf1d777f64e068fd3b9bf98ec1bdcee8305e37692c486a30365fa7c2192cf7d97b2db83cddf4f6b32ba3389778434f91577acd4079f54d91bd92ede0d72fbe8ddb87537eb7f78d2b3068f870d663fb4f5c77f008bf53df19444b1e0614ac06406bf04e30;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hca2b5ae09a09338fab11584cf2739e922492f460c6471f4d5b8db183558d344f64a7da4991e9b64efa720c77e184cf4d8516b724d067a29ea6b6445e5a27096d18472f5b45df7d67ca0832398122c775d1447946578ebdb12f7b9ac8eca128d9da1fe421ae9c488d7cfc9a6b6d643e9a1;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc907234eb599f2a24e561e055d4280970233c3cb871751df8c10a8b554e49f87008f13c3c5a40077ad8ce3576eba6dd70914af99a3e5ce12be8c96154243dd1064624613c6e4768a22fedc1b3165296480e3ecd97c4763bc49161960f8723b26840e7a1e991bb8d66aa19afe08be34ac2;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h64eb4b5bb0ccb46d6d00575dda28dcc029e8c85931b4a8585bc7c2a787444779e762a75e6941c5b6768afb451070a97b814506164f8b1e769dc7e67002c5e2dc139cc4932f565315ae5e9dd15f82df8b865fbc292ae96ce2b490de7119b65a18ec79e31fff7da72bd71f846e0c4aef20d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf0cf53bab231c3b03f3c49ab5259e05db8050cfc4d01d0d7c91f96c143816fb75e357a0c133f24e3227f7397cc923bb1595bc18f46d649299e072e4ba00533840b1ae6c4b49793636b9b0b877de7cdd3d2ffb78668c1b0076ee752aa3cf176eb78377e19c2d6c8dad1a6d86f4f4f95df6;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h313aa65fb1b2177edd67e22b1d01fcaa7510c5d90cef9d6d397ec64413dfc7ad516eb447a83bafc16ce4cfedc1aea65b8339d812bd1adeedff1515d9818a064fb0269464f7c89f728ef626c7220b84ddd33b4f6181c595da96147b05923d11e82abe3988a3ece622742c69fd436c133f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7671f41fa8d74467c9bf494cc111dcd42170a845d03398627446e004c72ac8dc1fb92dc0dfa71cd3e57cb22e805771fcfd7c09187ebc9bf1a937eca8345f8d0aa2a2aa2c3702331655f17f6c1ca17f41ef3f1450abbe2c7feda4f62513dbea647ae5fc7977d09d747628a010f24485437;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h74006deb6d65c06e1b23c617c3e230ff1640c8bf92dd745992bec25ecfd2282d33e5f3302ea645877e4d500bcd774e86cdb3eb2b9f1338eb155fe84c68bed0f831e26faecf01759f5411f7d35930cfde92264c596dbdb6e1212696fe33240c8c1ff17f60c2ec919a1a9eb02a9a55f644;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6c9922b23544f970de7058f952efa719e332d92427c015e467256c650475dad493d4ce587ff97b7ef4c2aa42b0d05f028516e80ec6aff52107660597c2c0272b93474df9fe00bb556b2aafd1d59cebf54eb88cbe8d41e0d094c8d86804d2cde48f3e9b82faa69c73178aa36cc667263f2;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h342c8ace10d2e610840886d96eea818a447a82b193f32b72a0793d204f70cba35380f61bc60209a2079da18fdc8d0beb6d6a96f4df7130ae4be57b28e41aab0e193e12d2e3cea82cef104f946d0c2e492eb234e28cc595b7c6d16881485c8c872791d70f4d8579026a4d8861a76f87d0a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha25076eaf43cb722dbd5e3fccfe4543923180f6c7e2fda141606548afccc2800733fbfdf37495fa79cf85299598b603d87d21ae2e91545ea9d3b31c338f9f18e7746a4fcd53a8136e247825042dbaa789224a8427c24a983ab5c66915bd55452cdcac1a4b70ef448873bb61a069233bab;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h36bff5faa81091de59e4d41e87e825a7a9220095ffd15acce28408fff1d26957fecbb8c2706cb03d6312d247a58e3f5d5149eec5d1205ba1f146b3ad91eb36d138e957edd5beec8fb76bbcf6276dae1c952de7d0c1637d73b56f87a38e80879232175a5987bda5453b145fb503bd1cda8;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1286bb170af8a98e9559ea8be75042a6a1b73f7202e0137508d5b295e5fb1af8a8f3a36adc6d0b806b2c56489253f311508fa2316898f10fd3156ef14ca33928911a502da97d29058e4af6b078b30aa3ec87fea1db5a29eb5406f3e47851d6de7045fbbf30ed62b5f3c77b99580be83e0;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he3bb5ba9baf4f39a9858cdec64fbeddb64d93db29807481e920b0b7802696ec36e97ee7b60b86f581a49219ced6e86c47e977c0bdb14b4a0212654d1a251dd6728cf8009178268d470514dfa36a5d6665f7486ba2ba2ae7731594daa9290e7c8c3d11e24afb778f9e282768c5e5176197;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h93a1831d96a7cd910380af11370fa801f31c7ba7e68e4f54f2f9ab4f519d7db5645a57d3c164ad845ceee3aa57d8e312e9d856da15aaf67c2b40b1a10800b0ffc4c3d02967c463ac94d3c0e3eef70f8c61cfe72711d1c3b0b098696b8af998a5bf8c2a3d185811181792a90938c1984b9;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hce22d917d7ca851e59ec621f24269ee0a1a97fc223605bb3bfcf023c58878033933a24672c2f02b51f90408d060a0eeeb9cca67b6e434f6f69f856e2345b755de82cb7ef406ca7fa39375b11d59daff1417eb8f388a3bc3433059f4ae93bf3f29b2cac02ab41a09f45c19745e5dd7f7b7;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h45414cf463a9fff8994f37c75c7e033f4faec94f9fd966cf24362946ab0e15d51a555bcca42d87748610dd770a000319c9f51e10f83771d83ecb867b0e91dc2da64850343515022164b3f7f6237339c8a95acaac109bfcf3db0cf61d4473e0cfbc45df3c0edbc0d66c2833fa4e172f752;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hcc2ef48dbcdf98d87f7d8abd9cb93f30a6e237b76c26eb959c516b95803eade251b216485ecb5b53a6aadecb8f5fc6f93bb4b34d9600a23118026947606b3d60ae7b8bdfa1f9264b6f2881dffb2078bf56b6f0078a3228c258022627fadf3b0df5a410144f918910d2507651961c8d261;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h65c9ad5df2224196140b12bae7d2ca8412d4cdcc601fd7d726b6b649f38f5a1089ed808baa611df2bf2b3ef0591d6d56c33e13b5f3d870b3158dd5719f9f42fae91197f062b32e057a4b2b1a0662abc560d97fce18bb881d5bfbd6d42d0059a5599857e87c30beb667ef70471a83951aa;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb3c55820966441006db96c7509c506bc2e5c88409a75832e276f1c770645262d047cf4d2c00b39d226b3bd7cdcab1b00d0b4a41492959dfb296967d6fe79022ac1993b7a75ce325bd10cf62d5743af4799053b0cb92f71432b9318b9dd8fbe835573eba40e18b5926441560def8e81d4;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4e315f638d1cc531bfd8e087cb6be0eba3d1e81b33a20d6b3e4efbaa54551273e0583138ae4436fa6e81260b41a3b12fb35db64864c830452e7094664f19615ce53cc6fac5bc1a99faf877b4ba7dfc4fb97049bc8c6f64f1c370171b467d4ab20156f3d9fac6948d10e51d5f570b45517;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1bf502372ff30355228752f8402f58c4dd92dcc99be971dfcf22bf5a109a093ef56e695a46a10b687f2f06d482a0c3024dd476bcb16bfb487a0e1b9e348c24678a89df4a2c7877a1d4e12f256a52bbdf88f0d1fde6135ae2df14109cebc6cdd3b718afb7d077d85a5c9e7564ff8cf7757;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb5c2396b3ff375b917a451bbeeea65a5d92e6bf9c7e4e2722c257d955d1a60ef3ae3302c303f55483ca01d592f0c94bf66daddb227e70608bd7429e2565b7921d35a14e424decc75a3ce5013a322da2b984ea07bf0400f93649f45fa986be95d132b9ba16d95dca6d6f1feb9793c7f454;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb69a835960e4c27557849620c983760de416d28423fd3b9f0750196a9d2da0f07030ea1f8ffba3f4ac40bd8025ae96c9815fac85037151f0841cb3b29b14482a1b827a54d6a1a738f289c9612ed21b238b2fe21b0f476afe99a9f06c955450060a563f2ac290770abd61488b512191eeb;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb8cc2202e25dc0fd7dc65de71ae3d7acc85136b5b2cbef6144e5c2679820868c6d10aeda585ca3b92b4580d57fb6b98111437e86c27ac216a2a44c4992dfbcf6c36011a7248ccdad5e17881496077d7187ba7e9b196fe79fe033dd5467f56f9923c4c7e89793a8276a16b24e38ed9aecc;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2cb57babf9e151be1876d54ad909d96ed58519d87529c803263be9295e51575d83c51a40833db5310d2039f64d633031a20e79cc0f71edb5e70763b8468478c5e9bf05caf4b05ad80accec977de8b731fede542cbc0d6d8663f107231053fd6291158b354f62bf42b327ecb41afe70e5e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h40699e6e9d6f07523f02579f352883a9ddde9fdaa82038be61555fe6849a9cacbb3b903b5fd817dcf44ca6c28d3ea8af2f4ca51db744b252377875f54ee8ab1f0a02c027d5f31171e7df2e3dd31796492a884fbc59ac1cb776984c1fcfd3eeae9885da864d941dacb8a620263a9c13d32;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h49158f46d28015cad5683e868566ed11e2808872d32185ba13cecdc2c5e27ea2a0a6f6293166766d9058ffbd5b9fb4c489884de56cfe2bf9fd7ebe7f9556fbda4651b45cded4265bb1613211a0b27cd5ab025cdc14621b1c38a6b4c3d49009e2d2505fc1b2b00994e26f50e374b67f3f2;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2cf0bedc6b11c08d33c40dc2ba526b40c6abc3248b6f061a9d82c3251d75f66f76403ea320c19bac516d10a103fe5343bcd338acea28b926f41c445c6d7bdb19e19996391fca2b09e5333707322279e37d8891318173d737353eea6b24376fce5145a28d8eb0ac71a762951bdb4d58030;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdaf071a365be00d4e241d1c1cee6a9b1bd0798f2ce0ff07fbf569822323b777da744b5a0a0fbc75cf00a3bd7bdc7c9228a719e6e048814da0e6141793e5133962805f3ba2afe8ba52a6bd0a9beca3825e39e88ea76a856bfc81e34f39cc9d9900ef28a191b0455c613e8efea82682d567;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdb3f2e669648a5a62f8202a712ee97ec8c6263a0237253984c018b99b5c0ee4fda21307f7e096110bb7405c0f1940978196d039c628705de262ba19ac8872c47d4e8d5c3f305aa82e1ec942ff76db413590335789999aa58e5074b846927da8ba19a42364375096e718ecac336d097616;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4ea701bb2f3c1ad216ba42f6e0cbefe0229a411e053a1605eb815e300ab22c1e6dbf5b50cfa6589d58e1201f5102830d5400cbfe36128f68ea9b49ef814feeaf71aca2378004c5d3085093060f8929a5812d0036d6e305d64344ce76208145a5194f2ff7e03353dcf7c86358a2a094e53;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd9e7c02eb8fe892d35ba9b3c8110beb179032c98ae9d2f788967e29f63572e23d13866a11f866d0c0efd1b8a7dcc964f85a62cd985c99ac1c97f3dba7d8828454c210bcc729d945677be80470d0b9978e512bd88eb0a06b48b90fe3c342b5b26196ad3d90ad2fbc4ae8b81e6996b0d3d5;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h82dd39b09d2fc0642b61d02807951b77349af0caa3e38212708d71c287c7416ec4a45303a234267d9e255dc4638cab135f78546643d2cd74f3d928991f7332eb23d78b56a8d4eb85d0748eec2eef45a85998d8435f5e9f2f3a32df5c07a0c2bdb408cb413f0a0b52fcae0f542b06edaca;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h420594071b065f0fcd240fac0d420d26a91ad17d5e74cdab0550631c2a58b7687ec03534f5d4f74ed609bb1a06a8dd3c715478165fe3b8243ade11083d0f05ccf710c26794a4a069d71d7de9b7b722d79d37f9a4df65f0800f80d7c767eb51d8a8373a2783e49495fa4755baabf3048a9;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7a6696ef7e9cf04cf5b2f53967cad4cbb714bd98d0f516f0b23f22b235e0a567fc53845d4f412c055c00001052d7443ad109128db98e211bffd33f2b10e9547d674ee4745cd99946e7c3087dc5a8f49761974513f40e95f2db5b43dd9956cac00e234c9d654e1a66a3e5aef8c61ea040e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h95d82f0a976669db442f7ead8a1fda3e57709a8c58518ca8b7e5c857c5745ba3ca90c01f223f25e9f79da6ff9a45bf95cf4a7b4ccf69bbbd2f9645cb13468ede9d49d4c6e9dd9a9a77b89ec4a196510e69579ff9d4df9ca05df19544af760fccbff2a3371a887c44503f86ba46350809b;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2aca365ef091d5d745d35ba2d3a0fd8a3d4f9133d65aaa167033231f96f339e9102dba27ffe332092eeb836431edd26e7def5f861c8ee9d95d9c89fa75bbc0de5807e9558bdd352fde8205f5a3fedb7a0ee6829514234f71889f5438de9a7c3077b0462adb9a5d7f6a8fa72d219a4017c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h185519bd8f3ce16c87e8062265f1f4678a5e5989047e18d1f500c36ed806767f570da1ceed631f61ad537a4a69f6aa862d16dfeba4ba575911d672ebce62a5cc3966c0754ab2912bb603a0029154ba3474ba493d10e98b56f877bba0f8331d95a4cb4433d8b5285aaa790ab00f7000353;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h28d291bd07d916589b6bab6780fb1282d8850dd00398b304572e095f08ebfd85388e67bc8bb1e620f41ba5d208948fbdf92899802a350d8ce1578e4efc64282e4f496b2fdde0446a74194ad1fc65d7dc9bb5de55063bf64230050f07c2ca46e54884e65e044fdd59cb3afa7e66e487135;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb6099f52919e7786a66d29909f90a929cf01a64eede772e445fb581a55084b3bbd79b6fc8aa55b0b31d33bc9d941450715e5ce777f93e6b10486ed08c89c057a8784df4f5d95a944d1adb877ac94cd0f95f4fc4bac9fd644af0c7f8618900dfdd8eb3489053749364ec5e1dd22f995aa9;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha183b7accf9e24858c1a6bae07f0c7d6dc44b7e27feaa3e8a71fb8c713f744ecef8540f647391e9d26890b76640211117231007175958744217891be6b2994f87b27353a14b0ed40c331adb3474cf689b43bf0a1cd2865ce3cef2c8ebfa93e450ea3d7df7cc6ebefb1818353dbdb290f4;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha229b8c5ee2871aa5fc9d852b953cdbdcdd2ca3781c66a3b4fd6a6b43c662fa6f75ed2652312f716f6b4f7710e00d2c3b7003f0f5f0e2a9fd71775a6eef7c2d77ffa449d0fb8f13293d1605372de28a94a474fa79a825cf17f6363291c6af14201e395f56cf0c3536f1407e7fd9c18cb5;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hef8f8f5479ccf40c46378b31ed3b48c76c18e083042401cb068af8c9fcc664a125110d029a6c8c04b179e095169951e863aa2c1a598449e6954aaeef1ce5e208df04f7983784fa80f077f0c4d1fd48e0fba0b5d42fb24c7abf059c355ed8d51d249e14a1b069625e8c0581ff5d515a743;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'habb0eadc9ab858348824383a4b84515e994161dbe04f6a6b3fdca87677f8ebd5303963c2f9c054d6d849ad958b32bbaa2c8e354deec67837ffff5dfe8f5224fb5121b3ae4da9345d4ff2abe1d7df5e011ab68aed385a4eaa926ce80146dfe73f21143b97e7591a7f49e9d53234b5535b6;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdbb56f31a28ae178706259c2b2c785a859273769ce42b206faf197cdc092cb29c3071adf7bc67336547fac1bd20ddc42981677353578c545462d391e6d805f441279fcfe812ad99b67d6e9d953981c6e71df50ba35c01cee9ef826d96bf876573554f38d82bbc4de95ec52b603272628;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6bdd2363a3ecbfcf65f9be20a1a054f9232c69729b1a3d0e1c3a408ad578aaa0416d8af37ea10c59c475fa4c02579bed40cac199d4b15373e7ff36add1acaff7abe59fa028fff1ab1a108f8209240952237f7d4badb240c5e6a53f43056aa54e45c601c6f62e25898e02d2a635b3fc047;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h80c569418123f36366649904b9e830005d7a0f274fc0c1ffa134dd778f2a1cb2b9c8b7abab96217df2eaed376754598e773dcde6e31ea555114b8650787d9ace0d65cf8d856132b2dc78b0e3290e9d84cf2185810e16b7a2bd0873b33279310dd65e4fcbf3736ddab1d080e396c17ade9;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h79518a0e5b250baa57aeb7e0ed3a658865b443571105e94263e53e91b390de939d981900bcb09be357bd1abfc476e5b44d41f560960c33bc4784cbf20bfbaa01bcca7e29fcf8c8c3ae22f767825cefa81b406931bf892691bdf66db85a53692678baf992b8f86a8b14a467aad586c99c2;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4d9fb8753d6f884cdb53654f99249e314bd525739ad9fd9efee60cd509e3c02aba27d7eb6804c0b1e213b704ea530c32a399a6a6d72e4e40dab4ae6663e775c3050662b2f8946a4728549c8f33027937e59426f8cad04918aeb6a5b111f264afef98a1aa234df0107ab0ef8b1773b1fb2;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hcd5833fbd54e1cd5455e32c737b6436d51ffbb32df9b20591d601091ecdc47a02d78f671a840173dc5164cb0b643693e4c43aecb92498ca73b107b8bab85df706c9cb2a7e8119e5f70be6f7b55cbca2f02ecf8660585a7d63504402919ee1cae04a372ef01fe34bc74dfb30ca2ceca5c6;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h75b7b748aba215df825f1659d8e534b1146ceacbe2fcae4f6ff3dc01709dfbcbf7636cd365a111457c2e5e038097fe16de0cc2aee8aa146e99b8dae6b266adf67d1b940bd7e835eefc1a2f683cfd7f51560a49ca7ebc24ff7694c41ba5d7ad3513701a3340617523ddfd91c8040b9b92d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'habdb26e11825079c18dd3ca03a44c96ed0cd37830015429228d92c21632c7d0d56a0f85b7818f35786523252ed7b90e97aaa2a0c9779dc3e26b7ad2f42199893b2e2dfecaece03fa3c5a498cb03fbdb6cdb99bac26fadff415aca603e0b1f6ae96741c49cce4b6df1affb1ad29a15d2c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hcb9eea439fa3b39ce6852d1b2b2e03f0b7ce877ce39827914cbaf66edb6d6f556aca6b3db78b2c11481b3402aad4b67f27920e94d99e9ed6aca98e1d5bdf1dd039be8a876ae893402b78743a837731234e5bd432a032d4bbd2706d6d3a225bcbb012368cb47d62e09f9b1206b95b175c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc765905d2c68b0d29c66adbddaea08c9fd5f9b188ee65bc81ae237d7f3e3666467effb965d8e1b8772e56092acb0c87029bdf30f778ee8526c65985cb033378e809edc8256e0ad6ede3f078c00d5549b9825ad86a9a5f0b0ce324975d6ea528332ec9e9aa2d37f0bf55bd00eee8c51ccc;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h673ee5dacdb2f70b7214cbd646f927cd11c57745b34577fd5d6cd01eec4e2ee1fd1545d87b50a0da414f4bf0dbbec8de796441e6a86350366d6d9159f909637a9af1fa6dcaf56c908119ef623fb5685851af2d9b4d9028cb1185cd6ffdeecf018ff540405cf2ee9da0d78036e0deb6b5a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb761b22deabadc82d658c246cdd0c2bb982888574f01a96a75aa9757b360522f6c9e8f896f98108d6b057f9950b0fdd9c1bdc2d3a44521796336acf8c9b1284252db15aefc99fe01c04eac1ccea5ac4636356bfe8c758b957224366956bb495734774debe2229bf40f7d96de5f958cb48;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he1294b68d15ffdbe4b83c6557adc4f7a9836b35efb24108f9d1e55dde3212401de10b4e3c9666237018b509fc4d97c4383ea9096c1f0bf88004ff6a8863a2da5b43b6dadbea34693cd125647c55fd1fdd8e6646eeee463734d9a4185ebbe5dc81a292556f8eab10985332b93465b2532;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3462c7490c30abb68af8f845374a4b7034ade6f0d68eaf6c7902cf8552defd203bf1b2de6274ad27aca6080ddc5cc296aa173e0e63d4a60d08f0f2284db4e72f259de3b4d96c1c17c051793fd121d4d28da669721a67dd7e08afc90c887fd52f0dd249b71e15d5aa00bd5c7264f9f00d3;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h920ce4c40c9388a44760760fa12bd7b1da554dad300ab4cb720003805cb8bc7b0d9f4118afd66cbc28c89cc8d98441ca9fa22808555a5705d30e40184768d691b49a8899c7e06170acd6dc9999b5a37be612a87b27f7316a30dbdb1befc811f50fefa3526140fe7f5b0df9b57680935f6;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h70026f333f8ec46020cd00335170f2e3873615e5a94c5611f325dc42f54573334439e14fc19b9b57c4512ce64053ff1f32856ec2c506c6e659fb8d88fe06ea8edae5f1d970d66a80ef3d5c48ce493ca8af8bc219fee7ec2d8bc5e76cb797526d5cc0cd5503cad7c4482fd35154f317361;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h70b519041a23478acf0a97d7cfe120befa0b8c84b432c4337d75789c9dcff30ab4837aa148d8a40dd50e9953b06b91876a0a7213545665d5359cac8a4497973c3d570a52d0e9c1f1a8ca0b0dd66000612e00c05f7258e6d43a6ecf991e87dabed46d02f5d6f8a886f23d343af0582abe5;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2602ef6d7a438688f1a7f1f5654163edf7698cfb0fe4781fa19963b41b0a7d8da3b38d150e38a069fe27d3e184b14de0e354c1c10b43d9b6eae37e4444491e6066787f4ce8bc7c3475dfb6dfafca9258d6fafca3daea9bd5f26fa6042666c3e1f27af09635aa28c39b17b5a5cf7a979cf;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfa93fc371f017b1be1a8b787390f754c806f9256b8c55e3fab8b672c6121dd710784b681450462056d539c5706d2b103cc7878ef3b735f0982ff98a69df3ea9037740c2d03fe01fc58b37f2fbd4afd2194ad3508e1538155481ec12ddf4aaa3756c369fcc6ddfb9c62eaf6a844d6168ee;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h195b2f3a70008e2e7975e1d3eacfceae4c6191c61225829c756988e2a964093b31d219ab85fa3654d646bfe715a6f15524ce1437bcac327d99d0d2291773f725d376d613d8e5bf04791264d73ec53744aab46d4ca78e6ee3d98e3e50bd03c6ea0d7af79855bf2473fb031f72d2619a14;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h129f656aa972beddd19af89aaa7166b62b6f71f5d31a2543166646b05869f552655211054ae291fde39817cf7ac428e15adbc944caa1d718a94569ac8f6b9e70f4b93ed8611f26e4f66564ea8812d21de3230cf163a69cd3565c2206fd68d7eb8e211ab47b155fcf2630bb8ba692dbeaa;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfa03438a6f497b04209371deb90cc0fb663d2a9d58d4e1ecfd9b1ec5ecd7dc9ea72a43a69043e50e18726749522475be3df3bc60bb5833fe320e078c65ee33535f5e6dca444fcf843d921197e214186b78dbd2a853beb1a94a044d66157bb6034d86e54b9d61485ba25a5b43fc74ae3ea;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h94f9cc3f96e91bc73e72834f025e18b929b99a0aecc5166efd12987f5d4abdb2e635d42eb5c6a213033550145b5af99b499602d714ee52c2fa9412faab7ade9b843c5de133b067449332f289ccdeeb92a91ea379cc59d83b6acde2f84feab00110321c3634a80bd568521eec459a199fa;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h49a421a05a9b235529cdee45532c8c6630a301df76d2bfc3e0bf36cf95fe79a4146386a20d62119c69b4c241968af6e471e882a00f45f5e99fcb71d6bc45aaab34a24958e2f0d8b2af58f60108e961397bf108a237e63440c0bb15236a650b4fd3235358406fe09bffe2fa3de440226b5;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc4475a00a7292e2d6fde637904ab26e10e7199654e73cc87611be8aaa6bf22cde02f2c510fae0337cd09b839484754ab54b8574651c46a19c0f649017b152b8c7b9a6cfff3f536d970f5c2c7c925622ea486b68ba5a1611e323b06baa7b7aed72e2ef63dc811fed6699eefb14f3437045;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc51e0f3f9e6af9c0dd208a11387c06d04ce231f3e128468044d86852ab1c5dfa1743c3e45b2d7c306dd76d7a4209a49e090ff3fcb14ee1d70e7e772c046e22bef949004e43a06b17a453f9b733cce7c7cce314847fe275e18a078e5e41d3a8cde4a55cd89cb4d0ad54b1067b9670507da;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdbefb2fafdb538534b0180caad200269ee3ff5e270f9dbfc94ee2848823c5cb24633859d5ef11532f99f421f311877f7cd4518f0bb37105ea454eaa3285fd1eb5a982cdb2bdcd506d53f394c89ec8cdc4b3a7f7626e96b3f89be715e05962b31adf241639bb19cbb33ab67ed45e628be3;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbf4d8cf7640da3f882bcb6e6be15bae1b5e07b2768b5814b12512ec39154a2d30e11762a962a4f4518f4f1ca8abeba8e9d4f66b8f6b55ef36329a0a4f90a555eb76182b0d47b10fba5814108f863f5ee5e913d1ae18764a6fc6fb2ecfcf68aa2950ca7a1f6727faf20726485d3d693089;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h38450fb6a0824cbad924cbcee44c1923f0ef2e78ad90acd64ae7755c641a3afe49bd9172f9d2bb872d92837e61f51ce572d44e1c39317d8cf1fd7d01d3362da8d855e344a4443e66828b7cd45a17b03f84e2423285adf571fb390fd1ee4d8fd4a0c93f7fe5d32261583b4003ce1eaf2d3;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h156402db17cdbd7a302dad0356a109ef8e8bace964640a7cbc42adc8e195945fddc85e76212245afda97c33f7cbce38f91b3f9bd7657e640eb858e4ba0b7c5e2487b02211fe0e40149df688e034dd016ef05a24cedfa6114d8068e5f1949647f8efe12948dd3a869bbfe79302c25177b3;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h125ce68f90f3eae6297f4ea6aa5fb5ca330af84bf1a5c1afb2a4d1ec181670cd52242466670157558e8b53dee256695238fd80ee4177b4f0e4cf256a0f89dddb75650df19656e7d02bd9bfecdfa462d6886de9d9ffa2725d82fb65da53a91b3a1fa0d9e135d87efc67874ddf5e3b18ab9;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1cddc76be11b5ef027fab13724068590c88d397667985f0cd331e030b4f73442c5bc1b799e0d694c7b4002edb95060e337a2a25a3418549b7bb5180b3a0d8bd0189122920cb0d0c2af41ea3b707cfc059f5f90231132a814b356b2e9f09df36423396d935047b419b9e565ef537d17e5c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h73088277cbdc8fa5e501a160765c2499b97a3069fad01f2b267aeaf3628b6e8e753d23e4bff83fc72f01ddcad12b64c91c7bce69b48499e5433a51f1b18f8be5ca41212a8c5871582555b08a01a882dd5e226e3666214f77109c5d72434ab99f52a00fa1c9ce4c418c945c8457c0d0637;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfc15b07c197716092009b8be3c3f2b6e7b6b291cd718138fd37958a0c3447f325ec457c5588108dbfbff46804a3079d156a1234a08dae666d203d7f6d096660a8b3ba988236024bca5edd52ed0510dea010d47af68adf9f7bc198ee469049b0cb39678ae2588863e55f697eed5f7f9719;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7819700565829ea3f028034422837606c499a5b611acf2a0bd112f7e232dbc1b61c33cad479370948f440778fd1dfddf328f1b2fd002986d3285b99a3e66c2e40741fdae85a5c14d0d583b118aa9659b4193aafe808ea716e61bacbdc7bcf7a148aa729db01149b70d08ea91fbfe4000b;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hefdfa47fc7cd82d10b06adfde275adb53337431993495fbda28ce9001033c6eefe5e0c4f61ed73d63b5df899664c2cc7360dfdc5c3dea3c818b8538c9ac3b37c729ef015792d0e5ded7090e3a27bc3f0e78b55307a4b5a0ab55940ea9f4e4b8c5af8a6af541089d8f1ce1bf5f59803e79;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h147e3d9037e16676400cc3a25236c900e24f2750a9c2a5c3c54bdbe593d6159f365e1304d4eefb63f5caef8bd473390d056f8807035df0f141d4e231d9cf0127cd355fff880b26655f4c1bffaa27414ddf8aafad6ed3c4590b8a64ca16e8ae16d8585c706e90cc0eedde6e7126771157f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h48fa239ddca6d5a57d2406c3da34d2ac454bf132b1ec4d46ea0601150c469f0b6a74b309105b781829757e84f109ce507d02b17213492d88f31c1586ab3953b441756f0f00da50b67bcd030abdc832e6ec0a1a1ea7332b35998440365b5fcebc776007e529bcaf74566ea0053bb99496f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1e370369f757c78357c7868157fbdb2b078982b341831f45ca69060e2e90fa128b35713220aeeee9afc1da049349f5b61d8441803c18b18ac7e5c2e2d07ef78400514a0596cd9bb1a1ac93124c36a342110fd32eb3c8b265f436c283206a85af499aefd613783cec8f2479f2a17b1f20a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4ea7817f9bb67840641a5f0d682b039f61bdb217ba59558e614923649246ceafe1ff800c162ef538b5a406bc0ca87fe88ebbb9d0905c5cf2004caa21ae58c5b66f84a1701021ca30c9671a66c13fde6a64f8072cd476cd2948fb63379f48f54c51db89825ae19bafc61111890944175c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9eb072c1ff41ffd865174161616c0f31c302b2b05b5e13d41fc46757b4096828f563d3ac6d1bade4250ac5b6579f0defdb67c928aaeb8719437e5cdbb0b936170b9db8950417d2bb77744347fe6a9b72d0ee7e3757472c48a1f8bce65d0a4642371f28c26fb773c1dfc5db28519d7f30f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1f2ed445d4a6fde044086124deb99128ddb80db6094185686adae615d1cf266823ad6f9596e33e14041d3c70b119eb8736868bba27629962e7dfc8d0157d3b0c3d4167d80f1f6595c4dc306770fd5e67b5900ccf14bfe2d61f437e04f85b7341b6fec789510e1a0f43d83d7e8c8a8a45d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6800ffa39f53cf0d9fd2a7b413b7f1dbeb6fd833f0a688c2ce9b909106df5959ef6feabc48eeba96a02bcd3fe7e177619ab35a8527c2519dd1b5baf81f0b842791b65b195776e8e017dae689bfd128deb75b30b3acc8a85fcef9aa796917c1e61aaf8c936dde6b0304ea63f5157ca72de;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd1493cd15b11e264a5ad01f4a411511ce6d2bfb54798004e32b8e6f609b07624aeaa836d4b8cf3311b0899c9bcb5a7dabfdffb1f10337696a43a76f0059a36df8cc238515731ea4b2cf8b71e0088c495b7c75e60b9f71d6ad67beb5d83f3ee8424e323c47adcae641d9239cc176593e96;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8fcaae4f81f514374434e8b60f9ecb08eed5dd11120dfb7a1b4a442b25f398d4b38a0df8bedf4532fcd8711bf515f2dbdc9c97d9e648771054b31f86b5238cea6baba18f0e2767381ff3e80096276e1ed765dee7a9881cf282b79a59a964a14a34133cecb8436cc5d1629204b8160df65;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6cca2b3777b71426123f793430e71a64e23e1941972c03904c1b38a59efa0a7a0df95593629c4cab5432dc2e62a72242ace6fd0fc9ab48229af77062225cdad7af25b44878adf40e611a1014b6c01edad848d2d2caac6e8d77fd3c18ce4c146cf7801ab952ab5e74594fc9bd927e6ad78;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5c6a4a042a482b418fcace2df3b2412a4e7a36c9c8eb71acbe37d7c2eec07bbacc2c344b15ba3775dab389f244f84bd68c5b4f7001844a58be646ede97504c17c0de09902ed31db1fc424dd60a717ddcb743e2f36b5d4fe44256a9e61ec6709f50d0c2899c459415295776060342a1b13;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he0e792bfec969cb4f489d20fe442a39a2b98314f48971ba746a785fa5f6815be8ad8921ce953dc973f192703f944c965fc80191f3c6cf3fe3bd27ab05bf9e6b0f57d51024354c65a3ffc72c5989b133528c8894e86a412a008a702f23e91af605025e42a74559e274f88362f8baaa010e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h924c7bb6a3a2303a59878b0d161b54fa28f6b39193d46c5c55a05da4754c553d7d650bd209b0c0af05d5486410d88a252404e80514a984f72af14ec1b63f4dc91c77e3f0a1b4ec9f1ba4bccc0caf730b26ab9a9dab47914dc63ba7ac0e78ac41ed07af812b092200d7fde20dfa48797b4;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf346d728d5de29126f857580a2adec4cbec7e4c5cc0f1e93680a3d6e25f23f680ae8e4424a09ab95853ff0a4b0da9f2fb0c61bd41d428933d731a7037313cb68e0f2cb90d04927403feb4b409085dee0388fe337defb251ba8db116365d39f2529c8faa079de411a02079fe4bbce07f68;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he18ec42012fa96dcc4be4b4899a34e33c28555f7f6bde5d1f5d6e87c20e097a17924858c1b2f2bbe7b4f537f9e3d41ca455fc597d8537ea3a3c374a99836bd2ada6f05725b774ebacde4f37dc46a9be57a8656776906110ad59e2fdff85410d5b301b231c82777b969fb0dd1a0081f244;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7ca3aa71baa8459982e85b8c8c23eb04ff4dcbc20b645dba32853f888681159c789dfd21ba5625f03b29cd23c0ee03081660f1bc4df3256a651eefa4d67efb708b43d213f1f75ff6b1c66aa262b27d08ce3ba912ec751946fea31e709c48be0b1faf3a49b2572f5f8a9dfa04478140033;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8ad1298c63d1d1a109e6000f4a45bba7adedcb701e1ad57eaa16a6b54ac24b94ec5a6c4a264dd5aba6966bc8168d2c090445eb6b307b908683234309d194dbee5ff7f6db0db1c7009b3bd6df86673c23790ce19d30a95dc6b9f929059e4d5eed7c834449b3cd329a3774f2af0529f737f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8519207568c76c4f1d9639212e2227ef794f6fada6ee577e58e1064bc0d3eb9527c57a123d2746b5bdb736632f0a07b823bc498b97a0e0270dd92e5e777e43d4d97806da5b0df2b7a29ad9a3241cf9180276199ddd2f2e58f62cd37c33aeddfc2c95cb070d0b3c75f628d80cdecdba237;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbbc3ec10a0a69f4d5ecdbeeea297729063ac0f5a5b6444b6bc94cafc75f23e538ab848e6b1bdc0311781655defd8a3fd4729302d22553bed2fae1b915b3943ccc9ca7a28f9c81f11b2192fb44af6062aa1842692835adbc3015338525590e1f6782633a3e015d0f8fb59ad949073a0d83;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h47ed0723a8c55ef655bcb501bde78e80e0ad62b9abd23ee933fc60b51deb4f8b11e9ebe2809cb441c503e0088e3826b3a4e4c18ec0d40d8a0ded16ad01d20a32ef17a94e18334ad78b5c15ff4af78dba76df6ea830fe67c933683ecca9b21ed2e73c63c3a741036072bcbfa72cdacb6cd;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h630ca4f59250706a7f7d786de59ac7656f25e2bea558507066146d94f9f281ea62466dc9cb3c0b414a0279bd98efbf2fe75860c39ce1963cde726b8cb9685d67894447537f68f174e30772f9f27a026e1cba95d9c17fe12c80cae1c3a1023109a95e36af659eb12ef1b01d3d446f94071;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc9fff26ea555cec5f4030089ae9f1a56c56728bfef02f21040d497875f64a1dac8ee3cece696956c1e63f05aef90579b04d322fd6477f5c34d39c0308fa899894c608dee28d71b2c43bf0435db0be3623412795633dee5d3eed8a77aaf13a737dacb858853d52b8af5d45ba9212630919;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc487dcfec4df2a72ebc562f93412c66f73df0ef593b6bd1f099e2866b5b9f29f946dd06d8f17b012e0abd984c4992eb9f52bcc5cdc31247db1356d1926f90a6920d9bd7dc094b2c53a93b4296595c7468f56341d9a415ce33cbbd4671d0ae7eeb80ebb95d79a1c583269cabee04a4f2dd;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd67fcaebee7c0b7e2497941f511d6b52d0478df854bac7362fa601d251c6f623249b4da730198f759c3f4636becc1281d034f59d3649fbb7b50369816fb8c462a88202721820ba42cbce7a3df3cb46ec949a7e624dd9a5f5ee418d41655557da50f8581a32dea505d2204e2363e9d2af4;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h42ba4ba68ba0375a81ba7670c2daae0ae856e792eee4b73f710d5147f4fad0f24ea916e0ca328225441f065a02d6b204d32f02c7cb3a3b8174180420ef0f1ec15324961414b9cb182d06c3c0ffba764dd9afaa2414bfb48d0ae8517937bfb797ace761c5e3708ef84a293ebfa223c7e95;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h62f437fbf6a8f5adf09f5361bf63ad9573642655d9b570bb2a5f6526823c29636693e3f591a1213b92fea40d3dae006635fc17de705b0614a7bb40ddb00305a80314cde7b276bfbea4fdc9d46f5746ec74dd66f77449f513bc3bf242e1c1255c7d33ff0273c62bc5aaa71fef006c66187;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h94defbc5652c4c4b8c51e56912d58361d26c4676a421e7bccce0c8c058a5a2ed1f9965c45fcd7589dc9122870dcfb1a945c5f79dde690cfeb9ea397fa6ddfc0cf5526ac3773eec4d0a839a6f2dc319952188b3c9e50019ff83e393479f6fa29ab2462da176c81884416c2a018359ac1ae;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h72c1f1b56076274ded721642ea7baebf4dbee388a98cabbd75ac27d2fe545d89bc6cc3979d9e43e4c59deddf6bf0334202c88b275ecd43567e81a62828fe024fbe4a4a6d15939fa7d608f71204bc587c9c8b95421795a582e78527493366d130fe04615954ffba4c412db648f41949098;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc95c09231133c8cba5f64748eba1dbed52f84e0bcdf42816fbdffd6dc03e8609128fa85af40d9f328ec80a10129a63757cd6cae6684f9e26d48883e012d4d07b0c77bd1f1378f05928c10413e640e8abbb230065d2058baa5e2030a763079973559d1997cd0e8674a0fc18e2a53765d85;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hee2111c396478c1c964b8e5193e901dbff1db3ff2f9db0e652ab94fadafd478a6de8b7b4e5099e09818c3febbf6a433fd2eaf4d2dc42eea0734ee9edbd9b5345126af14d3e98b43bca19370f64a65212c4d4c753b5c5d6ccf91e85f6569970cad9123f8999cc03503233b7347b15de242;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7634f048d68b9fbf565e27d0f935498baad6a89fff8f379a3bfad42ccc54366bcc664aaf07a031dbce12d6f36b1f7ed8865ef093d841d16fad80341a49f83b7cd1fd459d32eb968c65ceed30325a21d55cb51ee83f777a1d27e2a7e8c509bfd9d78bcbd83505cb77b18c4e7d489f4844;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h54d25395fc6d683e31516827d1eb0186a9f4b008b0b86ca19ae1abd5155a38d22b035332d23f9c1a11c12959daab5e3cd5095fe3e7940e9890e91cedd4eafb74de699e947bdeeed3b21748bbe9fbbe6a9e67b008cadd4133121dba2c19d66a8f7f3abff1a208895c52af0d592cfd07d79;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h902d329a76f23d69c9076e2b33727070b065660ba9f51e01d49fe81b2d7911fde01375d911ab613902df717f9bf955bef82bebc0031e01564aeb64e985761d5cf2746b391ba5d9a44911d153b6e7270d7c2d1ff80faac2f0f5b4fb6511a20c3aee1b5d99462006741cc88538dcdbf4001;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h98839542963678c5f22c76c62aa104e07be0eaf6f4ca7de3e7a717355534d0f73f65a854fa7876473036f831717fab7278b4b081a22ba848eda1641762f32a762cb9428d8be40832b3a0ad037f207bf90a0c2ae73b592b71aa292fbb80e4244d8f18d18b9830da1764b384a3e1b9cce98;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h447fe8b70bfb812f8e3c066fd4ed971cb352b9dc61c50e9b4e588e734105feaad38c547fee15725aa15aec613b390f42c5e8cdd312419d556bcc4a0460056cde9f801be4ce559972eacb0a3311629782e3db56da0be53149bd0c903ae42a559c38aa48745c685458be291dc63cb3fa39c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3ca8aeee5412865c038fc70bc17041db01014478309d9cd627733e7a8a2fa1a492bc872e113ab55cc7e936e97ed828122215bf0e0f86466ebfc6997ec294f11de5a9e2247b97fcce0f1b3e0337523495b29bfdea5d842a48e181e1227f92cb42d4865fe024f3dc6d95633b876e97948fa;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3c91c8866b73ee7bf518dc220e9014072e79fb49675e484fadb0c8f87111206046d5a20f6288cabdc917c27ec702f0b659ac0ef32c6b751e324d62f84f5a2562f27f86faf044ca543c3a52881b117d37e57bd024ec08ed2157d1b5c9c0e7583730c8ec32c50cfe23c3071891d99908120;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hddd95385a1dfac28194fc8662ea05a0d7426f22f5adb4515482763a8ad527b5cf5942388853a1121b539cfaf24f2b78a07942cb92937bb7447b3e67e601e682cadc174a81a5ae835809cd77ee810e6d44fc83cb84967d656b805e6bdc25722afa9c29bb707f3ab6fad1e9769e9662a591;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h30e8746c008eaf490fdb15bed7a519f627d03a870c13d450fb6cf01ee43d247ddaab0122bd307aef7da4cecb85f47edc1bc68684a0111cd782b405332d9a994ace15b48e33f736095106a2b9afeb6d63eaaf197eca73b1cc59071a70a0f4c36439eca9f2b31c8480500cd4db3e60a0ab3;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd7933b95645c17247d516f87b4b393008ebf5a63513d8a0b883a99a522b2647f12c4c1d8e5a3ed97400f3c00a0c7b3853bfa8afbd049be96d6fbe068972aab6f360676e9be7eaf7522630b051b53a4c08e3b0e2a22f9ffba4e7b317f1ba33473d105b85a1e3c87fbf9c60e9e761fa0689;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hca590d7bace035b3e9e257b5fc8c92d0e074ee1e2b28e00717181bd8b9a0bd8d10a676b5ac4c502abd11b7cd68dc479e431db59a529e502c6c05e44302e7a804cdc9072589a7182ffc5e14e389cf1ac8287f9c0d10bf7f896efd6d2a1b5b4aedd0a5e6d38030df5543e03689f63165916;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h253b6bac93d8212262dbaa0bfeff8190388a71de8799ca595eb170ec8f21af660b52dda7f7773fe80ca74847fc338ac53d2aa1e27cf4c1f70b92d6f2a2dac2338338e62f79237a96454d5a9d2403b36512f51e34583d5f2b584f88d9bb25637758299bedb20c77ac0c5055521d00d814e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hafb251b0322aae042861d8f7367018679c1b82b42ce0423c71ef5114e407ef3dbb915357763548558062e771b957849b16d66682658a9ecf073a37dced2b00390ef8d5a7c17be5ba1d4ac517ed302edcc6975b9937b86bd51e815d1b0c979ec42131ee2e40a4d7b552f8fecb5e7b327c8;
        #1
        $finish();
    end
endmodule
