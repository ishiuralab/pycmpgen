module testbench();
    reg [13:0] src0;
    reg [13:0] src1;
    reg [13:0] src2;
    reg [13:0] src3;
    reg [13:0] src4;
    reg [13:0] src5;
    reg [13:0] src6;
    reg [13:0] src7;
    reg [13:0] src8;
    reg [13:0] src9;
    reg [13:0] src10;
    reg [13:0] src11;
    reg [13:0] src12;
    reg [13:0] src13;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [17:0] srcsum;
    wire [17:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12] + src12[13])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13])<<13);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8660af667d84bafae09be3481ee7be90f2614662f473f37c4;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h317b078294a342e6bcee42e44cb2d0d0dd5d715b78c588222;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdc838cf4e98fe6b18133a8acf76249fd67215e8c63ae4d513;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hade78bb105be488c3c4621c68e5f5efd9799cb8132ccbcf67;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf8e6c2085456353a9144a701eb077499eb9437dd3409698db;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h46236bef030274c124511ac4d3e8c67ea7a944671767b2c8d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb7a1460ef51e72b855d7195f88473fa76af25cab456372839;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha12728f371f89b943015933058384781dc65de183df84bd75;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1ba561770e1a4bfc0b2f7862ae6924afff774ccf9f22a236e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hef29a4a2a4ad31bd99f40375bd85f3bac5801206c2d688adf;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbfe718eed1a6b329e50b50fc3fd1b025ff7f12be3f225cb6c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'heb0252845b8fc556a0d594465aff49322fb51c4673907c78e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h748e1779c33ead6e5c865241e019b29296076d1e817680b4f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbe1c546a11e9a33d56dc7e0b083738e52fa697456a057490f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h13c0c909d277708d167d40d091b116268414ac298a31b5b38;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd529c5e84ab3e49659e796d94907f701afffdebbee0a4621f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc03329b4d24bc9d74438c67f0d02cffdbd281f105b58c290e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h454d44228da55cbaeb3acd937c393769a887f503a0b01f4ad;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbfbdf83803e280c93f721e24dfeb9d9c82da1f7f116400fa4;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfa719f969a496907a02af2025ce9fd027a43eb65023667b03;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8d1bbd00e5c02092b7e89510165bebb44d7d08e195fbd4795;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4e28217df72f65430e9441199ce03b44684f8ac197fb807be;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hafe684c48ef72a7b1b7bfab5744034b71645793ab138c46c4;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2dac7a99058cab95d675c2e941ca6ac6df48c35a1b0019342;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h71833821ad752817846a98609b238cf56c8796833898d59a3;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he4d009312c1e0106dc5f5b938a2698d3ce20350f029ec6b99;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he6de172e0677616b9191addb9329e25012783d983d861609b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfb4dd7a103506f09fad25f6bf00e92f56778118033052370f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha623e82330f6d4821389a29cd2430b7f4d9113fee3a86bcf9;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1e58ca4d3ec35619fc745822ae39818030ba3648187bedb4f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5f7940261cb459f545f7fe04f8bd9734a10735d69d2fe92c4;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h533060719b70758fafb44f96663e4721d4555566e38059d19;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2ff3402d7c8bc3e3e31094ab7e8cb469de6284f34da8a1e3d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4f8099d02bf6337005d4f5f2d31befda4e9f1d01e3af0a49;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcb123ed1864e81bea5a823eee0cea8b47b3e1d278c33c3b92;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h42e82f160019020a5f9c6d720e45be70b7ce9b8cdd27c87eb;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hba7b17e357283e46ffa8fb24c8b28e053cdb005604490063f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb3ecb79b578df070ca6cdcff0b7a127ae847b31372ad2cf2f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hea93b432d96966b37323dadecc376b9d680a436020c1b22a7;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h918d9a3f22f49dee259d98ef049b1e506bb2cace9417a4084;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'haf5378b3bf575fd306d6de4082986529b1f67b47b5d2f2f2d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc914f0e1556d603acff5773ee3d932e3bd08445edc76877f1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h420e29b7592ead32a143c0032a116650ba61309378776c91b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h59e34b7e624e833cea59e954f7a77a5825090e968b0c1f7dc;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h90ca96b971718c359d4af55ec773e5963b6d48036efe421a5;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbc3cbd0dd8e2a9e3a374edf0aac4643c830c7eef8ca3e5ac9;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h818508334e8c365dec399cc075470cb464d3d8572d5d3e2b8;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6c59149c6c7f71854592976c79ec7c6480b0d6e61f6d584f4;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h89e3ba435a9bdc79cd9b75744a3f2a509b038291e7c616ea3;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9755fcf4e3e705e426f170937b8251caabb1eeccc1ac9be92;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h588796b384a799529b268f26d2eb8b541e6e33b2fbee61f1c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd1a7439c6f37f6b3fd513203564fdcc89e0f72de1140f1436;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha11a85f37b1ba970eea3596b134a687b9cd2144e23e697d56;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbe022a4f196c3c2aa51f30f0f4fdddf29620e19ef910b722;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7d17ba8e6bcbeea9380e99a819287a768f30a872d45f010f9;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8cb94bc51c84790695e532ccd0d18b2eb5743c955dc1d9cc8;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd9082710b9c8f189d9449b8f123bceecbe83750081d742dc2;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc8e0358507827491149d380f884b0d2626990c6fe20dc3edb;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdf4d1eba04b34ca44f122d4bd2d0dd5f1e85381a4b16c26eb;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7a6290f9dc81c97da8b7a903f717710574317e82a7d2eceeb;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h15fd77cf1206f2219a395805a4b23ead721aad789f3c03404;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h78b819db1e22540869c5da4a825ac902861749c687fc31cd7;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb28094ce760a795e22140285f1fcf6941a9fb4fc3b9f46580;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h19101d9e35efd56120d0be11fdb2faa3f97fb8dfdf4968dde;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h29cb35060eff266b5176f0805998697e8d37bcf57f10ac2ef;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4846457bd13d15ff66a66fbbe9c14d3203e12a32069775cdb;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3470ea4cfce20698bb60c5ee2466978081ec6b1a0d9727eef;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h59f32e06f3b58d118e275f5781392099f1a47d714c09c9070;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h252dd4068cc30164e7e4f55eeb8da4068efc963ed0da0ecf9;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha7163a3910c3733d7bf008e588a5e9b8005e9b24640345adb;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h11ea3fc0995dff2897e8642dab980e9f53e0572277ac260a5;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha576a2d3f09089d081d2e486fc8ffc5c4b2e21b496d62d37c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8bf519bfc5a7b94a902d04e0d16542098038559eebd1c6ef5;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc7545b04a54af1c2af9dde9e44eb8fc39debdde60f0f98e63;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4563d15871b5818f7165bec82a459d6b5517e17220b5e1c50;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha3f201198810b9af5343a03dfa5c0c6c20e9d1912dd61b8e3;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h57e6be58643a313892e4b73da6523d74e0211577edb69f095;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h685213b6693246c8fea440665d24178d601d6ee23b5372474;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hafd12d25c8c23881fc6fe7a16c08c0c3aeaefb30358891665;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3305f77769e52a9783fc6f74dbf4ba53b9c5d93cde4cfa0bc;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9b5bf94bc240fedee93815459f95003f8fb6381dd82a10a45;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h244f610138e968775548535144addfad39b586e553bbf6700;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9b4eeba10a91aeb0bd3c4d5271b332aa51adf24b828bd19c7;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h77d94028ef07c7ad86b88e1c7eafecd4be9d4296094e77ce1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfc0b5f6fea1e7621345853d8ae1960325426dab817a5a0fb9;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he4c5d3563affd1a5af0f28ade31d7b176da9b7b1f34b08155;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5f29d7bdefa4aeb54d089d94bfef260937c75357d3c5a6c82;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1f586decab5e7f311e1aac9d5403db8c6c033e4f2a18b826d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd732ebd9e7c38aa0a355c76d5dcadb3c6eb5e8c948090f7c8;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdb670a7330d94506eed7bc36edb5427123771cf408f24d0d0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1d1a957090cdc670bc6ce3ab1b65fdacd6dc24b1f1d36d5eb;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb0c05020d6f3bfa8f93bb6d5e22e025f9849ac6ed10588022;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he37e51c7167b7aaf088e5be9f24b64212f511bd130767cb36;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3f793a46d79022d8c71cb9938c16c8ca4c4d88ef92a12660f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h16acf33a05c8f8a33c7f99366ebaab2c1431151d51b020656;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7f4c9a13a41ff7cd81cc3791c00b51144a971b6ab06801ea5;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdcb51a09ff6ba1801b14917e18e3b7a13115deff9f0aa9fa5;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h89e2421aa11e6430a1f6cc06c9d2ddf8defe9986fdcd5c505;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc1ee72aa0900a989b10136e9bed5129e39d05d80a2056ed5c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he5d14baac43589ea74e2eb174a809dbf71f64229690334a1c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfdaec1612ea7140985414dc9cd5ab92b22f3b8c33e39ceb8f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha012d3c21e3330323873547cbf1c67d8ef92b1aa1d254e928;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6f207a35b24e2ce6acbe0302377693fdb3c68d3039cdb6847;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hed05ad2d356467186fc24c979877ea899b9cc1aaee40f74e3;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc4a315a8167a399a355c72663b8feae45c4ec3e148e8d550c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1a1e9650792c7e3d0a680536743eb737c26d05279593aa414;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8da6dc07033ab8e2f74cebab40ec7b415204a30230305fd9e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9ad7ca887db4b29026aaa0f1760a3607a3f49d009aaee44c1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h12bcfd78631979001182a9f5a2aac18037260fc1a924d817c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd938e140769da93fd4adc5a0ea46512dd0667e1d895120109;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8a82f223f68341ec332a484a8b41883e1285e96ea8f384dfb;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h85938ca6876fa340eae9f15514e9fabb98084e6faa9c6566f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h42e2c9afef187e80ecfd351b5f2dc7bbaf6d936ce08005cde;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7e3ba8f4176146c02e084d13b7127e2de259f80f48f49192a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbc81f909d608e3d5050bc0829c99afbb7824071dfc28ac515;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha703b64cc4fc8427e7e475c2b1afdb202dbe9357c2dacbf34;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha202157de9eed8cfff02b4346c92e5fc08df059fd31ad1e26;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf0010fbc1a3f29c299266d72379e3facf9b00906c1fcf43e4;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h401fb600e64e5d80833b8d8c8019d5dd9eec9d478d0d59564;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd6cf5f2fbae6faacecfd8cc2fc86fe11cbf0d8729e99f8ba1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hde26f1fadb0bf19960bef88f118e565ca40912ee6264baa32;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc0f2d7014d736093e95599c14b13dfe1483397e0f1c3ed43c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h28af47daa925d877c290c64501b71012f7a0fadfb790c69cd;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha47d162cb9df5d78f67c12fbdedfcd0ac5022c90d74dbde3a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h503979d60e44de4609882940358bbc12d4df9dab14396f980;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h928100a1ef7c141fce4527bc9b201b9416dbb3bf35140962a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'heb0f5febd53ed0981e0fba289ff45f8f5d053ea46b416c18e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdafd6bec7cb57801203ba964ee78bde2fb987d23cd49ead00;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbbb120b34d43d9814d66e8188148f06c2fecab15bb00a07b2;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4a4b20d6ceac44f4bb00e380edb523f4c2337ef1ac394244f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4ce019921ddef6854764fb1dcfcc32be9d85dcd7fb989c107;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2044136a9c01df2c76b8aeb057cc3508ead243fe841b077a5;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb1fa56b36bcb9b02e5f33d6eb787e4a8d420e76b0bb7181ef;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'haf4a577841f98b143cc6dd27e39566d87224dd3f67f5e63f5;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hea57afd710ed4b1ae28fa41679a53f0d6972de4bb1cde76c9;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h59141cb9e19a10135510dc3ed301a6acedc122ea9b94a3ba0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3eaaa6a280b58abb7688e82899e44146e2d17086c86c57afc;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hab690a99e01a8e16ccf3e6aaafa8320a9b28d9716a07976ef;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hade65ee2ef4a88ec07def0809fda9fc2f42f1ba615d31c697;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7ab672e7414ea1362db3c0f45314e71ded01845d31ac491af;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h39ee0c9ff8905d575af2e35c4c56945c72dc3e630466d8460;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd1151b2b80701f52764f1f01c0ab24e0749f5af5a3c252ecd;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4d52372f1e509d458a02a9788148abc0efbeaf717277ace4e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h633d8d5cc7eb62a53341bbcec2056309741a662b79e1c48e9;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha0dcd2aba458352ae526c3aaa6f4c1938399b6ee30235bb6a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd589b6e75c23009c29f14e1502184b8620b644e764efd2b3c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h41fdc93b42921b0d8b06a076c1eac4f12fbf284c585cf6df8;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd6297b62a5c6e707cccddbad0bd5c97e637bdff8e374fa367;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf005df8dc50a64050377c9281bbdb74879dc1ef761b0ed35c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd450d6b698f085572e8c156217d8979c0ee99d8788833492e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3571f52cfaf534dd308c916593128319aadcc20257de06323;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he9ac34f284132d59df4a10f24ecd44492b594858ef71830b4;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h304382afd581a32ff2ae93453b76e4aea24310590b5a5abc1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8ac4c9d1cdf6b5bbddd4f5375917196966dd34a39882a15ed;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h142a43d609dd53938ac2a0558b362219f75cf4acfc538b18b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5903e7d90a15fe704001b46f6170af582f60e67f04464295b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'haaf730ac1c520e346c18e839f8aaade927521c1cad9d5d72a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h367c88975a268df05d877d454265d821d63a46847081b76d3;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha0add9c03e10274c91b1a311c46eee6c981d9ee7ab5d65cde;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h134ea80f95b803b5d222bf953f5f32c6334bedf33a1edde24;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h35668238b171129813ec29746bf0d0406d4a83f4dc7ffd1a9;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfcf9fd7fc1c094963d0c28d2a507f41ed2237d70e345833f5;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h41f5518de9d8f2592d0197c516fa684353ae86f3f250d1710;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfc7af2fb02599d37236c50f086f0306d36ae0922ab4b33fa7;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9a2aac32926fffa53097ebca3675dc18222f2ee73114106c4;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb3a9eff80f6742660ffef5e7084b6ff7ba593a0d5e387764d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h67524afb4b3270bee2cc2ca74c75fe8b9d8e123e2b7a2af74;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfbcf74826c9137e2243cec8308d688007d9a2f96558686d58;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5dc42bab0384cb629462af855abb7fae01916dba0b1e77cf1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he02aea6cc14ab0a64f7c1d78ced2af815fa90ac6a6718eb9b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha334be12c40b27f31d1aa5d64286668633b2a7bf9652c26e9;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hae0c88ec4b6afc85a31fbf272f3e4f4f55fabfed17cd80a89;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h890be9acf0bbff2abcbd38c8264b7d14c2cc1283d44c0a09a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6f401008ea1df77f2b83b8d0dabd64014de40334af358331f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h861a3eabdb2610e248b04dfe65fe10634a4c278779c950832;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h65dbdbe88c45b8dc1544e10137a21b0157dcb62451b2d8457;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9df55bfaf2c362d37d7cd6fc5c9ca497358e41cb5c5ef1491;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h19e2de0a568e8aba808dd83f0833b103a1049a5dad50bc81b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc32cb3275c973a7e5dca12b0b92ced9a826e0fbe57f478ccb;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h11e830727a815d440f81688f4e2d90070872fb25885a87990;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3dd58132be3fffb0ac2a0ac4103089b344a121df44d78bedb;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3839ade76ccf601ee8863b119c27e89f2e28201e0f64de657;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h63c0eeeecd81347be4a12edf57d2f174d06fd2ba19d013a8e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha7f8958c111825b7f5e627d6f4c19768eb00a046b232d3b50;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h830b9071ee3df559e13ef470b14c9be5edc22384225776f16;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h92619a0d9f96026e65a2c651ef32c140718c54d083420973f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7aeadb849dc9c852c726b9219464c14171ee902bbd8af4ee6;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h512847240c34c1b15c4628e7fcfbf38b5cf1ce2b3d42f9d06;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9626ff2c2bfdb31ae305df83aba2f600915198926a2cd9a75;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5d7e5df6ac6eedce6adbb72c61d88aa78b9cc9fd59733ec52;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h96c702f129f55d99102226023be2d11473217df40d7d39833;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h113137ea66736d61eb7cd80e4f4ad5142788dbce1cebb8881;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd3229be0a6547c3146b3ae35ff84de6fb359e392c093e08e4;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hda4021e88b853d1748ab3a0e5580140fef70755ec6282c083;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6708e8c2b100719671f6a3683e2e0631f7dee32cf317a7b9e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf7be7a698e15b419f4e26ebd9c2d2e8450578007c97909ae6;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8762e8d7142a5e49c09c132b4008bc51177822afdfd5bc7c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc127c73ccc252fcd1ada19cc2a14384f19518c042c747e09b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h18e9622e157f231169ee315aec8b5d272af8839f91120fb0d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha1b615c31f9ea95f96d79726f6568760ab526f3db5176f5f1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h911ad47365d72f3b292960e81146ce451708d7b4f26abb409;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2b798049214bb98a663d4fa17cb440d715ea837cf3e47eec0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h49f2c00d7e38b39947629fcf5e11864103fa6eb8467df78f5;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdfb67090fe1a28b5e0bddb1de53990f8d8ea620ab762bc57c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf9ae04e806fdc920ea9a9a3e9711872b3314d6b4bb73c0aa8;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcaaa82bea7bc2b19fbcc783dd8dc1fb249af19f434384c03c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h794b214fce93a60ae7ba01612cfcf3966adf5607efa53740d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcc1c339afbcb30fa4933d332c13a74346d53a39db9a626e99;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8e3c990aae600f790fb98afbd09e887e2aa859aefc6ce9994;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc9a6e4a696664ec8c97c16c38253d0e23abf33cb7fd975ec9;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha3935e5116bf3cda3522f5a7069f06c90dab102cd9dbca9ab;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hff093048fd13be6239707f89395a779a7ba84dc6b3a134ce6;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdffbfdb0ee82a53060071dcbc74a6bd67d5d61b6debfc8a6;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf0b34aeab1ebb90ed56205a90b68b287342d7f1d48d492a25;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha55d7ad68b4e399506843871dfde7f97852e4133b1a9c4f6c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h63c60cb215fe06700071214f382f561a8f652800670c316c8;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc1f29e42665affe6858009f3ca7b3ca112f168f1fce85370e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h391f7f7524f223bc4c8822005969c1e84bf0ca8984b007ba3;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7f3c933caaeb2897da396387850c6e54ed5b4c32b01a1533;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha620dcc61490c41d91bb93f4c9ce1477ac48e1442dba88bb;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha42de48e07e975b812122c70b33a52e2961f909c1a301592d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h56fe7834207668ed4f26efa58677d2329f942a17e8e30e9b6;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdc9b2157f7aad49d64bf6a628a91e494e3490d7a775232220;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9bb8bc85dbdf0d82103ba5d24643a6cc196007da35bdf4bd3;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha667a235e8170b3f76ef6bcdf7f054f98ec7e34d21fa71666;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h871b02ded24ceb72e8ad5c4e9f40c52dc94cd209f824ca14f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9f28f132cb4ada12c937ec892a548a3c0575eac2e41731e3b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb7db396a3165940081695c2d81b644014f194d85313d892a2;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbb258dbf9d898cc25f63bf472ae738c9fee35da762cdeeedf;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he836af294571c1276aeddae157a5373d96b3ba007d1efbf74;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc56605fc092f1312fd15c8a79603ff96abc42c1090d002d84;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8374614d16825e0d5bf12fb4b62c6f2784536fb9a93761282;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he0aff205e719316a511626ae32a118c898cfeeb7bf76f5a9a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3ca9c55c912bcf7bb58bf236e80d5ab1af7d18500ba327356;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h282dbdbe1184634a8444a159090e845e52cbb51f36390d4e3;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h856d3a8a99920adba023f20e4fedad90dbad0173fefc9c999;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb65fba0d30336ecc6dffee5c1f219d3ceebd1abeace0e769a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcb062c9e1c649a9a352ef3c3febc5833173a1dd0e9d365223;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1a9655428a97fb6ad043d351455d6dfa9053d99806e784cd6;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha1cee11c47bdd88f26ea43c52c847eb44e2569f6e157599a5;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h77fd92d642d8f700a28b91c4ef1cb24db3f0f2a4fd1912e21;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h576816fac26a1ba14ff8876b014a2becf48a5867aad6df310;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h246a1876b064bb8c59d97e1b7ecad854fcf2f73bc7a451712;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h86a8203147be64e71c217929bcf0658b3a44ab66e2a800b00;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h50023a3069d38c0c83753ab154659513586e5e5542b549dba;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8d999a5e09ca3207758fff41c17c3786e74205a96a2bfb063;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h75c7c2680c6bd23184becc2bbd2d6f131c70ee4f8589b207e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h32f67d1c9758a71c0581542c845d833977142785dc917ec92;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd301f60edd643c4aea8b8687a50f0dee3953d825171130787;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3607d3ebe4e601260fce95c5203ea78215eb99b017e18a790;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4f1aa38a47da35796e3da329a6b3694db684e951b38a8f537;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h543023be31591d59c63bbd0da691f3649340b6d9ee4d75990;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h215612c1748336f707a8907fbddd4ed11960e593c4c05ef18;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4945adb91e5c6db7e961457e1438504506827747c7a25330;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h47dbeef39d7fd05343d2814ab8f95054edd492d06ca9562d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hde349797f1cd3a0d1d1cb0a1d2746b92c6760085b3745ec79;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbb883166dbdaa4a31deef44fe47822d19095cc0a6243602e4;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h42d8512183cf71e8739527b880cde36dca9722535b6745e46;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd02ded3ca8d3a064df09941b620aa4b686c0f2ea838d77a74;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h413a365d39622bc8d60859100910c99a1ccf283f41891a118;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h22a318487f701bc288204ff09beec98f45bda2926e532664a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc4c813789834c8e99380c13d580a6788dbee774013f736649;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf515711307e9d6381e02703837d204b13c8eb4020f8679f23;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h48c132de2800c5373b112881c07bd30ba507646c39e16945e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdb24f37e29b240c204b446fc5149643ed4730fccf432b2860;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdb42aed409092af50a36361d79f2aa1b51d5d92f9cabe34b1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8986e544e4794148dee9b9bc9d0667fc9c66a96f0cc80f049;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h92fc7428f492d87c872ee9a3c4a5bd7f708305c6f4cf468a0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd18cbbfded9790c58c4b6fa4b8dc6d9f9cecd657f6d8c9ccf;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hda36a0c24067057a9ab539bb9de2bbe0252d1d83e3f306d45;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'habc2cf4a1122c2f322145e50ef19cdf9396c5b729b82c71;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbcce325febed4f8182576e2255e251a6c6c04207461282904;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdd38b4c65d21ab58aa4f7cf52d971e40f992b091261c2d9d8;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hea0a2df6379466b01194bfee9c4203c69275e38e7f5a865b1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he200fbb1cd8c9d14ec85ca0b82c77048d46e7375a371f1d14;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h66378ab6a231888d3c4b777841dab7f18b740a07f7d5eac0a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7b706eeab0c60582d507ce94a81298fe7fb4fbdb32926500d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h22ad5630990062201c933a3aee31a66f192f0535fee2a28c7;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbe0e810914f461e820d674b4cae634b00d95503540b8f4710;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'heb715f7def60f9b3ca9edc780bb01946662618adef12dd61d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h92a27fca621576d12d468723ffff248c9c8069aea1de8ca8;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h60c8b18c87f20329e67f603966761593d2e6e681a20a73c9a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd194751bf3a892690ecf852c11ebe77f08117628860e77471;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h80d1171391e5cfe0c626b1a18b2c091924eade5679aba0ce2;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'haa17c39fa31fcc96566f49728af520a1aa39be454c1e7c0e1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h94ec5b212bd577babd3be3f8452cca501d2e97053447b25d6;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hadee70e754458d88d69e34c113936144e43fb8d9e751ac84d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd9c885295a94276c2ea96d1cb2ec2609942dd45812afb24aa;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h182a8c15e3543f2cc88d5448c81314dfe4e7bf0f55eb5a6ed;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5f3d0bac2ef6b9724a2e9717fdbe7c5792d50656c72750253;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h606ef720bd9f04c1f3b0c88a10626229481ea71614ff98cf1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbc4ffd6c2bb93da190ab05702ba83dbdd7d210bddb41bc711;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4b2f2049adee8246605074cfcf93a0703c71ed6299c80e2cd;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1dbb85e4ecf2fe3390a6394ff25b857676362ad814dd3def2;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf6dd33a443fe681c982a87f5c573038f59451746d112d091f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h26263b758a8f5c017e7a606372cc4909cc8e7c619fb68b59b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1ee3db4549b94b25825ff49483814be27bb8e43044e76f9ba;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdd686e4931f1c2f282ce3b44e16bfccb10afc77009053efac;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfb0844099437e973dc80aafd17f7b396a13f18754493abe99;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc74235e5db776973ed766fd2262d6c8ad959340365be13d59;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb98469eb73a4b67b916039d980bea2639a1c7303883aaa437;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h902fb9a94c2e03e717b44dd66a7c4c2817e010082828acf16;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9f5a26037eeedfb2ba62c9847870cb2ed30018c4ca3c97445;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfe6211347a90e03cd8257ab89622daad163779c2785ee3573;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he7f7c527aafd6988c6dab933999d73aebfd99fcf54a7bcea4;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3851ccca11be221abd619351133181d557647c43e71d82d13;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hef1ec73e322fa85f5a7467c4f5f3b69c4c9af71ef01c60526;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h14d943c12882829a507d2a2450185e6e29f927fae089c6264;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h540b71c6fecffa5ab743260d1bf1914549bbd42ae46b51340;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he565b62b1a1ccda9be2d2b7abc2d22fa3533d6a60e8d0566f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h695f9a52668fd4f245906bbc0c3dc1518fd6ee20a969fda2a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf099947955efd4740c1b7f7ce2aad27504d3c6d0a0c46db37;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd8cf26184c83b7110ee4f52a0f3a724a04ec1c2e31de63477;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8f7271edddd159d1db9dd88e644e48bd8dd0167a1f9d3245a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf90b008981335870fe277959c3f885e494ee81c30d35d105d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1eb10e28bd4899468280bd814b156f4c5ea8808e2071d1a8c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h218cde3020481096dcf43343f0dace41fdc51e7635876e2e8;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hade5644bfed205175aa5ad9a22e8f2db000cab9712fb3f262;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h90d441d239c6eefb351127c356aa184113635e6aa8efe4e80;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h21733d09fd8532b18e9d34c737fd0da7633e72bdcff7023b0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8b90c9fa86fcdb53f3f95643988dac31475575637856b00c5;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hba384a39eefefee1d9178c1b5880cf59957045cee1055b5df;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha2280dc3502c26a356ca9048c51adf53dac02f4a3280fc39a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcbd72a175ca7d2e449ef425fca4e10f6c3c6fc4ec46614801;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc7290d1c47ba82d9568d31f50aa2a620e22ab744974e520ad;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf402848f3fb18efbd32f8f7cd98bca703d61afa876d9c0f4d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h623a5b1c90f298ecbbd3bb5624a0bff3d5f3339ff8ef1bd76;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc557afa55efd8c7aa3e0808eeb3f9fdb7c0b387aa970ccae0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h577efc7749a86d942eadb003a964d1a0b9c70bf5883e2eb21;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc03de457507c1204fe3f41b7ae2e9d575d4831ec9fe81cd99;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6a9aed8209e530e131370aed4dfc506aa9a893beb89945308;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfef7e7cb5fffa585d2873deea7646d79a1b249247c07407e2;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h348dbb84a5eaaee30dec70e9def49e4394550c67670800504;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h93ff3d027ce2bc3f0650f7ec2d3918122314742ae657b6718;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc7f9cb2ae16937b8fbfc63d67d48edc5a44bacc2e60008edf;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc815abbbae6387ed0ce3877d01474d47e7f4639f98fdb5b3f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h191c2891a05a669a39c49ef74fe73af1bbd740892f06efd23;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h30b7b1c9224f4afccf97417ed198b00b63d92356e64387bce;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb0b51299eda0330074b7597891cf25a8f9b68f4451bbbe8f3;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf616c70fc817a7e5fbd996ce7b25e15b5b2c0e6febb035776;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h10607b44ef61f02ab912b08f844ac726cac8c2fb13e412df9;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcc2da5aa3e296bcbfd266c76705ecaed60adf83047a7f195a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h46873dd5449dd9a6838a697d8e338fd4395f670f3547b6741;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h356bcdc09bb41d81d2b6716283ef7fd3903b4fa42bd28a2a4;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h284e3428c709ec37f5878e050888996fc791beffda691de4;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hccbd8bff1510d1475dfdc182355abeada4209a320c6de997a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7b17e0405b9d912bb48e11953137e266bc713c2f947023b20;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4e1561577ee32c6efe1de6b55ece8d16902bcc2a56c95077a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha6abb4542399c69bfa1d0f23e674ac9a30b4136ee32039fb9;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'heb192e6bb722d649e610adaadf9e4cf38829c018126c32687;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4a595e294ac30ff36736cbc6a8e55be8db5642507dc6e28c2;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hea3339629b5ea8f2ec69c86dfb449947099663b2ac66b92ba;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8321c5c1c40a21d410709df0726bc2ebf07ec2ae7e8b1634a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2e2ca8fb3faaaba1574a81b4582913692f27311bf311d564;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2bce6d5c5b3949274619c118e4b9afab303f34955f40163cd;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcecd12c9866ce255e452460aa9db66967183e62338ddfecb;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h31b47226e2b06111320256871b100ea48f89c2f163194114f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8f1bd60b9495a0e84b52d009ff4bdeeef0178ea4b765d0d3a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he33f218112e825d928b0fff65342cd56e5c05b418a8828497;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'heef91ed33e0b417de20739b479c03f452e15880b4be38e837;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb58e6d1227b54b46dbc08fda555b21a308ec58815a8873b94;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5f8acb6eef1d72abc295d2e76759f443f46c0646e8f36b926;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h14302a6e7e2bc1137769b419057691bb209d6f409283b035a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc33261dce06c5405a3b067edf848e0a332c2c9f3092b520f0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3491641b9b31f5bc0b550423d87a688d485f829e4688ead90;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7aed3ba5ea38b574c9a115da94e34ba3749df5c53d70d8a67;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h60f429ab24114f57a21d29d8fcbcc9ed0ba8764bd240af2f1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h68caa29f6d5c34428ac80c8383d9ee38597f815f3d59e5a44;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3ccf4b220d558bb5685187d1a78c85b5cfd5cb9f186425dcf;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf7e975e0df3628d3e996855040b159eb897ea3ef001eae1d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h40def8436dc05611b44dabfa23a95166c17389d3b541c1078;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h27c2cc2bd90d6cedbaf362091cc582cd4b223e671c698cf85;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h94c900c07f11ff0e31c3278a288bdce4c337f5b98c3d405a4;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7759e9ab1a71f7335a9407c915be05d51d3012fdaac524b10;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h24eb6258adb2f4f1df8b52da49f81048beb5d29fade0c6324;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4cb5fa983f71b2336793bde13e8b55c993cf1a72d48b0a7c5;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8711bdc7b9c746e5016aebb01e496a9057363f828605ed3d9;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd3bec447fb667d4c24fa25164c9df9ea9ddd414335b7ca500;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'haa16e64729dc4d95b8a37ae933dbbf82f923c4b1b0bfdfddd;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h27371d4d1fce02e79b8a4bf297b5644f2e68d26c069237931;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h93624df30d959578f8af27c45beaccee71278eb7d0891d770;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hff567e90b9642ffe874e8b93e90e0330e6ca7d0dae0c4dc36;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h32efc0d8ef50a98bd7eadf97e8298e7314e0c6385ec081a91;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb4439601821a69cd0f42ea1b9e78e3cf11a20d134e512cf00;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc12c08beede5cee664d13802bc0fe8c08a066802c9a5a0f3e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdb7568d7468b811b94d6684934d65db9edab6df676fcdba40;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hab3222fa006e1afc19e9a224ef7788a5ff55f7c1ecb0aa42b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h806823b14601e2ed9fadb7d11d8a0706e10a40a6b9283971f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'heb5325ee0ace20a6e68b19e110f2c651598ca404d8048e4c9;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6965800cce89078d828e0eec7d522a940fc21b85cdfc41692;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he54d7d1bfe20752d4aafd8f11757092abe51ad24fb6a4333f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9fd92ab811c38ce2891f360868701148122ea0dc793ebed60;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h25821ae7b05ffc8cb78352549679460c2d0ac72585916dd0a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2cc6d9f3e6e052537cf6db54ee2406561199bf8c18276d97c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h989dabf2839f05c1dcc14a46293b51c15fca0a8d1b9e868db;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc43c5c6cd68d364d75c5764c9bc0166536d7a37894d21f664;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb0c2dbdccefbd30caf48fcccedd2e7c75d571c468654f5be;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc713f1879647e000d008bd703db2b967a3648203ee2d97d73;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8d96627384871f0bff29a609007fc4860911db2c31268ae77;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h98926867f1bda89a123e820185370bcfcd335aa3cdfc5b5ac;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb7dea1e2d863d57162adc53cd45ce3dd07fac187ac9b27522;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4ddb5df066eee6564782b65066a63438cb1eae7af15d67e37;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5a4ca29cccb4b89ab5f6e1e96648ab37492b69ba4a9459884;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdc77047100922155ecea30c5c86e2953a7c53dd0094ea2bf0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h769ba15f26dcebe173b1aaa004cf70734005d6a220c5ec117;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2284f84d6181616f2ad815090172867ddf9a40d5543c9433;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbfab8047d64c44d1916833ffc58dc94fb0eecc609513793e9;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf75a7e702d1fbba15527b9bad606cf1a260e8133e82faede9;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd4fbb33a1946f0254a8354278e7d8d76be61513a1152f7fe1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he791aae2c7ae00ad091e9527a284430a13958bfda48179c16;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h380aa865dc5793191bd9f75640f8e4bf45e9e013b434e4024;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf79b42b59c3d31f2743e3b8e047a6fc8b374e44c92a6e9ac8;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h83fdf1050e08bad16a49960bfc0c75f81ed2d5f6d013d169c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'heff90fe2048af657e5b670a88a77d514419e29fca2b341b6a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2a78e2615ac24d4007a671e9f2e336f069d77dcfb6fd7f72a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h195892c0f862261196fbeb2c6a7375205f6d1f351e2ab695b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6a83b552fc0e0d638fa94e5a5d6e8628b2480e7fd6ad508e4;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd756242588078e4323751a8977803d4a026b79d1e5d69246a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h87247e57d930d808fffd02b91da7c29ad084403da576420e9;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h790cdba058634d611c0b1c6c5cae4ff09c487f0c59cbd4365;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1e99e69a08eaebb3d4dd841dd83d2703b286c5bab1e61a755;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h781f7d562a0f04f6d28a75e3879746d6d2cbb0634aa79bc40;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf14137268ed1e74803a0f42aaf83ee02f952e9297f27c62d8;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha2f69b0306f2610f29a419685acaed50a36d79ec3843e7784;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdf005fbba3f0ff85322dee47d1399228616bab11b7a74e2f8;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h998a730509293e4da566d68aa706274538f093fbbe1e8858f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9aa85ac11e047923ede5e5e45aae937fb1cea245120653a64;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h21b5268a624df8364d308647884481688a528a7abdb935c83;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h103e10e66d9f02a03459a6a45ce0e27d43cc3a0515c46f4c0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1cee5632ea1e26bcbcf10c807b7a5638bbd3b8b8211235de5;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h27bc95560eab40fee95a049c364df64189909eb5c5ea07cbe;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7e5c20261d9c5a3eebe4160b8540c0c7c8db5f7e4a0778262;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4d9707a4ca4b57dfc526ad6968e3f9861be562407f0b1a42e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h38a1e0e60751ca1c26ac82c67f1fa1565af19dae717a7b4b5;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbb1fe897ffac1d48f3830ba33211d231478444577e6424fc;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hab90e3f41b3a277db83cc2ad2d6e1cb48cafd0a2138219ddc;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h38d0cdc715446ba000a0df4bb9a8ee4cf6d33c29fe22ed0e4;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h695093aae9c7b61c940f1afcfed2a197aab00c8d0545c9fd0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h367204f606630ad4c410e083c2fd3ee4c8f7c44188decf938;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5c226cc22ec427e032603c9c77b36a6e7c246a8aad6ba6fd4;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha5353830d694bf3fe580413142a934abd9b75a40d5ac3cfde;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1ab9df6ca2c0193975ff91b6cc20864503256cdfa7af61451;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd4905d19b294a43b8892d75198fd3787e394944cb7faae7e2;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he3d1411162149261c1a91a178221c72cc3cff174889bad77a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd337710f440630a1f8d48128329b04988d1ca350b9930b162;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfac4373e593af32b789411bcb9059232363c8c6df35df3b74;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8fe087aa7098f68e01594b14d56a245b07d4ea4d8d49d9bd6;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7e0dd9c4d7eb1b1f8dca46b93e3ecedf7e6573ddcfa7a30ce;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2440da8bfa58d8b12402a326cd1cf4a43f871d2bb5a20735b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he8cd59582ab14f824b98822ed40988bca4677d5269db8dfe4;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9416b33274f45acfb43414376ad5ef26b1f737a8f5eada1d6;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7a461064858cf8ef64fcc88af732aa7c1d527914b3771e4;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfeffdb3a747e36512b47eac949cfa787eb3946a0493338c98;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbf5030ef44b30533b4f3488e6a86d0831c76047b2901aa866;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc4e784959ccb18e13b53f16194bef7340fda33fb0f71d3947;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc7bcf08e76fd8129b84ca8ae766d8165187b1a6e86bac069e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4564f771675e738142e2fef0565926c6a931c6dfd9d0f1bdf;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb0309035a9104f89458b7c196cef0a297e44d94bc64f54d0f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf7d4c08d0197247a525940007476996aabc5fb3b1a281115a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc933429680ca384f92ca03bfc0ab483f27593ef2b0715841f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb32ce5e2f80a4a914946c1587ab4aafb1399348342d8fe5be;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4481473d1c953b05d01888c34bd79ade568a4f16a45ba7e33;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdd67e2b5fbc9420e9f5215d92ca36cd9f55a93a33d54a414c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h91e57ce38aa6d8c55a657e4b8c688c5c61e1a95580c96781c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha887b20c2b0888e228b95d47c4c0f441810c0f672a1f9ff95;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hebce3236424a9a6ebc470b6506154be625a9129894f6cc312;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h86595c28b96029377b85a734eb58f78d1ffebf120187578ec;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3e2eee728c39a6228a90a6fece79b7c590be8f63fb1e3515;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h30551f9396c8d349d9032561e53de0701d7b693fce56c05a0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h96f5df8e16e9b52cb9e25ac6ee8be480a53d7786ec058798c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb923147b141dcfa3a45ab95aa2b46549dd4d4f296b361569c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hff87cc1635eadb669513abdaa1d3a5797ceefff3bf74d5d56;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdf0e42ebc56f37a342766e809bb0303f5538ea6bf4c9cc138;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf3dfb6e6a25f96ef96cfb54c2ce3760c9f39ef4f444da9b6b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3e6a32dc795522ff880d3fcc0e2b8d3bf678224fdfd4a1fa0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha8e8b0a7679cc5f828d566bdcc778fff6a37836ce26958ce9;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6bdccf560dd8834d9a13d877f2afa496528174b0b685e8141;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h152973b91be618b51c1f463090db5765216d25a051756abd6;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfc461c425e49c34d298bd1c23329391decc5cf5f68b374dc1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h946ae967b4b3385c5ab07a6b7dccb71b97f8f48185be6a42f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcb49dcd43f287115732a39c4d4835ee30541a7d801204ae0f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hed9c7b4e01086c8b942d2e73102b3312e2898863401aca9e0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfd6579fb51d289f222af2ea42ebf03bba1680ef6161ba6a68;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h308c59c2fd680c2ca6bc5e33d1b65fa195a1b630159f1bf29;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf31b4aef71d55d01e7dfb5fa75623d0ebc6d3affa951f3b3d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha63802dd698597e3606276e555f9dcb5f5a4f218a7f25f818;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf6621638977fdb966d3401a805700451fbb0d1ecfcd6f8147;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbe7a437925e1d1f87ff643af6a6926a4a58cdd8dd3acb2e43;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h47324e7e1c8113f7121cceb9391575feaf624759feeae12c1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he2224076be3412496f344c6c7a35797177caeb83adfefbc87;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he56e1be8d3152b8754680ce7b5beb84c24c0ca388761edd4f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6f44b72c9be752db582b6ad81948a7cc65e1de9c1b4e7f7b0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdcd351655b52c2148ce717b25b039417b1ffcc3424f0b267a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4b848432a6bcbe00ca642d232f69b0907f12e8b470c2f0a9e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h87f983ae59e5292ad8d0ff137787e88b873b6283353e9258;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf10b0e12f002c122f59446206b3a0142aeea2602d3cf325a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd32bf383a7a21b65614a62146dee384af2f4cf3bf92c69120;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9f8fb2b7134c2118b977feee99366c1e0408737bcf4fae58a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfedab4a26b2e0618f0b8f95aaa7e4c7fbbff7ec372769da83;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc4db7659b57cef1ff8c70a6c55ffb95384e3512baf146901c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1b50f9b5328a62c7b0eb67c867a6a923fac8a7ebf39a1dbed;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4d500efbb76c3b675dd643340fa9ad88fd6bb17e680f70645;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf326f1436ada54d381921261340e33263c2ebd985819531ad;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8be304b3adead7f86812a18737f9a7517c085c62d081a5cec;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfed70b41bc2ac39d9d5601939f18e8d966c497f2d83a85e4f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'haeb91258f2ecd370115c72cc46029fcf63321cc38666c231;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he4886f1c02cae8368a04edde6da959ed754b40930589d9561;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9037c61c343a71e70a004771b19d54df4b85579346c0b0286;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7ad3ae209af0c34c143d34c9f4b5ae0e0bc165256f8aabb6d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4ad23ac147885ac7a8860460416542bd23a89a295a592c18a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcae262e2744cf9b3ec7f128c8139e30728935efbd7e050ee0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2b5d7c2948fc83c9fdde61941c3152622a49ab086bbe959c3;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'heca4258975de45c02ee1aa961040a2dc7340b6c5e6656c7c4;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4c62f49cb8e6cc86253ec4c2686b1fb0cef5d4b8fcb854e0e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3b313be163c0931fa72e497355f508e299c409bb12ce3fece;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h84a81c6d4e3eae9bdf9ece161bdfecf69c776cc0873aa64d7;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbd452cdae9ca87ba9568d26bf02786b948c82a257352ebaca;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha78787c91aa1a3ca10b56abd77fef87512468eaa5b173a017;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5cb2a39d6a1953b93c7cafc9e8e7facb1f7913ba2eec24340;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h43a09e65ae920f56e3d685e0c9255db748e2b7112b76c65b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hecef1af0500926ee6986ce6b222b3a35876929bbec72ce065;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha4bc0d75647ca31edeaebe35a54a16ab751d9239e60197366;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4f211ff357fae5f25568c206f443119b9d3b2e51f8da81b09;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h777ce06b2fe4bc1a08f0ade5deda437de16b5fc07e36d46a1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1eee9231b9ad7e0bebf8e7c457b1fa118e44a53c5abc79d2d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc61c6bfd0f41b36766ded39ce1f39efa760cb7a7db6e20885;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha6133a2026910e2c4a9c66621a6a6c5c9b7f63b2e93930a89;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h24f657b4ee8e01ac368fcd24163f03146d5ded085380c18;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h945de27d4698263a6c4b6ebb0aa67f324aed6d64db4ecd9c6;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6f29cf7505eb30f717f5525135031fc2c1abad4835bdd5be5;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7cfc5f704b76a264e832727ec43a9aa2d019f83d7676ef244;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4e74900ab388a29e6313598de4f48f26cffa5990e77b2b0e1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1a14ab3db6038544858f74b8f43b8158b8c3a32689de1f663;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha9df51b6cc7bc14885592600b6993a725dd3a1cf6bb6c5834;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he97f52017ed05dbbb8fd5ac967d1c720f81dd41cb1e25524d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he75c68e1f7062f6ae6afac7a1403baa4ad7532563d86b194f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd752dd9fc8ca874d2d6fb77888b918bcbd090f29bf8349100;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7f712b2e705f55fae0e98c6d05fcc8c191cf8f8e04d9f99ed;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h209dbd6f39c713ea5b2f9859b0a2722faaadc46bb7ec2a3fc;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h75485928d28130f8ed06c20ad332bd241120fc835cf50120c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h81699ff3664ba8470287be09baa92f7e463523e20dd6a7a7b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h96a88b9a7ae48941c2176ec92d0e4935d31869142c8d29706;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h79a0361b99a4ef32d2c1459411ae13413ed7afb0e4146239b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3079f10a055d556836ce73a8e589e117172243c2273a20fde;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd483666bc5b565c138e2c7cf01f22bf7b3b2c1f8fc3233ee0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h881b5b8f7d25cbaad0059a0171368030af2a0490b84eeb888;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4da22616f1a5414f8a91030f321ff39c2caa1b91b29809cd5;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h98c58b6a7f9fbb7a6cb375c3211f8295fc201721823fd036;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcc152571abe10cdc94c8da9e11fe72b20de3fa2c13137bb2e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcc328f91688e5e1e185780db94ab3a2e951e6e26d56a65827;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8b733d1e0df6cc2d69c85b251e58f258be201964100cbd32e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1b5fdb072449400e95321759cc090b4f4b227c5b5cf7184c7;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2178cbdc50d4a805b873e4de75156c1dab070996a41cfdd8b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc1f9aee10489aa4decbc0de40940bf9a12b2d3733ba8a7c77;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd23adc2175882cc2eb9d0fa760a591e6d8036dced4ea3529c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd55d818ad0a7a4083009a8967af2c18bed925a747654204b0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h23c6d62ea5cda9521d1b60d139c695080002888ab0ccd7966;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he71936278d68d043fab083eb78def80a53d21bb44c47061fa;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha76264cf126ad7b2381949ab36df3b31e522c4e3d17dfce3c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5d94b66c2c0207042d0ac171c7bcab22a7e7209a50d331d61;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h831e81e4ffb77843e6416498f8c91b298bd3b8c40a079c943;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3c8158bcb7de35bd494197d2f3b458e38e0aad66373db7389;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h40233c0912e9c8266126557630ba88dc67a2f9a8703191069;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6b1c66b0e8cfacc49cd2e55c889cd9e55967e697b5b4ae5c1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5111a47b6d74c3b1fc084fb57483505014866480b802b7290;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h40c3778444e21998c8eadc30ecb61a932f6c28690acf36115;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9e904ea9b31f4709cae5ed3b09562263cfce186f1109b9d2d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd6a37adaaff65954cd99d33b1f60c20e3eb29c561b60a7a95;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc0e2b7a227d345982344827f30e5ad82446b0ccc0fa8ae44d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6a723df36b3dda59249cafa3e628cf617145d89cdb51f7adc;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc0175da5f0b894eed6d2ddfb12334ed3856dd2c550bf46411;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc74051676cffa746b53b5aa4d8f3b3036de75ce396c3a3aa4;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7ffe941036e3c080c8a47b0e6cdca676942c529b8606cd97a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h354aa216c9dcba0b7f7549b9ccd6bfc8c19e0f0ffae8a1e11;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8828986eb3b0585d1baeb6ae7104bcac68907d0875867f661;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5a29cda443b9ef297e693b1f9d88a10ee65c1f9679c2fc144;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he3d16540d204fbacdc7f7b6a4312bb1fbf7c2a9657a2db767;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h58d8373590ce8f932354920149450db8cf03d78cedb56ed82;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1f0c961a7fd55021438aced440c7d22db01da6284fcb22e35;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hba8d56c04f3889fc8ae80f99823184d038d8947522d666527;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6efa6d5a6219ba5920c41d207eecc16c262504d96272c6203;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1dcb07cd0fb543b4a8345ba18bfa9bd82d4607b9666b0e693;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb3e9e91860f8c4f0316fde8d0f89a3b550096392d1f6a3189;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hae1aff1106f1b8412ca6d7cfd67ba946e21e536dabdaa37e3;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6dbff616c03773ab432c2869f11cecf33990e8e165976530;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6e9637a93c181bf455e1c004f095e22442c10392b4711473;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hddb23284748d05baf8b8bc8bb0d3672bc612a0d9c1b00ba02;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h73e862535df15096928a9d5bf76fcc3c176c61abc66da7c35;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfdce71412c73f0ef828d235b84c534a28846f50dda49028c4;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9c76e3ae415b562b98beac38f272ee0a3e1c109899c1c2578;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7612ee72b6b37247086ef7f754f20f50ba7bd7e707186fc61;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2fcbcf4ed008987fd8294d503937a6eb3ecd5d05b514bc04d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h93fe4f735c2d803da6237ab88f2188fc4243564e9c44fec8b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h18d0eed421f81ac6ac2332683216aac0493a9f0b29db4ac64;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h404359652b27bd703d1ec03751049d1bebd0660de3eafbf07;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h30cbc3b0e6f99d5d07557deb1b2e97e2a5142c975a66882a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h895dbacca977fb610d56395f1fe6a94cb4d1c745b69c45cb3;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb461ca1b057f740b587d648721af21ccd7533e16abcdcfb04;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h13d527bc47ffa7ae856d74cc138c22eac840d88e07ca74ce2;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h555cb79f6bf59bcc46d5bf9aff9b5f3794bc23d9d12e3491;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc10c2186ff4ef4a8ebc418b013dca7c8bfdc712134ecdd3f8;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdd8883b78d4f02a5b9d38d49ad25613aee928599ae250d92f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9609735a789a4b9c83fb507564de163612e0f61ffebd4c39d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb2342dd6a092a8a0e631ee03c9e8384a574aa9afc322e1833;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8784ed2c3f0ec350a15eada60d35579f3d1c9fa826f82347f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9b27cdee158bf5a76426d77f03ff6cf63304208674535882c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9dd479a331cbbd11d41864785afd7f6ee55f4140823de2c71;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8bf9fdb21f64189f58d5004fcdeb02dc020b4b45af059290b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h68567aed7084156de1b136a1899a93cde2461238baead92e9;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'haaffd78cee186f3cafa9fb88e0074833f789e36585fac8090;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h589f3dcf53e562c3585b071e79f6ddcf4c957d2010e006150;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc6045b7b27899296532fb3240164d2dd2b2b821a9096c2846;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h17278484fd8ce7df004dd8f90ef7c7cdac192b24c525dc0e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6469d001cca3c755ee7a61090b5e22390d10d2316f681830b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hec4aeda3c4b3b4e497fd509b39ff83aae2751d844b08082d5;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h91021d40b3b5f1d7cfe65682cd546b4c95cdf15d092663536;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hca512b66f2917e6a6aa8729fe541af5b940822232fb16353d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3acc4df236fa561cb53e00cbb8d4f24999ea12a6641e47c6a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbbb93d4b931070713699e5ab6cad0d01109262c25834a0da6;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h99890c1abfbd22c3fb8701a268347d3037dd1707203a7848c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5c2212345a6eb4e918d8b8e45b2696a8ca67efb6417bc43b8;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3e3737cc86df7b4f750300f39b579931e1d780d78b1df58db;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h900196e274657199094b6532e9aee79bccee4a69878503b4c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbf2f6450dd589562c35fe720d8b0bcb6008da9a82c0340777;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2c31dc67435795de811c50a7e6f20079bc193e11ea2fc18fb;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h639c1b2da2212be80da20e3604da62c870af125093ad65542;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7415790a5720c374990576e7c08018e30d5d7e7167accf2df;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha0ae918c13bea1af3029e7a473079a665706ea7a8b5ff305b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc4004a225db3281e628d7bfe874b0c4f9dd631428c1805df6;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6baec8dc36d058cf324b5ccac239efe099d0f202d1d52f04;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd943e35aaff78e42358a8a9c4f505352e3df451b5c4d4431b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7b076a81dcdbf95d2e7117082d3a767ea552355d9ad3a2251;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h97cade4e7d0d1b16a0a5f8da29c2f77738daa33818c2d51ac;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbcc88afacc949a0360f853382235bf042490844d517967355;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8a823b9b09d332a12f9c8cbab289a495d0a99ef02816f5603;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf3588ebf44c3acc5185e5992c5dc9b017f515f93e3088b05a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h87f8b0e65467ac36161d92f35780145f43cc3057984fdd196;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7d4373e69a5b236916d8a3e1c9072abbead543ab9344b4dad;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3944d07e37865cfbb0044691ea5ffef377f9edbbc2fa3287d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2d3dbbf7023777e66e7089e57683b7b59fc10dd9178ad00f8;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdad7b9cd2abbe319a2e344847e789f89d01555689334314bd;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h84712f17fa9611428e514c1c56781243b7a3db41846db19d3;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1015eb157ecc01fbc9620927707bcb428e75f886f509708db;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfdb8635b78a183b0312877df7b60916042b7a08e6dc2fb996;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h888af2062689c4f94d64a65d27d86d56416d0afaf8884fdab;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3cafa78d8b3ed2ff56eccf8f1ce8f0f664d5af1e5086dcdc5;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8622327ba00716e19c3a4a3c0c50480495f0141d94ce57a69;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfe481f87d97c426cc5bd7849fe76acf9aa026406a4900f211;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfe588b2bf10c838ba097ddc56875be3195d80ae3bd4176295;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8b3bf74e972fc65c5ac862892a618e4802150d1420bdbc171;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6a974796a32e672d409b97c44dfcc50c005bc5e05dea7c3b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4593b631dca87906112d0c86797f8ef6039f78edd7cfd909;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc1b1002fef55fa982d90f7b19360f27f24bec6cd8c07e66c9;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h34294cc35d1779d2e92f30db6ad8b8c429fa751de7ed929bd;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7292f377ec60ede5de5f3babe81e1de17efeca01440f13f20;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h85698308a8463c05235bff826455b6ddf704c2c4a065412db;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4a9b126f074a807a9f1331bc41e9353575efb525dde1c3d35;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h14473b3d2522a017a4efdc135f335a20c1321320c57aaeef5;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h737fe792f3687a3e40f8554ac4a5db5f3e92bbf06032d813b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h954f903c87963eeff61ace67098a3ff67bba221b97fc2a1d4;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcbed7bd5a5be73fc4ecfbdad3f7ca734d11d39d8bf1fdeca0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8547913cc15a2cb9bc6520ef8d737d2941985ec9f0a510375;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hec4b951bef4e398104fa701cf48ea318337198afa4bce3163;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9ecbbb013b51e25b5f3d7b935d8bc0e92f37813ef73e91a91;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9ae6e772937556b20fef0e88872b60c4a336ecd69b8d15b51;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h65002275d41ee5120d1326e144f08aafe3b11ce58c011c583;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'had46bdf49cd96d18b0ed2e1159a7fcb12d067d7702b355bf8;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h858f62d5456800d72dbfa33ac29f99b06ddb49d39b705a5a7;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc51ef37a9a6d1a8a238468782c3e632a5381c722dea823f36;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdd38baf1a3ceac94cb10a26a482daba2a4a2cfd1a1946d9eb;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h798e5a6de1aa4c88e513d441f133652ef70b03aaf0982dd81;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h90a6df3ea1dc9b7d5db1f6ce4cdbf229d80ae6572d2ad7d20;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he864bae8fe386ab27b6245ab8baf80aa946ee111ec62338d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2adab35dac81e8636b3532043e9a47b2e950accc3db091527;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf5e1ed954d75810071ddba68e0a3a9664cd1b272b3f074609;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h914f833c8dd07e470af0bc3576b1496edbc712f20fa410fd1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h18115f818b80911ed65cd8120c87cfc0e08b9bcd326234213;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3b9484cea7103f1f6f9d9d834aaec736cb8d49ccb4f298222;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8141d0fca5830f8fa964c3b886ed99908417da7425e4c7657;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h85d5000d11c998f6cdf0961b8a3ab77a66478296f8664bca;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf8e2db4470744ed497b3ee4cb35e86d4b1298099be3536b8c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfa6305e562944bb0b9b206bcc187dae276bcb505ac630cf5f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he04a06a1b2582905c1ab925b7863fed788d6528bbfe84d567;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h78caa6a8c1543c85af67aa63f5032f040079a519292d72a6;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he26f9faf8cac79c335cafcc58f43572a56d91f03b34268bdb;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcd4e5a7e68d7455587df9886c92526e40084d9c297c83b16d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc460dbfff8054b1683c16327164f2f030221d669f195aeafd;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h611835796f31339d6784b71f720698b5cf80e5f12e6957358;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5d4f87f2d31cd0f3db31ab1bedad7814593abb61115f896eb;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf23663ad6e18a78f8d4a007a0bbad98eacf905be3438cacbd;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1a620a3455f409f08fb126baffd7edb4e76a434d85f56e38;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1ec6dfb9393ec7d4e9d03234fb7f3505f0e9e08901bc11d76;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h37956ae2a618be2f8fbd5162f85df060fa7fc590106dd5729;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h926aa99dadc3a4d18f93746fb3ac9edc004a432a2ef36b756;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb452523958f77e7112e79f90c5df62abb6f7a099f042d241b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h320e6d0d8502691a3366fcaa964e8ae7ff7086b61290834e6;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4a80a3ec6716cc3727b772cc957b19e660804dee5af771e83;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9b9a9c354be6fd4a15fc92f381985f99fe1ca1bb455938ed8;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he669ec23cef1b8a31ab1294783c593f272ca7f52905faf252;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h61c89706bfb7fb435382db6e89fc22f870a1c90ebb0fe8215;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h74d8bbe2834660ee63b3d12030b10607de69d7fa6c4a62dd7;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h59848f270489573686dd41d96df29d2ab18fff703c82eb65e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'heea1ed69b91c532a4347a323633222ed6880a0a6b43947332;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h31801d0f5b9bc091b25fbde98660e718fe3ffa67d6cb90d99;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfb8a765cbb2ff2235dbc8c6ad0f47c78948bb571fd735842;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb1c92eb42cef5d42ac118fc7ea3087ff8757e9cac85e3769e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h84f78ccd3e6fa610e4dfab852e29cf1a26046dbe4dba98c92;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9f0d5bbbd0ba2f21762fcb733bb2fd2f10e7c1ee858f27f7f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5d83f04a98854fb3372cb9a326bbf73449a5e3bdf57b4fd1e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9f02715a5a4d4cb1d6e6415157e5af9125a2aa5eab1a623ce;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h85858cc340a0e330de96dafb1da9fe3c8092431c92343c138;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h714b6aac2ce088558340c3e937f2f9d1ec8a0c80b9ee0ee8d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc7402029b77797384f973b218dd430fd825dcf33b0678e792;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha175562e94446a9b2f2eacabd34beb70f5f552f925638167b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h49cfd01d5ffdd5d687e581ca5e625088252497405f0b507ee;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'had09bed390dec2c325b12e344fbb34bb7956660088dbd7164;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf0e0ea91ba5a37ae0eaa268641c176b340203a04642f4e30;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf999a5b913802fb16b7d066603e8fd655ba92198824253cbc;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h46bdff7d2d0c70788299223d22b8dd0a650c53752934f5f6e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hba5f74320f36a5c3ec1e7098a6f2f1adf031a0d69d7581af3;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2269895eb3ff0fef6ea41d47e226565786e1856d582c7a724;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdac8f82f0b7e416bd90875da20733dfbb05d37583dbf8403d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h51739643c5c9611d2fd9d07046b8ae06f8b66d52b12d90c8c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc83ea5841f3468ebd1207e56a6fa61f74f230367b979eae33;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h545364c7d8ad31beba34e4ee147c4ea733170868a3f4bef8b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9d8389d4ab5a472df2ba79f9f7cff5427348e969b5fdf97b1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha14cb085525bc6d807fc9ed4c804f5b3058129e498b89ec88;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc6a0b82303764e48d704099a6cdb55e7f9ddb620da733957a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3789a09820b5eddb1255fa6ffdc41757e65622a97f3ab8a7c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc534652ee0e8d054354a322b58cfbaf53d3f2d3afff1e25c4;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9fa85064c1bf27c29c6b2502fd7218ed05bd16ce29ef9f846;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6e505536d2b797a71cbaef6133a600b292a7a4a31efaa27e0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdcdccf51efcfd8f1f7c19b22644a4e0b4ab87727f8d06617f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h30bb318ed2d0449b8a68024935411efa0118ce02d99cde0a5;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h19061159048b57898e1f2e5240e7955d721e18b6031e6a4a8;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h40dd5d532a1c9303ffa11ec840c39f6b5d60c36e6dc6d0241;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha484de117713087ec9c4a84539b62198158a2282eed51c29d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4f47cabd2f4923e1382e3eed7534bc1f2c31e3b0f5522335a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h91ea010b314709b817404e5ce94f4241b9759c44c1174f6be;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h98b47506d7ea0e1203481dda3652b3719fd63694a40e3842a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbc18c36aa082670c059cf6c1783dab9c18cc1e403bd48b7ab;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd98a44ba005ec0ff440c97de0bf33e48d8ecd2e71c660cde8;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4b83802c665b5285393a468c693c0af3bb3738457f1133117;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he864739e5bccf3dfd9f7a18fe06a9efcec71ce064a5116998;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1f3be1d1c05c59dde1e0da2f2423c3c99452c00aca9558aa;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9b2b966324e1e2faee9b10e1163ac9fc5f8eb99a618432026;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hab414b6982b64551215f5c86721024f51a122e0faa0abd8aa;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd913c696d240a3dae76cd5038727534e11cfc7b882cb48b56;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h67fe97d6802749cda527b40b8963c1f18a30d468ebec4ae06;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7b98228a942e30949fc7c256af3c1322610fa661644aa63f0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he02cdde1ca05463dd13bf9eb93f38110b44060ab079abc7c9;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb8d6a7f1ebb65d70f1f20c4933312f0f14252e196d97f1603;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha77738259f320572060f07583360e66fa09607a35293b5f76;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2b1aabdb6340857b0c432dfb797e18cb9a089ce393539bd6;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h42c1f95f0459fcb15cd978d1db98eb726e826ab620ad127ef;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h61c29810df4bf7f244c164442869d258058c01e82970f20d0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4fce5253101eeaa6d9589959d82a957c01713dd2422f949a4;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hce21bd810242c5058f7fc9b4c7108bd5246e26fdb1d1f2934;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h619c6264f6a77d3d07c637f12a4937b2bc9d1b7990b2db8c9;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he3ba3329104233ae3367e666bb71a09563208d2eb9f732512;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7d2be4d199df59f844a85024040a8845ba03da3dcf25212a9;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h176a7ecca05def6ce32fb69bd3b873b507ea6a916b30583f7;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he697986a1cacbbae1f55c222838f42b109ef35e9b61e833a2;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h580a7bcece5961548d60d8767479c745fbb63ce5ea6716ad;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h977ae3112021d9bf098bd9a06d4e406039c26abd61aaa3c8f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc3d4db12ce41fc117a080e747b9e36e9624027da71a19b157;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha2f04a2942fa3b648855128408d73603bdea92ceaf619bf78;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h564340d00df656deed0dc19f971ecb4d01458dc6896bbaee8;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h56b82cb2f9cb1fb1bf1f82f6b27727945066205277d494695;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha573427dd47a3849b1ccac3bc50ef8b822123dec23e25cf4f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h94cb5ef0c9f642b0c3c16b3bf211f6ec53893fd45539e7c10;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd0bee1261c8f96a6004f5bbfe5547bb621782b3afca9fde04;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h67ecc44ac3e9c635ae489d79e0979715320e41df3649697b3;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8b12261c1d3bb697035590481e06241b2d9c56de5b16678b7;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5613ba99690b8bd41e20c96e843f3577636fb252f8123d5b3;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h11ff4da14c80126747daf0e1f84c91473999af8765130fb1a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h414146981bb3ce5b1a9a264a3e491f2dccadd3c6f92255c4e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf6957aa0c9b7b0556722b7adbbc64c8ed4dd85332fb343aa0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbe78529463bab87325c7af7120512ff9f03c81985269d5374;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6d92127c9ec8c0ef78d2030fd78e0b62a299b537b2648856c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7eeea074f61029e7acaa3516f6007449aabfef96ae5a99f0a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1b20ea8d1fd9635a6ae2cb1a4d117dcd048093d3ff1df7db0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2f9c554fc8502352bb66dae179d4886c19d556dbaf5177a42;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha73a1ad008c32060ca1f40ff90538bb16d38d221d6803092c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf52028a9590bd02b65c66803d5609123f1368ae8f1a11c58;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb0a96408fd7c44a1fb1a568d01787b038fec6facd3004c3d2;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5f4eb6bd3bed3289e438393b079b6ef8903feb31c25bd1d28;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h828412cf3af12d74078c2c2a650b10d454f0136c9b120c47f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h173d835776d05a2c6044a33c7afc7a03f050394dd0247aefa;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h598752bf9df026e92358fc6670383bd2a90f5823a32458223;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9992282fe4b8867d227b00c756127c0c3a152a9983d91947d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdef2aa83d4ca631948ca52968c49204727f075003a40456d3;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcbb4397df9c2d039c6ad20774c9a88319fccb819f0e49ce01;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2d640dd8724517e407bfad5e9e2c2c37ef3561db74ffe09de;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h32297f2ed1cf642d882986b34591dd2d4537964a60b2c4709;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd95071be2039737aae46d5ea57a934bf1b64ff4173504548d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd069b33bee0121ff24f7b5043d2e3d46761e9d84b5310a3ef;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcb88df952499dd5d3d704518901b038106b02342d5e23ecf4;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3f0647c5c10d0b8b3bc49b80af49a98fc123fe3f883404a82;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb4711dda4f17edf72e757cebd6488dc453c2f9c4b7241c766;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6db4e739d78f7dc2ef0c6d99bea0c0631af488d9345f2b98c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4f71a4ac17466059d4d5f6c292790a06b4b53627ac5d2f791;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h48dbf6ed8193231f8a45a99bc0432361b413fb4d160ecc26b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he850fbbc14f2c187a30ed9dfaaef6c530af6bf9a470005411;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9267e4d4037f865f8c30bba235d776b665a40380b73f95e52;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc4657d78926709cee724402f26cd4c3da4ce85bd6731f8032;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6999bc7bedc3e38cc0dd7f4c955f56eb196d5f4b5925274d5;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h47377cc83410d28e3f2e424a9b5cdcde803ca2d88c8fb7135;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h51092fd444f1124d8cc3e699ca1d2c64b29af91234fdeda5b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h56e2f086293b1ffd194c47b343a7c28997f798a5751a92030;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2618d0983bf168717631703cdb2b20b57bcb06fa4851c617;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha6ecc3cfed8a544b80d6aa691649f6e65cdbf0284bd1c16c5;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb57176a80952839614b4b2ffc5c813da86a27e9ab0c9d78b3;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hae56616b1cce7a4b4031490bbe4c965de55d2119385e0120f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf7ee2fcbeba92724ca1d925797879f99586fad215cc0ab14e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h48aa3bf1616e802b84e7913ac244f219abbd840c7e4e491ff;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfd1c3ba4996efeffcffb4aea098c0d189441ad72e7185f5fc;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h61bc948d33e62eeb590816417bad15d7805fdde9466cc9c7;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h269310ade770da3f19df2d97a046482e97f5f33ef903a3da2;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h370f9af5b76377c2477213ee14d7ab058379ffd36d12a35c4;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5a92eca28ea6281e00e4f8d6f88d4e5904687bcb5a9018f3f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'had6a2f775ebb394b45ccc112bf571c014fdb33f2f8d34bb7b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h85e3bae0f0db2d62d3b22e3f15349e31983a95acbc53110a7;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha48a637150a1cd8939009f07be10661254c6713bafde5c355;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdb9523546941344a902ab86caa90dabb8fa83e0aa9e1f8c36;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb8daaf628f82d7e66079c3158fa7035468db85b47e3102640;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc6978741192bc4f230035d256e33bbad957d75e17cc76a1f2;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7fd1d66cb0fedf0382dc4625d818a34bc34d1d11fa2337ed3;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8042030cdb4a5bb1638c6b693b1c388e6d2b8bb4857fa619a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h60f22753328a04f3331827ead6fe894ddb9a1b2240b6c74fd;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7b57c20bac000739adfe70d216bdb651f6daa8871db169220;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha95e7ca9a44049d597ad222d6b0b4d4f227956b7f8890e8c9;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdb24d7550069cfc3d3099f7a3d93002dca223ad4e2302e7c7;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8be4d2988408e93d4e0aa7491a7965c76ab92d9dfd54d32c7;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he3ee29b318dc5353c66faf64518316f58f5da9af7a2298f13;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb833be2f89e1a4513f01ede9bde46bed5cff0217f4e444783;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he30e38af702aa41d63e7f9abb8f5a727b4bd96ad939aef77b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h404ba703610e31ed1c95e0bee090846c610699501a1796661;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb008653c8e6736defe21f3cd48b48a9de48468a2d26d59f6e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6308b98eb458e28e5aec9ddcae35182fe9899abef0d841eea;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9e2fb9b4dc94df1668f9cb3f9b49c358ea0410853da5d1ed7;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5fb2e06db6f0581736398aba251a16616afb2103217560488;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8f0182176ed4763d50f769cdf25510f7edb85920f3349b3d9;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h47af2e4c60c7dccccbb7124fd0012fdfdecfc05c6a4c342d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf8cf1de85005669015b5dbfd22a68d2840ed1b75e7e5f90cd;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'haa05b6a99d17dbaac0b8d65bf915335cbb8688e08f24205d4;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h93dcd8f8cebe2c4e3b647dc29e47c4efe963a3be6e8d5f1f9;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h18eee468e084905bcdf6c4e02740ebc32832ab2e047ad85d3;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h764666c21a316f2886da214e95cdc96e1b8636a503d83aa03;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1186bc81ca2515d650d768a73b227e3d1e665e4fef1e369d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h59176ccb3823ea61c47c20b46ac5d50fc13851c6c6f85c76d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha1f31ec6eae96842ed1a6b71784a697e93b43bf725b145f5f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he09fa1366f5600dc2be6e2ad62671e334c6bc861a8fdf27a2;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h72d37d0d7574a70e4f6850a679e1efff6d3ed9691fb849793;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcddbe4c7f7feb7a9837892c2f23453aa9c58ede5015586419;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5d72eb577d49124c6882c49798b959d6aa8bdb0881bffdd34;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3bb2397ce30d61af6606beb33fddd6ba5370b67678deb5f9e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h899afaaf30565d1ae53f873791021c33025c0a13c507924e9;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd7ed1a7efb1eaf4adf44a39cf961f28f76cd063d5e475b495;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4a6ebeec7e5a5e5e42154071e4a5e98f924b8b99a5a9c9f0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h71ab99d3cdc129256c166a065018bc03bccf9b3006e56d2c0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd51e28c0b81b067d2ba6f37cd1bfd33987dfee9c965a16ed5;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'haa33da630aaa1d57ff8e057546206f2249204f7d00a779633;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h319b2a3e5c7e26c38c568e97e29ad9c114b0607b4ee2b767a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8a7de1970fd9ee0123ee839f9742afd413458b39ee507e624;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb1e0c3587ea15b9b80b858a66a7948d02b6cff56699ac0e6b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdb91ed2992253b2e660adc7f769ed0e1da3c9100304afcc23;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha02676d01703fbb9bfa5e1602b32ac088b7ec896caf658f04;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5aface7aea9967a4631b512d3966cd86355384668c91bfc2d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3b3fc0394f7c8d967c4a93f454a23c598ffbee65d16dedf14;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7246722a59130d8e6f8387937f7797ce2c958ee1123e06391;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3dd23bd7c74fc1935edac0bf3eb99efc8ca84b9ba65a469d1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h73291226644fa68fae2bd46275918cc024542369930b2348e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb9a192e0c04f388a7fd5b92545d1c819dce11539e38333597;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h78b6401ebb3f04d3416313dd4de460fe4c4c48e1668e0789e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf60c0ef2bcbc80efdfad9f60a8133a817d25eae5271f819d9;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h463dc82a16e456a42c90a434ee286db56900968450584c3a0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb5eb98c4243115cfb736baf4577bf94c13f02f7fe9ab8e8bd;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h651ed52899fc8b960199bdeddbd08ba95b78fd645eab15933;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc70fc5443317fe08013b1adeb59480e65050869f61aa111fb;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h546ca023a5901530f96aebe785154ad988f345157f6e35344;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h65626c6d590eb416bd4b8aa29d31dd4ef825e7004ca3fd76b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb0d7c89aa4ade6c006e8916165ba6563d1b4c14f596cce946;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hacc38028e81933fc2326bff9e33cc0fc47b95c6ade64c2b7a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4377b8cebb6ba795c921dffd0f52ab5000fd383bbae5b066c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h742e36023e2c331e6790772e89604db35446c69e4f4f45dc2;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4f9335b2cafd29100a97a52d7cf166825c9fd6ce93ff11886;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7deb79704cdd7b39842292077965b686bd69cc5a511b0d599;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9f759df584cf42d01eda353f59aff995d63fbb6764c995cfb;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h16705547a223c6c11d933b24442b965d498e1e32a40c216e5;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb85fee431c7d95b5d9cc8a8788bae44583ee54179e11cb938;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h349e9545cc2243e12994efb6252a111956f946b7f39cffad9;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h349251d81a3e83cf4715a25074c2f4f4a65a9c2a94dbfa4a0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8740a61a699bf4d21e4c0ffd947736bb3d6eb9ef66fa8e710;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h849118d2de3a79b99b4a43123651e07b374ccfdf284dacc36;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7f99abb00151eafbf5e971cc96d86f385d926a7b98c4ed94a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3f2944b7d281220079d19d4974cf6b690e236777b79f074a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'haec63511e6ca3bb95c741bb60ac235f8a4ef3671ad75d7a83;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdf5137749b4201054a310c6066d814904c539f9272aa91393;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'haed4a427e56b8fefe0667d204acddf42dd440705f1ee33f99;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h50d97ddea0d221ba290b8214ca2bc1a1899d6537c0199c7f2;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha680e4dfe48896cf4787deeb7a88f021c55b6cb0c22f47e8d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbab5aac035e9207fbc863970883ec581497b22307b818d5ba;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf009e7c2d5ba335765ecebddbf01c4b54be3bcf2ee2e5942e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h340fe112f430361a965cadaefb55335d4546ba14f5511dde6;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he97673277636e02a156ee389a713217c7c094d226e5802e9f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h78a860facad7f558b640d4726364989c1c3fd66ee01c07845;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf72d99032daa49e8aed57842d42e18bd6b1b663b84022fdf;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4c2942e05eddf5d3a0c6fa66df9e97c350ee1d4c78dd95441;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h61105a8343dcbc915fd7aea4631e652ded0dc125e36cf728;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf04eb7819a73c276d519928e59f1f01d1afd66409a92b3070;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h901fed672118f898214fdbc187faac636e0198d37d6b0b2eb;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6f09e705ae4a57bd45c9f06832e77244a4f2029784fccd2a1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfb2ffda1e258641056fee94c31ec3d4fb543fcb8436c3a149;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h98c2e6488e3a3679cea9826447113f613d80403e93fe301dc;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7eebc6ce538980b8d6b627f9cefc4316cca2f68445030a8de;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hac519a5c84697804c963b3798632350ba71cf40a9154fc6e8;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h18197b899e25061876f1c45036261e92759f9f081a765f2c2;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7deda779d68aa971f480da327abb5258357d1fe1d147957a0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1ebbb2a85781e293e700ff47573ac94c23682c7dcd0c4e5af;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5251ecdda9b8432537dc807a3de83b29a0d1edd1dca4bcb2b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd860b91a548e5f5aae7c059b11e55179b974e266a407b4872;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2cee3553a327f8e0ae862cc5d4deeccfb26d3aae4941aaa13;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h837ef6fb42bc2eedd2e8ed03c34bb7463896b9cbe670b8f73;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc83bb4713437e4dc4dcd67b3c843886d37b2bf0a4dd6f739a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h37fc91a29fc35785deecaa3950b99f5867eba2c4d091269fb;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc5244e5ae3452803da9a205b398e2cd012cd127a773bc3bed;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcdff7a66a0ba3439140be1984c73e4c0ef4f2d1225a6d15c3;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hde9fc022d5303a4de94559d0c929a5bc7cd9fe3261bf5e195;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6ae5ab20bce291b7edc9b605576ed7d371df55570c5672c0b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5f25e66eb6227f08748acd4ed88898431b2bfdb1d05177452;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hba20616e29283262ea361c2f4eb2de6ae308b9bf9a3575fad;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2a9e4d9c7e05937724904edd4d685b8b3db170ab253966350;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc6b5a086570e71c00ef2d5fcdbb5dc11417dee14396b825ec;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4ee0c444e4ca80798a560456702d926ea3bcb26b1bab429bf;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf04c3c9cc58a021bfa9cf27f990b7e5b2b77ac3754362f719;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2e4b5502dbfcfd68a1b628d773a18dbb899e29dfa00419959;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcf238f5a92662c58943331af44afe91fc0bb94029cc115cfd;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7e257a9a7a79bc54263fce477f4c5d728abfa1dd393451531;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2d449fc8e1be134c58895e9f494d736f1b02cf851f4a498a7;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4ad70e0bea24b25cd47dcca8e857e1d7ce4673b5dcc1280d7;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h17129a0e5d6e0d623a42188d41665323954a4a39297632738;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb503bc4a39594583c6329bd89d097e4d0a29ec890314853f2;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h440d2a67d44a7e4d20be2539e6be5a6764bc2c1fe72b7d827;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdb6a8d325847d46accd9fd30ef423131294ae735de0a14d6a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf6011b159cbd81298d3e15d767fa9e2f7dfbe36328e39d7fc;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h58e9db4fa52aeecb2c2944b112bf11edb777b2c7d5d2b13d0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h98e05ac0d6959bb256fb412fdfa1f0f4799449a65f214c2ef;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2f1c0f08323af3c5537b4b95276387f1a2aebcf108a745486;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h92993ce6f57ba2c1093ce887815667ec9acefbd00394a5854;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1a46fd4f75dcce5e196f55854f4f54a5f8e05ce120ce1b879;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8d94babf67a9f4cee3d1a0f3c2df42b0a6d41e55b180dfeb0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3b81ec382ff8afd2e89b05b9b1e1277111c7f7275b8379e36;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hce7f5c67c4b2d3f2b92488034983a9c938d23eeaacc760833;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfa3e5c3f8a81e32fb9c745d356455a68f66e35f280cae9bee;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7fd04908209b8ede4c001a61facb190ac01ee0c6191d75214;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he6bd97f38009decbc9b58f4097ab236756752cc952bae8399;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h27612b0fee585f43b2c1bdd70d1a257644af681e93885d2c8;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h57b22fb57231eac0d72bb7e007b4ad3e591690dc96bacf61a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9ef7fe2ece1ce49e8a2d8d0ce1fa546d0224f2fe01a3d2023;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he0eb00ffaaaec264592bd916851a5d9e099e000cad0fb06c7;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd189a369b56c24653eec33f4ad9d6461ef78d0c6be576ac05;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf0c8f7c57410470cf9de084b7b2c0fe9dda333dec0f9dc2a8;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h13d30fb13e95f450135f5260b8cb9109b16e1dbd0cd362d84;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5f817eae4a150aed76ead5e007fc22296adda97ab8b2d7d0f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h86abb2f86bb452b4784ad4ffc9e1c9515ca20aa5a69d698b2;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6abc74bd73bf45ee8bed8c63a284af8c6cfbc116ee2fe6364;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha6ebb3379dabd4a70931d0da0e01574ed23b2ad20392eb802;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8be8a9d966d4f0b3e25fd1f54a5a21d14fdeedfd76ed7a784;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h582cd27ffaf40132618af4a0a45492325198425354766cdd6;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb37dfc5f883b585bfd2dc1dbedb0511661c70b1ab2e31b531;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcf6dca0a8cc17f88c2e641e81e1be87b6a22b23721bbde5db;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb36c6293cfb14ace1217a86e292d9cad37e9b13c323e395c6;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha06d09d325be4816c4b3a2e6be39385103546ff21b34e1911;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h67b1d699443d15d12ce87008b842bf9170485c71406eb9bbb;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he61b96b3932c9df0e321286076293c153c1db7e255278ae5c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb5e71352ff3ffb456ee4343bade5e4b8cef7c1a17594b6129;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h17307e6172af0de5fba55c6af857cba5e47cfbf862b528ae1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf0db9be03aeed33695a035582e7e8305bee4ba525bdb57a57;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h20f3170404511792e290715180d7eaf8ef697ab6b49c22f93;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9d334826e74e181a1a10d643bec62cb8e259f6ab1c1d83005;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2e9e4417e2a9a1d62416eef98a2407b62974c1918f41e2313;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'haddfbb01cd84497d24d2cd3e1aa0a5fef0f607c833ae3e688;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h321d85aefdabd87c13b18ddc227a71ff50e090b1ba7fde4eb;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdc4ce0fd57ce9565356be5733db6aabda34818d3a90a9be1d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb879a4dd0b39c4f681d4ed39ac613e1395754935c01cd9fd5;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc7a517175a4f5f9ceda1bb62d9f2d45c0b93447f1b3ff916;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h276c7e1f56a8bdc285a806e24f1bad714bb9e435b487063ea;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5ecc6ce28dc0517c43f7a17fe16e9157c51df34b5e43d6baa;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc9657714d36eab4c88e163a21eb89ce47165cf326a2a3d270;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hef63c1130db3a5cc6963855b9e8d83dac715a7728775d9ed1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2a9b359bf0358ecb30a1b85ba02765a311847d2d7d1962228;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h28b1d482265be0b2ba7f1190919662816ed01a64e69076af6;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h17be818585cc1546edcdc17d30798d222aa6044ca4a849c7c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h59111c441cd32bcdf60a677ee9f411e1559f8697fe26c49d7;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h328442afb788eff5aa05b8bfe009e570fd49c0956b6d8253f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h710854bc510d8ab86dfc6282b7c6287c6b7de0e2e7af4b546;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he99c3a47dbacf0148509108ea461f743c20b70dfaa764e4c1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfa209bf2405b3fb1863db44b496a076103b9c429c46ea27ea;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h727517d0f7792c3250e27d1a009de2f5e335ea8d6dd1b6c26;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbbadd535b140acefb393719aaf1c36504bd22e50bff0c1d4;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8476f5d8081cc8d2e9bc994fcf26cd90e6529d1a48bf5a535;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h67cef47e66a6be1d278fe2924af974b573ac20ef46884175d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h50e2664593fa53c2524da521088bfc170f5e785906a9d3198;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7caf9196f257798882c5307777ea1bde1ce8f0f59b3c22f48;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3c542930f79ac57a39dc77d74aa60c7fa182b3ea43bec3c43;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2266a7791f0d925c9f0a2150a6b993e6c1bf40617802ddc4e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h41ca2b904adbda3acdb2d349335f135850c7d7f7f0823937;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3fae650d60f42a92cf9f5c6059024c5dec664a069616fee5c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he167c66b2775dbaa0da21dad0418412b89c577e5bf697692;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb1b8bcb2fbdd3db2006e2dd9dee33ac28546cbb2c8f90132c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h94df9799099a1937969d25b9abde50df8c63f84cf6e880e47;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3a9bfc5f28a066c1e7c8662d430dd433e65358a40f0466ac7;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfce8534fb2f2239552b3fd1ec11a22b56d4f61ec8d9b79394;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he7bfc4a08773512439648d163426042bf4b85f63516af22cd;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3eee421c1a192e072e72559b18ce3d3cbc89e0256ad5d6f18;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha6642a769a0ae4bb9e96a7e2be16736afa6f4611e020a9085;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1183555fd37624a2addc6e5e145619377de5392866dd734b8;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd919a8f203cc707ab125baf053c337b0c206f93593eec9bf;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h973db79606d849620391bb9e346c86a510a39e52149756a0a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h28ef49bd4ea9b0c66f849ecbffa3fdd0f799cd6d5ca080d8d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2cbe679e3f75df1357d1ea551c9b75c5d635821a3dde3e39a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb0404d26f4aa833000dcf5e62cbf49f04c8049ef5e3c47410;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5963e682d03802c88c27c923b9952a5f61f8fce8689faa804;
        #1
        $finish();
    end
endmodule
