module shift_register(
        input wire clk,
        input wire src0_,
        input wire src1_,
        input wire src2_,
        input wire src3_,
        input wire src4_,
        input wire src5_,
        input wire src6_,
        input wire src7_,
        input wire src8_,
        input wire src9_,
        input wire src10_,
        input wire src11_,
        input wire src12_,
        input wire src13_,
        input wire src14_,
        input wire src15_,
        output wire [0:0] dst0,
        output wire [0:0] dst1,
        output wire [0:0] dst2,
        output wire [0:0] dst3,
        output wire [0:0] dst4,
        output wire [0:0] dst5,
        output wire [0:0] dst6,
        output wire [0:0] dst7,
        output wire [0:0] dst8,
        output wire [0:0] dst9,
        output wire [0:0] dst10,
        output wire [0:0] dst11,
        output wire [0:0] dst12,
        output wire [0:0] dst13,
        output wire [0:0] dst14,
        output wire [0:0] dst15,
        output wire [0:0] dst16,
        output wire [0:0] dst17,
        output wire [0:0] dst18,
        output wire [0:0] dst19,
        output wire [0:0] dst20,
        output wire [0:0] dst21);
    reg [53:0] src0;
    reg [53:0] src1;
    reg [53:0] src2;
    reg [53:0] src3;
    reg [53:0] src4;
    reg [53:0] src5;
    reg [53:0] src6;
    reg [53:0] src7;
    reg [53:0] src8;
    reg [53:0] src9;
    reg [53:0] src10;
    reg [53:0] src11;
    reg [53:0] src12;
    reg [53:0] src13;
    reg [53:0] src14;
    reg [53:0] src15;
    compressor2_1_54_16 compressor2_1_54_16(
            .src0(src0),
            .src1(src1),
            .src2(src2),
            .src3(src3),
            .src4(src4),
            .src5(src5),
            .src6(src6),
            .src7(src7),
            .src8(src8),
            .src9(src9),
            .src10(src10),
            .src11(src11),
            .src12(src12),
            .src13(src13),
            .src14(src14),
            .src15(src15),
            .dst0(dst0),
            .dst1(dst1),
            .dst2(dst2),
            .dst3(dst3),
            .dst4(dst4),
            .dst5(dst5),
            .dst6(dst6),
            .dst7(dst7),
            .dst8(dst8),
            .dst9(dst9),
            .dst10(dst10),
            .dst11(dst11),
            .dst12(dst12),
            .dst13(dst13),
            .dst14(dst14),
            .dst15(dst15),
            .dst16(dst16),
            .dst17(dst17),
            .dst18(dst18),
            .dst19(dst19),
            .dst20(dst20),
            .dst21(dst21));
    initial begin
        src0 <= 54'h0;
        src1 <= 54'h0;
        src2 <= 54'h0;
        src3 <= 54'h0;
        src4 <= 54'h0;
        src5 <= 54'h0;
        src6 <= 54'h0;
        src7 <= 54'h0;
        src8 <= 54'h0;
        src9 <= 54'h0;
        src10 <= 54'h0;
        src11 <= 54'h0;
        src12 <= 54'h0;
        src13 <= 54'h0;
        src14 <= 54'h0;
        src15 <= 54'h0;
    end
    always @(posedge clk) begin
        src0 <= {src0, src0_};
        src1 <= {src1, src1_};
        src2 <= {src2, src2_};
        src3 <= {src3, src3_};
        src4 <= {src4, src4_};
        src5 <= {src5, src5_};
        src6 <= {src6, src6_};
        src7 <= {src7, src7_};
        src8 <= {src8, src8_};
        src9 <= {src9, src9_};
        src10 <= {src10, src10_};
        src11 <= {src11, src11_};
        src12 <= {src12, src12_};
        src13 <= {src13, src13_};
        src14 <= {src14, src14_};
        src15 <= {src15, src15_};
    end
endmodule
module compressor2_1_54_16(
    input [53:0]src0,
    input [53:0]src1,
    input [53:0]src2,
    input [53:0]src3,
    input [53:0]src4,
    input [53:0]src5,
    input [53:0]src6,
    input [53:0]src7,
    input [53:0]src8,
    input [53:0]src9,
    input [53:0]src10,
    input [53:0]src11,
    input [53:0]src12,
    input [53:0]src13,
    input [53:0]src14,
    input [53:0]src15,
    output dst0,
    output dst1,
    output dst2,
    output dst3,
    output dst4,
    output dst5,
    output dst6,
    output dst7,
    output dst8,
    output dst9,
    output dst10,
    output dst11,
    output dst12,
    output dst13,
    output dst14,
    output dst15,
    output dst16,
    output dst17,
    output dst18,
    output dst19,
    output dst20,
    output dst21);

    wire [1:0] comp_out0;
    wire [1:0] comp_out1;
    wire [1:0] comp_out2;
    wire [1:0] comp_out3;
    wire [1:0] comp_out4;
    wire [1:0] comp_out5;
    wire [1:0] comp_out6;
    wire [1:0] comp_out7;
    wire [1:0] comp_out8;
    wire [1:0] comp_out9;
    wire [1:0] comp_out10;
    wire [1:0] comp_out11;
    wire [1:0] comp_out12;
    wire [1:0] comp_out13;
    wire [1:0] comp_out14;
    wire [1:0] comp_out15;
    wire [1:0] comp_out16;
    wire [1:0] comp_out17;
    wire [1:0] comp_out18;
    wire [1:0] comp_out19;
    wire [0:0] comp_out20;
    wire [1:0] comp_out21;
    compressor compressor_inst(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .dst0(comp_out0),
        .dst1(comp_out1),
        .dst2(comp_out2),
        .dst3(comp_out3),
        .dst4(comp_out4),
        .dst5(comp_out5),
        .dst6(comp_out6),
        .dst7(comp_out7),
        .dst8(comp_out8),
        .dst9(comp_out9),
        .dst10(comp_out10),
        .dst11(comp_out11),
        .dst12(comp_out12),
        .dst13(comp_out13),
        .dst14(comp_out14),
        .dst15(comp_out15),
        .dst16(comp_out16),
        .dst17(comp_out17),
        .dst18(comp_out18),
        .dst19(comp_out19),
        .dst20(comp_out20),
        .dst21(comp_out21)
    );
    rowadder2_1_22 rowadder2_1inst(
        .src0({comp_out21[0], comp_out20[0], comp_out19[0], comp_out18[0], comp_out17[0], comp_out16[0], comp_out15[0], comp_out14[0], comp_out13[0], comp_out12[0], comp_out11[0], comp_out10[0], comp_out9[0], comp_out8[0], comp_out7[0], comp_out6[0], comp_out5[0], comp_out4[0], comp_out3[0], comp_out2[0], comp_out1[0], comp_out0[0]}),
        .src1({comp_out21[1], 1'h0, comp_out19[1], comp_out18[1], comp_out17[1], comp_out16[1], comp_out15[1], comp_out14[1], comp_out13[1], comp_out12[1], comp_out11[1], comp_out10[1], comp_out9[1], comp_out8[1], comp_out7[1], comp_out6[1], comp_out5[1], comp_out4[1], comp_out3[1], comp_out2[1], comp_out1[1], comp_out0[1]}),
        .dst0({dst21, dst20, dst19, dst18, dst17, dst16, dst15, dst14, dst13, dst12, dst11, dst10, dst9, dst8, dst7, dst6, dst5, dst4, dst3, dst2, dst1, dst0})
    );
endmodule
module compressor (
      input wire [53:0] src0,
      input wire [53:0] src1,
      input wire [53:0] src2,
      input wire [53:0] src3,
      input wire [53:0] src4,
      input wire [53:0] src5,
      input wire [53:0] src6,
      input wire [53:0] src7,
      input wire [53:0] src8,
      input wire [53:0] src9,
      input wire [53:0] src10,
      input wire [53:0] src11,
      input wire [53:0] src12,
      input wire [53:0] src13,
      input wire [53:0] src14,
      input wire [53:0] src15,
      output wire [1:0] dst0,
      output wire [1:0] dst1,
      output wire [1:0] dst2,
      output wire [1:0] dst3,
      output wire [1:0] dst4,
      output wire [1:0] dst5,
      output wire [1:0] dst6,
      output wire [1:0] dst7,
      output wire [1:0] dst8,
      output wire [1:0] dst9,
      output wire [1:0] dst10,
      output wire [1:0] dst11,
      output wire [1:0] dst12,
      output wire [1:0] dst13,
      output wire [1:0] dst14,
      output wire [1:0] dst15,
      output wire [1:0] dst16,
      output wire [1:0] dst17,
      output wire [1:0] dst18,
      output wire [1:0] dst19,
      output wire [0:0] dst20,
      output wire [1:0] dst21);

   wire [53:0] stage0_0;
   wire [53:0] stage0_1;
   wire [53:0] stage0_2;
   wire [53:0] stage0_3;
   wire [53:0] stage0_4;
   wire [53:0] stage0_5;
   wire [53:0] stage0_6;
   wire [53:0] stage0_7;
   wire [53:0] stage0_8;
   wire [53:0] stage0_9;
   wire [53:0] stage0_10;
   wire [53:0] stage0_11;
   wire [53:0] stage0_12;
   wire [53:0] stage0_13;
   wire [53:0] stage0_14;
   wire [53:0] stage0_15;
   wire [13:0] stage1_0;
   wire [16:0] stage1_1;
   wire [22:0] stage1_2;
   wire [17:0] stage1_3;
   wire [34:0] stage1_4;
   wire [24:0] stage1_5;
   wire [18:0] stage1_6;
   wire [18:0] stage1_7;
   wire [25:0] stage1_8;
   wire [26:0] stage1_9;
   wire [18:0] stage1_10;
   wire [17:0] stage1_11;
   wire [25:0] stage1_12;
   wire [25:0] stage1_13;
   wire [17:0] stage1_14;
   wire [23:0] stage1_15;
   wire [16:0] stage1_16;
   wire [7:0] stage1_17;
   wire [7:0] stage2_0;
   wire [2:0] stage2_1;
   wire [7:0] stage2_2;
   wire [8:0] stage2_3;
   wire [11:0] stage2_4;
   wire [9:0] stage2_5;
   wire [11:0] stage2_6;
   wire [10:0] stage2_7;
   wire [7:0] stage2_8;
   wire [11:0] stage2_9;
   wire [12:0] stage2_10;
   wire [6:0] stage2_11;
   wire [8:0] stage2_12;
   wire [10:0] stage2_13;
   wire [8:0] stage2_14;
   wire [7:0] stage2_15;
   wire [9:0] stage2_16;
   wire [6:0] stage2_17;
   wire [2:0] stage2_18;
   wire [2:0] stage2_19;
   wire [0:0] stage2_20;
   wire [1:0] stage3_0;
   wire [1:0] stage3_1;
   wire [1:0] stage3_2;
   wire [5:0] stage3_3;
   wire [3:0] stage3_4;
   wire [5:0] stage3_5;
   wire [2:0] stage3_6;
   wire [5:0] stage3_7;
   wire [4:0] stage3_8;
   wire [2:0] stage3_9;
   wire [3:0] stage3_10;
   wire [5:0] stage3_11;
   wire [5:0] stage3_12;
   wire [2:0] stage3_13;
   wire [2:0] stage3_14;
   wire [3:0] stage3_15;
   wire [5:0] stage3_16;
   wire [3:0] stage3_17;
   wire [3:0] stage3_18;
   wire [0:0] stage3_19;
   wire [0:0] stage3_20;
   wire [0:0] stage3_21;
   wire [1:0] stage4_0;
   wire [1:0] stage4_1;
   wire [1:0] stage4_2;
   wire [1:0] stage4_3;
   wire [1:0] stage4_4;
   wire [1:0] stage4_5;
   wire [1:0] stage4_6;
   wire [1:0] stage4_7;
   wire [1:0] stage4_8;
   wire [1:0] stage4_9;
   wire [1:0] stage4_10;
   wire [1:0] stage4_11;
   wire [1:0] stage4_12;
   wire [1:0] stage4_13;
   wire [1:0] stage4_14;
   wire [1:0] stage4_15;
   wire [1:0] stage4_16;
   wire [1:0] stage4_17;
   wire [1:0] stage4_18;
   wire [1:0] stage4_19;
   wire [0:0] stage4_20;
   wire [1:0] stage4_21;

   assign stage0_0 = src0;
   assign stage0_1 = src1;
   assign stage0_2 = src2;
   assign stage0_3 = src3;
   assign stage0_4 = src4;
   assign stage0_5 = src5;
   assign stage0_6 = src6;
   assign stage0_7 = src7;
   assign stage0_8 = src8;
   assign stage0_9 = src9;
   assign stage0_10 = src10;
   assign stage0_11 = src11;
   assign stage0_12 = src12;
   assign stage0_13 = src13;
   assign stage0_14 = src14;
   assign stage0_15 = src15;
   assign dst0 = stage4_0;
   assign dst1 = stage4_1;
   assign dst2 = stage4_2;
   assign dst3 = stage4_3;
   assign dst4 = stage4_4;
   assign dst5 = stage4_5;
   assign dst6 = stage4_6;
   assign dst7 = stage4_7;
   assign dst8 = stage4_8;
   assign dst9 = stage4_9;
   assign dst10 = stage4_10;
   assign dst11 = stage4_11;
   assign dst12 = stage4_12;
   assign dst13 = stage4_13;
   assign dst14 = stage4_14;
   assign dst15 = stage4_15;
   assign dst16 = stage4_16;
   assign dst17 = stage4_17;
   assign dst18 = stage4_18;
   assign dst19 = stage4_19;
   assign dst20 = stage4_20;
   assign dst21 = stage4_21;

   gpc606_5 gpc0 (
      {stage0_0[0], stage0_0[1], stage0_0[2], stage0_0[3], stage0_0[4], stage0_0[5]},
      {stage0_2[0], stage0_2[1], stage0_2[2], stage0_2[3], stage0_2[4], stage0_2[5]},
      {stage1_4[0],stage1_3[0],stage1_2[0],stage1_1[0],stage1_0[0]}
   );
   gpc606_5 gpc1 (
      {stage0_0[6], stage0_0[7], stage0_0[8], stage0_0[9], stage0_0[10], stage0_0[11]},
      {stage0_2[6], stage0_2[7], stage0_2[8], stage0_2[9], stage0_2[10], stage0_2[11]},
      {stage1_4[1],stage1_3[1],stage1_2[1],stage1_1[1],stage1_0[1]}
   );
   gpc606_5 gpc2 (
      {stage0_0[12], stage0_0[13], stage0_0[14], stage0_0[15], stage0_0[16], stage0_0[17]},
      {stage0_2[12], stage0_2[13], stage0_2[14], stage0_2[15], stage0_2[16], stage0_2[17]},
      {stage1_4[2],stage1_3[2],stage1_2[2],stage1_1[2],stage1_0[2]}
   );
   gpc606_5 gpc3 (
      {stage0_0[18], stage0_0[19], stage0_0[20], stage0_0[21], stage0_0[22], stage0_0[23]},
      {stage0_2[18], stage0_2[19], stage0_2[20], stage0_2[21], stage0_2[22], stage0_2[23]},
      {stage1_4[3],stage1_3[3],stage1_2[3],stage1_1[3],stage1_0[3]}
   );
   gpc606_5 gpc4 (
      {stage0_0[24], stage0_0[25], stage0_0[26], stage0_0[27], stage0_0[28], stage0_0[29]},
      {stage0_2[24], stage0_2[25], stage0_2[26], stage0_2[27], stage0_2[28], stage0_2[29]},
      {stage1_4[4],stage1_3[4],stage1_2[4],stage1_1[4],stage1_0[4]}
   );
   gpc606_5 gpc5 (
      {stage0_0[30], stage0_0[31], stage0_0[32], stage0_0[33], stage0_0[34], stage0_0[35]},
      {stage0_2[30], stage0_2[31], stage0_2[32], stage0_2[33], stage0_2[34], stage0_2[35]},
      {stage1_4[5],stage1_3[5],stage1_2[5],stage1_1[5],stage1_0[5]}
   );
   gpc606_5 gpc6 (
      {stage0_0[36], stage0_0[37], stage0_0[38], stage0_0[39], stage0_0[40], stage0_0[41]},
      {stage0_2[36], stage0_2[37], stage0_2[38], stage0_2[39], stage0_2[40], stage0_2[41]},
      {stage1_4[6],stage1_3[6],stage1_2[6],stage1_1[6],stage1_0[6]}
   );
   gpc606_5 gpc7 (
      {stage0_0[42], stage0_0[43], stage0_0[44], stage0_0[45], stage0_0[46], stage0_0[47]},
      {stage0_2[42], stage0_2[43], stage0_2[44], stage0_2[45], stage0_2[46], stage0_2[47]},
      {stage1_4[7],stage1_3[7],stage1_2[7],stage1_1[7],stage1_0[7]}
   );
   gpc1406_5 gpc8 (
      {stage0_1[0], stage0_1[1], stage0_1[2], stage0_1[3], stage0_1[4], stage0_1[5]},
      {stage0_3[0], stage0_3[1], stage0_3[2], stage0_3[3]},
      {stage0_4[0]},
      {stage1_5[0],stage1_4[8],stage1_3[8],stage1_2[8],stage1_1[8]}
   );
   gpc1406_5 gpc9 (
      {stage0_1[6], stage0_1[7], stage0_1[8], stage0_1[9], stage0_1[10], stage0_1[11]},
      {stage0_3[4], stage0_3[5], stage0_3[6], stage0_3[7]},
      {stage0_4[1]},
      {stage1_5[1],stage1_4[9],stage1_3[9],stage1_2[9],stage1_1[9]}
   );
   gpc606_5 gpc10 (
      {stage0_1[12], stage0_1[13], stage0_1[14], stage0_1[15], stage0_1[16], stage0_1[17]},
      {stage0_3[8], stage0_3[9], stage0_3[10], stage0_3[11], stage0_3[12], stage0_3[13]},
      {stage1_5[2],stage1_4[10],stage1_3[10],stage1_2[10],stage1_1[10]}
   );
   gpc606_5 gpc11 (
      {stage0_1[18], stage0_1[19], stage0_1[20], stage0_1[21], stage0_1[22], stage0_1[23]},
      {stage0_3[14], stage0_3[15], stage0_3[16], stage0_3[17], stage0_3[18], stage0_3[19]},
      {stage1_5[3],stage1_4[11],stage1_3[11],stage1_2[11],stage1_1[11]}
   );
   gpc606_5 gpc12 (
      {stage0_1[24], stage0_1[25], stage0_1[26], stage0_1[27], stage0_1[28], stage0_1[29]},
      {stage0_3[20], stage0_3[21], stage0_3[22], stage0_3[23], stage0_3[24], stage0_3[25]},
      {stage1_5[4],stage1_4[12],stage1_3[12],stage1_2[12],stage1_1[12]}
   );
   gpc606_5 gpc13 (
      {stage0_1[30], stage0_1[31], stage0_1[32], stage0_1[33], stage0_1[34], stage0_1[35]},
      {stage0_3[26], stage0_3[27], stage0_3[28], stage0_3[29], stage0_3[30], stage0_3[31]},
      {stage1_5[5],stage1_4[13],stage1_3[13],stage1_2[13],stage1_1[13]}
   );
   gpc606_5 gpc14 (
      {stage0_1[36], stage0_1[37], stage0_1[38], stage0_1[39], stage0_1[40], stage0_1[41]},
      {stage0_3[32], stage0_3[33], stage0_3[34], stage0_3[35], stage0_3[36], stage0_3[37]},
      {stage1_5[6],stage1_4[14],stage1_3[14],stage1_2[14],stage1_1[14]}
   );
   gpc606_5 gpc15 (
      {stage0_1[42], stage0_1[43], stage0_1[44], stage0_1[45], stage0_1[46], stage0_1[47]},
      {stage0_3[38], stage0_3[39], stage0_3[40], stage0_3[41], stage0_3[42], stage0_3[43]},
      {stage1_5[7],stage1_4[15],stage1_3[15],stage1_2[15],stage1_1[15]}
   );
   gpc606_5 gpc16 (
      {stage0_1[48], stage0_1[49], stage0_1[50], stage0_1[51], stage0_1[52], stage0_1[53]},
      {stage0_3[44], stage0_3[45], stage0_3[46], stage0_3[47], stage0_3[48], stage0_3[49]},
      {stage1_5[8],stage1_4[16],stage1_3[16],stage1_2[16],stage1_1[16]}
   );
   gpc615_5 gpc17 (
      {stage0_3[50], stage0_3[51], stage0_3[52], stage0_3[53], 1'b0},
      {stage0_4[2]},
      {stage0_5[0], stage0_5[1], stage0_5[2], stage0_5[3], stage0_5[4], stage0_5[5]},
      {stage1_7[0],stage1_6[0],stage1_5[9],stage1_4[17],stage1_3[17]}
   );
   gpc606_5 gpc18 (
      {stage0_4[3], stage0_4[4], stage0_4[5], stage0_4[6], stage0_4[7], stage0_4[8]},
      {stage0_6[0], stage0_6[1], stage0_6[2], stage0_6[3], stage0_6[4], stage0_6[5]},
      {stage1_8[0],stage1_7[1],stage1_6[1],stage1_5[10],stage1_4[18]}
   );
   gpc606_5 gpc19 (
      {stage0_4[9], stage0_4[10], stage0_4[11], stage0_4[12], stage0_4[13], stage0_4[14]},
      {stage0_6[6], stage0_6[7], stage0_6[8], stage0_6[9], stage0_6[10], stage0_6[11]},
      {stage1_8[1],stage1_7[2],stage1_6[2],stage1_5[11],stage1_4[19]}
   );
   gpc606_5 gpc20 (
      {stage0_4[15], stage0_4[16], stage0_4[17], stage0_4[18], stage0_4[19], stage0_4[20]},
      {stage0_6[12], stage0_6[13], stage0_6[14], stage0_6[15], stage0_6[16], stage0_6[17]},
      {stage1_8[2],stage1_7[3],stage1_6[3],stage1_5[12],stage1_4[20]}
   );
   gpc606_5 gpc21 (
      {stage0_4[21], stage0_4[22], stage0_4[23], stage0_4[24], stage0_4[25], stage0_4[26]},
      {stage0_6[18], stage0_6[19], stage0_6[20], stage0_6[21], stage0_6[22], stage0_6[23]},
      {stage1_8[3],stage1_7[4],stage1_6[4],stage1_5[13],stage1_4[21]}
   );
   gpc606_5 gpc22 (
      {stage0_4[27], stage0_4[28], stage0_4[29], stage0_4[30], stage0_4[31], stage0_4[32]},
      {stage0_6[24], stage0_6[25], stage0_6[26], stage0_6[27], stage0_6[28], stage0_6[29]},
      {stage1_8[4],stage1_7[5],stage1_6[5],stage1_5[14],stage1_4[22]}
   );
   gpc606_5 gpc23 (
      {stage0_4[33], stage0_4[34], stage0_4[35], stage0_4[36], stage0_4[37], stage0_4[38]},
      {stage0_6[30], stage0_6[31], stage0_6[32], stage0_6[33], stage0_6[34], stage0_6[35]},
      {stage1_8[5],stage1_7[6],stage1_6[6],stage1_5[15],stage1_4[23]}
   );
   gpc615_5 gpc24 (
      {stage0_4[39], stage0_4[40], stage0_4[41], stage0_4[42], stage0_4[43]},
      {stage0_5[6]},
      {stage0_6[36], stage0_6[37], stage0_6[38], stage0_6[39], stage0_6[40], stage0_6[41]},
      {stage1_8[6],stage1_7[7],stage1_6[7],stage1_5[16],stage1_4[24]}
   );
   gpc606_5 gpc25 (
      {stage0_5[7], stage0_5[8], stage0_5[9], stage0_5[10], stage0_5[11], stage0_5[12]},
      {stage0_7[0], stage0_7[1], stage0_7[2], stage0_7[3], stage0_7[4], stage0_7[5]},
      {stage1_9[0],stage1_8[7],stage1_7[8],stage1_6[8],stage1_5[17]}
   );
   gpc606_5 gpc26 (
      {stage0_5[13], stage0_5[14], stage0_5[15], stage0_5[16], stage0_5[17], stage0_5[18]},
      {stage0_7[6], stage0_7[7], stage0_7[8], stage0_7[9], stage0_7[10], stage0_7[11]},
      {stage1_9[1],stage1_8[8],stage1_7[9],stage1_6[9],stage1_5[18]}
   );
   gpc606_5 gpc27 (
      {stage0_5[19], stage0_5[20], stage0_5[21], stage0_5[22], stage0_5[23], stage0_5[24]},
      {stage0_7[12], stage0_7[13], stage0_7[14], stage0_7[15], stage0_7[16], stage0_7[17]},
      {stage1_9[2],stage1_8[9],stage1_7[10],stage1_6[10],stage1_5[19]}
   );
   gpc606_5 gpc28 (
      {stage0_5[25], stage0_5[26], stage0_5[27], stage0_5[28], stage0_5[29], stage0_5[30]},
      {stage0_7[18], stage0_7[19], stage0_7[20], stage0_7[21], stage0_7[22], stage0_7[23]},
      {stage1_9[3],stage1_8[10],stage1_7[11],stage1_6[11],stage1_5[20]}
   );
   gpc606_5 gpc29 (
      {stage0_5[31], stage0_5[32], stage0_5[33], stage0_5[34], stage0_5[35], stage0_5[36]},
      {stage0_7[24], stage0_7[25], stage0_7[26], stage0_7[27], stage0_7[28], stage0_7[29]},
      {stage1_9[4],stage1_8[11],stage1_7[12],stage1_6[12],stage1_5[21]}
   );
   gpc606_5 gpc30 (
      {stage0_5[37], stage0_5[38], stage0_5[39], stage0_5[40], stage0_5[41], stage0_5[42]},
      {stage0_7[30], stage0_7[31], stage0_7[32], stage0_7[33], stage0_7[34], stage0_7[35]},
      {stage1_9[5],stage1_8[12],stage1_7[13],stage1_6[13],stage1_5[22]}
   );
   gpc606_5 gpc31 (
      {stage0_5[43], stage0_5[44], stage0_5[45], stage0_5[46], stage0_5[47], stage0_5[48]},
      {stage0_7[36], stage0_7[37], stage0_7[38], stage0_7[39], stage0_7[40], stage0_7[41]},
      {stage1_9[6],stage1_8[13],stage1_7[14],stage1_6[14],stage1_5[23]}
   );
   gpc615_5 gpc32 (
      {stage0_5[49], stage0_5[50], stage0_5[51], stage0_5[52], stage0_5[53]},
      {stage0_6[42]},
      {stage0_7[42], stage0_7[43], stage0_7[44], stage0_7[45], stage0_7[46], stage0_7[47]},
      {stage1_9[7],stage1_8[14],stage1_7[15],stage1_6[15],stage1_5[24]}
   );
   gpc615_5 gpc33 (
      {stage0_6[43], stage0_6[44], stage0_6[45], stage0_6[46], stage0_6[47]},
      {stage0_7[48]},
      {stage0_8[0], stage0_8[1], stage0_8[2], stage0_8[3], stage0_8[4], stage0_8[5]},
      {stage1_10[0],stage1_9[8],stage1_8[15],stage1_7[16],stage1_6[16]}
   );
   gpc615_5 gpc34 (
      {stage0_6[48], stage0_6[49], stage0_6[50], stage0_6[51], stage0_6[52]},
      {stage0_7[49]},
      {stage0_8[6], stage0_8[7], stage0_8[8], stage0_8[9], stage0_8[10], stage0_8[11]},
      {stage1_10[1],stage1_9[9],stage1_8[16],stage1_7[17],stage1_6[17]}
   );
   gpc615_5 gpc35 (
      {stage0_7[50], stage0_7[51], stage0_7[52], stage0_7[53], 1'b0},
      {stage0_8[12]},
      {stage0_9[0], stage0_9[1], stage0_9[2], stage0_9[3], stage0_9[4], stage0_9[5]},
      {stage1_11[0],stage1_10[2],stage1_9[10],stage1_8[17],stage1_7[18]}
   );
   gpc606_5 gpc36 (
      {stage0_8[13], stage0_8[14], stage0_8[15], stage0_8[16], stage0_8[17], stage0_8[18]},
      {stage0_10[0], stage0_10[1], stage0_10[2], stage0_10[3], stage0_10[4], stage0_10[5]},
      {stage1_12[0],stage1_11[1],stage1_10[3],stage1_9[11],stage1_8[18]}
   );
   gpc615_5 gpc37 (
      {stage0_8[19], stage0_8[20], stage0_8[21], stage0_8[22], stage0_8[23]},
      {stage0_9[6]},
      {stage0_10[6], stage0_10[7], stage0_10[8], stage0_10[9], stage0_10[10], stage0_10[11]},
      {stage1_12[1],stage1_11[2],stage1_10[4],stage1_9[12],stage1_8[19]}
   );
   gpc615_5 gpc38 (
      {stage0_8[24], stage0_8[25], stage0_8[26], stage0_8[27], stage0_8[28]},
      {stage0_9[7]},
      {stage0_10[12], stage0_10[13], stage0_10[14], stage0_10[15], stage0_10[16], stage0_10[17]},
      {stage1_12[2],stage1_11[3],stage1_10[5],stage1_9[13],stage1_8[20]}
   );
   gpc615_5 gpc39 (
      {stage0_8[29], stage0_8[30], stage0_8[31], stage0_8[32], stage0_8[33]},
      {stage0_9[8]},
      {stage0_10[18], stage0_10[19], stage0_10[20], stage0_10[21], stage0_10[22], stage0_10[23]},
      {stage1_12[3],stage1_11[4],stage1_10[6],stage1_9[14],stage1_8[21]}
   );
   gpc615_5 gpc40 (
      {stage0_8[34], stage0_8[35], stage0_8[36], stage0_8[37], stage0_8[38]},
      {stage0_9[9]},
      {stage0_10[24], stage0_10[25], stage0_10[26], stage0_10[27], stage0_10[28], stage0_10[29]},
      {stage1_12[4],stage1_11[5],stage1_10[7],stage1_9[15],stage1_8[22]}
   );
   gpc615_5 gpc41 (
      {stage0_8[39], stage0_8[40], stage0_8[41], stage0_8[42], stage0_8[43]},
      {stage0_9[10]},
      {stage0_10[30], stage0_10[31], stage0_10[32], stage0_10[33], stage0_10[34], stage0_10[35]},
      {stage1_12[5],stage1_11[6],stage1_10[8],stage1_9[16],stage1_8[23]}
   );
   gpc615_5 gpc42 (
      {stage0_8[44], stage0_8[45], stage0_8[46], stage0_8[47], stage0_8[48]},
      {stage0_9[11]},
      {stage0_10[36], stage0_10[37], stage0_10[38], stage0_10[39], stage0_10[40], stage0_10[41]},
      {stage1_12[6],stage1_11[7],stage1_10[9],stage1_9[17],stage1_8[24]}
   );
   gpc615_5 gpc43 (
      {stage0_8[49], stage0_8[50], stage0_8[51], stage0_8[52], stage0_8[53]},
      {stage0_9[12]},
      {stage0_10[42], stage0_10[43], stage0_10[44], stage0_10[45], stage0_10[46], stage0_10[47]},
      {stage1_12[7],stage1_11[8],stage1_10[10],stage1_9[18],stage1_8[25]}
   );
   gpc606_5 gpc44 (
      {stage0_9[13], stage0_9[14], stage0_9[15], stage0_9[16], stage0_9[17], stage0_9[18]},
      {stage0_11[0], stage0_11[1], stage0_11[2], stage0_11[3], stage0_11[4], stage0_11[5]},
      {stage1_13[0],stage1_12[8],stage1_11[9],stage1_10[11],stage1_9[19]}
   );
   gpc606_5 gpc45 (
      {stage0_9[19], stage0_9[20], stage0_9[21], stage0_9[22], stage0_9[23], stage0_9[24]},
      {stage0_11[6], stage0_11[7], stage0_11[8], stage0_11[9], stage0_11[10], stage0_11[11]},
      {stage1_13[1],stage1_12[9],stage1_11[10],stage1_10[12],stage1_9[20]}
   );
   gpc615_5 gpc46 (
      {stage0_9[25], stage0_9[26], stage0_9[27], stage0_9[28], stage0_9[29]},
      {stage0_10[48]},
      {stage0_11[12], stage0_11[13], stage0_11[14], stage0_11[15], stage0_11[16], stage0_11[17]},
      {stage1_13[2],stage1_12[10],stage1_11[11],stage1_10[13],stage1_9[21]}
   );
   gpc615_5 gpc47 (
      {stage0_9[30], stage0_9[31], stage0_9[32], stage0_9[33], stage0_9[34]},
      {stage0_10[49]},
      {stage0_11[18], stage0_11[19], stage0_11[20], stage0_11[21], stage0_11[22], stage0_11[23]},
      {stage1_13[3],stage1_12[11],stage1_11[12],stage1_10[14],stage1_9[22]}
   );
   gpc615_5 gpc48 (
      {stage0_9[35], stage0_9[36], stage0_9[37], stage0_9[38], stage0_9[39]},
      {stage0_10[50]},
      {stage0_11[24], stage0_11[25], stage0_11[26], stage0_11[27], stage0_11[28], stage0_11[29]},
      {stage1_13[4],stage1_12[12],stage1_11[13],stage1_10[15],stage1_9[23]}
   );
   gpc615_5 gpc49 (
      {stage0_9[40], stage0_9[41], stage0_9[42], stage0_9[43], stage0_9[44]},
      {stage0_10[51]},
      {stage0_11[30], stage0_11[31], stage0_11[32], stage0_11[33], stage0_11[34], stage0_11[35]},
      {stage1_13[5],stage1_12[13],stage1_11[14],stage1_10[16],stage1_9[24]}
   );
   gpc615_5 gpc50 (
      {stage0_9[45], stage0_9[46], stage0_9[47], stage0_9[48], stage0_9[49]},
      {stage0_10[52]},
      {stage0_11[36], stage0_11[37], stage0_11[38], stage0_11[39], stage0_11[40], stage0_11[41]},
      {stage1_13[6],stage1_12[14],stage1_11[15],stage1_10[17],stage1_9[25]}
   );
   gpc615_5 gpc51 (
      {stage0_9[50], stage0_9[51], stage0_9[52], stage0_9[53], 1'b0},
      {stage0_10[53]},
      {stage0_11[42], stage0_11[43], stage0_11[44], stage0_11[45], stage0_11[46], stage0_11[47]},
      {stage1_13[7],stage1_12[15],stage1_11[16],stage1_10[18],stage1_9[26]}
   );
   gpc606_5 gpc52 (
      {stage0_11[48], stage0_11[49], stage0_11[50], stage0_11[51], stage0_11[52], stage0_11[53]},
      {stage0_13[0], stage0_13[1], stage0_13[2], stage0_13[3], stage0_13[4], stage0_13[5]},
      {stage1_15[0],stage1_14[0],stage1_13[8],stage1_12[16],stage1_11[17]}
   );
   gpc606_5 gpc53 (
      {stage0_12[0], stage0_12[1], stage0_12[2], stage0_12[3], stage0_12[4], stage0_12[5]},
      {stage0_14[0], stage0_14[1], stage0_14[2], stage0_14[3], stage0_14[4], stage0_14[5]},
      {stage1_16[0],stage1_15[1],stage1_14[1],stage1_13[9],stage1_12[17]}
   );
   gpc606_5 gpc54 (
      {stage0_12[6], stage0_12[7], stage0_12[8], stage0_12[9], stage0_12[10], stage0_12[11]},
      {stage0_14[6], stage0_14[7], stage0_14[8], stage0_14[9], stage0_14[10], stage0_14[11]},
      {stage1_16[1],stage1_15[2],stage1_14[2],stage1_13[10],stage1_12[18]}
   );
   gpc606_5 gpc55 (
      {stage0_12[12], stage0_12[13], stage0_12[14], stage0_12[15], stage0_12[16], stage0_12[17]},
      {stage0_14[12], stage0_14[13], stage0_14[14], stage0_14[15], stage0_14[16], stage0_14[17]},
      {stage1_16[2],stage1_15[3],stage1_14[3],stage1_13[11],stage1_12[19]}
   );
   gpc606_5 gpc56 (
      {stage0_12[18], stage0_12[19], stage0_12[20], stage0_12[21], stage0_12[22], stage0_12[23]},
      {stage0_14[18], stage0_14[19], stage0_14[20], stage0_14[21], stage0_14[22], stage0_14[23]},
      {stage1_16[3],stage1_15[4],stage1_14[4],stage1_13[12],stage1_12[20]}
   );
   gpc606_5 gpc57 (
      {stage0_12[24], stage0_12[25], stage0_12[26], stage0_12[27], stage0_12[28], stage0_12[29]},
      {stage0_14[24], stage0_14[25], stage0_14[26], stage0_14[27], stage0_14[28], stage0_14[29]},
      {stage1_16[4],stage1_15[5],stage1_14[5],stage1_13[13],stage1_12[21]}
   );
   gpc606_5 gpc58 (
      {stage0_12[30], stage0_12[31], stage0_12[32], stage0_12[33], stage0_12[34], stage0_12[35]},
      {stage0_14[30], stage0_14[31], stage0_14[32], stage0_14[33], stage0_14[34], stage0_14[35]},
      {stage1_16[5],stage1_15[6],stage1_14[6],stage1_13[14],stage1_12[22]}
   );
   gpc606_5 gpc59 (
      {stage0_12[36], stage0_12[37], stage0_12[38], stage0_12[39], stage0_12[40], stage0_12[41]},
      {stage0_14[36], stage0_14[37], stage0_14[38], stage0_14[39], stage0_14[40], stage0_14[41]},
      {stage1_16[6],stage1_15[7],stage1_14[7],stage1_13[15],stage1_12[23]}
   );
   gpc606_5 gpc60 (
      {stage0_12[42], stage0_12[43], stage0_12[44], stage0_12[45], stage0_12[46], stage0_12[47]},
      {stage0_14[42], stage0_14[43], stage0_14[44], stage0_14[45], stage0_14[46], stage0_14[47]},
      {stage1_16[7],stage1_15[8],stage1_14[8],stage1_13[16],stage1_12[24]}
   );
   gpc606_5 gpc61 (
      {stage0_12[48], stage0_12[49], stage0_12[50], stage0_12[51], stage0_12[52], stage0_12[53]},
      {stage0_14[48], stage0_14[49], stage0_14[50], stage0_14[51], stage0_14[52], stage0_14[53]},
      {stage1_16[8],stage1_15[9],stage1_14[9],stage1_13[17],stage1_12[25]}
   );
   gpc606_5 gpc62 (
      {stage0_13[6], stage0_13[7], stage0_13[8], stage0_13[9], stage0_13[10], stage0_13[11]},
      {stage0_15[0], stage0_15[1], stage0_15[2], stage0_15[3], stage0_15[4], stage0_15[5]},
      {stage1_17[0],stage1_16[9],stage1_15[10],stage1_14[10],stage1_13[18]}
   );
   gpc606_5 gpc63 (
      {stage0_13[12], stage0_13[13], stage0_13[14], stage0_13[15], stage0_13[16], stage0_13[17]},
      {stage0_15[6], stage0_15[7], stage0_15[8], stage0_15[9], stage0_15[10], stage0_15[11]},
      {stage1_17[1],stage1_16[10],stage1_15[11],stage1_14[11],stage1_13[19]}
   );
   gpc606_5 gpc64 (
      {stage0_13[18], stage0_13[19], stage0_13[20], stage0_13[21], stage0_13[22], stage0_13[23]},
      {stage0_15[12], stage0_15[13], stage0_15[14], stage0_15[15], stage0_15[16], stage0_15[17]},
      {stage1_17[2],stage1_16[11],stage1_15[12],stage1_14[12],stage1_13[20]}
   );
   gpc606_5 gpc65 (
      {stage0_13[24], stage0_13[25], stage0_13[26], stage0_13[27], stage0_13[28], stage0_13[29]},
      {stage0_15[18], stage0_15[19], stage0_15[20], stage0_15[21], stage0_15[22], stage0_15[23]},
      {stage1_17[3],stage1_16[12],stage1_15[13],stage1_14[13],stage1_13[21]}
   );
   gpc606_5 gpc66 (
      {stage0_13[30], stage0_13[31], stage0_13[32], stage0_13[33], stage0_13[34], stage0_13[35]},
      {stage0_15[24], stage0_15[25], stage0_15[26], stage0_15[27], stage0_15[28], stage0_15[29]},
      {stage1_17[4],stage1_16[13],stage1_15[14],stage1_14[14],stage1_13[22]}
   );
   gpc606_5 gpc67 (
      {stage0_13[36], stage0_13[37], stage0_13[38], stage0_13[39], stage0_13[40], stage0_13[41]},
      {stage0_15[30], stage0_15[31], stage0_15[32], stage0_15[33], stage0_15[34], stage0_15[35]},
      {stage1_17[5],stage1_16[14],stage1_15[15],stage1_14[15],stage1_13[23]}
   );
   gpc606_5 gpc68 (
      {stage0_13[42], stage0_13[43], stage0_13[44], stage0_13[45], stage0_13[46], stage0_13[47]},
      {stage0_15[36], stage0_15[37], stage0_15[38], stage0_15[39], stage0_15[40], stage0_15[41]},
      {stage1_17[6],stage1_16[15],stage1_15[16],stage1_14[16],stage1_13[24]}
   );
   gpc606_5 gpc69 (
      {stage0_13[48], stage0_13[49], stage0_13[50], stage0_13[51], stage0_13[52], stage0_13[53]},
      {stage0_15[42], stage0_15[43], stage0_15[44], stage0_15[45], stage0_15[46], stage0_15[47]},
      {stage1_17[7],stage1_16[16],stage1_15[17],stage1_14[17],stage1_13[25]}
   );
   gpc1_1 gpc70 (
      {stage0_0[48]},
      {stage1_0[8]}
   );
   gpc1_1 gpc71 (
      {stage0_0[49]},
      {stage1_0[9]}
   );
   gpc1_1 gpc72 (
      {stage0_0[50]},
      {stage1_0[10]}
   );
   gpc1_1 gpc73 (
      {stage0_0[51]},
      {stage1_0[11]}
   );
   gpc1_1 gpc74 (
      {stage0_0[52]},
      {stage1_0[12]}
   );
   gpc1_1 gpc75 (
      {stage0_0[53]},
      {stage1_0[13]}
   );
   gpc1_1 gpc76 (
      {stage0_2[48]},
      {stage1_2[17]}
   );
   gpc1_1 gpc77 (
      {stage0_2[49]},
      {stage1_2[18]}
   );
   gpc1_1 gpc78 (
      {stage0_2[50]},
      {stage1_2[19]}
   );
   gpc1_1 gpc79 (
      {stage0_2[51]},
      {stage1_2[20]}
   );
   gpc1_1 gpc80 (
      {stage0_2[52]},
      {stage1_2[21]}
   );
   gpc1_1 gpc81 (
      {stage0_2[53]},
      {stage1_2[22]}
   );
   gpc1_1 gpc82 (
      {stage0_4[44]},
      {stage1_4[25]}
   );
   gpc1_1 gpc83 (
      {stage0_4[45]},
      {stage1_4[26]}
   );
   gpc1_1 gpc84 (
      {stage0_4[46]},
      {stage1_4[27]}
   );
   gpc1_1 gpc85 (
      {stage0_4[47]},
      {stage1_4[28]}
   );
   gpc1_1 gpc86 (
      {stage0_4[48]},
      {stage1_4[29]}
   );
   gpc1_1 gpc87 (
      {stage0_4[49]},
      {stage1_4[30]}
   );
   gpc1_1 gpc88 (
      {stage0_4[50]},
      {stage1_4[31]}
   );
   gpc1_1 gpc89 (
      {stage0_4[51]},
      {stage1_4[32]}
   );
   gpc1_1 gpc90 (
      {stage0_4[52]},
      {stage1_4[33]}
   );
   gpc1_1 gpc91 (
      {stage0_4[53]},
      {stage1_4[34]}
   );
   gpc1_1 gpc92 (
      {stage0_6[53]},
      {stage1_6[18]}
   );
   gpc1_1 gpc93 (
      {stage0_15[48]},
      {stage1_15[18]}
   );
   gpc1_1 gpc94 (
      {stage0_15[49]},
      {stage1_15[19]}
   );
   gpc1_1 gpc95 (
      {stage0_15[50]},
      {stage1_15[20]}
   );
   gpc1_1 gpc96 (
      {stage0_15[51]},
      {stage1_15[21]}
   );
   gpc1_1 gpc97 (
      {stage0_15[52]},
      {stage1_15[22]}
   );
   gpc1_1 gpc98 (
      {stage0_15[53]},
      {stage1_15[23]}
   );
   gpc1163_5 gpc99 (
      {stage1_0[0], stage1_0[1], stage1_0[2]},
      {stage1_1[0], stage1_1[1], stage1_1[2], stage1_1[3], stage1_1[4], stage1_1[5]},
      {stage1_2[0]},
      {stage1_3[0]},
      {stage2_4[0],stage2_3[0],stage2_2[0],stage2_1[0],stage2_0[0]}
   );
   gpc1163_5 gpc100 (
      {stage1_0[3], stage1_0[4], stage1_0[5]},
      {stage1_1[6], stage1_1[7], stage1_1[8], stage1_1[9], stage1_1[10], stage1_1[11]},
      {stage1_2[1]},
      {stage1_3[1]},
      {stage2_4[1],stage2_3[1],stage2_2[1],stage2_1[1],stage2_0[1]}
   );
   gpc1163_5 gpc101 (
      {stage1_0[6], stage1_0[7], stage1_0[8]},
      {stage1_1[12], stage1_1[13], stage1_1[14], stage1_1[15], stage1_1[16], 1'b0},
      {stage1_2[2]},
      {stage1_3[2]},
      {stage2_4[2],stage2_3[2],stage2_2[2],stage2_1[2],stage2_0[2]}
   );
   gpc606_5 gpc102 (
      {stage1_2[3], stage1_2[4], stage1_2[5], stage1_2[6], stage1_2[7], stage1_2[8]},
      {stage1_4[0], stage1_4[1], stage1_4[2], stage1_4[3], stage1_4[4], stage1_4[5]},
      {stage2_6[0],stage2_5[0],stage2_4[3],stage2_3[3],stage2_2[3]}
   );
   gpc606_5 gpc103 (
      {stage1_2[9], stage1_2[10], stage1_2[11], stage1_2[12], stage1_2[13], stage1_2[14]},
      {stage1_4[6], stage1_4[7], stage1_4[8], stage1_4[9], stage1_4[10], stage1_4[11]},
      {stage2_6[1],stage2_5[1],stage2_4[4],stage2_3[4],stage2_2[4]}
   );
   gpc606_5 gpc104 (
      {stage1_2[15], stage1_2[16], stage1_2[17], stage1_2[18], stage1_2[19], stage1_2[20]},
      {stage1_4[12], stage1_4[13], stage1_4[14], stage1_4[15], stage1_4[16], stage1_4[17]},
      {stage2_6[2],stage2_5[2],stage2_4[5],stage2_3[5],stage2_2[5]}
   );
   gpc615_5 gpc105 (
      {stage1_3[3], stage1_3[4], stage1_3[5], stage1_3[6], stage1_3[7]},
      {stage1_4[18]},
      {stage1_5[0], stage1_5[1], stage1_5[2], stage1_5[3], stage1_5[4], stage1_5[5]},
      {stage2_7[0],stage2_6[3],stage2_5[3],stage2_4[6],stage2_3[6]}
   );
   gpc615_5 gpc106 (
      {stage1_3[8], stage1_3[9], stage1_3[10], stage1_3[11], stage1_3[12]},
      {stage1_4[19]},
      {stage1_5[6], stage1_5[7], stage1_5[8], stage1_5[9], stage1_5[10], stage1_5[11]},
      {stage2_7[1],stage2_6[4],stage2_5[4],stage2_4[7],stage2_3[7]}
   );
   gpc615_5 gpc107 (
      {stage1_3[13], stage1_3[14], stage1_3[15], stage1_3[16], stage1_3[17]},
      {stage1_4[20]},
      {stage1_5[12], stage1_5[13], stage1_5[14], stage1_5[15], stage1_5[16], stage1_5[17]},
      {stage2_7[2],stage2_6[5],stage2_5[5],stage2_4[8],stage2_3[8]}
   );
   gpc207_4 gpc108 (
      {stage1_4[21], stage1_4[22], stage1_4[23], stage1_4[24], stage1_4[25], stage1_4[26], stage1_4[27]},
      {stage1_6[0], stage1_6[1]},
      {stage2_7[3],stage2_6[6],stage2_5[6],stage2_4[9]}
   );
   gpc606_5 gpc109 (
      {stage1_4[28], stage1_4[29], stage1_4[30], stage1_4[31], stage1_4[32], stage1_4[33]},
      {stage1_6[2], stage1_6[3], stage1_6[4], stage1_6[5], stage1_6[6], stage1_6[7]},
      {stage2_8[0],stage2_7[4],stage2_6[7],stage2_5[7],stage2_4[10]}
   );
   gpc606_5 gpc110 (
      {stage1_5[18], stage1_5[19], stage1_5[20], stage1_5[21], stage1_5[22], stage1_5[23]},
      {stage1_7[0], stage1_7[1], stage1_7[2], stage1_7[3], stage1_7[4], stage1_7[5]},
      {stage2_9[0],stage2_8[1],stage2_7[5],stage2_6[8],stage2_5[8]}
   );
   gpc615_5 gpc111 (
      {stage1_6[8], stage1_6[9], stage1_6[10], stage1_6[11], stage1_6[12]},
      {stage1_7[6]},
      {stage1_8[0], stage1_8[1], stage1_8[2], stage1_8[3], stage1_8[4], stage1_8[5]},
      {stage2_10[0],stage2_9[1],stage2_8[2],stage2_7[6],stage2_6[9]}
   );
   gpc615_5 gpc112 (
      {stage1_6[13], stage1_6[14], stage1_6[15], stage1_6[16], stage1_6[17]},
      {stage1_7[7]},
      {stage1_8[6], stage1_8[7], stage1_8[8], stage1_8[9], stage1_8[10], stage1_8[11]},
      {stage2_10[1],stage2_9[2],stage2_8[3],stage2_7[7],stage2_6[10]}
   );
   gpc615_5 gpc113 (
      {stage1_7[8], stage1_7[9], stage1_7[10], stage1_7[11], stage1_7[12]},
      {stage1_8[12]},
      {stage1_9[0], stage1_9[1], stage1_9[2], stage1_9[3], stage1_9[4], stage1_9[5]},
      {stage2_11[0],stage2_10[2],stage2_9[3],stage2_8[4],stage2_7[8]}
   );
   gpc615_5 gpc114 (
      {stage1_7[13], stage1_7[14], stage1_7[15], stage1_7[16], stage1_7[17]},
      {stage1_8[13]},
      {stage1_9[6], stage1_9[7], stage1_9[8], stage1_9[9], stage1_9[10], stage1_9[11]},
      {stage2_11[1],stage2_10[3],stage2_9[4],stage2_8[5],stage2_7[9]}
   );
   gpc606_5 gpc115 (
      {stage1_8[14], stage1_8[15], stage1_8[16], stage1_8[17], stage1_8[18], stage1_8[19]},
      {stage1_10[0], stage1_10[1], stage1_10[2], stage1_10[3], stage1_10[4], stage1_10[5]},
      {stage2_12[0],stage2_11[2],stage2_10[4],stage2_9[5],stage2_8[6]}
   );
   gpc606_5 gpc116 (
      {stage1_8[20], stage1_8[21], stage1_8[22], stage1_8[23], stage1_8[24], stage1_8[25]},
      {stage1_10[6], stage1_10[7], stage1_10[8], stage1_10[9], stage1_10[10], stage1_10[11]},
      {stage2_12[1],stage2_11[3],stage2_10[5],stage2_9[6],stage2_8[7]}
   );
   gpc606_5 gpc117 (
      {stage1_9[12], stage1_9[13], stage1_9[14], stage1_9[15], stage1_9[16], stage1_9[17]},
      {stage1_11[0], stage1_11[1], stage1_11[2], stage1_11[3], stage1_11[4], stage1_11[5]},
      {stage2_13[0],stage2_12[2],stage2_11[4],stage2_10[6],stage2_9[7]}
   );
   gpc606_5 gpc118 (
      {stage1_9[18], stage1_9[19], stage1_9[20], stage1_9[21], stage1_9[22], stage1_9[23]},
      {stage1_11[6], stage1_11[7], stage1_11[8], stage1_11[9], stage1_11[10], stage1_11[11]},
      {stage2_13[1],stage2_12[3],stage2_11[5],stage2_10[7],stage2_9[8]}
   );
   gpc1163_5 gpc119 (
      {stage1_10[12], stage1_10[13], stage1_10[14]},
      {stage1_11[12], stage1_11[13], stage1_11[14], stage1_11[15], stage1_11[16], stage1_11[17]},
      {stage1_12[0]},
      {stage1_13[0]},
      {stage2_14[0],stage2_13[2],stage2_12[4],stage2_11[6],stage2_10[8]}
   );
   gpc117_4 gpc120 (
      {stage1_12[1], stage1_12[2], stage1_12[3], stage1_12[4], stage1_12[5], stage1_12[6], stage1_12[7]},
      {stage1_13[1]},
      {stage1_14[0]},
      {stage2_15[0],stage2_14[1],stage2_13[3],stage2_12[5]}
   );
   gpc606_5 gpc121 (
      {stage1_12[8], stage1_12[9], stage1_12[10], stage1_12[11], stage1_12[12], stage1_12[13]},
      {stage1_14[1], stage1_14[2], stage1_14[3], stage1_14[4], stage1_14[5], stage1_14[6]},
      {stage2_16[0],stage2_15[1],stage2_14[2],stage2_13[4],stage2_12[6]}
   );
   gpc606_5 gpc122 (
      {stage1_12[14], stage1_12[15], stage1_12[16], stage1_12[17], stage1_12[18], stage1_12[19]},
      {stage1_14[7], stage1_14[8], stage1_14[9], stage1_14[10], stage1_14[11], stage1_14[12]},
      {stage2_16[1],stage2_15[2],stage2_14[3],stage2_13[5],stage2_12[7]}
   );
   gpc606_5 gpc123 (
      {stage1_12[20], stage1_12[21], stage1_12[22], stage1_12[23], stage1_12[24], stage1_12[25]},
      {stage1_14[13], stage1_14[14], stage1_14[15], stage1_14[16], stage1_14[17], 1'b0},
      {stage2_16[2],stage2_15[3],stage2_14[4],stage2_13[6],stage2_12[8]}
   );
   gpc606_5 gpc124 (
      {stage1_13[2], stage1_13[3], stage1_13[4], stage1_13[5], stage1_13[6], stage1_13[7]},
      {stage1_15[0], stage1_15[1], stage1_15[2], stage1_15[3], stage1_15[4], stage1_15[5]},
      {stage2_17[0],stage2_16[3],stage2_15[4],stage2_14[5],stage2_13[7]}
   );
   gpc606_5 gpc125 (
      {stage1_13[8], stage1_13[9], stage1_13[10], stage1_13[11], stage1_13[12], stage1_13[13]},
      {stage1_15[6], stage1_15[7], stage1_15[8], stage1_15[9], stage1_15[10], stage1_15[11]},
      {stage2_17[1],stage2_16[4],stage2_15[5],stage2_14[6],stage2_13[8]}
   );
   gpc606_5 gpc126 (
      {stage1_13[14], stage1_13[15], stage1_13[16], stage1_13[17], stage1_13[18], stage1_13[19]},
      {stage1_15[12], stage1_15[13], stage1_15[14], stage1_15[15], stage1_15[16], stage1_15[17]},
      {stage2_17[2],stage2_16[5],stage2_15[6],stage2_14[7],stage2_13[9]}
   );
   gpc606_5 gpc127 (
      {stage1_13[20], stage1_13[21], stage1_13[22], stage1_13[23], stage1_13[24], stage1_13[25]},
      {stage1_15[18], stage1_15[19], stage1_15[20], stage1_15[21], stage1_15[22], stage1_15[23]},
      {stage2_17[3],stage2_16[6],stage2_15[7],stage2_14[8],stage2_13[10]}
   );
   gpc117_4 gpc128 (
      {stage1_16[0], stage1_16[1], stage1_16[2], stage1_16[3], stage1_16[4], stage1_16[5], stage1_16[6]},
      {stage1_17[0]},
      {1'b0},
      {stage2_19[0],stage2_18[0],stage2_17[4],stage2_16[7]}
   );
   gpc117_4 gpc129 (
      {stage1_16[7], stage1_16[8], stage1_16[9], stage1_16[10], stage1_16[11], stage1_16[12], stage1_16[13]},
      {stage1_17[1]},
      {1'b0},
      {stage2_19[1],stage2_18[1],stage2_17[5],stage2_16[8]}
   );
   gpc1163_5 gpc130 (
      {stage1_16[14], stage1_16[15], stage1_16[16]},
      {stage1_17[2], stage1_17[3], stage1_17[4], stage1_17[5], stage1_17[6], stage1_17[7]},
      {1'b0},
      {1'b0},
      {stage2_20[0],stage2_19[2],stage2_18[2],stage2_17[6],stage2_16[9]}
   );
   gpc1_1 gpc131 (
      {stage1_0[9]},
      {stage2_0[3]}
   );
   gpc1_1 gpc132 (
      {stage1_0[10]},
      {stage2_0[4]}
   );
   gpc1_1 gpc133 (
      {stage1_0[11]},
      {stage2_0[5]}
   );
   gpc1_1 gpc134 (
      {stage1_0[12]},
      {stage2_0[6]}
   );
   gpc1_1 gpc135 (
      {stage1_0[13]},
      {stage2_0[7]}
   );
   gpc1_1 gpc136 (
      {stage1_2[21]},
      {stage2_2[6]}
   );
   gpc1_1 gpc137 (
      {stage1_2[22]},
      {stage2_2[7]}
   );
   gpc1_1 gpc138 (
      {stage1_4[34]},
      {stage2_4[11]}
   );
   gpc1_1 gpc139 (
      {stage1_5[24]},
      {stage2_5[9]}
   );
   gpc1_1 gpc140 (
      {stage1_6[18]},
      {stage2_6[11]}
   );
   gpc1_1 gpc141 (
      {stage1_7[18]},
      {stage2_7[10]}
   );
   gpc1_1 gpc142 (
      {stage1_9[24]},
      {stage2_9[9]}
   );
   gpc1_1 gpc143 (
      {stage1_9[25]},
      {stage2_9[10]}
   );
   gpc1_1 gpc144 (
      {stage1_9[26]},
      {stage2_9[11]}
   );
   gpc1_1 gpc145 (
      {stage1_10[15]},
      {stage2_10[9]}
   );
   gpc1_1 gpc146 (
      {stage1_10[16]},
      {stage2_10[10]}
   );
   gpc1_1 gpc147 (
      {stage1_10[17]},
      {stage2_10[11]}
   );
   gpc1_1 gpc148 (
      {stage1_10[18]},
      {stage2_10[12]}
   );
   gpc207_4 gpc149 (
      {stage2_0[0], stage2_0[1], stage2_0[2], stage2_0[3], stage2_0[4], stage2_0[5], stage2_0[6]},
      {stage2_2[0], stage2_2[1]},
      {stage3_3[0],stage3_2[0],stage3_1[0],stage3_0[0]}
   );
   gpc1163_5 gpc150 (
      {stage2_1[0], stage2_1[1], stage2_1[2]},
      {stage2_2[2], stage2_2[3], stage2_2[4], stage2_2[5], stage2_2[6], stage2_2[7]},
      {stage2_3[0]},
      {stage2_4[0]},
      {stage3_5[0],stage3_4[0],stage3_3[1],stage3_2[1],stage3_1[1]}
   );
   gpc615_5 gpc151 (
      {stage2_3[1], stage2_3[2], stage2_3[3], stage2_3[4], stage2_3[5]},
      {stage2_4[1]},
      {stage2_5[0], stage2_5[1], stage2_5[2], stage2_5[3], stage2_5[4], stage2_5[5]},
      {stage3_7[0],stage3_6[0],stage3_5[1],stage3_4[1],stage3_3[2]}
   );
   gpc615_5 gpc152 (
      {stage2_4[2], stage2_4[3], stage2_4[4], stage2_4[5], stage2_4[6]},
      {stage2_5[6]},
      {stage2_6[0], stage2_6[1], stage2_6[2], stage2_6[3], stage2_6[4], stage2_6[5]},
      {stage3_8[0],stage3_7[1],stage3_6[1],stage3_5[2],stage3_4[2]}
   );
   gpc615_5 gpc153 (
      {stage2_4[7], stage2_4[8], stage2_4[9], stage2_4[10], stage2_4[11]},
      {stage2_5[7]},
      {stage2_6[6], stage2_6[7], stage2_6[8], stage2_6[9], stage2_6[10], stage2_6[11]},
      {stage3_8[1],stage3_7[2],stage3_6[2],stage3_5[3],stage3_4[3]}
   );
   gpc615_5 gpc154 (
      {stage2_7[0], stage2_7[1], stage2_7[2], stage2_7[3], stage2_7[4]},
      {stage2_8[0]},
      {stage2_9[0], stage2_9[1], stage2_9[2], stage2_9[3], stage2_9[4], stage2_9[5]},
      {stage3_11[0],stage3_10[0],stage3_9[0],stage3_8[2],stage3_7[3]}
   );
   gpc615_5 gpc155 (
      {stage2_7[5], stage2_7[6], stage2_7[7], stage2_7[8], stage2_7[9]},
      {stage2_8[1]},
      {stage2_9[6], stage2_9[7], stage2_9[8], stage2_9[9], stage2_9[10], stage2_9[11]},
      {stage3_11[1],stage3_10[1],stage3_9[1],stage3_8[3],stage3_7[4]}
   );
   gpc606_5 gpc156 (
      {stage2_8[2], stage2_8[3], stage2_8[4], stage2_8[5], stage2_8[6], stage2_8[7]},
      {stage2_10[0], stage2_10[1], stage2_10[2], stage2_10[3], stage2_10[4], stage2_10[5]},
      {stage3_12[0],stage3_11[2],stage3_10[2],stage3_9[2],stage3_8[4]}
   );
   gpc7_3 gpc157 (
      {stage2_10[6], stage2_10[7], stage2_10[8], stage2_10[9], stage2_10[10], stage2_10[11], stage2_10[12]},
      {stage3_12[1],stage3_11[3],stage3_10[3]}
   );
   gpc606_5 gpc158 (
      {stage2_11[0], stage2_11[1], stage2_11[2], stage2_11[3], stage2_11[4], stage2_11[5]},
      {stage2_13[0], stage2_13[1], stage2_13[2], stage2_13[3], stage2_13[4], stage2_13[5]},
      {stage3_15[0],stage3_14[0],stage3_13[0],stage3_12[2],stage3_11[4]}
   );
   gpc1343_5 gpc159 (
      {stage2_12[0], stage2_12[1], stage2_12[2]},
      {stage2_13[6], stage2_13[7], stage2_13[8], stage2_13[9]},
      {stage2_14[0], stage2_14[1], stage2_14[2]},
      {stage2_15[0]},
      {stage3_16[0],stage3_15[1],stage3_14[1],stage3_13[1],stage3_12[3]}
   );
   gpc615_5 gpc160 (
      {stage2_12[3], stage2_12[4], stage2_12[5], stage2_12[6], stage2_12[7]},
      {stage2_13[10]},
      {stage2_14[3], stage2_14[4], stage2_14[5], stage2_14[6], stage2_14[7], stage2_14[8]},
      {stage3_16[1],stage3_15[2],stage3_14[2],stage3_13[2],stage3_12[4]}
   );
   gpc117_4 gpc161 (
      {stage2_15[1], stage2_15[2], stage2_15[3], stage2_15[4], stage2_15[5], stage2_15[6], stage2_15[7]},
      {stage2_16[0]},
      {stage2_17[0]},
      {stage3_18[0],stage3_17[0],stage3_16[2],stage3_15[3]}
   );
   gpc7_3 gpc162 (
      {stage2_16[1], stage2_16[2], stage2_16[3], stage2_16[4], stage2_16[5], stage2_16[6], stage2_16[7]},
      {stage3_18[1],stage3_17[1],stage3_16[3]}
   );
   gpc1325_5 gpc163 (
      {stage2_17[1], stage2_17[2], stage2_17[3], stage2_17[4], stage2_17[5]},
      {stage2_18[0], stage2_18[1]},
      {stage2_19[0], stage2_19[1], stage2_19[2]},
      {stage2_20[0]},
      {stage3_21[0],stage3_20[0],stage3_19[0],stage3_18[2],stage3_17[2]}
   );
   gpc1_1 gpc164 (
      {stage2_0[7]},
      {stage3_0[1]}
   );
   gpc1_1 gpc165 (
      {stage2_3[6]},
      {stage3_3[3]}
   );
   gpc1_1 gpc166 (
      {stage2_3[7]},
      {stage3_3[4]}
   );
   gpc1_1 gpc167 (
      {stage2_3[8]},
      {stage3_3[5]}
   );
   gpc1_1 gpc168 (
      {stage2_5[8]},
      {stage3_5[4]}
   );
   gpc1_1 gpc169 (
      {stage2_5[9]},
      {stage3_5[5]}
   );
   gpc1_1 gpc170 (
      {stage2_7[10]},
      {stage3_7[5]}
   );
   gpc1_1 gpc171 (
      {stage2_11[6]},
      {stage3_11[5]}
   );
   gpc1_1 gpc172 (
      {stage2_12[8]},
      {stage3_12[5]}
   );
   gpc1_1 gpc173 (
      {stage2_16[8]},
      {stage3_16[4]}
   );
   gpc1_1 gpc174 (
      {stage2_16[9]},
      {stage3_16[5]}
   );
   gpc1_1 gpc175 (
      {stage2_17[6]},
      {stage3_17[3]}
   );
   gpc1_1 gpc176 (
      {stage2_18[2]},
      {stage3_18[3]}
   );
   gpc2135_5 gpc177 (
      {stage3_3[0], stage3_3[1], stage3_3[2], stage3_3[3], stage3_3[4]},
      {stage3_4[0], stage3_4[1], stage3_4[2]},
      {stage3_5[0]},
      {stage3_6[0], stage3_6[1]},
      {stage4_7[0],stage4_6[0],stage4_5[0],stage4_4[0],stage4_3[0]}
   );
   gpc615_5 gpc178 (
      {stage3_5[1], stage3_5[2], stage3_5[3], stage3_5[4], stage3_5[5]},
      {stage3_6[2]},
      {stage3_7[0], stage3_7[1], stage3_7[2], stage3_7[3], stage3_7[4], stage3_7[5]},
      {stage4_9[0],stage4_8[0],stage4_7[1],stage4_6[1],stage4_5[1]}
   );
   gpc135_4 gpc179 (
      {stage3_8[0], stage3_8[1], stage3_8[2], stage3_8[3], stage3_8[4]},
      {stage3_9[0], stage3_9[1], stage3_9[2]},
      {stage3_10[0]},
      {stage4_11[0],stage4_10[0],stage4_9[1],stage4_8[1]}
   );
   gpc1163_5 gpc180 (
      {stage3_10[1], stage3_10[2], stage3_10[3]},
      {stage3_11[0], stage3_11[1], stage3_11[2], stage3_11[3], stage3_11[4], stage3_11[5]},
      {stage3_12[0]},
      {stage3_13[0]},
      {stage4_14[0],stage4_13[0],stage4_12[0],stage4_11[1],stage4_10[1]}
   );
   gpc1325_5 gpc181 (
      {stage3_12[1], stage3_12[2], stage3_12[3], stage3_12[4], stage3_12[5]},
      {stage3_13[1], stage3_13[2]},
      {stage3_14[0], stage3_14[1], stage3_14[2]},
      {stage3_15[0]},
      {stage4_16[0],stage4_15[0],stage4_14[1],stage4_13[1],stage4_12[1]}
   );
   gpc1163_5 gpc182 (
      {stage3_15[1], stage3_15[2], stage3_15[3]},
      {stage3_16[0], stage3_16[1], stage3_16[2], stage3_16[3], stage3_16[4], stage3_16[5]},
      {stage3_17[0]},
      {stage3_18[0]},
      {stage4_19[0],stage4_18[0],stage4_17[0],stage4_16[1],stage4_15[1]}
   );
   gpc1163_5 gpc183 (
      {stage3_17[1], stage3_17[2], stage3_17[3]},
      {stage3_18[1], stage3_18[2], stage3_18[3], 1'b0, 1'b0, 1'b0},
      {stage3_19[0]},
      {stage3_20[0]},
      {stage4_21[0],stage4_20[0],stage4_19[1],stage4_18[1],stage4_17[1]}
   );
   gpc1_1 gpc184 (
      {stage3_0[0]},
      {stage4_0[0]}
   );
   gpc1_1 gpc185 (
      {stage3_0[1]},
      {stage4_0[1]}
   );
   gpc1_1 gpc186 (
      {stage3_1[0]},
      {stage4_1[0]}
   );
   gpc1_1 gpc187 (
      {stage3_1[1]},
      {stage4_1[1]}
   );
   gpc1_1 gpc188 (
      {stage3_2[0]},
      {stage4_2[0]}
   );
   gpc1_1 gpc189 (
      {stage3_2[1]},
      {stage4_2[1]}
   );
   gpc1_1 gpc190 (
      {stage3_3[5]},
      {stage4_3[1]}
   );
   gpc1_1 gpc191 (
      {stage3_4[3]},
      {stage4_4[1]}
   );
   gpc1_1 gpc192 (
      {stage3_21[0]},
      {stage4_21[1]}
   );
endmodule
module rowadder2_1_22(input [21:0] src0, input [21:0] src1, output [22:0] dst0);
    wire [21:0] gene;
    wire [21:0] prop;
    wire [23:0] out;
    wire [23:0] carryout;
    LUT2 #(
        .INIT(4'h8)
    ) lut_0_gene (
        .I0(src0[0]),
        .I1(src1[0]),
        .O(gene[0])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_0_prop (
        .I0(src0[0]),
        .I1(src1[0]),
        .O(prop[0])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_1_gene (
        .I0(src0[1]),
        .I1(src1[1]),
        .O(gene[1])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_1_prop (
        .I0(src0[1]),
        .I1(src1[1]),
        .O(prop[1])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_2_gene (
        .I0(src0[2]),
        .I1(src1[2]),
        .O(gene[2])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_2_prop (
        .I0(src0[2]),
        .I1(src1[2]),
        .O(prop[2])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_3_gene (
        .I0(src0[3]),
        .I1(src1[3]),
        .O(gene[3])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_3_prop (
        .I0(src0[3]),
        .I1(src1[3]),
        .O(prop[3])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_4_gene (
        .I0(src0[4]),
        .I1(src1[4]),
        .O(gene[4])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_4_prop (
        .I0(src0[4]),
        .I1(src1[4]),
        .O(prop[4])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_5_gene (
        .I0(src0[5]),
        .I1(src1[5]),
        .O(gene[5])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_5_prop (
        .I0(src0[5]),
        .I1(src1[5]),
        .O(prop[5])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_6_gene (
        .I0(src0[6]),
        .I1(src1[6]),
        .O(gene[6])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_6_prop (
        .I0(src0[6]),
        .I1(src1[6]),
        .O(prop[6])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_7_gene (
        .I0(src0[7]),
        .I1(src1[7]),
        .O(gene[7])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_7_prop (
        .I0(src0[7]),
        .I1(src1[7]),
        .O(prop[7])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_8_gene (
        .I0(src0[8]),
        .I1(src1[8]),
        .O(gene[8])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_8_prop (
        .I0(src0[8]),
        .I1(src1[8]),
        .O(prop[8])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_9_gene (
        .I0(src0[9]),
        .I1(src1[9]),
        .O(gene[9])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_9_prop (
        .I0(src0[9]),
        .I1(src1[9]),
        .O(prop[9])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_10_gene (
        .I0(src0[10]),
        .I1(src1[10]),
        .O(gene[10])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_10_prop (
        .I0(src0[10]),
        .I1(src1[10]),
        .O(prop[10])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_11_gene (
        .I0(src0[11]),
        .I1(src1[11]),
        .O(gene[11])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_11_prop (
        .I0(src0[11]),
        .I1(src1[11]),
        .O(prop[11])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_12_gene (
        .I0(src0[12]),
        .I1(src1[12]),
        .O(gene[12])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_12_prop (
        .I0(src0[12]),
        .I1(src1[12]),
        .O(prop[12])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_13_gene (
        .I0(src0[13]),
        .I1(src1[13]),
        .O(gene[13])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_13_prop (
        .I0(src0[13]),
        .I1(src1[13]),
        .O(prop[13])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_14_gene (
        .I0(src0[14]),
        .I1(src1[14]),
        .O(gene[14])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_14_prop (
        .I0(src0[14]),
        .I1(src1[14]),
        .O(prop[14])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_15_gene (
        .I0(src0[15]),
        .I1(src1[15]),
        .O(gene[15])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_15_prop (
        .I0(src0[15]),
        .I1(src1[15]),
        .O(prop[15])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_16_gene (
        .I0(src0[16]),
        .I1(src1[16]),
        .O(gene[16])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_16_prop (
        .I0(src0[16]),
        .I1(src1[16]),
        .O(prop[16])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_17_gene (
        .I0(src0[17]),
        .I1(src1[17]),
        .O(gene[17])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_17_prop (
        .I0(src0[17]),
        .I1(src1[17]),
        .O(prop[17])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_18_gene (
        .I0(src0[18]),
        .I1(src1[18]),
        .O(gene[18])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_18_prop (
        .I0(src0[18]),
        .I1(src1[18]),
        .O(prop[18])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_19_gene (
        .I0(src0[19]),
        .I1(src1[19]),
        .O(gene[19])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_19_prop (
        .I0(src0[19]),
        .I1(src1[19]),
        .O(prop[19])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_20_gene (
        .I0(src0[20]),
        .I1(src1[20]),
        .O(gene[20])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_20_prop (
        .I0(src0[20]),
        .I1(src1[20]),
        .O(prop[20])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_21_gene (
        .I0(src0[21]),
        .I1(src1[21]),
        .O(gene[21])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_21_prop (
        .I0(src0[21]),
        .I1(src1[21]),
        .O(prop[21])
    );
    CARRY4 carry4_3_0 (
        .CO(carryout[3:0]),
        .O(out[3:0]),
        .CI(1'h0),
        .CYINIT(1'h0),
        .DI(gene[3:0]),
        .S(prop[3:0])
    );
    CARRY4 carry4_7_4 (
        .CO(carryout[7:4]),
        .O(out[7:4]),
        .CI(carryout[3]),
        .CYINIT(1'h0),
        .DI(gene[7:4]),
        .S(prop[7:4])
    );
    CARRY4 carry4_11_8 (
        .CO(carryout[11:8]),
        .O(out[11:8]),
        .CI(carryout[7]),
        .CYINIT(1'h0),
        .DI(gene[11:8]),
        .S(prop[11:8])
    );
    CARRY4 carry4_15_12 (
        .CO(carryout[15:12]),
        .O(out[15:12]),
        .CI(carryout[11]),
        .CYINIT(1'h0),
        .DI(gene[15:12]),
        .S(prop[15:12])
    );
    CARRY4 carry4_19_16 (
        .CO(carryout[19:16]),
        .O(out[19:16]),
        .CI(carryout[15]),
        .CYINIT(1'h0),
        .DI(gene[19:16]),
        .S(prop[19:16])
    );
    CARRY4 carry4_23_20 (
        .CO(carryout[23:20]),
        .O(out[23:20]),
        .CI(carryout[19]),
        .CYINIT(1'h0),
        .DI({2'h0, gene[21:20]}),
        .S({2'h0, prop[21:20]})
    );
    assign dst0 = {carryout[21], out[21:0]};
endmodule


module testbench();
    reg [53:0] src0;
    reg [53:0] src1;
    reg [53:0] src2;
    reg [53:0] src3;
    reg [53:0] src4;
    reg [53:0] src5;
    reg [53:0] src6;
    reg [53:0] src7;
    reg [53:0] src8;
    reg [53:0] src9;
    reg [53:0] src10;
    reg [53:0] src11;
    reg [53:0] src12;
    reg [53:0] src13;
    reg [53:0] src14;
    reg [53:0] src15;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [21:0] srcsum;
    wire [21:0] dstsum;
    wire test;
    compressor2_1_54_16 compressor2_1_54_16(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13] + src0[14] + src0[15] + src0[16] + src0[17] + src0[18] + src0[19] + src0[20] + src0[21] + src0[22] + src0[23] + src0[24] + src0[25] + src0[26] + src0[27] + src0[28] + src0[29] + src0[30] + src0[31] + src0[32] + src0[33] + src0[34] + src0[35] + src0[36] + src0[37] + src0[38] + src0[39] + src0[40] + src0[41] + src0[42] + src0[43] + src0[44] + src0[45] + src0[46] + src0[47] + src0[48] + src0[49] + src0[50] + src0[51] + src0[52] + src0[53])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13] + src1[14] + src1[15] + src1[16] + src1[17] + src1[18] + src1[19] + src1[20] + src1[21] + src1[22] + src1[23] + src1[24] + src1[25] + src1[26] + src1[27] + src1[28] + src1[29] + src1[30] + src1[31] + src1[32] + src1[33] + src1[34] + src1[35] + src1[36] + src1[37] + src1[38] + src1[39] + src1[40] + src1[41] + src1[42] + src1[43] + src1[44] + src1[45] + src1[46] + src1[47] + src1[48] + src1[49] + src1[50] + src1[51] + src1[52] + src1[53])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13] + src2[14] + src2[15] + src2[16] + src2[17] + src2[18] + src2[19] + src2[20] + src2[21] + src2[22] + src2[23] + src2[24] + src2[25] + src2[26] + src2[27] + src2[28] + src2[29] + src2[30] + src2[31] + src2[32] + src2[33] + src2[34] + src2[35] + src2[36] + src2[37] + src2[38] + src2[39] + src2[40] + src2[41] + src2[42] + src2[43] + src2[44] + src2[45] + src2[46] + src2[47] + src2[48] + src2[49] + src2[50] + src2[51] + src2[52] + src2[53])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13] + src3[14] + src3[15] + src3[16] + src3[17] + src3[18] + src3[19] + src3[20] + src3[21] + src3[22] + src3[23] + src3[24] + src3[25] + src3[26] + src3[27] + src3[28] + src3[29] + src3[30] + src3[31] + src3[32] + src3[33] + src3[34] + src3[35] + src3[36] + src3[37] + src3[38] + src3[39] + src3[40] + src3[41] + src3[42] + src3[43] + src3[44] + src3[45] + src3[46] + src3[47] + src3[48] + src3[49] + src3[50] + src3[51] + src3[52] + src3[53])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13] + src4[14] + src4[15] + src4[16] + src4[17] + src4[18] + src4[19] + src4[20] + src4[21] + src4[22] + src4[23] + src4[24] + src4[25] + src4[26] + src4[27] + src4[28] + src4[29] + src4[30] + src4[31] + src4[32] + src4[33] + src4[34] + src4[35] + src4[36] + src4[37] + src4[38] + src4[39] + src4[40] + src4[41] + src4[42] + src4[43] + src4[44] + src4[45] + src4[46] + src4[47] + src4[48] + src4[49] + src4[50] + src4[51] + src4[52] + src4[53])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13] + src5[14] + src5[15] + src5[16] + src5[17] + src5[18] + src5[19] + src5[20] + src5[21] + src5[22] + src5[23] + src5[24] + src5[25] + src5[26] + src5[27] + src5[28] + src5[29] + src5[30] + src5[31] + src5[32] + src5[33] + src5[34] + src5[35] + src5[36] + src5[37] + src5[38] + src5[39] + src5[40] + src5[41] + src5[42] + src5[43] + src5[44] + src5[45] + src5[46] + src5[47] + src5[48] + src5[49] + src5[50] + src5[51] + src5[52] + src5[53])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13] + src6[14] + src6[15] + src6[16] + src6[17] + src6[18] + src6[19] + src6[20] + src6[21] + src6[22] + src6[23] + src6[24] + src6[25] + src6[26] + src6[27] + src6[28] + src6[29] + src6[30] + src6[31] + src6[32] + src6[33] + src6[34] + src6[35] + src6[36] + src6[37] + src6[38] + src6[39] + src6[40] + src6[41] + src6[42] + src6[43] + src6[44] + src6[45] + src6[46] + src6[47] + src6[48] + src6[49] + src6[50] + src6[51] + src6[52] + src6[53])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13] + src7[14] + src7[15] + src7[16] + src7[17] + src7[18] + src7[19] + src7[20] + src7[21] + src7[22] + src7[23] + src7[24] + src7[25] + src7[26] + src7[27] + src7[28] + src7[29] + src7[30] + src7[31] + src7[32] + src7[33] + src7[34] + src7[35] + src7[36] + src7[37] + src7[38] + src7[39] + src7[40] + src7[41] + src7[42] + src7[43] + src7[44] + src7[45] + src7[46] + src7[47] + src7[48] + src7[49] + src7[50] + src7[51] + src7[52] + src7[53])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13] + src8[14] + src8[15] + src8[16] + src8[17] + src8[18] + src8[19] + src8[20] + src8[21] + src8[22] + src8[23] + src8[24] + src8[25] + src8[26] + src8[27] + src8[28] + src8[29] + src8[30] + src8[31] + src8[32] + src8[33] + src8[34] + src8[35] + src8[36] + src8[37] + src8[38] + src8[39] + src8[40] + src8[41] + src8[42] + src8[43] + src8[44] + src8[45] + src8[46] + src8[47] + src8[48] + src8[49] + src8[50] + src8[51] + src8[52] + src8[53])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13] + src9[14] + src9[15] + src9[16] + src9[17] + src9[18] + src9[19] + src9[20] + src9[21] + src9[22] + src9[23] + src9[24] + src9[25] + src9[26] + src9[27] + src9[28] + src9[29] + src9[30] + src9[31] + src9[32] + src9[33] + src9[34] + src9[35] + src9[36] + src9[37] + src9[38] + src9[39] + src9[40] + src9[41] + src9[42] + src9[43] + src9[44] + src9[45] + src9[46] + src9[47] + src9[48] + src9[49] + src9[50] + src9[51] + src9[52] + src9[53])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13] + src10[14] + src10[15] + src10[16] + src10[17] + src10[18] + src10[19] + src10[20] + src10[21] + src10[22] + src10[23] + src10[24] + src10[25] + src10[26] + src10[27] + src10[28] + src10[29] + src10[30] + src10[31] + src10[32] + src10[33] + src10[34] + src10[35] + src10[36] + src10[37] + src10[38] + src10[39] + src10[40] + src10[41] + src10[42] + src10[43] + src10[44] + src10[45] + src10[46] + src10[47] + src10[48] + src10[49] + src10[50] + src10[51] + src10[52] + src10[53])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13] + src11[14] + src11[15] + src11[16] + src11[17] + src11[18] + src11[19] + src11[20] + src11[21] + src11[22] + src11[23] + src11[24] + src11[25] + src11[26] + src11[27] + src11[28] + src11[29] + src11[30] + src11[31] + src11[32] + src11[33] + src11[34] + src11[35] + src11[36] + src11[37] + src11[38] + src11[39] + src11[40] + src11[41] + src11[42] + src11[43] + src11[44] + src11[45] + src11[46] + src11[47] + src11[48] + src11[49] + src11[50] + src11[51] + src11[52] + src11[53])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12] + src12[13] + src12[14] + src12[15] + src12[16] + src12[17] + src12[18] + src12[19] + src12[20] + src12[21] + src12[22] + src12[23] + src12[24] + src12[25] + src12[26] + src12[27] + src12[28] + src12[29] + src12[30] + src12[31] + src12[32] + src12[33] + src12[34] + src12[35] + src12[36] + src12[37] + src12[38] + src12[39] + src12[40] + src12[41] + src12[42] + src12[43] + src12[44] + src12[45] + src12[46] + src12[47] + src12[48] + src12[49] + src12[50] + src12[51] + src12[52] + src12[53])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13] + src13[14] + src13[15] + src13[16] + src13[17] + src13[18] + src13[19] + src13[20] + src13[21] + src13[22] + src13[23] + src13[24] + src13[25] + src13[26] + src13[27] + src13[28] + src13[29] + src13[30] + src13[31] + src13[32] + src13[33] + src13[34] + src13[35] + src13[36] + src13[37] + src13[38] + src13[39] + src13[40] + src13[41] + src13[42] + src13[43] + src13[44] + src13[45] + src13[46] + src13[47] + src13[48] + src13[49] + src13[50] + src13[51] + src13[52] + src13[53])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14] + src14[15] + src14[16] + src14[17] + src14[18] + src14[19] + src14[20] + src14[21] + src14[22] + src14[23] + src14[24] + src14[25] + src14[26] + src14[27] + src14[28] + src14[29] + src14[30] + src14[31] + src14[32] + src14[33] + src14[34] + src14[35] + src14[36] + src14[37] + src14[38] + src14[39] + src14[40] + src14[41] + src14[42] + src14[43] + src14[44] + src14[45] + src14[46] + src14[47] + src14[48] + src14[49] + src14[50] + src14[51] + src14[52] + src14[53])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15] + src15[16] + src15[17] + src15[18] + src15[19] + src15[20] + src15[21] + src15[22] + src15[23] + src15[24] + src15[25] + src15[26] + src15[27] + src15[28] + src15[29] + src15[30] + src15[31] + src15[32] + src15[33] + src15[34] + src15[35] + src15[36] + src15[37] + src15[38] + src15[39] + src15[40] + src15[41] + src15[42] + src15[43] + src15[44] + src15[45] + src15[46] + src15[47] + src15[48] + src15[49] + src15[50] + src15[51] + src15[52] + src15[53])<<15);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'h0;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'h88f53284c68b8c6211d19c49e62d463695f4f2751783100d797ede9c2ddcbf4dbedeecad10c66c4fb2952467d69d28b0ba825d1f667d420d637037260144a10c249b5719f5b9c9a5c69f89193b1c1107b170cff5d51198a3c3deab39d4f01f99a54e6510d322b69323dda37d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'h9e74f072c794d39128b7cd69543a59d0c007f5b1aa6d4bc08788e66abfc77841422b8dd03a3224b3798da5014331880a10a3563eb79b9dfe37afcc0576a2d0317e9206587cd4f1fca7ce68c08fff514f121c8339f394b373696e00170d76a8e2e675a050976c76cbc243c80a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'h38fe5a67e0c449bdec53eaced600c7fa8fff5f14eb0608a04083decf7b9c7f2a55f361e127f61f7cc3cb76f714f91c75f2e180ea0cf1dbd73db6d63ecb9aec387a2108e4dfdd722a296fc015dc3f5aad3a4718742c099c24f16486ed7e59bd2d06109790e6b3d2a8d0f33a15;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'ha62a9a0f1a55980dea4546531e5e7b3fe53a5cfc0abca142600d2f097d750d4be2c5c7c26bdbbda114fe77322182dba243ee71efbf823a486f37db3b3202b039306e6063150b5d18490b085297f34a6d61e1c7ebe1f49555b83e3577ff968af3e07bcf3ba529701bbf27c29e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'hfcf8466866b9642aa1288c44d356259fb17511febcb7e912733df3d397222d061ebc0b64173e497a39146365ee75d19a0490f53b3038dcc7e6237d729cccba92e5aca3267bfa56ff64e481a842a285ce29da86097038d0560f33236e14cae76df030e05d7dc01a61ebc757f0;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'h562a29b84cd640fdc10a33bbbc06810c38c2dd00a1941f225810277f23d12be97d86c276eeca3b8ac67027659278e087f0eb207f62b4a2633c7c1cc53ca7250f0516b574ee21cf30168eea4ab415aa86d9ebfa9da5e07d9aa91f3af9002e406cfc308b674da0c9f385776ac9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'hecba213ac7a7a45ce868b19a6891d1a307622582eac90ec091b24e1fad6ab79cfc8b5c0ad76bc0f7b9e37ad21ef0635387e83b362140754fe1990b794ff6a2a96c9537681598a585cc7732bcd36ab49df42a40fbfefb90d1b1b7982b0f5380a776be3e9b488c2e5dd226d53a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'h5e05ee99652fc32c198c52b027f8864e7fb3992630379559362f9d384c590a02ec868466ba43bf22e9caf949bec0e28b2497d65e2aca22e74db5f7a8c2ac5dddfcd6bddada3d1ec98db7334f751ebc386fe3fb8e174cf72bb38d5300a5112bc77b191f36d956af77ee7cc38c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'hf44cc1ba195dc1fe08916dfdc11a9b167279c9f32673cb4f2120b37d0834190cfa0150f010e7781fc392542a6e8544132cf94061ec84e8a2b88a59f27b9380644c78c5d6c8572855f89a1dece1a429a4a928d159c15a7bd6fbe30b4c4c4e567599859512973ec36b72f37380;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'ha8cdab0cea6a9e490d03a369b00395df6c212fc13a90b93a06f8a2b89f6f5cb35aa34c456adfba46ca858f739d491b9432c300e516f429b665b89e8b910a513594f7dd4155ba4e6a57a33c2e225d5f591394d7aa216a5423c3bd8844de7eb975c4eab67473c4b18d46ed87c4;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'h5e5c42a43973884a2754adda1e1b7c134b7835dae0a5d1f9c503d2f25a861bbde71c9725cdd741704ab0459180a506ec1169692961c24873c60ae2ae5dd856ed88de7f685baf81680b7f397b5119eb877819f9f953a98dd9cef0da38057f955adba3be889225cd4604c26582;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'h7ccd49744ed13fec4d95b5bbbce9b5b3f3739408f98f35787eaa8ce2ea51f4a043e3d73d3027e8f5fe77a6028f92da05a57f8a5e595f7ec132bb25448346a61eccee2a46e931e5c63128ac85eaed15379f160b95fced237303a3a168290191d00f0c5988c1f950c4c66cda1f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'h34efe93cb5618467c374b5e0f0dcb8732856f9ca6c881820ec8baf6c56b7906dec43b7031c60111917abe171033e0d7805adf1fc58198df9f6c5041677412dcc73f6ea9261a725e59e691d48812ba0b6053806dfd864b221cef8c304bc5ff7ebbb7ed2b70491a083ecc5c41f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'ha08d85d2814e273499851df7a1abccc8642bf9e38758703b5cdba2e92666cf23e8a5bb62cfb1ab4b6d5a9087f8f505e550353f30931097085a9d3e82e996514076d95c350d0febef7e2943a5ab211f307aa3fa9ef072ae007bcfa178472a724cd0a08fdde7fcf49d241a9e61;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'hedd7bbb844ad43b386756e625fd3048d0296dd7806b33c524f6e62953c098f90e4b054264971f25e9c8881e9d2ef06ba997af073e6a6cf8ad631aed0480957fb0351ba1b1b2b8017c86655b0dd7e911cfc9be48bae5c3fa4ff8950ff26e971a04652a1ba0d9f141284e44b98;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'h7f02b3dca4f65eedd0ff1da5089743d3af8a70938f706cf1e42b16e151562d1013e6c2d7f5d314eee8f48060ae883fc4cf4a1d7ffbb2f9cbfc823ac58da12f5e54e8471c36bc71083b49b73409894c0a920bd685547e9d01c6e3576703334b68f8a089d595a3aa076a855f2a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'hf4134744f4f5e3a1c06596294abfb1fb82a8e4bd8a5860ebeafad210ed79ef5bdbb717ea89b67b505cd8e19557212091c0a6ef9d33fed3d3ff8a00c7c4b722a74b607759ec548e46072682dbd67cc1bbce1a649d84dfff855a0b2baa3b946aba18285ad59c0df3b186b8aeef;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'h40257f37ffecb13c3140ec9116b6c02874ea7f2749d022219fe4b3e1e8b6e0306b738f4ba92dd90f49e1dbc3a929ce0f0bec8623439756dee7768a60014a3e9be8b25ae76f4b361cfb171b02b2fee91ec1566db09a922dd5cd30e91d0bbb7e3c737a90cdaec2b151b037088e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'hf6552b11da7b77108a9cd77b18cbf6a066836c2da8e70d30e73346f44ee7b8dc46f99e067961a97e0e01da7dbfdf9e752b14ca497e4d17f5bf01033cfb6e5969aa7a1b599f8b80a4528c1546fa8b7c343d15a15957e1d51cd7dc68661438ba773a71ef2dee7177df9361b063;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'h93a4b81beeb772e1513b1865a7fe668b83599e148fd9cec639caf74c9fe8c69f43f603e3ecd4e468b9ea49a969139ad760968309bcd6860cb98c67e115909a9da11fefa5fa43578f5900569cf1af0f8a6a9a9f6fb6c2dc14a160b4f5e1560e194a1235cb88fd253952f9c6ce;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'ha56005723d103ff6a0c0b82e856c5e7fc4a8616726f27fdb0c9849af72d8058c58850b7cc31c9e350615cddf7471faedad0df33bf5337f28ffc29f702d3692a52b20dbba07e8117e6154ab443dc3b9af3fccdc9e16bf1bb7fa52a8b83178c9dfb05cc33fc8f7b491fb4a5edf;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'hac5be2567cae744ebeaeb3273fa0e61d110f5557f894fa37b1e6f599514bf9e509cb253eaa0ac2889a869a478e9be1cf29db4a39eeadc3721eb3ce91e501d1c6320acb8982c764c4c1927e66b2f969889f35437f1dc2da9c7413597b25b526ae747da31d5a32581be55a53a6;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'h5bd4ebce9a3ddc966b3e0dffabc9ad3ee2403ca1e912067e233a72bb1bf334fbb80527cf41aa7b17e75da316d0f00a7aed77c64beacea272ef9b444fb92c1f13a7e15670179211535f30c0a132fc39ff6428801f909f798b943f4328367f83c19d063332667e0bc6545f27dc;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'hfe086308797140b04145cdb5b32be2385344e849c7fcc4f5f58634b3e4ddd66f62865e0d9aa66705b9a54ebe84e10b206a86c6013e7a37f3a70ea3eac8a53f283e3f981aee41a4bd5f7b054fe3491e10cfea22fe279e7284834e93dca869b5ab7476343fb6a71b8c2ad8ec50;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'h816a2fc247236eb1f0a6145c2e474448fc1f0ba0bcf956da17ebebdcdfa7b5663a7f471992779de23c1612997cac809fb276f9bff3845258b8305f995df0a6f3c9f0cbd349617496c0e8925329ab6ee5ce5e1d5de9559460d445d2adf8a92d4806304d61debc237de1abdaa3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'h70ed15b07fb4e2b8f6d20f90ac71d09cd1c9d9cd133e509a2ff175ff17633c5895bc1157a9ff2f01b928aefcbd1501ef32d7bdbfa68edbfb00e2711c8a5c97a4a8eee0f71180a93574a390b30c09e571062cfc83d0f5a8839042f9488f9243c43fd5b466e1d1207de409e8fd;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'h2c3ec31e40f57120211624a5fc1154d9f82030aa7908ef5285acb7b9c20017139ab04438def4ffe3a1c26de742c4e8cf65171ba8c245b082c099bdd68b1d6aaf011fb00d01e84c9ccb1b515bd25cb58ab9eb8219752692b7df3250a15ff228416a59d3effe424ad332e11f11;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'h43ecef8923d9572255abc5a8688a5055d03a6216a99a2e9cce82f49440053d314bd9c6526d6d0b5c2a6ae4d9471a3532b1ea429ad876d057ac3b92fad8b0f6733e6b91d5cbb5a737365b5546db0eb8dc2db2df0428a17cfb4bd15ea2da6d28368d89b135e8512f1b183758eb;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'h9b7b9af06b7b5c1b9ce895df2e39870a28da3ef3471e814ef5620fd9bf16cef8e66a7f75bb4e7a979793561e2079c24cd0a3f972a6de490b47eba6d8c13b621a84887fd2de76fad94477d94db88142de5893f7117af09d16448abb6d4e8847e2ec4a6d40aac4b7ab0d0a6045;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'h705fe32fa54acfd40e4a6f68d01d584a09f632dc39ed228281b8e1cc85902bbdbe0a4f04adb046cbd677dc0283340c9fe92834c51652234b98774e13e2811dd8255c2afd37b43bb9eaf6a5bbcb018cfeffa75e4ac0230c0c8e97c2f0ffa3aaebcb7ccfb51d31b8f454d4dea9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'hb4dbfd3f89ff01e9603d7fca0614ae03439cbfb966db164be5c765853d40a5d25884df16f20b4c643994058ce4e014dae4650eeccaf216d680a13b8d6542f51c8eb63c60196aa26f650e372ab2091dd7d726b6346ece5fce9f7c3fd13a3e1ce3236ea3014213dbfb3ef1003f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'hd06a3cf96ae1587ccb7b127b4ad0aab95cfb0681a7b7af203169c68307a33178734e5cbbec8418cca46363f1acc166a69c4b9d406d74bd8200e49e504e97395fac180c936f0e002b6b6b3a264f4f59af0a95960a38ebe665e452d1c2cf25351aa4729218d5cf334ea1ca53fa;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'h6c0987c4c8817af21ca4ff51de342ad4bad872145cd00b3fdd036ee9caec5b0c3a1c8b94d7e90fd5071347ad9c329df28b95103f0fdb6f80b4f77dd25c7cdddebd58641ceaaf582911551a3f67afe25292aa1a14daada450bc12e479dd19f31235ffbff171ec9c387893295;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'h8b0906293dc3aba081970e36ca7eaa672b49a1407be7d644a7243af527ed4e518646860c692373abecfd188abf65842eff86e519e03c707c48995b51575e8650ab108a1712590bb7f460c92fa3a79049464a8867bfa943723bf04d7252d7b1c9415b0c5fa4e14b5ae0a4f4c8;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'hbfc941628141c4f917ade5c7e10f1d48f5f1c0184eafebc16005c18bea274bbd176ced169ac45e7adeaa7308a1959f4d76af631631ac09485b71f3604cbbde72cd6389759ea1781269101e496e5aa7ec73ed9e8371eeae5864fe08e9d73023b611c443be5bd46c36823356cd;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'h6e434f039debf6431375adb7ff20ae88fed2433e3958ff843c9ade4b64333cb58297f7367ea59af99ff6c6660ff24db78c81be8083342c0eec560f8a17fdb658e5d305ff61b753b26adbeb747e21cfc83a93ece52633efce67d52a1ca4a4debb2476a78faa6cfb8794654aa0;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'h361d6406aec4df6ff4164751b52aa2244e40237378616d91704447c6c8a1ea7e97caadfec2ea187c5493f5ce8100454d1919e5944287dbe8e155d998ec7925eba768268f25087a80f8d50fff8bf6eb489cd474a9d8e5b2166746a33692dd94c14d3bdb7a9fa19ee3163cc10c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'h5a74684e1d0ff6b904e2d4d26c12ef6071b3f9093f9575bb397cb99859ae9825aea33afc834c0328ea9b11837508cf679b93d010eb29ccc5ade50bf1641ba8a956d2e851e13b15feac7d9599ea4220c8035c045c7c43283d98ebe1d49af6f09110fd4cdc74204a25fe5a601f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'h617853d50349c5ab404bba30ccd6b0f093828e1dd58ccdabc83bd2c5d02cafb7965ae35ab4075f355377d40750601114dea4c2fb7a4949bbc72389a44f0f8d14db91d9c3b4e68327eb0a39691122e3df4711aeb525a6f5fc5e84d02e2cbf55a2c3ff3c14a80bfd8f12c340fb;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'hcfbf5b096d3dd680ea2250ca97a382fe00ea48d976034c35ea3183b94f4d3325a85d5e3ebc75ef2044ce931867b8dfbb42859eb0852c2ed83f350b9282c9ac6b044f8fa9fc55651dc0cb08a14db81f601226e3119704201df1c336963a317caecf0625ba857d14aae37d2c3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'h1abd185be14117115be377d634920e135d56928cfb3ab10d8ba6e0df90452259af387be769ac8c28b029aa4cde4df525755bf92c927c3ed75022ba9525ac325bac409a82730e52336c2856b410b5cb811c760356a6401d4a2ebc5b006464d86bcb8a3db5eecd18953b4f9526;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'h3a0df25c218e4b649abc9aee23e10facb76ff53f09cfdb04100014f6201853556d808d4d46f8ed5b6edc3ad2a545a2fd76f67314a59c868a14d7c7c10a0b17a802e00abe6db1b303e28d9c6791ae3266c3044dabb4b8ff64905962fc3acbe4841acaaefca7812363fd53a5ec;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'hbcbec2b325a21bf2e0062e00f6bff411f765bd44fb5cb17e130e6156fd203db2db9d3de5bdc542b4322c3e0af7f42869549453862310fa7a448967cd4da673831506831bf18b54fa51e2ac56a625bd55d637eb42a2fefcb4af345018903417983e3f60dcaf2ace7da19ea950;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'h13534fdf653bed27bb5df704a0a0c2f035e202ce0ba2592a30b1f70c11735131d54c9ee263c78276dc58f275a2c5c77ffd092661f743ca9430053588f2a45dc0a8409cadda18432f2c6b3ce900bc6f4f0aaf866079206d3032221cbf6681922f7014d1330aa152437ec95827;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'hc17764b1ed9ed7593eee215fa00b1738363b38f8052b03edcf6acfdda57713a3c31a85c51df47a663921871ddaf83942a195a169c5ccd0289cd115faf2808fa139dc0419c9aac2c5a1ad8739e6f139535b28875f056cfa24bc4c2afdd106b47c5ab7ab3041d9bcae751c63a5;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'hb1a2c8b0ea124dfcafc8de330bf1a438bd7735d2c50816da46506e6a3f9a0975bf1be01fecf1de6261b47b6bfdd3cbe0d8125ce652d529a79403d64336e45510eb5cad0ee3cdb7440d47054068f1414dd8135f4d1c3ac3a18101038645ecb792aa7f42a3204aa1a704cd2a77;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'h8752d603a14cdb8a7fc39b4aec61ccc83fcf7af99d4810b0344ee137a7456728df032baa3d7d4a8c4c31fe6f356c637af08327ab283c0610ea85e1a10617ce6beda611ea0f3a2c56615b185043481ffd8ab8012d7fb6e55b95d089af2a206246abf27c32777050f6e4a500ce;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'hebd3eb226a0f4e62409af966e3fd5106b8f5afa5f4a8894c64803d97ac819890d337be672c9d4a7bfef5a3a97299f0d67600f6d2f64b4abe2bccc2da38e8ca0ce4d4518f0180ad4d14ba57b3a4dc48cb73f405fe6b31b7527b26d5d35e0454b26a0555f01e8b6102404569d2;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'h26ef0bf1636a08f607581a91616c2be75ba7cb8413747fe03e6cf550dc84459c11190c80301636914502de026583346fe5d4b426b4e30fceac3d75463cd9725b2794117740b494c0c026e71eb8d6dcc76c052e34bb1ef2bc6b0db181a2b8b2a03a176c462b2ebd577d8f7908;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'hd73e46911b17e49de035f12147289f8d38af4fdf64a29da9bbb0d527edf82ba138f724edda38051f3650e1638e11172c9cd4ef731e2e9206697798146597718c830824a5eb91f8834450e4bfaf81287f43909513d7613795942acdca7511f0c4e3da0a06d89166416b7ed8fa;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'h20667e68b49900b090d5866088caa682d33d7cec1aaa672f8ac115fc4bab0bd6297dc8e63800f6e2e9ee90e5cc29531d81332f3d3aa32e53ce9e848a9c3dbeed0efc743731d78f013e42c037ce3d24db9a811f0baf1d94a6605b7043d00c29170fae56269d0f829a122f3d7b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'h7a9b0b251d77a7410a290855e7d64c06b9b68e63d8504c2a83080ddf9c2d8444b00b7dab2fc19fd8928d996c667048d37b7ce982a6e20e57d2feb097653748745dac3771d4fcbeb047025e12d7be48c5027e297617dca85f34c93be97f2440a1a868919bb340efc41a6724eb;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'h81196f53d0f1a8afe7e07f5bd209e7d80f9e480ae72ee02b5ef37f4379251cbb8e1a4d5986e64c1f262281e62371354cfb3e435b80c55f0d41746cd1776fe1ad4ff5e2bd5d55b4b6166c8a84fb6dffd3d316d6e5808dcdd9d5c90b1191b45ba13287acfa66c67241ef930cd3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'h88b712bd35933be300cfd36726f744f8a3afe2c477f6a843f5cfa7d0a91b6a28905c0a72223be75f46e88b617704e3c34a3129b50e9bd86046a4c521c5fef817764684f6ec7a67ba130cf9957986e16eb46719fcbf64d2d221a65c6038f25ba15c6e2b7efc67cba4e5fa5fca;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'hb817f50d6abcd78a39a592f6fe52dc5f064b1ce5fc231c5f90449f13243764f87f27ef7ae1bbe2900080b29ad8273dd749494518bdc31c0cd12bfa624d1c79b349e1bc0087dcd7ab8256c3f5a2a07bf8f59e38be1ad95a93b2b70e3b74e31533580b13d9d478e4f3b8903ef7;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'h51e5dae767241b0a86566b550243d77fce78c6ac585ccbcedaf21ce2db13c5380e4b3614fe0215fa2783166d7639ddb2de56bb781ab3231a8f02bc652a5e19c79a00e8fe98db9d4f28604ce8848e96f5da137476140a243ce52391a9a27214b0f413bca4e5c72b7c3bc61149;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'h29fa5d389795745ea98a87640c852e1c111d4e5574a33bc0db87b1e83451ae47fde4c2d32489850478974c4a02d0a5e9d2e617a2d16b91773a5be85e1b1939f333a94af0286bcde3273d061b119d5ff19f92b1e16c6fa762925e3fa2a32ac605eef4aa69389e652c3a4ad805;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'h56c8382f3783144cf0b0b36674ea9158a063b825f737929e1693bcc8f8ec81715e7b42bc9ba7bfb06aefbb3a72349d0402e7d039f3b4718f184cb13e4b49cb51da0a0f2d85b61bed6f59e4be56e117fe046f56e60e8584105e20cda0c34e38a013efab68e8795866068e2caf;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'h6407646da03608f904961c3ced59f84db73d13ec559148e69b8f9f9b1de2e19e046ddf1657f89c8be0f11b75072bff01a11b81f45fae5ac3fcb6d9320b9e31894ddb6a27740d74c8e76e697f26db85db174f9c406772ff4336541507a1f4b6cf267b4cdae8c5a4386e3c375c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'h74e41e37805f4345daeb6b2e7b5524d67348618491664af84d41663d3d1c5a0952176809eac133fe26d427c99096c44c02fb703a6a7dc598dec1d79a8e15924f30df03c5a22f30d43fe57508f4312fe1350a996384fd4c06b9ec069d25251ecea129afac00776aba934c0cf2;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'h3c078d25a4583327a0f42054106298e24f055676de1819c593c8af9530947bad5f250677449cdb11f9a00bfc0c67143a7eaab7a24c80a5d2be07e94ac1144930d57d0a4cc8347c7ab48e79c6916861f12abdf5c921b30ae9fd6564030347bd8a38f836dc29b4e32e689acff;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'hb237b7849b571096e5450c7fd02310ea0a0c6428c2316fd7e31221a94beca5e4a2b8be510a9ffb868de7c95e9070c0522385ed79530439900b4db5766a64057ca4a2c42aeb00e892db5bb5ea945c611dabfaee6187db35fcfe76edd5a572a19479f91a313236aaf2ad408796;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'h9391a890b7db0884b2f03f84dd3c80cd4ccbf0c1210cee7278aa0e1a8fa6dc4e0fd2d2cbd686cd6115a18cc88c4ba32fa15d176d96ffbdf884e1af34f2cfe540609f6686a3eadddd77684abb9c0ed1522cce579f284eb8399ef9404b9fb628db543b9e77019f77fd939451a3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'ha0b85d7b25d0949c4769927578ef1c9963cd42f2c210f94dc5ace258457a28a204446dbe486d587511485db6875189092569ed9d3bd8ab44cec8bcff84dfbb72d9ee65679dfc9e79a3a194a4fab45a7082708f722cdf77b5f34b957f5e42a5906b616fc3005a469aadb1512a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'h8b920a336929e922065110bd0d3d4f1853376931b87306e289e72e9a8fb63c475e51c2b698e1708b8666f74d01fc775c6cfc17ae105e89807078b64e4b73364595eb61734cf4ebdcd81deb47c998437ed5115c9f343691bc03a1e7379d65337f35cf64538a8c1b6a7b98f11c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'h4b1e0f6b4d6a4483b4b8b50367f0326212053a010d95b9f85dfc084a908459390574465b66178274d02b9b3b9c0fd2ad3ce119c6fa33fa0b3e83f333f2937568806fab311a4bb857cb080810b71402f1277d86f0e7a54022f8d9be5c2bba6ccd0d3bb382f57cffdbec7a68b7;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'h3ab6bd77a3fa699677bcf360739b431141a7f06e14985f045b2bc0dc88d520df6ff04f717bd684062722a311742e0a7ae61ae5a3c081cc47c5fa2a715da1ee17e7d4aeba12bacd070b240f11fc679ce8b9bae3789471b7a435ce97aa046b8ee751d7acf78cb63da458834a75;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'h21a364df4d338502c09062d17c97d8c70b1a9ce1f816b00ea8f75cca27ed39dba0b6184a958d34980f176c98674e3af18df9ff06c9ceb2166753514a5aef810b23f21b28f3a3aa13b81d419d16659b69a9f5d1da27939fd639ce8e3980a09a9eb89387b1dd0d5623b793b9da;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'hc0ac0cbf4e1367f226a86e03d13508a99df3af6c35bda11c170c6a5e2d721e6053a40fd6ea516cefb3cb112e7da18e4fb32455b4081da311472f6199903d04a1e68faff23d201e64dd8d1050eecc257e462d3dfa8635f38ad7ad1057ead02d92e6361423b1010b738d5e669b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'hdfd543a0d8a719889839ab5e9b7a34465388a9ae2c1e8f3bd6d57b74682341f884387a7507adfedf9c6a0abf5d2342bf102d47fbec7e7d2d799ec6ae338e8d3940d28abc22e4606f964607a644a921b5c3d02135264d9a4c6ef46eeba36a4bdc0068624b450713d976fbf948;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'hd1808031a0a02f262710ce606c5eb0d78a6de0f38ac68177126262050ddb2d72ca2706d09ecaa35c83b157d93eacf9e19ce38250986767ac9feef12a9f742eb51b1d7c05661836d616031c419f2b2a55b6aacbc785f2aec7a2220da91d7851a1084b5b47f104893a8f31cec2;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'hf0e883e36b34020bcceba61299ccd2974fd32f04895ee1026c1c48476be0258347656a7a8170116f456e182b29073e91efa2237acfc5b3b221e8cccaf8cb9aa0908c76dc5b6ef3d74f315ff8968b8b3d826f90eaf1c00ddf85b0ad352587c3e435a10657d26e92bbf4fe5e6c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'h8549c1d782817115664d1e21a63f3d55fe886d8b0707c552d5025b26d52f738a0a7cd5a1037c6e594b972f539ee62ed2959d8e52727104d47a6e5e28fa5dd49d5c3e2686f4da31a55c89a87de104e078a1998ab7c4d1e3244d217468a81b1f5fb31745c577295522b56de6b7;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'h356a0d1ec73ac4f4e18a7978ae7cdf2ddeb6cbe3bb5e40dc47e4c3bd0f478de4e0f819883a63f42ee5b801f495abca48e2853bf84256f7bf44bdd73ce996c2831f1b9c0954a5d394e929bae1fdc4fbdbe9241797d8004e1a6f0f800edf4f5512880b4746198b14a0fa56e4e0;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'h9d90a8ca8e1432dcbc89c2c429d37027aecbfe80c31839c3f0c929fc8365a0cc52fba248344a46e53c70744e95e8f85217c5928cb1c4480f094dbf23fd5e51b6d781c53dddb1e6795d76e926f20b094114c0bf101e88e9bd4b012283f6f3034632feea8f5d4988ccd5221eab;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'h2c69cada09550f2283e434ba710e1287defc63564ec027665c887baeb567c189682ec6b3af9d7b78bb5b31f696ccc989259b09cae693f218434bc4b7e7b53e2ade3ec38ef0259328acf657bd656f51f352cbc3ad679d750e35f001b92c990d23e3b29d7f82b82bbfc5fa3b37;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'he82d9724e0de9451742a88202e82f1a37833fa7c6ed28bd83657a4e0e72ebd7342519880580e8751e129d9df40c2226fdf7585264b8bd529f9f6d7b2c9e0d40b49be50e8fd3fb4166fbf13b2f8e7c2732e755fc3590e52323a17d409fddf3fa4b1ef944f2bd3d798f9316606;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'h17d30d33dbf05af7010ca20bd73c12f17fb19dfd39a785685896ee22f7586e220b2c297fac45cd5e14cfd750d887d3858e8614b1ab898a14e11e676c25eac836db809b665780069f59f7f21a15e879880d3de08554f9db1f03179353b5f110ed7559e64731c7a50bac3bc4f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'h1b063c83dc343e13f73fe0b4c9bcee5aaa6d0af6ddeb2ae08dae086d537fa182c9b0bf071f3b173a352e86e192ced17d7a23bcf61fe7d24a8fe946ea29145929d74567d128085e32be6e08cb5853b1505166f16bf62ad719c9092c164e5710b7f7a2d1e35cfca61e189bbfb1;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'h8a762e2069d02313da5cd3e2449429da6bddb53932eb27a7a242fa3ddb0b1038f29822bace020d36becdfacddad11c5334a98498ddf67993d8cda51740f565a698c312862977a667629574d4abd964386834a6e8dcaff6c1b454737690f0c01edc6904469a2c0104d7124396;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'hdb57525f9c9b3948c0d44efacb3dabdcfa0bb743deaf662b51eec026bcfcd81264e99cb36377f22f824ad3930bac36ac69be8b0a7731440c5896dc9b340390783416d5a56843acd4a7b8688e31504ed2437a912f0d5529ac2ed60a7dde577a3d8d677e2214eddbd1c3b30ad0;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'hc87c5bc88f4973b350e0b0a43acb70fa77dab1373a8cb4f7959112491446cb3c732bf4e185316e3d2bdca0a6e837914dd9402dd92f6e6bc8e7aa357c34b9c0ddc9b2502b1441049d8207a301054eb66c2b1ce239d885029ca0dd562954528e8f1cb5360452e6bbd81e6586cd;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'h9ebb0bc8a036a3829015ec223ad557d4ebdf24945701ee0b2cc91d51b567b8ae24dd853f1128de66a9ece0a75bffb21335884defd83fb2e078f89de42a0242ea0876139b516dd76ad17bf4e61d4de738e2055ab618e212edcf912cd1f9c94a02fc4287face27ab15f41cd090;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'h62b6bead640aed98e2c66ca33d44e3c1754480244520b464123300228fe7c2787fa46e5d2067d0125976a1833d4a0d79d8a9e18773fba731e28a63a2d72b3d45b7d01b1bb5e64f2a27f74fac27c58d0afb953a1aef4542e177902694d3e9e19f3df834cd98adfe8be987e58f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'h6e6d9f565627fb1432a8ffff686a95cdc3f9f8c07dc349ae5159ae8e3d7ad8ea42f079559236b2847a79d8ae8aa6f87cd4f6a9fda20012d3a3a2b87a1742e409289dd53388ca10ca23499a2211cc81f4cb6df3e0b1a0ca0aa38d1c7c5d1f43740d532a0d1d68d93eb061f0fa;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'h56e193091c1d6f828910ec4315d1bda6aa3a4ec5781b892e4dc2c040dc2251fd07c640604d91c8e970674e4520561156f44703d510b35d491a0844579a039ebbcd29a7744474a2137a41efbd264386cf50e9809960260777436f161f6162167fa6334189e647220c6d6fe5b8;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'hac17389b19fc749b519c2b77b63f807c4f187810dfbe297685113cddbb14b788e0ecfb49f2c6cd05f42316f3c053d0a1d59cd1d993052f8774d7dd73f5bcdcbac6391963ad549008b648c9847a97c78f693ea56fe6802f8a5289e4a61b4d1896852aa6feb6eeab1ab5bbbe98;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'ha6eab35967325700d5828f8ff1b92b761f2d078a7be4d16f68037813eb5d5397346a7ba8047714594f2a53b84ffc36ea819c5923072f1e463a265894b199bdbee4ea6f06124ad44e7b419196299079e410ace0dd6dbe2c71c7a452a8ab9c0df21a15943cff54b2a996b0df3b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'haa6f7505fb156e0431b65a58966869f657d7fe1200725e4a6b01a025f9bbc022815404543d743e883a55b1dd6b02f45cedf75c12a0b0edd0e95a1bfc6aa73bee2691fd42ec49b98342523a633cbac8e1c4597caf24958dc17c298819f07ae1e5d53a7600491e77a0605ec0f0;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'h98e0b53541a7093bb412d71e3d44ed957cd933c2414229fe4d4ad2eb28110d535d56b2afb45ade1304d43653b032fe5704beaa9c2de1ec9b740569ff5a945c90d7d316bd46e9688465a8c2812e844d8af8390a1e71fc29f6da4a35ba7da8a98c5fa9d8be1e51d5cdfc40dacb;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'hf2d1ebf30eccb722a34804908c9d5cc8951f30b9cdee5850b941145a95fb5b5ee2caf343530847a79a50f74f51935e5a84a4835258bfacb9955cd3369abf0001060877700e98a56155f75150e9dce5da8a7eef9c70fc4363c52423ae37ca0c79803ff337a955c1be593ef82a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'h7bd12ba7d825deab847e42b7405317cbb362327cecb316f75c9310673c6a4e6d3f685348f58375114ca4e10b884e2cb327307ae709dee7b0d23ead923a50489249031ad6081d76e4d67e6ef1e0ec70a23cdebbeb77caab867cf65b11d2bbde7120494aa0843541bd068156c3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'hf5f03b8c9233cbd8aab8b5e0287777f4eccc454524d3b9edb35f83858e5498b977f8d43387e4af44edd19ba66b19cdda5a0c5713751d0afe768a8f62c18c025089d1646c1e159637a191684696c8a4ee1b8655ec3e419dcac6cb6afdcf2d6c13f925a0d412081d3c5ee3da1a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'h6068f9f660a2249865de02828f3e52d342e12e99cf2a42653240291cb46726f796d70faa0cf2daf76ba06df729bc618985fe4a90d779c68484fd8b492a43a79dd2761f3873134041ca3d87f56644551cfbdf78122f82c33b97d2036e622d319dd8b9030225929a1ddeac3b2d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'h7099c5954eed644fe549fd8ec7ca613bb0bcb80b4faad081269c4409853a2e032a0d4c18d17490be4e7de18ffe51f671cf96f780892f80a5c1761980396b08852f4d88595e702a71c6a5e80298a9a23b2ca0e968c1860bc78b46ab6316f7ee4ac292c96b17b8a4b8c966ef93;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'h45aad152e5b04eea291044749ca7579996c1e2bcc994e7fec8572976966557f61795dc6b73077ccffd5a571f02b33d8220bd506f6b63c8003e270936f212ec9fa6027263e3f10ec9804ef07f610c795ed892f102a67b6fe6e9be663ab0dcf33ab169dd094534787e57236382;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'hc0af523d5d0a8975c1f5042a94fd0c13b31744673025f20d6cb5df7bf2e476528ba77c874726b51c90e1c4160a410ce59b616b2aeca4ac00d5a9b111b42fe2942739d2a50f4ce6163d9e7d43e1feea241287b5b0f6c43a653e17e5799e91540576f5fa89e61058a0e3a96e98;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'hb9c4f4776cce7ca2a877e3b8e5b400a8465637bdf1bf0163d63ef70a8143877af7bc686f80ab72e17c69fd07e1239697b795f29fb7febcd92a82e1ea9b93afb440b23562ad8ee613aed15dfabaa8e390147704b6b87babd29c7389ee670673a82245d8d381d3f3949194d751;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'he6c882c58eb87ca76e95b6c0bb6d8e6cf60415e48b398f168b744e28b7f35881ac848c7178957b51619dd6455b04094d7843af634e5f2806e403c8b4e899225e324e287f8d664657edac710f4450e9c916ddd08f68c69efd28aa73df4b0899a35dd15b7e993526922d0dbfe5;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 864'he5b8cdeee1372b82fd78bd60e85ce2fa82c6c75a8878b98bed85e635b5c0df2411b366cac23121fc6eda46f2a16c11814ff5914099c6eb3ef35b1303e23c504e6e57a3503576962ec4f528c2daf18be18b5b905b830d4655fb1b1e5a2c770ab93de7b9bc72728544480bbbb3;
        #1
        $finish();
    end
endmodule
