module testbench();
    reg [11:0] src0;
    reg [11:0] src1;
    reg [11:0] src2;
    reg [11:0] src3;
    reg [11:0] src4;
    reg [11:0] src5;
    reg [11:0] src6;
    reg [11:0] src7;
    reg [11:0] src8;
    reg [11:0] src9;
    reg [11:0] src10;
    reg [11:0] src11;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [15:0] srcsum;
    wire [15:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11])<<11);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hffffffffffffffffffffffffffffffffffff;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h53f76f3f539c3df44034d375631d4c201424;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6a84c87e34138a677cb5a889a80e674734a7;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf68c8a7f078c6157ba2e6e6446baef8d4067;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc21547115d3ac7926caa1b583b8637b97fe9;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h62deb92760d489910164c7e461f598bc2f8e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4ee9106715ff0214ef6dcbb1119ce90581aa;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h40f0162b5ac2fb213af794459e237e4ae67b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hba5b046855749248d5afd1826b329de81133;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hdbafd0ad09a57672be736e8b5b4d412be9cd;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb2ca86452b72c4053de8fdf8b507fdc3cb3a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h56c2fa092b4c5e2e7bbc95091cff6c919043;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he3989f1184b5e9488acbd5098ae8967c88fe;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf8aa36accd0860b0cc7a0f105f8f5c35be20;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd3446c8e29a444c3891c932c6d41cc02e0c3;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h44520229511d35f3a5edf086fc0438bfca56;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6f2a1a148a8c7c46d23f05452fc3e2889d24;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h73635e2fc3e04095fe3db4db25ee47061a5b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd8b39e185ee0f5a162e9ef72282aafabcca2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha613dd6030507878f07d437b0bd38113d975;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc73909aed89225bf9aca1150c9c1f3a86c1b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hcff2a8175b98c9f67ee7d75a2671be5915d1;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h74938856d1a60cfa922f7299ed9fe923ec5;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hca0543ec9fb4e524cf31d553f09c54d1f40f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1263f6508ef7df7dfafb8bc88e44cfc0019a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1e4da16e5a1656dc0a4db5c5cf5d9e0b2e0e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hdcf8c6ecdb6a5067792e3bc5dbff8926ce5c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc55618aa41c9587e7a78a5d0846a988692ee;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb3f4ddd905e9d808bd61a3c8434fbf6d01fd;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hedaa6f8cea8ebd55ad8c8185cfff22c5b2c2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7ca72b864e510b36ac51aa07ae6c59123577;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he924a50bf8f22bbf8611f6356bfcb79f3589;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf66271fbe0fbd9676f2b456e23081b653f9a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2a7e89e926950ef054ac6657650ccd2e19d6;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha88e9a06b00ad1fc75993817b4be4a0d1ef;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha75bdca4e14f19fe16601492a2008e04cd81;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h44431a87de73f1cad09760951560f7c47a4e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h10921e10aa034f9faf395617b31789dfbbdd;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hfff97b10734b923793290fdfa11f1e70fd7e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hde040a6b961d85d9cf7fff2ba53fc3e9d277;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hcac04b7708f2093397154a6fb9356150cf48;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7f3748137e343100f152ab396aa6f0f0ffd;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h229fb1f5071d7e3693768cf8d4a658123572;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9671d83b9e33f01a08ae1b607e82a8c4883d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbcd8f9a74309cfc066ea0784c55260209852;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h12f5c33a0594614df6ebb7a7186f5793c841;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1b89c5f96b5a028c054b62278ef0e7285f9b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbddaa5e041295feebb7d4601923177e1c662;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h104acf40f785d18cfbe0e60e592674b18fde;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha34c243219b5c27777f677006ba4ad3bce17;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h70e60ae6c9f604850e91b3f63ea31a48a5e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd5b8db7aab89ed17f6f8c228c3ce161a0790;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha29a1b7a9bd6b7ebc99cdd59db94b5ee8bc2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5c21d571520ade88ed7d9dfd2aca67544827;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2adf1f0eff70d40d0387309b3102b9dece46;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc204b7a3ea64f04276e46c4a08766b2992c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hfbba14a841e901d2438280c47904ec0968f0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h370e8f491b7b744c5cfddee042474419fe99;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9e89a4f4f9555210c6b14d87bec7ba4f7280;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h999ac57f1f61db8acd8eef84e5e41f689649;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb47c350fa65ffcd45b932c40a249e2db687e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6bc4c83f6766eec27ec1d18c899757c4174c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5380e8b83ce25715543f868356c49b909776;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9fca309ce13bfd9e7f5350f917793773adc5;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc9d1fe536d629afa67b9d18b3412db037a4;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h979f63040087ab40d1fa85b6e769ab8eb4f5;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h73d51f45cfa0c28a4ff1245dfa91fbabf47d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1a2f4b44f16e759ef0ee9f80534538cd311f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3d4b04e00eb0fb6648919513deaf09123b3b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h704cdf25ec3aeeb19c8af1915a49276dd17c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc73a1f3aa2ac97dc974de6230d8f667ce9d5;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9df024edf0476332f123d804001091efa6e3;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h747c85f140f1dea96fd2996784ae7882c37;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd717a5b3da9a0f41b6027464fcb5063a1ec3;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3d9a442181a792574f4ed006f2e2a6633567;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hcc7ae5c657c78b5ba9c3a313fe03506d2123;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6ee5f82824ed271200301066e95323cf3560;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h275675f186726e5f5a956c67d9d7ffd10213;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2267e2ba4a75e93f87817bf1d8bff91d7e6e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9ba5a7b24c73d73c70ffe0d40b56cecbb1f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h89b7f500fbdde1dfcdf7a6bbba288adf1c5b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'had8cc3ed3c1b099e2395004caf2fde31467a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h80e331906133a89c1f6dc1e755a23575b06;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc1d1ecc926ddb15d220bb18a4c0258193d90;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf0ca71b0218e9ca4a229f2183b1f332a9abe;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1d4a00989750dedd084ba3f592ae9aa579de;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h64b9b73ea79309742774e3a794a6c8ff7e0e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h52c6b75c86d696e5ec66a5454af1d391c79d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8120f5ab172ab3a0c048896d58213745bc6;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc2555ade84bcc3da2a9fb48bfce3ffcbf335;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h34b7ce22df8eac7c81a11efa5690a98ec165;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hac2060380f9bf7258fc33f0d8cb16f2ba645;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha6dbde0ba3ca52d43b03762f3ed93ce5868b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h15517000167b8e2fd0ffc8704d43e27d9f9b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbe1305905a5b8dc6f9a40d5cf64341b59280;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7d1cde143fdf1b6b33a0d17c5d43fb476f05;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf41ca9ca6c2ae361b889d2527e7edfe2c197;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h24159b39593ab84a55f3f3c723a511a3d3fe;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hecece89dd1a3f23700b7bdecac4eb0d739e4;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he12501bc27802f4f468b7d0bfaea46a3470b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7dd559be5e0327580489e2c54d604e32c5ad;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hade86c544e0654a35a545a172d1a250f5ad4;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4b8c22bc1b2fd9720e3171fff6a5a7b8cf67;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h93afde56539f73c260265e631326401eadcf;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hca54cb05f6a1513b7d7c6210b813bc907030;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h21051952e6079d02e61e6bb739727b1dbfc1;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb0a170650bf3e7fb7d9900a44ba1250d4853;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h367addd87109f9789e6242e125e9f39fda14;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4f4aeb31cca44c2671a319b512d69a663979;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7a98364742353c958b726e3c4291c5cf92b6;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he12c48a6def31ff1f91ff7ef9a56f7fffb3b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1c688657751b21663280f88f62a84942a2db;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h14913412e082ce86136803883c78c7f444eb;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h51ec15dcc9bcc9dc119239c93b41194446c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf3f1b5a2eaa6c97ff7a894bf80147205a106;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb4b64c73a8215fccc25c12b06ab5ee889b49;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5cfb13750a0aa620812edf69ad3c59fdb198;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb3af0cc1696a2af9622e7a01b8fd44f1d8f9;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he58614ffa1f91c48724af8776f08892f2179;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hfcc4b6c3cc930069c8a13b13ed741827b782;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc643f2ce8ef713cba53a6af6717eee0ab534;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h17a0709b27468100c2c92da14c764a34bf1d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1dc55015d3a26bb9a2e50bf51d867c47100f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2480903350680187a8826598d53a5549e64e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h77450632746d5bcd312a9ef599da8db544df;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8aa861f367ff2fe88224d75f2392eeca1668;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4414b9de5ef62aafc8ac6da1748b3b79747e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb4b9e65ac8dff77f24fc518005622fffde79;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4e49202ef988bc122ea24525129ef515686f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h53d0f6dc8d127b0562c92e7d3c7e3b48a614;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6c83b34630427e5c228250a8859a5019a0d6;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h543b31e08c12beee17ab6760b0013819e98b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3e0aea6c47ae117fe45783b70466278d8a0c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9e8a253fb951e7576f947ada2e4bca990634;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3bd8ee3798d5dac193513d9fccf464b94ae1;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hcad97ebbee4b86bf0f32c048234aa66f90bf;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4c20962ab573018d59c4d4254b82572623a3;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb4b5169e86eafdb99f9200e393f16729956d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h70503b8cd9a67a3c846601180708ee8d35f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3d747530dc61ef558161d785332077944231;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h42ff92b803a483eb25f465086a7dd14a157c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6af1b66a6eabc6afbd19c100a77590cf5f39;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd6eb1a621b649b8cfa15ea962258611c8a63;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7f26e1a9fac0f73ace695a40d19a59f75568;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hdd36a5980de502ec7146e9ca4afaad33c461;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1bb40a5e226fb832cdb1b6f9c4431cabd341;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd41b7f3ef857f222522cf4c64effd1d7b76b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h513d478bbd60da3a18eb5d802c80dd0e80a7;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6d45f7b651a9b565686f333935393751bef3;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf50dd672e9f26137aab03777a9db5d7a4a39;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hee4b7e9c7a7605cf877c9267081e819f239d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2b79dabc8b371b341acd77413a255f938e9d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2b00d746a802d422aabadd009f945783e13e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5f2de41e3f70b1b8cac006217804afecb937;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha11592b11b96a4d46454bf7e3c902e3dd881;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h97e78debdba20576da17ae6e73d2ed7422e3;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h68a7c009d8c969ee3b757bc4dfe901110770;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h509c6b42a335287c3b95bbca08483f43c7e4;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4ce3a5060ca8fefa5eca4a19c16375b2137a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3d93a2f5cfc7bfedd14170ed556c81a8d017;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf5a9a9fb105b1c2edfda1bdec1bf773d4e21;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2047a74219885eb9951bbc5de6619a60f1b5;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9fd918e28d7b909cca929e2b1b05f39f96c1;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9b06d9cd4d078b5fb444c52e87f59f81806d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h50603326b96a1bd8fd73c2ebc814bbb5fd4e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h787dc2177cb04916200e4ec23396b8ddaf76;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf8fc995ee1be92536f59a8fd6a9fc9f8df23;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf8ff1d11cdad2efd34e3fe717e3bb97790da;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha55ae689e1b27e20e3b5f4c3cba4a70ec082;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h855cabac366673ae3a7461890cd5a37c3aae;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h18c4319b35ec7bb7403caa2d6e354b335955;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2946687cd9214044cf7d60838b3bb3fd16ed;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hfb97bd7e55e995f9438a3b82684d0b5b202a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h886ebbe672ada84519df7a157fdd89ec5819;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9c11e474959cf34051af2a1fcbfe217deb0c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he835e4f4534273a93dc5a0a4e2e21e2df563;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc1ca9cac09d827f8c5dae4d6547e869dc34a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h267b793300ccbe71bdf4e85a91497a0338f3;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb10179f25a2d120cce308024ccd1ed24c5e5;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1ff1ebfe457452b36b16e210808496c22c82;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf08125d4a5bf4965037418232699ea783978;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h51ea1ab244baa526a01c26477fc3d7c35518;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc3036ee30f14131f645d34b6afc78cebed7b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2c5808a55239a0e66a4689ca317eba59703;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2df055ffc7cc6272270025aa7e5af528e58f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h16d94cc2678133fa78262ebceede1572ff1b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h852b50f38fef7f52284cb0b89a581fb0abb7;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h899a2ab17a6da9ab3973467941eee2b78107;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb987d375c25ea6f3d71172d07c512165dade;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h54a3b39cd08b4e8db208377c14a5dc2519c6;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h620c50283ba7acf5acd622bcbc43892773c6;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5d1a2329b9dd09afc618603637a49517a34e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h47ec40c741c0335977c6d7fe9fc93200a73e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h50eca844c7354caf2019d527417b4e358484;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5cfb22a55d2bc86bfa2ca624358714c7a530;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7bab4b10aa3580f683533df48effe08d517c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h45360337b785a43343c212eb536d4a14d5f2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h26ef74a1a2ce3702e468edd63091b2ae70c3;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9be72b77e5b0c5d8721934c3ca6eff969bfc;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hfaaba508c4e26e543510a19c89c21d07c7f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha7bc9ca003fffe458d925499762db8a06994;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hcb6763a2e21c94e93d86fc085373c01e5597;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hea1c8c59282f4ba84c96fd4435ab494e084e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3e42f474301c5a8db2cb0c2bc9d9b9855576;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd51a886400b6c4283fdcd32537c3f0543496;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf11612e22d097f0150743059006dd10a730c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1633ce80432cf27da83d1d87dfc4c15ad1d2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc6d3da53e6011ad91bdaa87e004a9ffb72a9;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9730666debcc2dc2382754aaf76d613ca0db;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha648e4cfc32b290902a50aa2e7f96319084;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h573f720bb5048ad3924206b9e238076b159e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hac0b97165eb1e8a8ef2c7c1185ef469b3683;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha9f6b39f73d6bc45fbf42511a9ee2dbb22aa;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2e9db0fc60fd4dafc25e102511a5308f976e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hae4da0562a8fef8ca12606b1ea975b64da30;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h63ef86e165edafcc3c9a7daf3a1e48c2cbcc;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hba126415187033c7b29e85f4d511989adcee;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h34b3e9e4e5571f0bdbd78c7f0718c9f3243;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf8503dbf5012cd48f0b34dcf44f99144902c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb4a0bae276eda273494f7a12b7297097b84f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h61b6a2bf8fd45aeac1868ade42a1b89b300b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha2bca6e336e642a2490980d9e64ec92cf8a7;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha5cb5efedf1ae3d2e868588b87cc80bad22d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6cc8d5abe3b2ce9bcca526c4cae20464faf9;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h85ca91afcc438fbce0ebb8464e7dd95470a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha58354180bb3caf6b428afa7aa41299f9651;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h141a5cbfe3fab05e40a9cfffa3877b6560be;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hfe933a9ef407277c918075c198e35f0e48a0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5593ce4185578cf4746ae9a0726ad5d511f0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha0592638c16bc9ae1b94cc5b00cc4df6687b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h875ada85905aa5f41de4c21a581f2df63ffb;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8f6e72e9a9fb8676ede4595959e93e23eddc;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc031972a097ba0db7548961d5b221c5c9570;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hfa721bf495b536fc932449372e100185e015;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h83a636b4fbe851b8bded5e96a98895ee12f5;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h45b51fd8998b253fe788f769c07340673c25;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf92dc9df027018650aae6c8db97218947298;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he12839f2aefd3ce89c219812c2ab30b35a15;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hdb783702227f72b7596c7c38f4c59bb7e02;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h187371e4a4d55209f9c07472fc7857f203f1;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hffa8338bfc79f0cf3f1fc9aa1508acf0512d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h51d743602ec897889cab04aa5c0cadc30f9e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc406dc2fc357b2b04dd9c41faf3ad7853605;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6614f3f3231b5ac6627dcb949326cadaa456;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h941ebfbf2dbc8c5513c4e1c3af7722265e45;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h67563282773eb57f8a25ec068d44ad68d9d1;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h75477c8a69a4cb530932cd09a309b8bed4e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha44b5f3dfb6898009beae8a2da5634d1dc88;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb1adb0c068cc7a3cce30127251d2093dddf4;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7c02d7f29b8abd7005eb068b3cc706b127df;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h593fd727ef132bb59bcc110e1dcf10ee84da;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb6d6033c2115cd08d0345900a83422ec08c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'haa735bf4512aed003ba04dd4c7f07df165ce;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5e1d0aab90ed8d670a3991f36a972fad2b2f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hdbdb9ab3f2844c941d1a3a81615bd91f5ee6;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1bb26129e56e2d6eaff31f82799792bb682e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha1dde8c9bd0d25e6710b3941ebd1ca07317;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd95a0322c8f397835678c7deb20233e218a6;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbb97bc9dd09195739d7bdb23cdb42b9a33bd;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h60e1818b3a21467a6ef7f3d8007ea0e8a2d5;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h55239364d26f0783ee4d3bac7d308c19838e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1a080cdbc97429aa47b2cf5a9b8efff5f3e1;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h45172ba204bf560f8e2661e3954224374162;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9229a6f3486bd9b1279278913de2316808c7;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2ae33b3e334f5696abb105f0a8b8701fc94a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4f5dce5af4e9b6f682179d85f865262be59;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hfb9714427ef06e9abf54ec07969f733a1289;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc0de5012a0db81622b5fedc1153ce1761e5;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5cda755cacf13b7b115fee3d3705c4dceadc;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8bec8994faecc98c1aae25888eb8d80ae95d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7e24c0ad42ce49e6c1cc73166d9e7a826a1b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1ca722464910f3536fdfe7468623061325ac;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb427bb6bcfb3140db4d599288c1e89c494fd;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6f97d9fa3cdd956b2542f7732dfb9d9a792e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1eb466dff9eae2f13e844b28f2709f670cd4;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5172d249b4f4a583dcd91428ba0c58cda947;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h537063e0674e9595c46f4e112f31ccb095c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf03f521797b9d6ad54915e72d11f550b2590;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5668080a34daa2b53b9e99d9db3959ce27c2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb6fdcd5ca5d6788547c7cbf85fbaa15d6fc5;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3ef9ed2548ef7d237589b5df0b27f97faced;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7322c477cd774f8545d7a585fea82a67ed4f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h788dab9d99bca1565fcfd5c886db215bb00a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h37ab782ff690711d59cfa077efc6d03c758c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7ec20515184c1a6405acc00d2022fd1acb01;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9ecf0a0dd7fca8b3189dae81ae588102319d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h36b279bac63bf7b757cc2f6f0f4f47d68ce6;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hed932293c9e018329419ef151151963861f5;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h661d4b359b119242a09bc8606f613db3f112;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc7b09f0bc58750cd058ff05a295c3109809b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h41acadeb56f4b26a660279409002274d8afe;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc8913f8876665afdef43112cb95427019a79;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hfba8444e0ba3d9b10911917da3477700a638;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1dd1f86c495cdd493a5096ca60dd9674709e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8eb8cf39c76aa9cd0523cd76bde19caa64d4;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd0d339c41b3fb350a0cf97d932df7b30be5d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7bb4bdba5230451a09969d82fd8126d5fbfa;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he7f1fcc39af57ed41c82abc43d90985efbcc;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd16948c006322d68edec56332cd67fca6bdd;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h954bb80589968dc839aab3ad82cc58a6c809;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h16a3d3916a0be12f5bb522eb6cb60ecdf879;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h242a3a2f4f756c9591e668e3449f884357d5;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9cfd6a274ce5471ea532befe12beeafbd317;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc0a41808c5074620ee3b7f597ddb5e4c4d71;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf4eb6deb0f723900d372cc29d4a53fe613e9;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'haa60c56d1850a131905f04cee0fb76faa4b7;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h723d212f232a8f85023683a97474d3dec010;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h773482e027ea485485bdeb90abb90c6a932;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd2d382e1978a757f0aba4a71c4ca29439aa2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd0b6b7474d1d9bb62cc9f9db7d7beff53907;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3f957db1945392b32f482c6269d2bb03a956;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf03109c8d40062bfa49122dcc516bc63012;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h68ce9a2d700a47e81c11d67517068562522e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd4c924050408ad5007a1448253053b0eabe0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1bc28481f871e66b8b8998e222cca842cb27;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbf53705054232bd7382bbe9a72062244fca4;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1eb46df4590ccdaa474599c7c10eaf0864f8;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc17c70ef43043bcfee6300ffc89e71e57578;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h185ac4183b7a4a4e3f33eafa5e4dc98e8757;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h387436cfd2f6e6fba1763dde3550dcf8e24c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1342628ada8fa7abcdc16d0c25ea99e40d0f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8e4faa649bef7a7266dcdf793d187d66f15c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4d311a6c8e0aa2d400eb3ecda7e258342ef8;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8f05f4d22184938408c1bb1407d02218c37d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4182fdb4c27be910ad07381680aa5e1ba831;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h90cb03fb318c37b637203dd30a3ffef15fa9;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8bd59e57334cdbcaec81d4b8176894a739a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd87ce9af73f87219f25abad3ba7982850831;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h20f19133a02c99bb52b5e81c1f835266baa4;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h299e3edf3e91135bb81e85b54624734ae690;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5a328fe1643fb69869d019eceedb3023bb07;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd2d1875bbddd58631c37cd3dd035ea74da7d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h87ff9fa59885802df1116fc60c9733df07f3;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h210cd2b17912514a07502a6129c5fd363817;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he130893b6f1850610a2b8b49842bfd7ebd15;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'habe45156f96b656be79aabcb979555d4ed3e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6384df3924839e20c978b7ce500d933ca073;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd99388b39017a4f4d0c7216d1f66ea2afd41;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb8ef59c9ffc8cccd0f04b8c61b3d9da19e8c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbea9e7f8222a8c18e60a2c0343133d849344;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he246578988bd48b4f3e2fa587dec1ccc818e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h686601b928b1514da8dddb1a0422ccf04c94;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8e2d3ca5422ebec13cb9bc98b765b71f35e3;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hfd6c83093a666fada42f5b0e58bcef130dfb;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he9d74202ab7615cf3823730439d535a9a1ba;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha407f2a5f898e4478598a6e760a6942746f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha4bf906fff6b2b1ed88dc52aa13b8da21f6e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb0028b10415256d7a69941d7870ac1194ebe;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hfba06f49ff7a412c6a9afc2be66132f5ba67;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he54831abc43ab0f674082b069ec14879b651;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1833d9224b8f16d394332dc6a8d23e559089;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hcc5cde0c12cbdbe5789bd15aae254fc76b66;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7535407f6d48804666b64f8555f225fca532;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbcdc40a3d2aed6ed011b153868ee48e1a311;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h11f3f546973a52c4a6801e80ca35024379fd;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h69e8b7c981cd047234750784406a72519282;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd12b6cdde9c60338e3c23c4e0d99d65e5232;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h94e9fb7f1aab9cce4ce0a8ac8c2e7c72e5ce;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h358ea69e7d813ee74b3bca1699067f81c489;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf40ced8cd42315ab5d353e5c22c831888631;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1afd810900313342aed497edcac80f6b75aa;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3ad13ab889fb8293807194b0511e04de34d1;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h41c609b52b6fb9dd48306e070887bb6caab2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h986ed2fdbacfc5c3eefe81232f425de7cd36;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hfa6f02606d9ef65ffcb43ac7f8fca7499ca;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc8d7052a358e30cf85a73c3f77f7c7389088;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha7525c7bf8567a4f4a9199cd64ee9aefc4d6;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4b95aeaecf92c9f5248bc4ab634614a34290;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9adcb131375710578cc68c1a2baa250f3496;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha5b6851ae31f6e8b627f92be013d2bc08bc5;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha1b4f590c0f9b211f8f4ead60938496a4042;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8971611f2be979794ad758f31751f50b53e5;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf9a54b0c0ad75c9789077259403bf035661f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1185e52b6f2ea333657492f6436fda1bf3b5;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h16d0bf14968efe37c3061607643bd7e69bae;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h102499673f4a00fc8f3afac253d779e7608b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h54148f3f1935dda38db6dce543befafd1418;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hec29c14a2836d9fe3c66641bc5b9244ce7aa;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2e6fe35babdf94da362e76c8c218e0edce81;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h87800102d73f31e4679d9d8da8881785d531;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h619137e915aba3d3d2f770d8302a715acacc;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hff14ce36704da43060fa718aec11bcf4cdd7;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5ee91642a2e66f88760adec37fe2cec3c34d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7070ec27ac4ba680d743eab1280ff7803b1e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8186a2c46d82aaff903ed433bc43bbc8808a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbb870f45efed9386e27b7e98efad391f28d9;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2ed9a28ed3e8abe6b88aa27ac711be75e5a8;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha8e942f3275f5d6d9678b28335b4fdf93f53;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hebacb5edea4f6ee1d64416ac569689e056a3;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h72f4fa2399e721d15d1c7fc6fa4f407a9049;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h84838bf63f04ea1dbcbbdd21dcf74086f648;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h508bbc98e3e5ec584f4d0bcf531195b8834c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h480b84cdcc1d7e83f53c5591582c1488f2a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he90db7ee65c54d67999624c642a5a5ac435a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9dae66dd26eeee2a3f4dc28a11ece9836f5a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha0fd51a5cfdd035b3c8e99baae7ee3213cd0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb035b04d491e69d6c48cbf59075a63be8322;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf4c3708c71c1be740d8c9414920d7d14f05f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8f6d8f31b1776096835d7f134b26016fbb9c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h55805b2f663121888d895610e74c9e6c4ae;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h899dbcf115ae67460edf7aeb58b677eb3842;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he2e5987276745659ae59fd8ee02e92ac2696;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h36406b56a1d194b62ea679f8eee73a808df0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3728fdfeb48a56b843b0860b93157509eb0e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3ea0a65d081d6a64dd8d159aafc89e89d000;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h38737eeaa45747b925ca10b258c8c8040308;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he09ff94833245bb05debe2d0a17e72b82ba4;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2b2b2a7cafdc861440865593bc3b6246b295;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he2db17380864935924971a9ed5743d58785c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h681f217bf895be444cf65bae00993b989792;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb79ce020fcb80e7cc3982360b71975cab372;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h830ca8a692003a4736e34e6f06399bc50469;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h45ba2eb0cb263d98608d4a48b6e9cfb24f08;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf87daa6422c1c33fa7d153d68d956214438b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h33af485c9df71720e105ec7b5d80d3f75ec0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h13981614ef07defa94f3630a118baacc7d5b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9f0588bbb5ed69dc138d63a7b843f7ccf3bb;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf7a6fe536a3ea224c3bb6811e8397ce83b54;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb3848d5c248b3c362fe0555f7a709a1f3b77;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hdbb7120d6f4cce6804de1cab79a73c96ba22;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1d67b3a394e4f9a00b5a71e4d7bb12e9d613;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'heb0a4d04bd131c3324d31473aaeafc28ec3c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd6e5a9196b8ea13deab4031f452093f57285;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h18f4fc223f42219527deafd785c424379b65;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h19c11f63d528970caf37fd38d7a2e02dae88;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5711603a9c13b05f52a5b847cc8990e7d773;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7fee955f8bf3dc2c999538d0e9c0573531b5;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6770f20299d4c1d5aee047ee3623197d8c5d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9fcc0591a02fa8d728a668aaea32cbaf40a0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha63376598ff43bb2b333455d013af7d949e2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h591af1a2e5c20558073a6931c54aa8399201;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6f69c452decc8e9d8e7ad69b7c41fa3abe0d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf046fcb31d83bdaf127c9d5408592c13a803;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1b043b1f24cc23a2b6c39de00f28e40de3f9;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha5df9eb30718150985a354cb303be520b751;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb22889a6692d519a2eeaa7eb48654ab2ad4e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha600047bac57df365f71386165926739aac9;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3af356f8a6157198c33ef975afdb4aca5c07;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb1670d6faa76943e1018d00c6d30aec64234;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8a257c5b76a36cbdc6990d55f3281108b9dc;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h44c7110412c32b9c05b7a3c76ef023a12f0c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h170e2f76e199377c81408f13efbfceaf31b8;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hcf1d359ce253b93bebb58038a9439f9584eb;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1f384393f3f77165ced384e9fff593d238b6;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hedba1881f9be7ebaa05017a6b924f6995ee1;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hddb4168e81a8ae7b8d618fe87ad7e04dceeb;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h25a98574c529b37887d92881cca5429d26a1;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha25de53570722a1cc76573853948efbdf9e0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd34126f604fe40d6ac55a14b6863bb9a0a5e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb0b71f64d8636c537b9aa79b434a1c897c07;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc3590c58d77b46656e0393396feb88e4e4d2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4f88443a16692c0279a94fd79c91a31e1cf6;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h716595aad8b815e0c582ac97d4265804e30c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7641ab14f66d895be5b72f890c7678f79c7e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7c85c1d19b3d5eb79143cf2f3075cc2fdc45;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5163464395890fcbaa644d95f102b66a3d3a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2d5eeb9fdc0473543954bd69420557717028;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8c9192e19173fa7063904a0cf4a4d3c66562;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hcd2b6d560c2aacb72fa61ed6304c69042f0c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hca9d841f4cae1fd8f3ca1250650fa4e9438e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6e48579bdd9769dad69d52c4681766a1ce84;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3bf3260e1fef7d32e16c752f62d1ccd22c9e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf9f32740b488bba30cb6b3c880de7398623f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4d2b0d44c17ceb46c675a7c189fb2632ff1f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h56cf24bbb353d15c725b94533ef44cae713f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3cfadc4701b1b0e2404c5162cc1d805a672c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8e8b9438be2ab2b1139505ce20d1aa5d46d4;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7a4baf45d792ddadc410fb9dd673f8d9bba6;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h171717a9e9687f51873d01174081847c8b87;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha990d4fdb0f5fe337fd1ab122c143361a4a2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h70e48df3237626c82f9e4c7f4e221f08a092;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9bb14da6835cacaf778611342743c13a0425;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd5a5549c3791acf2fb65844d09eb16022ae6;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h18456ccdf2a3a73cfe1e1652d4a15e9d5297;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4c93edd9eb85cff4d5bec2b3d7e1cebf67c9;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h58f16989807c76705a5feabfcc9530f464c4;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h497f6993bf43ddc671d4080c3f5b0ca0a1f3;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4047f15d90af6515a2afe25459e5a6bccb27;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5712b83e3eea2943b9ac3e613c9dfcc75540;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1535059525be0a91da0c29741ae1e42ce45;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h46ddf701a6216bc026e4b28ea3c7d6d04669;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8985c097b69a66a1f7df8fb7a44f47ae731;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8b41a0617852bf359372839fa056cbca4055;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h74138911b5d5a432b463b90aca4b5d159cea;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h35f0ef59a6a4c3ab62acbb49f2b8cb23a6e7;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4dcc6ccba893bde99cab28c5d73b8097b3ae;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5c9f367a2ef2c7c4b751d86ea956fc6c35a8;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7ee0eff19de3ed3d95526e905ce73c5fc9f6;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7b38ae3d75f939a93b85a03e11407259a256;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc0ab260cd62f32db5c9adf23602ed43abbe3;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2b4c045e44554e34ba2415652d550b5c78c9;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb874de4e278e11902a9ce72d337c674fa1df;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h77837e375698ce93bfcd7c59d5971ceca78f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8a977a028f10d3d9efd7c39498c63395ab60;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd122ba108df57efcf090c913939a4bac9b6c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2ac28732b59aced1ec6df0f5cee495dd14f7;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h54518f7e4700d534d283039d9e82f32afc27;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h956df5060209c8671c65af5d140ac5daf6fc;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd81a39061758fb02664bd415940d339c979;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf544de7212ec887e18565df0b0f55834808;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h171d1e0f6bf80eecf9334da2c1de4a554c48;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h94554c8a31b156774ca8d9d578dbd31abbdd;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5783a18e45950a639a235fa232e2beb5165e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h75a7f53a7bac36adda51abf23322d561f70a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb4d5f1787808e16e7790547af40b041d56a0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h197fdc6f15d7bf9a8ba980f2fb9ec6736291;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4ae3076a56c140016b09b15f84710499cbf8;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h22d511bc77eb9e590115fc30bb04146f669c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h819571489de784ffc27985b99586b4e06b3a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hfc6b0620eda09e4bcf6d12f46532c97a03c6;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h794e19812f10b0c184b959a8817e803dcf1d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h53645c4b6b1e4f5ee796ddfe0c6b60bf8b2b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'had989853a2bc1d05c43e7aead4e9f9e01b3c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h97a5ae917bda4cbd569810cc7ffe0afcd59f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2c9afac13d5bb31289c2da7bc3ec10cd84e3;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd301f37eadaaae7d8fcaa1426eb8dbf54a94;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h387fe65d219efa933edb7c262c99a38caf45;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h61edfd848909d0acab87976302ba26a5deeb;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5f9c13c4b30d4af2df21729339c87c21678d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hfdbd35618d79a8c7a73fc09e2528e9e9463d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hae1bbe21fb6332d1ffaa2331e3765f3669a3;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h89bcd05e81f8d307b132438b324c095cd76d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h90f2468f702f5850f7ca2fad9bc537219ae;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h81375e246c9b9cf00d39d424c4f353d86a19;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2007127ae75ea3c709b0f0dd08149b5520a9;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6929cae29ad2df0c284a2df071b226f4c6cd;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc8d5bfec53a093e99b6c63323adfb91ac70e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hef23c278c999e628d6acce4f201f5dc1dac;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h62cdabdf59e60c3e5757232ef759e79bec95;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbf20be9044e74eed4e4d228a8aea52d21288;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha67cb72f7238fa074049edbda52b73f8373f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h99436479e5a8b0e57ffebc4acb66919b5e5f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6a6fdac37afbdf9791f2715fcc0a45bdbefd;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h59d07e5e403c530896533fe33cccce33ff38;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3ac32dff536460348d2dec7e2ac1f96e3c05;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9d5d3890bf708c4db258ae83ae346f35427e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha28ee7b937468498562b27927cf9805c52b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h72518f39ea3435cd5b9dd52f7af8edf3e1f6;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hcc8f3aafd6380b3d197dc009b8c7c106b981;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h806ee611687901f0ddfb89b601b93a1216c0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h15452d64c9ea03950bea3e9cd6a0abeb81c9;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'heb49cb38e77df456f06bc9519207ee4a8e1d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h57a632e175e599127ee6d7df91f8dc1d0773;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc3b32c25f7bd78256d466c70027e20f81b3c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h13b7302028ad83ad1867a11f9cf4428f2f33;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb46381c29340fa95b869037316820c088cfc;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hcd46064b5d75b601c7e5ba9899de7f1d7dd2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hac2cfb5f4467e6f4f4f440c6032fa2fda10c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h106f85a489356ada6e417190ecd191c38a6a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5a9db82f4caaa6e75a0b3c7053299d6c5999;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h503fdadeb8c42fc2e48914a5e87954622046;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hdfd126af71543fa43bf2c5d15f2e7022b0ae;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hdd2794d071839c475ea90020190832808430;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5c1d2b3ba3a280c2a0a48efb64e9348346a6;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h422d9153da48cd9431ab9467e2989b8f2ee7;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1bb68215d932c42bc555761b3f8f8dfa84ce;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hcfb7e3e1c7eae0c089a588dcd927732144a5;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h215f5606cb3e0bc3abfbd20cd45e536381ef;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h59ecce6b551e615f542e92262c3ed99863d3;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8940407c3992aab66a311c4a1185a851ce4b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h19720bfe0b73c48cbfe17efba1569c024713;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hdb344ff805913f761919cb6ac0ac31830c76;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h679cd9b4e209a2797c63271145b9feca6806;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h95c5c1d6437107686c1c7df2266337ca0358;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb6f63ff0e9f81643aa2b9597565791dded54;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h95448324700003646970119c5f7083555872;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf64705b7540bda8ff15829a32314446f69ff;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h698140b2220fe1696aaf6081b698b621c5ae;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1ab727f8af2750595b6763ae2f525953f518;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc8996bd524daccb970dfb33c1afead8c4314;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'heca94b7c7d8c9ec3e522ef6513c0a4fd4558;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9b4aa17e428990ad795ef1c268be06bc8a61;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h15b84d06f8530175d84bac317ca431eaa3cc;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h444458869764c225c8ad1b3d9325ffcc521e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'haefc08c7ed9bb301c6c834b3b5f8c9320dd9;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h930c92f20c62718d411f56e178417c55120b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h98814ee1b5267d2057d5e17843d1a01bd62;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h407cc2179175abd6d00a394e7d7be0b84108;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3b9924bb968600c20d9ca39a224a47224699;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc23096c347ef13d993294ef7281a7d9af284;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc90d4c8ad184703097972982c2008f59be2d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9fe8935304357b0071bef7784d9a2361a5d2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7d4eaf00062e71e40739bbf6b22456d45e26;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h61824cb6227556fc120690b9f8b0214aeca1;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf92bd37e206a01cb48eb4ecd1c1c19c22538;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5019cf063a71a31597d0d9f2052f8cfd68d1;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8c9d916a2936d8beee51ccbb7821c9f5dc9b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h11c15d0874a216e437531d06fe09330041b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h53ae72f9ffe2651de7c6b008d3a59e937276;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h36947f69778cb4c7e862788604703404543;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6ef15d1e124d54ded811a8068b7338275de1;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbc52816b5f0bddcb2ada9f37d46613541578;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h54b1e8865732f43865c1d473c2220848ad53;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc03434d01f1181fe2ecb41db32f386700042;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1bba3e6c8ca493bb004cf81801c62f507cb3;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8ab945eb7ea4970c414022d2c3ddb33c7a6;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8eebc8e84d0e0a19fa5134cf13600aac0526;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbccff8c6e273e9a0b29e4d07fbb8a32218c2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3908f2cbda81951ff307bb3fa41831a0172;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h190a6ed704e0e1c9131c7ea5f79b213306ed;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h971329ad5c2aad99f9c7ad54ca30a493d335;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hda10a691ebcdfcde7e2ca742f20e8ad9c9aa;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h67026e16f51b8f7051831243537219b81972;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha61efd5b9d9a7a18e8eb439363ee724b202b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h626be3c69a5a6065e3da732e525c766f00db;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbc5e65e9c8816dfbe7c9cde9d08dc627a57f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd7d7e64cd10f865e42fbb3ceb51e013d99d5;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h72d8fb336a93e22b138472cc330f092e4667;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf29cde58831203fe11226978d1c1f62b7048;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4d266d3e0e8ffe2b1e2cfb65c0a2f31deb5f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb39f7fc1986f52a0ac41ddb20d64c4aaffa;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8fcd217627cd5314fab54dace26cab87aea9;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7a0ea5249d0b2a322b88219b492635a10304;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h98fe55760f05635ad3cacb1813f218592320;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb5fcfa38501e382b73020f56aefa5a1c5adb;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h266b1ea66c329f7877ea93b8337842ace47b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h242c9011563d7eb60c6507aa8b481e340cad;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'heabce96f82f44eb4d618cf36b4341c6099cc;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h411b6819d141b1f7fc5ded5cd094155f159e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd308da7e75b25e68f9ddfcc54f8663677a1b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf84a88fee515797a1ec9785e3aaa8f51f1e5;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he2809c0b3f51eeea0fac2869e077b06bfc4f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he221de315a392b482d7b9cb248f1eae4c6db;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h36fb1b003db4c29939b898e3ad0a6c27a790;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd4b2e76a983a530ac6d4d54450834b31492;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he038630a99efe5254ae691b585711d441856;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9c344127d86b8e9dc06ded0b4d4222bf5b7b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9c9827980e4f91244e0326a16936e4659e3a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf47ac725d9dd56210a2f5867487bfafd49b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbb03fb3da51770681a9fb8a0c152b32c3317;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h63537e3d13ffc8768080c9ce20c172eade4f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf90e7c2c62569731b4996529b8b6f299bde3;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he06f525078672885f64a95543e3c04b01328;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hab721dbb40c32f79d3bc78d773075251e7af;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd5ab357b24a2f2768f77c76f5e90d2b187fc;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2e4dbd89c86c4ecd0a0427702dbfe1077d56;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h25ef9159fbf247e0991c28ffe96136d9b367;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf7bc17cfeab965269e49e4a0cda18401ead;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he9c46698c2bbd6168a4ef270cadec3b7eeaf;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc5e5a31dde933425bd1e6ce35d5e9e306f62;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf94c5be01cdf22bcee5ec348ce850f48e4a3;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5c2c44f9cac0ab5ba359138f07663eb14002;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf773163462ccb77b7c5c445190c6674d2777;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h681b6b07e81fce0a532212c832c4b8ae205f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h64ab6913f67b5a07c6bf605ecbd695f98552;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hba6d0087d18b16d319dbc37dacde702b17a8;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h68b947528a6716413d70afc9fdd180e67213;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf694002dd9c44d3a9cd765f4de2e2cb84414;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h89433184c4b5416a0b52b7bcc54cf21a8a4e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h54196bfad36cb4488916889b6a1c9455b869;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hac4c88d7011cda2dfb433cfe296870125699;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4b9974991751cbdb93be65e67760b200736f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h50f22507eefe00e4585439c0da617cd9818c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb64fb5fff0301595e5830eb4d3df068020b2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha54a62a842f185dfc08468c05893edd95045;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hfa5d95d0b7b63d59a828f7912930357fda94;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h37e2b4f15f629a0969751e4fa59b41b1cef3;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8be9d07fee91170432ce59f618bb93274c77;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9e657ed5ad88e3ab174dce9cd81959749398;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3a473bb46ba1394e19816458caf93d8bce70;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h58f86d35728310ba41b1eaca7002c04641d8;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha1f882ef767f6a703d00c70c064eb7004487;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1de0854d5d48a042351482e5b03a35d8c504;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2c95d564a87ed1d27e817d5142e8822788;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h79ca0524bffa442502d02dd26ff2f0d2b9f1;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4f5ba4786f040b0da448ec019cdfafad09da;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h750f7fcfe2c6015b7dca677aaeec7c3519d1;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h397e8bf569eafa7ab792ee97e6b666138379;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4532d3a559ae02940859987738dc15e05450;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h40856adf2030dfb19e1fbe0c78a6a1786bfb;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he29a98d9954e418ded80843b59f0f2a74a0c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he993ecdca08d2b571b9a9d3995c4bee8c6a6;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9a386f6893a4dbbd6068878290d9879a5c62;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8bb5a10567717cee45cedee03fb11a8979c2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8725193b4ee5c90c3ba5425b8f60254cec7a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hfcf8d104f00d0b563f5ef6bcca490a8b7340;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf35b8b097b7bade69b8d5be667b0d9114f28;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb623987aed808b95cd4be140b3e2c67e3d5a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h279c36c803379cdd348ed113df03fc2c315c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2540b244355dbfa741df36a37b5eeb7fe0e4;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h616ec69de6c2a984c4559ea04ba9c17dce68;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf68668ff01dd0d5d5507ebf7ef995a010e1f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'haea3e3d03d45f9d5438756b3fd6631d3ea11;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he3a8a72daaa1553207fdc6afbc735f8200e6;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hba4dcbb84e9cbd285b28f1a0db60ea89cab3;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h292c0b79ef124ad928d5bf901ec066191e3d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h281abc243f7eb98c2f07059134c57539073e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h489a7191ae6e630660e68ef3a8e80e61d356;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hfe3c13dbc543fca1e45eda37aff64f778f81;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hcf96ef9f97a7995bb7b10256e072632a80bf;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf89944b0e67d3d3c51478573234619e93b92;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h764ac0b2998d96b46d7fb62aa04200912474;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1fd2f1e0092135ebd4de23db9aa4e8dd0688;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha09234dbdb17b342aec7154c9c92c5e9010d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3bb1ed76e37eb54be7a67dd8eb4435eefe62;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h58b718a49b7d6418a816ddc79fbf2518cb2d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h77292a11f85888beecc54b703106b514b6ae;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'heb787fc865bcfcdb649ef8485d94c07fc251;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1e7cc5e69a0c92be44aacd4bdf7943fc8512;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2f119ffcb9e4b9cf32dfaa4482d5554e7249;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4fe70384ba80c4f38700900df0e33ab5a4b9;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h17a1fbe359b0ca321e63348a6db4692a1a9b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h12e97246e070f3e0e01e8d75a13088da117a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h515786caf20f949bae571d71276a677ecd0a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hba2245130e0b1a68287a4b1a13f46a7d1b37;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h84dd66bcf86e07ca2330d892353dea8d152;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha3cb0c07108341e5d2cea16c465a0f1f7de9;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h31a395cb04ca7cfe737ad9b6f3dbdf5b84f3;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1d1d5004ad276a36af1f505799cd08398d88;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4daa8a9d803df00baa3b99fa52d42a94c390;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8544f4b326f023830ef3ee3ae76cb1eb47fd;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7ccd4a7d8440cdcb20810b96fe246f9e731a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5bb9c69e8b7de5fbdff9e51ecf1650fe51a5;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha91888bab06633158814bae40e4d08a83474;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h70ff5bc26f700bdbd7d31744478fbff1ad70;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc91f733bd1bc36e5885a40eb05607cab9b21;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h83a8a563c5affd7d20133295501024c7d43e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha5958f3d15541995e071c8d17ae7a033fd3c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf31043e45e566c3e4db1c11a31cfb76a2b1b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5103bf23d3f6f3db156bd484d79edbd5e3af;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h39174df4c6b32f16c31691232e260f36d710;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2a8acf6a053a112bb6e59d8f7743c94ba379;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h59d9ab442e21942bd06b5ecb41fbdcb0ceaa;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hefa04e9dfae7a74610c8c41594c7495d6e75;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h697fd53d9736a2a0368316802da7a522adab;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1d82f22f20963e282a3360520d47d5e65bee;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha5f5a1b497ba65d693afa2089d85c464d5b5;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1253020c005bee723b0e351d15a5a2cde3fc;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1b45cc0fdc2fd3fbc20296948ab8d7db50a5;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hff1bb115f327b008c1183028df278586ab7;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hea1ddcef4884fbc3882f86dfb646f76ff89a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5cf967feff250be7220d0244415ff3674466;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h950873127dc7b60b738666d541bc85515a5;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9a714706b750f36bb075781200c057c1d5f7;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hef852c3546e0d05b3dffb50efe51d5561a6a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he913aa58630c59b9f9861231237ef7e656cf;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h715c0a4d3290993fe3ce56e594a15d3d1a25;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h365365f8ba7dcd7a2404af0dd30c1bc9e449;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hedd07a250c842e8e144fd226594c16ed871c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h12626bebbd4a35c42ef1756f03424f2aa138;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he6cfb7097411208a1a7449fcdb1bb10ddf81;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h10412d6f1f2cfc82745f451666c67166e22b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf345081777b0288a45ab33ac8ab9ae4db2d7;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1fe2ce7c384303684cdff96c1ed78123c5b3;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hda51560d1d10e49456dcf5adee0058ca21d2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8ab2d2f9941905b77b3e5194889d987d004;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h80ca0adbb3e033d4cfe8d1764bd54d9ebaf5;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd5b0e2eefe4e146ee80016478cb5675f14fd;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h87aa1c47cbbbbf473570f743f8eb2e40b6cd;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hfd249953bb1a6096dfa14d284947ab2b8551;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3b920421ecf9f11a020cb45db7f0e8919cd6;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h994eb6ed699fbe28503f96c70feb7cb60c62;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6afbafd5bcd35168cdbc7e1f1cd6bf29d597;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc8808ac438bba4d5d79735f389dec48b0f0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hfc479720bb3844480e6dbb5d6e70934f0f4a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5b4180d15060c07f1ef1852553be9403d5bf;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3eb86c2de7d73c8456e28550901556df92aa;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf96190a9231a9a09157c918f822ed8068a91;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h18fe04c18f016c3d850972ba58e92cfc0631;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd9369be08bd5f9ce7577a802913f260d0706;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6b7ecb219c249d1659c3c309ca2a276b5739;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hab422521687cb782fd33d500b5df5cbec65;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd71916af1c983cbb4d4f3ca87829276eccfb;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1d7837274cbdc674fdaa913c557a35b7d653;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf68004aa81d2a7b76ddc355d2addf26fe195;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h183d3f431575dde838c11bf2b84b7bc2c7ae;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf25d2deb4c27ec11127427187eefdaf772f4;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he91baff7c09f59222c15bc9dd69b213d9e22;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5b6997f8ff5565d62c05a9feb0caf48eab2c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h86de4410930d11f13d179bb23d206238c7c2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf140a223ae7ccc8bf8cfe6150a0e4aa71fb6;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd633d426d6c3847ab0ab3493ea8846489b14;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hafcef39a091e9cb02def7582788c8f7a4dc3;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1a58fe0d5fa76deef2b1ed9bc47d592051a9;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb6c7593a8c9d4ce244af8a162a9c23650c49;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3b42f3789a59fb084056a6abd53f0e4a00ec;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb7ae58e90aeae7a70633980be7dd1e245ffc;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc3bf21c8ca2195b71c07aec3a52b40537120;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5d8e3efcbb99e5b98dc75e2c1bb934013cee;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he88ccca476a11888ec969710b8b2d5a6e630;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hddddbd435bb8c7b2ea645e17a6935b514aa;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd215a54c52714018647f66cbabad5c59aae1;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf32a94db5de8ba1b9bb2f6befbb7a08758e5;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2a50560e3720403bd46171e2f5001fa16aaa;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7f997d2c80d236fe0a99d0a54f6232ab0c2a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h482e207980767304bfc0ee02b898577f13c0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc452205e0c0fde2397c1d95659c7efb001e7;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1267ce08484c7120d9b707c982f3cadb42e6;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6470e2f1280cf536303edf1c7382b811b05d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he5cc93b2440bc70f67455e4a802d9acc0930;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3b20a9d555298e11e6ec2c6c712c58e5f37d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h44594ff35b59c0dce6bbb9704ff57fcc9ef7;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9e1cbc54fa498affb519940696bdb2af9b87;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h473acdb2608488c5b4c51903f280d64addcf;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'haa40fd4650b37da6e6afa89aa1fad2a8fc48;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5f2ca41ec46c8d1a5dd7af41a7a960c1d6eb;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc38603e995f6980acb6560208a1c482b6eac;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7b6ef4a4c0ccc36667fc0e4c0b86926ab67c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6859e5dfc164df5e949b3df41a35aabfd69;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hdaa88eb12d5c82df374f18ccd148993ddc6c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h383d5f6a467b94fe864b44fd0a96d927fc1f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8503763d8b376c7ba1584422a4869bb58598;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha1398cd45eaee6962ed1037b6f64998cb524;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hab431e68791204d0340665f43efd9ee6f054;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf927e76aa734467736b685a2ccb2564b9f29;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he8f55ba8923a7fc38534cd7c2a9bdd488318;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf1ee361ee0c9911bdb5412d30d077da2d019;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8729f1d019a24b7b260c16eb9c8a0b6cf217;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha2995dd5130e5ff9e2ccd860912e641f3881;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h319ff943e84c35a36de5273f556e32be7c70;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h692cb3e5a30aa7478975e49f7cf72d88a7fb;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf650d88ef866e1632f900e770b7cd5b00460;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hec250fc876a6830dedf81617ee81c5811069;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hedaa3c63542cd01720abdf377a75f57fe8b2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2c21205df0f7534134d078d73bd139eaaff2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h55e3aee0152a0b263b79859f3cd0a9f36ce7;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h69296fb0f7895e3b318cb9734fceba105997;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h179766c94dc9f1de549891374d85a6e5ad31;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'heb2db8f4de79f52e815470c324682f31db09;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h978d9728c89e539506683084a7ffb8617363;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd612715a12379a8042df8d641cd1e0034b0e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7265c24084846cd672d78d1c6b7914a7a7db;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'habe830cb886763269f32add363d0db0dac1b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4b67055219b37a099f60e0cb39f383c571cf;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hec86511e73f1d9ea718969649919f2112404;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h883674533004adec17ab4cbbc381ea390713;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6ba0e2c0360aa2fe292cd7b7396311e4e99f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h68d716a7b835cf0b1818a0f1cfc6e72c2d08;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6b4ec343d43512dd400ca7c8aabc902bcb2b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h667c75b9e787996332e914b46bf873fe3ca3;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8a25e2e8f41cfa9a4712a95ef53f0fa0c408;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1ed60f2df0090a174eb9d5a27f9a140b56d7;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd1b80410d8c7255cb8b5ce674074fe0ac4ea;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h47e2a285ff7200a6dc3e89830a8d4dfcd012;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2f90da5de4fece9cd95102f7522215fc92a0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h35662460dbd5091c88c823310a7530157ecf;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h435dd069050cf419a590ace52c8e8d2fc4cd;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h73322f0bc01680295a70a031a3c1ff187689;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h622811a212ffd05135c1a8aba55bd2d867f5;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd942d4ff95b850410c77c6ffe51b5b5f4f8a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h76aaba496ad0e04a1d7343af4ba9e612975b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h481d479a0d3a1e0401fca99aae16983ca9fa;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7358d773e52806978f15846a895f298e910c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbc7a3c4a3af100af6167085d915d10fe748d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5de3ee9c2e234c1a6060addedf7e5361d739;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc0dae1cb145033ebf00fdccbaa4b0c47a005;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h221e351517806f353e885d1cf6a99bceffb2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6cb570e61e740c4604b1fca79da2f6ff71a7;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd27c7de5acb173381bbe3a558ee6938dafc8;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h60afa6188a845b964795e6b0f6666686e78d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf3422564fc6943b3c5587eb266033b41a984;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9b84992eb04cd7e541971d633cf6181a9645;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha6278825d31b67c3938bf6abfccd86fe16e6;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc457e8521007ba31981a0a07e1001d9ed31d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h468f2be9faaeb29119a8ebb160cff0033e8d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hffd325e7d13ce86689c67c0a27b5301069bc;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf2cdbb52327b3bddc49e7a32bd26a51e71d6;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h625f266ee01bfd0e265e1df2aafa5461dea4;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9ca9efccb0006c7117ee247cd4f80816dd9b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1408bc43645ff50e32f11bd7e2de5e130ec6;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hdbb7d9ea8f74b131f69030fc0665ed9701b9;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9b358cc396bf22040fe7726d244447720524;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h95b601f718a7f2c601ffca32c9a3ac8d92e0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4846f2c562adb50abed62f564b2575381b73;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2a3b0a04f3c793d0736f84547571aa9819af;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9e15296f55485df7b5e78b33bbb617ba7c9a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1c866df7e3885122b2dc2f2fbd08c6b451a9;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h843a01f0db63ec812b30407e7746f704af4a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha5779bc30ff84296e4d0da86385dc217e657;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9bbcf6fe249cf016aeee115ac0076f535e80;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h789bb201732eebcd4b51718511b6b1a42055;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb2986a20d4f1f4e3c74a68afb649541cec54;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hba2ed51e3cd72eda252e851a00aed9c69c3c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h808ddd01614232f81cb7ce03dc40e1bf70e2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he3808c1a814a63958d339c4ffe9bfe352708;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7997fb2ba494e7730b9b608f0e8e570f47db;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha8bef61c93ef409d09d1c5dda383f06565ff;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h499c99ee895830c7b879ffc11090ddc1a9a8;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf673c326613b329cd24ce05fbf46d781b0a4;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2c770e52bd23da29c95fb245070b4107904;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h333bd97c990cd2d6a9ff5a50485d42f7a6fe;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h292755e96455b6e27a98fa03920a0d6d30e4;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4cf6c608cc5ab943f161ae201495e02ab351;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd73e29c8bfc16702b012c4e348a28c07bbb;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h33da76d7a4678ee9d4a222de955ade5a1241;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6880f4c6e9f23bf2784745f7c01143ad3538;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he0b2981dd7ad609b8cdf973488fc0ea1ebc0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha89447e10ebeaaabe09aa14fe2fe40c43443;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hdbb0ff9609a94bb710b79dbdf29223620971;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9787a3c215cd1ae2f5af512965aca5d59945;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha97565ea58865859d128cd0eb95b3ba908f4;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h75f9585b6b17a4fd7c1cb535f4bda0bfb165;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc40e53ed75027caca7a6a471d58ae3aaa22b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8386ea8475599430976fc03d56d20229c8a6;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hfccc69d31855b7111b39a291e9e292c5936;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb48e028865dea6e5542720b9fdc086b645a4;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2c6c52999813604b08465f5bac0673347e4a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he3159104d1168f83f59e3cf3ab65f05cac03;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1a44e62ead140f712b400b607f118d0006d0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h13ca19442728b51ea016de83d9ace6c4ae46;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h26e708d244c994ec6cd75eee143149eb15a2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1d116f6f32ae85a045daf49049642166982d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc24195114a228e1aefc3e2059cfbf9ecbc46;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h171cee5835cdafd8bcda6db94eca747a7386;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h92fe257bd76e2198e9d9506576b9e4b68bab;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h92b8c39b52f81fa93e2ca705a3d6fbb46ffc;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1603662c47e74bc0f0369e42e90a7b014991;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbbe7853fb9b2709a01765566e15f7c7dc381;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hff253fbb242a4f1c7e5aa1af1416c234aafa;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9ab8d09c63ae6b34e00742c38351ad627d1c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h78daa92a1aa94aafeb5e012ac69ea561a6ce;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h14cfa8c48854f103a111d1daa259cb05e4b2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h566e57e7d6d7fdcc7f920cc2fb6e562f0173;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb57e5a088fd9ffa272bedb74bc262e3dff01;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he9719692f1d1c0d80bc132167dcf0525e91;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha64b5b2244dbd3173129eddea76d77b528a9;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2332b56b822f9edec6cd6039a6bea1220636;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h14128a52150e435405122516962cea2609e3;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h91dbbe5fe4e299cd185ec7e0363c05a7d26e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4cb42fc25c0884c9c3e4363ab0d3bfb016ea;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h51edd9ea3d4581142200e6a274c71114c967;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he42a20d7ef5181b9e8d9c377cc7ea57a6455;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h235f63a2955a59ba3baa098c6645dff1abf1;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6c55f52231844f6e4074f96f5c952f46bcda;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8a3cdcc19fc58d33732e7c141899e0f87942;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h48c61b414c7dd649eda1074a5919398deeac;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hceaa4b640b132f257f6b83e7bf08820b8b23;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6f85430ee25fbefa74e8bb2a32def3c98735;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6842f8ac83a8c12c699f4298fdf590a05e60;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hffd0f3ff0a225301605507f33bf1f37b282b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6c22038ace35889f5f820af94567f7ca8405;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h588ae17b0bc073e7287212c310080038a2e3;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf173494c572699dddcccda04636a6b2bdf55;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h371675f090e7868688245b4528b2529ba9f7;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hfe538db2bd2a0a570bf5b9167910baabd056;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h22f3899d43e4d131f7832759e356554b568e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha7e6d6ae75718004ff0b5e39f90bc7c92b81;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h940780742ad41194fea538facb5cd57603ca;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h414bfa94fb1c59f18e83dcafef2f9d750d25;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6de0d9a95ed91b79760be03ab8fcc2d9f739;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb70b1ba66c98491c4804954cd280737aaf7;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7f83fe0ddccc912affc5f6d9a0b6023e1f51;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf6d46624dea0cfb073925c34748410c23644;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb3d905b5141b3b6e3be18575f4fe00f351c8;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5ddf9c646a4cddf32e535ec54d13c934bb41;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he49d34ab9bacbe9f45592d7400086d63aa23;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h60f9bd3c11d707069e23f7a056a00302db59;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc6338b7db6feca539e00213cd13ed5193c5e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h873c16d2a92082d3b1e81abdc30cbce0107;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5d40bb0fa104677412625fd046a55f1d0594;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he478a4f71fccd35ae0e9b3977ec9f4548700;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h908f1ee9fe55fbeef15a04144d0d1951f830;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hcd2913f89a1caad2feee61e9f5d819e18548;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb5fca769894ace339102cd7ec933a4e284d2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h89d450da54c78b53a0b80d5b639af8fcc30d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd423c85e76162094b35506f1e312b7568180;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h63958b7d850fada4b2dbe686ac7b18cc6117;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h54a3ce52a1a386c88f6ea3f0dd3be616eb19;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6edd8d85956b3d733d72c389dafaf87ab93a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hff88216f9dd4718b37817ede475f6c3a1eda;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2a5d1b8fb347c866c65f71c216f3020df70d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb16706152c08db5e6e86992728711b5362e5;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hed516ad2c4b266459bc8e720afec991f49c2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6df130a08a30e63cdfc2d7e439012f3c3d70;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'had79b5a635d8099910163848324510fe0f91;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9c012fb6b2107418e1efb849ec30acaa46a4;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4f40a8c3c5e633b0255c9aa882ff1d134550;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf8c161955d0d482e307d5c84de2b81fc46e6;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3a697a7c7b26dd0004fb57d36fcba0081130;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9f9f5174247f503a6241df012ec5b5d25436;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9653a01635721d75c40a8427eddd31095cdb;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8c2498f204ebf74d14834f32b2d10477ed64;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h10ad85bc7ed835b21aaf9a52e8da90d9b400;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf6a948a5913ed36dbeb1c79b65a2e090ef51;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h608f892a4036f58d4bee988314319c3ef36c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4c154bcd936814f80c95c3b9526545e5eb60;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h374bd5a00ae814805158acadd329ac17f2f2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h12a1c746aa850b7416dc1dea5be162f065c2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7c429fd18b2d8216484b6b8d6e835e40ccb;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8913f9c6c5e058fc821a6b298a2eb21930ae;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1d646b0d031ec107787524f3d1885a8159de;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf5ffa6f69121b296a44d71952e7113b1fab;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'haf35487e6e0bdc03120b5a31a426b2edfa00;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6eeafff1666eb9db227cb59558b4555b05ac;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9d7d50444aec378ed1c3795db1545886f77b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha4e28ec5cff1d7692be2a8ee121fe509a1e1;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h93f311ad04c712c39b5a0853936fec9b58fd;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3b84ae8a81837967d1581aad09ed7326e593;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h15bc7b72985eba60ecddc0cdf2acb9a1466c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h59be8b0fe1a030fccd7730faf0154f7cd054;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hdb0fff1dc7eaec0218560862e89781bba4e5;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h33cd77f382ec7250f0288e0ff25db4d8f329;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf30a39b1b38ce67080768582236ac7126b4c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb411481f6a4431a1f6ee16b4ccda4ed48840;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1aaf24f23d855bd0c24ee4166838d4e6736b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h53ced004897985f56ba6fed379a491df591b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha0154960ecf4b0d84fcbe1d56895b6005a66;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h16f372e5a4ffcb55e319a3ea964d4dfa50a2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he1644d67212a4e19e1cde743b621fd975609;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc592d0b9824b6f712ad147e27aa9b68b936e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h87a15da99630dd72d32009bc20b1ca04033d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h11444783f64addc3170fac1b5fccdf48f6e1;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9c80be61d10f4173dd7399b4e6e25cd894c4;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2adfe9f927306421e23e56bfb7ab409a3b67;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb299bae5ed1570f495b6060dff2175b2c56c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h818eb5084f370b0caf7904a4904688d7e5ba;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5334dee11f27d8a3639fab169ed5e4852446;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf431b31be659583ea3e3350432d8773eda71;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1f2891e17411ccac112a02d5160e9861e1f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9874c125c3ca598da25139e2fa14890daa10;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4a1905ee8286165a19c771d2a92c5740f6fc;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5ffd91d06aa23c9fba96b936908342c3ffbd;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h57dc522f96a472b838ff454bc5bb650623e8;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3636a05375c1c5270b6fb05ca807a9c09a42;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hde44dd08984bf02cecb65a48bf406bc78860;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1b72716787f3bdd6bbbad2c53f2215f9ff41;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb7021dfac01f0d3516ad9c7fdb5d42a91a98;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2321a3b8028abf9a0cd557fe337152d36aa9;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8cf29f635e4ccef02cf37a66b33fab461aad;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha6b6d5bf573f4beae205ba901010ee256631;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h16b58ed7be3a8d36fe99dc3341f6ede83125;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h220ed3d528e16db46af2d8a8157df08f8751;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd587111f055298d98132227703f049076905;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hebb9f784e2d8f11bea2e477fe31031bf6e0b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd85f3f00c2142276ccbb6d38c8e2f8ea7e66;
        #1
        $finish();
    end
endmodule
