module shift_register(
        input wire clk,
        input wire src0_,
        input wire src1_,
        input wire src2_,
        input wire src3_,
        input wire src4_,
        input wire src5_,
        input wire src6_,
        input wire src7_,
        input wire src8_,
        input wire src9_,
        input wire src10_,
        input wire src11_,
        output wire [0:0] dst0,
        output wire [0:0] dst1,
        output wire [0:0] dst2,
        output wire [0:0] dst3,
        output wire [0:0] dst4,
        output wire [0:0] dst5,
        output wire [0:0] dst6,
        output wire [0:0] dst7,
        output wire [0:0] dst8,
        output wire [0:0] dst9,
        output wire [0:0] dst10,
        output wire [0:0] dst11,
        output wire [0:0] dst12,
        output wire [0:0] dst13,
        output wire [0:0] dst14,
        output wire [0:0] dst15,
        output wire [0:0] dst16,
        output wire [0:0] dst17,
        output wire [0:0] dst18);
    reg [127:0] src0;
    reg [127:0] src1;
    reg [127:0] src2;
    reg [127:0] src3;
    reg [127:0] src4;
    reg [127:0] src5;
    reg [127:0] src6;
    reg [127:0] src7;
    reg [127:0] src8;
    reg [127:0] src9;
    reg [127:0] src10;
    reg [127:0] src11;
    compressor2_1_128_12 compressor2_1_128_12(
            .src0(src0),
            .src1(src1),
            .src2(src2),
            .src3(src3),
            .src4(src4),
            .src5(src5),
            .src6(src6),
            .src7(src7),
            .src8(src8),
            .src9(src9),
            .src10(src10),
            .src11(src11),
            .dst0(dst0),
            .dst1(dst1),
            .dst2(dst2),
            .dst3(dst3),
            .dst4(dst4),
            .dst5(dst5),
            .dst6(dst6),
            .dst7(dst7),
            .dst8(dst8),
            .dst9(dst9),
            .dst10(dst10),
            .dst11(dst11),
            .dst12(dst12),
            .dst13(dst13),
            .dst14(dst14),
            .dst15(dst15),
            .dst16(dst16),
            .dst17(dst17),
            .dst18(dst18));
    initial begin
        src0 <= 128'h0;
        src1 <= 128'h0;
        src2 <= 128'h0;
        src3 <= 128'h0;
        src4 <= 128'h0;
        src5 <= 128'h0;
        src6 <= 128'h0;
        src7 <= 128'h0;
        src8 <= 128'h0;
        src9 <= 128'h0;
        src10 <= 128'h0;
        src11 <= 128'h0;
    end
    always @(posedge clk) begin
        src0 <= {src0, src0_};
        src1 <= {src1, src1_};
        src2 <= {src2, src2_};
        src3 <= {src3, src3_};
        src4 <= {src4, src4_};
        src5 <= {src5, src5_};
        src6 <= {src6, src6_};
        src7 <= {src7, src7_};
        src8 <= {src8, src8_};
        src9 <= {src9, src9_};
        src10 <= {src10, src10_};
        src11 <= {src11, src11_};
    end
endmodule
module compressor2_1_128_12(
    input [127:0]src0,
    input [127:0]src1,
    input [127:0]src2,
    input [127:0]src3,
    input [127:0]src4,
    input [127:0]src5,
    input [127:0]src6,
    input [127:0]src7,
    input [127:0]src8,
    input [127:0]src9,
    input [127:0]src10,
    input [127:0]src11,
    output dst0,
    output dst1,
    output dst2,
    output dst3,
    output dst4,
    output dst5,
    output dst6,
    output dst7,
    output dst8,
    output dst9,
    output dst10,
    output dst11,
    output dst12,
    output dst13,
    output dst14,
    output dst15,
    output dst16,
    output dst17,
    output dst18);

    wire [1:0] comp_out0;
    wire [1:0] comp_out1;
    wire [1:0] comp_out2;
    wire [1:0] comp_out3;
    wire [1:0] comp_out4;
    wire [1:0] comp_out5;
    wire [1:0] comp_out6;
    wire [1:0] comp_out7;
    wire [1:0] comp_out8;
    wire [1:0] comp_out9;
    wire [1:0] comp_out10;
    wire [1:0] comp_out11;
    wire [1:0] comp_out12;
    wire [1:0] comp_out13;
    wire [1:0] comp_out14;
    wire [1:0] comp_out15;
    wire [1:0] comp_out16;
    wire [0:0] comp_out17;
    wire [1:0] comp_out18;
    compressor compressor_inst(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .dst0(comp_out0),
        .dst1(comp_out1),
        .dst2(comp_out2),
        .dst3(comp_out3),
        .dst4(comp_out4),
        .dst5(comp_out5),
        .dst6(comp_out6),
        .dst7(comp_out7),
        .dst8(comp_out8),
        .dst9(comp_out9),
        .dst10(comp_out10),
        .dst11(comp_out11),
        .dst12(comp_out12),
        .dst13(comp_out13),
        .dst14(comp_out14),
        .dst15(comp_out15),
        .dst16(comp_out16),
        .dst17(comp_out17),
        .dst18(comp_out18)
    );
    rowadder2_1_19 rowadder2_1inst(
        .src0({comp_out18[0], comp_out17[0], comp_out16[0], comp_out15[0], comp_out14[0], comp_out13[0], comp_out12[0], comp_out11[0], comp_out10[0], comp_out9[0], comp_out8[0], comp_out7[0], comp_out6[0], comp_out5[0], comp_out4[0], comp_out3[0], comp_out2[0], comp_out1[0], comp_out0[0]}),
        .src1({comp_out18[1], 1'h0, comp_out16[1], comp_out15[1], comp_out14[1], comp_out13[1], comp_out12[1], comp_out11[1], comp_out10[1], comp_out9[1], comp_out8[1], comp_out7[1], comp_out6[1], comp_out5[1], comp_out4[1], comp_out3[1], comp_out2[1], comp_out1[1], comp_out0[1]}),
        .dst0({dst18, dst17, dst16, dst15, dst14, dst13, dst12, dst11, dst10, dst9, dst8, dst7, dst6, dst5, dst4, dst3, dst2, dst1, dst0})
    );
endmodule
module compressor (
      input wire [127:0] src0,
      input wire [127:0] src1,
      input wire [127:0] src2,
      input wire [127:0] src3,
      input wire [127:0] src4,
      input wire [127:0] src5,
      input wire [127:0] src6,
      input wire [127:0] src7,
      input wire [127:0] src8,
      input wire [127:0] src9,
      input wire [127:0] src10,
      input wire [127:0] src11,
      output wire [1:0] dst0,
      output wire [1:0] dst1,
      output wire [1:0] dst2,
      output wire [1:0] dst3,
      output wire [1:0] dst4,
      output wire [1:0] dst5,
      output wire [1:0] dst6,
      output wire [1:0] dst7,
      output wire [1:0] dst8,
      output wire [1:0] dst9,
      output wire [1:0] dst10,
      output wire [1:0] dst11,
      output wire [1:0] dst12,
      output wire [1:0] dst13,
      output wire [1:0] dst14,
      output wire [1:0] dst15,
      output wire [1:0] dst16,
      output wire [0:0] dst17,
      output wire [1:0] dst18);

   wire [127:0] stage0_0;
   wire [127:0] stage0_1;
   wire [127:0] stage0_2;
   wire [127:0] stage0_3;
   wire [127:0] stage0_4;
   wire [127:0] stage0_5;
   wire [127:0] stage0_6;
   wire [127:0] stage0_7;
   wire [127:0] stage0_8;
   wire [127:0] stage0_9;
   wire [127:0] stage0_10;
   wire [127:0] stage0_11;
   wire [23:0] stage1_0;
   wire [40:0] stage1_1;
   wire [41:0] stage1_2;
   wire [57:0] stage1_3;
   wire [63:0] stage1_4;
   wire [61:0] stage1_5;
   wire [44:0] stage1_6;
   wire [43:0] stage1_7;
   wire [62:0] stage1_8;
   wire [63:0] stage1_9;
   wire [42:0] stage1_10;
   wire [43:0] stage1_11;
   wire [41:0] stage1_12;
   wire [20:0] stage1_13;
   wire [11:0] stage2_0;
   wire [8:0] stage2_1;
   wire [13:0] stage2_2;
   wire [20:0] stage2_3;
   wire [25:0] stage2_4;
   wire [22:0] stage2_5;
   wire [27:0] stage2_6;
   wire [21:0] stage2_7;
   wire [26:0] stage2_8;
   wire [24:0] stage2_9;
   wire [23:0] stage2_10;
   wire [19:0] stage2_11;
   wire [16:0] stage2_12;
   wire [15:0] stage2_13;
   wire [8:0] stage2_14;
   wire [3:0] stage2_15;
   wire [6:0] stage3_0;
   wire [4:0] stage3_1;
   wire [5:0] stage3_2;
   wire [5:0] stage3_3;
   wire [8:0] stage3_4;
   wire [11:0] stage3_5;
   wire [8:0] stage3_6;
   wire [11:0] stage3_7;
   wire [10:0] stage3_8;
   wire [7:0] stage3_9;
   wire [11:0] stage3_10;
   wire [10:0] stage3_11;
   wire [7:0] stage3_12;
   wire [5:0] stage3_13;
   wire [8:0] stage3_14;
   wire [7:0] stage3_15;
   wire [0:0] stage3_16;
   wire [6:0] stage4_0;
   wire [0:0] stage4_1;
   wire [6:0] stage4_2;
   wire [0:0] stage4_3;
   wire [4:0] stage4_4;
   wire [3:0] stage4_5;
   wire [5:0] stage4_6;
   wire [2:0] stage4_7;
   wire [5:0] stage4_8;
   wire [4:0] stage4_9;
   wire [2:0] stage4_10;
   wire [3:0] stage4_11;
   wire [5:0] stage4_12;
   wire [2:0] stage4_13;
   wire [2:0] stage4_14;
   wire [4:0] stage4_15;
   wire [1:0] stage4_16;
   wire [0:0] stage4_17;
   wire [0:0] stage4_18;
   wire [1:0] stage5_0;
   wire [1:0] stage5_1;
   wire [1:0] stage5_2;
   wire [1:0] stage5_3;
   wire [1:0] stage5_4;
   wire [1:0] stage5_5;
   wire [1:0] stage5_6;
   wire [1:0] stage5_7;
   wire [1:0] stage5_8;
   wire [1:0] stage5_9;
   wire [1:0] stage5_10;
   wire [1:0] stage5_11;
   wire [1:0] stage5_12;
   wire [1:0] stage5_13;
   wire [1:0] stage5_14;
   wire [1:0] stage5_15;
   wire [1:0] stage5_16;
   wire [0:0] stage5_17;
   wire [1:0] stage5_18;

   assign stage0_0 = src0;
   assign stage0_1 = src1;
   assign stage0_2 = src2;
   assign stage0_3 = src3;
   assign stage0_4 = src4;
   assign stage0_5 = src5;
   assign stage0_6 = src6;
   assign stage0_7 = src7;
   assign stage0_8 = src8;
   assign stage0_9 = src9;
   assign stage0_10 = src10;
   assign stage0_11 = src11;
   assign dst0 = stage5_0;
   assign dst1 = stage5_1;
   assign dst2 = stage5_2;
   assign dst3 = stage5_3;
   assign dst4 = stage5_4;
   assign dst5 = stage5_5;
   assign dst6 = stage5_6;
   assign dst7 = stage5_7;
   assign dst8 = stage5_8;
   assign dst9 = stage5_9;
   assign dst10 = stage5_10;
   assign dst11 = stage5_11;
   assign dst12 = stage5_12;
   assign dst13 = stage5_13;
   assign dst14 = stage5_14;
   assign dst15 = stage5_15;
   assign dst16 = stage5_16;
   assign dst17 = stage5_17;
   assign dst18 = stage5_18;

   gpc1163_5 gpc0 (
      {stage0_0[0], stage0_0[1], stage0_0[2]},
      {stage0_1[0], stage0_1[1], stage0_1[2], stage0_1[3], stage0_1[4], stage0_1[5]},
      {stage0_2[0]},
      {stage0_3[0]},
      {stage1_4[0],stage1_3[0],stage1_2[0],stage1_1[0],stage1_0[0]}
   );
   gpc1163_5 gpc1 (
      {stage0_0[3], stage0_0[4], stage0_0[5]},
      {stage0_1[6], stage0_1[7], stage0_1[8], stage0_1[9], stage0_1[10], stage0_1[11]},
      {stage0_2[1]},
      {stage0_3[1]},
      {stage1_4[1],stage1_3[1],stage1_2[1],stage1_1[1],stage1_0[1]}
   );
   gpc1163_5 gpc2 (
      {stage0_0[6], stage0_0[7], stage0_0[8]},
      {stage0_1[12], stage0_1[13], stage0_1[14], stage0_1[15], stage0_1[16], stage0_1[17]},
      {stage0_2[2]},
      {stage0_3[2]},
      {stage1_4[2],stage1_3[2],stage1_2[2],stage1_1[2],stage1_0[2]}
   );
   gpc606_5 gpc3 (
      {stage0_0[9], stage0_0[10], stage0_0[11], stage0_0[12], stage0_0[13], stage0_0[14]},
      {stage0_2[3], stage0_2[4], stage0_2[5], stage0_2[6], stage0_2[7], stage0_2[8]},
      {stage1_4[3],stage1_3[3],stage1_2[3],stage1_1[3],stage1_0[3]}
   );
   gpc606_5 gpc4 (
      {stage0_0[15], stage0_0[16], stage0_0[17], stage0_0[18], stage0_0[19], stage0_0[20]},
      {stage0_2[9], stage0_2[10], stage0_2[11], stage0_2[12], stage0_2[13], stage0_2[14]},
      {stage1_4[4],stage1_3[4],stage1_2[4],stage1_1[4],stage1_0[4]}
   );
   gpc606_5 gpc5 (
      {stage0_0[21], stage0_0[22], stage0_0[23], stage0_0[24], stage0_0[25], stage0_0[26]},
      {stage0_2[15], stage0_2[16], stage0_2[17], stage0_2[18], stage0_2[19], stage0_2[20]},
      {stage1_4[5],stage1_3[5],stage1_2[5],stage1_1[5],stage1_0[5]}
   );
   gpc606_5 gpc6 (
      {stage0_0[27], stage0_0[28], stage0_0[29], stage0_0[30], stage0_0[31], stage0_0[32]},
      {stage0_2[21], stage0_2[22], stage0_2[23], stage0_2[24], stage0_2[25], stage0_2[26]},
      {stage1_4[6],stage1_3[6],stage1_2[6],stage1_1[6],stage1_0[6]}
   );
   gpc606_5 gpc7 (
      {stage0_0[33], stage0_0[34], stage0_0[35], stage0_0[36], stage0_0[37], stage0_0[38]},
      {stage0_2[27], stage0_2[28], stage0_2[29], stage0_2[30], stage0_2[31], stage0_2[32]},
      {stage1_4[7],stage1_3[7],stage1_2[7],stage1_1[7],stage1_0[7]}
   );
   gpc606_5 gpc8 (
      {stage0_0[39], stage0_0[40], stage0_0[41], stage0_0[42], stage0_0[43], stage0_0[44]},
      {stage0_2[33], stage0_2[34], stage0_2[35], stage0_2[36], stage0_2[37], stage0_2[38]},
      {stage1_4[8],stage1_3[8],stage1_2[8],stage1_1[8],stage1_0[8]}
   );
   gpc606_5 gpc9 (
      {stage0_0[45], stage0_0[46], stage0_0[47], stage0_0[48], stage0_0[49], stage0_0[50]},
      {stage0_2[39], stage0_2[40], stage0_2[41], stage0_2[42], stage0_2[43], stage0_2[44]},
      {stage1_4[9],stage1_3[9],stage1_2[9],stage1_1[9],stage1_0[9]}
   );
   gpc606_5 gpc10 (
      {stage0_0[51], stage0_0[52], stage0_0[53], stage0_0[54], stage0_0[55], stage0_0[56]},
      {stage0_2[45], stage0_2[46], stage0_2[47], stage0_2[48], stage0_2[49], stage0_2[50]},
      {stage1_4[10],stage1_3[10],stage1_2[10],stage1_1[10],stage1_0[10]}
   );
   gpc606_5 gpc11 (
      {stage0_0[57], stage0_0[58], stage0_0[59], stage0_0[60], stage0_0[61], stage0_0[62]},
      {stage0_2[51], stage0_2[52], stage0_2[53], stage0_2[54], stage0_2[55], stage0_2[56]},
      {stage1_4[11],stage1_3[11],stage1_2[11],stage1_1[11],stage1_0[11]}
   );
   gpc606_5 gpc12 (
      {stage0_0[63], stage0_0[64], stage0_0[65], stage0_0[66], stage0_0[67], stage0_0[68]},
      {stage0_2[57], stage0_2[58], stage0_2[59], stage0_2[60], stage0_2[61], stage0_2[62]},
      {stage1_4[12],stage1_3[12],stage1_2[12],stage1_1[12],stage1_0[12]}
   );
   gpc606_5 gpc13 (
      {stage0_0[69], stage0_0[70], stage0_0[71], stage0_0[72], stage0_0[73], stage0_0[74]},
      {stage0_2[63], stage0_2[64], stage0_2[65], stage0_2[66], stage0_2[67], stage0_2[68]},
      {stage1_4[13],stage1_3[13],stage1_2[13],stage1_1[13],stage1_0[13]}
   );
   gpc606_5 gpc14 (
      {stage0_0[75], stage0_0[76], stage0_0[77], stage0_0[78], stage0_0[79], stage0_0[80]},
      {stage0_2[69], stage0_2[70], stage0_2[71], stage0_2[72], stage0_2[73], stage0_2[74]},
      {stage1_4[14],stage1_3[14],stage1_2[14],stage1_1[14],stage1_0[14]}
   );
   gpc606_5 gpc15 (
      {stage0_0[81], stage0_0[82], stage0_0[83], stage0_0[84], stage0_0[85], stage0_0[86]},
      {stage0_2[75], stage0_2[76], stage0_2[77], stage0_2[78], stage0_2[79], stage0_2[80]},
      {stage1_4[15],stage1_3[15],stage1_2[15],stage1_1[15],stage1_0[15]}
   );
   gpc606_5 gpc16 (
      {stage0_0[87], stage0_0[88], stage0_0[89], stage0_0[90], stage0_0[91], stage0_0[92]},
      {stage0_2[81], stage0_2[82], stage0_2[83], stage0_2[84], stage0_2[85], stage0_2[86]},
      {stage1_4[16],stage1_3[16],stage1_2[16],stage1_1[16],stage1_0[16]}
   );
   gpc606_5 gpc17 (
      {stage0_0[93], stage0_0[94], stage0_0[95], stage0_0[96], stage0_0[97], stage0_0[98]},
      {stage0_2[87], stage0_2[88], stage0_2[89], stage0_2[90], stage0_2[91], stage0_2[92]},
      {stage1_4[17],stage1_3[17],stage1_2[17],stage1_1[17],stage1_0[17]}
   );
   gpc606_5 gpc18 (
      {stage0_0[99], stage0_0[100], stage0_0[101], stage0_0[102], stage0_0[103], stage0_0[104]},
      {stage0_2[93], stage0_2[94], stage0_2[95], stage0_2[96], stage0_2[97], stage0_2[98]},
      {stage1_4[18],stage1_3[18],stage1_2[18],stage1_1[18],stage1_0[18]}
   );
   gpc606_5 gpc19 (
      {stage0_0[105], stage0_0[106], stage0_0[107], stage0_0[108], stage0_0[109], stage0_0[110]},
      {stage0_2[99], stage0_2[100], stage0_2[101], stage0_2[102], stage0_2[103], stage0_2[104]},
      {stage1_4[19],stage1_3[19],stage1_2[19],stage1_1[19],stage1_0[19]}
   );
   gpc606_5 gpc20 (
      {stage0_0[111], stage0_0[112], stage0_0[113], stage0_0[114], stage0_0[115], stage0_0[116]},
      {stage0_2[105], stage0_2[106], stage0_2[107], stage0_2[108], stage0_2[109], stage0_2[110]},
      {stage1_4[20],stage1_3[20],stage1_2[20],stage1_1[20],stage1_0[20]}
   );
   gpc615_5 gpc21 (
      {stage0_0[117], stage0_0[118], stage0_0[119], stage0_0[120], stage0_0[121]},
      {stage0_1[18]},
      {stage0_2[111], stage0_2[112], stage0_2[113], stage0_2[114], stage0_2[115], stage0_2[116]},
      {stage1_4[21],stage1_3[21],stage1_2[21],stage1_1[21],stage1_0[21]}
   );
   gpc615_5 gpc22 (
      {stage0_0[122], stage0_0[123], stage0_0[124], stage0_0[125], stage0_0[126]},
      {stage0_1[19]},
      {stage0_2[117], stage0_2[118], stage0_2[119], stage0_2[120], stage0_2[121], stage0_2[122]},
      {stage1_4[22],stage1_3[22],stage1_2[22],stage1_1[22],stage1_0[22]}
   );
   gpc606_5 gpc23 (
      {stage0_1[20], stage0_1[21], stage0_1[22], stage0_1[23], stage0_1[24], stage0_1[25]},
      {stage0_3[3], stage0_3[4], stage0_3[5], stage0_3[6], stage0_3[7], stage0_3[8]},
      {stage1_5[0],stage1_4[23],stage1_3[23],stage1_2[23],stage1_1[23]}
   );
   gpc606_5 gpc24 (
      {stage0_1[26], stage0_1[27], stage0_1[28], stage0_1[29], stage0_1[30], stage0_1[31]},
      {stage0_3[9], stage0_3[10], stage0_3[11], stage0_3[12], stage0_3[13], stage0_3[14]},
      {stage1_5[1],stage1_4[24],stage1_3[24],stage1_2[24],stage1_1[24]}
   );
   gpc606_5 gpc25 (
      {stage0_1[32], stage0_1[33], stage0_1[34], stage0_1[35], stage0_1[36], stage0_1[37]},
      {stage0_3[15], stage0_3[16], stage0_3[17], stage0_3[18], stage0_3[19], stage0_3[20]},
      {stage1_5[2],stage1_4[25],stage1_3[25],stage1_2[25],stage1_1[25]}
   );
   gpc606_5 gpc26 (
      {stage0_1[38], stage0_1[39], stage0_1[40], stage0_1[41], stage0_1[42], stage0_1[43]},
      {stage0_3[21], stage0_3[22], stage0_3[23], stage0_3[24], stage0_3[25], stage0_3[26]},
      {stage1_5[3],stage1_4[26],stage1_3[26],stage1_2[26],stage1_1[26]}
   );
   gpc606_5 gpc27 (
      {stage0_1[44], stage0_1[45], stage0_1[46], stage0_1[47], stage0_1[48], stage0_1[49]},
      {stage0_3[27], stage0_3[28], stage0_3[29], stage0_3[30], stage0_3[31], stage0_3[32]},
      {stage1_5[4],stage1_4[27],stage1_3[27],stage1_2[27],stage1_1[27]}
   );
   gpc606_5 gpc28 (
      {stage0_1[50], stage0_1[51], stage0_1[52], stage0_1[53], stage0_1[54], stage0_1[55]},
      {stage0_3[33], stage0_3[34], stage0_3[35], stage0_3[36], stage0_3[37], stage0_3[38]},
      {stage1_5[5],stage1_4[28],stage1_3[28],stage1_2[28],stage1_1[28]}
   );
   gpc606_5 gpc29 (
      {stage0_1[56], stage0_1[57], stage0_1[58], stage0_1[59], stage0_1[60], stage0_1[61]},
      {stage0_3[39], stage0_3[40], stage0_3[41], stage0_3[42], stage0_3[43], stage0_3[44]},
      {stage1_5[6],stage1_4[29],stage1_3[29],stage1_2[29],stage1_1[29]}
   );
   gpc606_5 gpc30 (
      {stage0_1[62], stage0_1[63], stage0_1[64], stage0_1[65], stage0_1[66], stage0_1[67]},
      {stage0_3[45], stage0_3[46], stage0_3[47], stage0_3[48], stage0_3[49], stage0_3[50]},
      {stage1_5[7],stage1_4[30],stage1_3[30],stage1_2[30],stage1_1[30]}
   );
   gpc606_5 gpc31 (
      {stage0_1[68], stage0_1[69], stage0_1[70], stage0_1[71], stage0_1[72], stage0_1[73]},
      {stage0_3[51], stage0_3[52], stage0_3[53], stage0_3[54], stage0_3[55], stage0_3[56]},
      {stage1_5[8],stage1_4[31],stage1_3[31],stage1_2[31],stage1_1[31]}
   );
   gpc606_5 gpc32 (
      {stage0_1[74], stage0_1[75], stage0_1[76], stage0_1[77], stage0_1[78], stage0_1[79]},
      {stage0_3[57], stage0_3[58], stage0_3[59], stage0_3[60], stage0_3[61], stage0_3[62]},
      {stage1_5[9],stage1_4[32],stage1_3[32],stage1_2[32],stage1_1[32]}
   );
   gpc606_5 gpc33 (
      {stage0_1[80], stage0_1[81], stage0_1[82], stage0_1[83], stage0_1[84], stage0_1[85]},
      {stage0_3[63], stage0_3[64], stage0_3[65], stage0_3[66], stage0_3[67], stage0_3[68]},
      {stage1_5[10],stage1_4[33],stage1_3[33],stage1_2[33],stage1_1[33]}
   );
   gpc606_5 gpc34 (
      {stage0_1[86], stage0_1[87], stage0_1[88], stage0_1[89], stage0_1[90], stage0_1[91]},
      {stage0_3[69], stage0_3[70], stage0_3[71], stage0_3[72], stage0_3[73], stage0_3[74]},
      {stage1_5[11],stage1_4[34],stage1_3[34],stage1_2[34],stage1_1[34]}
   );
   gpc606_5 gpc35 (
      {stage0_1[92], stage0_1[93], stage0_1[94], stage0_1[95], stage0_1[96], stage0_1[97]},
      {stage0_3[75], stage0_3[76], stage0_3[77], stage0_3[78], stage0_3[79], stage0_3[80]},
      {stage1_5[12],stage1_4[35],stage1_3[35],stage1_2[35],stage1_1[35]}
   );
   gpc606_5 gpc36 (
      {stage0_1[98], stage0_1[99], stage0_1[100], stage0_1[101], stage0_1[102], stage0_1[103]},
      {stage0_3[81], stage0_3[82], stage0_3[83], stage0_3[84], stage0_3[85], stage0_3[86]},
      {stage1_5[13],stage1_4[36],stage1_3[36],stage1_2[36],stage1_1[36]}
   );
   gpc606_5 gpc37 (
      {stage0_1[104], stage0_1[105], stage0_1[106], stage0_1[107], stage0_1[108], stage0_1[109]},
      {stage0_3[87], stage0_3[88], stage0_3[89], stage0_3[90], stage0_3[91], stage0_3[92]},
      {stage1_5[14],stage1_4[37],stage1_3[37],stage1_2[37],stage1_1[37]}
   );
   gpc606_5 gpc38 (
      {stage0_1[110], stage0_1[111], stage0_1[112], stage0_1[113], stage0_1[114], stage0_1[115]},
      {stage0_3[93], stage0_3[94], stage0_3[95], stage0_3[96], stage0_3[97], stage0_3[98]},
      {stage1_5[15],stage1_4[38],stage1_3[38],stage1_2[38],stage1_1[38]}
   );
   gpc606_5 gpc39 (
      {stage0_1[116], stage0_1[117], stage0_1[118], stage0_1[119], stage0_1[120], stage0_1[121]},
      {stage0_3[99], stage0_3[100], stage0_3[101], stage0_3[102], stage0_3[103], stage0_3[104]},
      {stage1_5[16],stage1_4[39],stage1_3[39],stage1_2[39],stage1_1[39]}
   );
   gpc606_5 gpc40 (
      {stage0_1[122], stage0_1[123], stage0_1[124], stage0_1[125], stage0_1[126], stage0_1[127]},
      {stage0_3[105], stage0_3[106], stage0_3[107], stage0_3[108], stage0_3[109], stage0_3[110]},
      {stage1_5[17],stage1_4[40],stage1_3[40],stage1_2[40],stage1_1[40]}
   );
   gpc615_5 gpc41 (
      {stage0_2[123], stage0_2[124], stage0_2[125], stage0_2[126], stage0_2[127]},
      {stage0_3[111]},
      {stage0_4[0], stage0_4[1], stage0_4[2], stage0_4[3], stage0_4[4], stage0_4[5]},
      {stage1_6[0],stage1_5[18],stage1_4[41],stage1_3[41],stage1_2[41]}
   );
   gpc606_5 gpc42 (
      {stage0_4[6], stage0_4[7], stage0_4[8], stage0_4[9], stage0_4[10], stage0_4[11]},
      {stage0_6[0], stage0_6[1], stage0_6[2], stage0_6[3], stage0_6[4], stage0_6[5]},
      {stage1_8[0],stage1_7[0],stage1_6[1],stage1_5[19],stage1_4[42]}
   );
   gpc606_5 gpc43 (
      {stage0_4[12], stage0_4[13], stage0_4[14], stage0_4[15], stage0_4[16], stage0_4[17]},
      {stage0_6[6], stage0_6[7], stage0_6[8], stage0_6[9], stage0_6[10], stage0_6[11]},
      {stage1_8[1],stage1_7[1],stage1_6[2],stage1_5[20],stage1_4[43]}
   );
   gpc606_5 gpc44 (
      {stage0_4[18], stage0_4[19], stage0_4[20], stage0_4[21], stage0_4[22], stage0_4[23]},
      {stage0_6[12], stage0_6[13], stage0_6[14], stage0_6[15], stage0_6[16], stage0_6[17]},
      {stage1_8[2],stage1_7[2],stage1_6[3],stage1_5[21],stage1_4[44]}
   );
   gpc606_5 gpc45 (
      {stage0_4[24], stage0_4[25], stage0_4[26], stage0_4[27], stage0_4[28], stage0_4[29]},
      {stage0_6[18], stage0_6[19], stage0_6[20], stage0_6[21], stage0_6[22], stage0_6[23]},
      {stage1_8[3],stage1_7[3],stage1_6[4],stage1_5[22],stage1_4[45]}
   );
   gpc606_5 gpc46 (
      {stage0_4[30], stage0_4[31], stage0_4[32], stage0_4[33], stage0_4[34], stage0_4[35]},
      {stage0_6[24], stage0_6[25], stage0_6[26], stage0_6[27], stage0_6[28], stage0_6[29]},
      {stage1_8[4],stage1_7[4],stage1_6[5],stage1_5[23],stage1_4[46]}
   );
   gpc606_5 gpc47 (
      {stage0_4[36], stage0_4[37], stage0_4[38], stage0_4[39], stage0_4[40], stage0_4[41]},
      {stage0_6[30], stage0_6[31], stage0_6[32], stage0_6[33], stage0_6[34], stage0_6[35]},
      {stage1_8[5],stage1_7[5],stage1_6[6],stage1_5[24],stage1_4[47]}
   );
   gpc606_5 gpc48 (
      {stage0_4[42], stage0_4[43], stage0_4[44], stage0_4[45], stage0_4[46], stage0_4[47]},
      {stage0_6[36], stage0_6[37], stage0_6[38], stage0_6[39], stage0_6[40], stage0_6[41]},
      {stage1_8[6],stage1_7[6],stage1_6[7],stage1_5[25],stage1_4[48]}
   );
   gpc606_5 gpc49 (
      {stage0_4[48], stage0_4[49], stage0_4[50], stage0_4[51], stage0_4[52], stage0_4[53]},
      {stage0_6[42], stage0_6[43], stage0_6[44], stage0_6[45], stage0_6[46], stage0_6[47]},
      {stage1_8[7],stage1_7[7],stage1_6[8],stage1_5[26],stage1_4[49]}
   );
   gpc606_5 gpc50 (
      {stage0_4[54], stage0_4[55], stage0_4[56], stage0_4[57], stage0_4[58], stage0_4[59]},
      {stage0_6[48], stage0_6[49], stage0_6[50], stage0_6[51], stage0_6[52], stage0_6[53]},
      {stage1_8[8],stage1_7[8],stage1_6[9],stage1_5[27],stage1_4[50]}
   );
   gpc606_5 gpc51 (
      {stage0_4[60], stage0_4[61], stage0_4[62], stage0_4[63], stage0_4[64], stage0_4[65]},
      {stage0_6[54], stage0_6[55], stage0_6[56], stage0_6[57], stage0_6[58], stage0_6[59]},
      {stage1_8[9],stage1_7[9],stage1_6[10],stage1_5[28],stage1_4[51]}
   );
   gpc606_5 gpc52 (
      {stage0_4[66], stage0_4[67], stage0_4[68], stage0_4[69], stage0_4[70], stage0_4[71]},
      {stage0_6[60], stage0_6[61], stage0_6[62], stage0_6[63], stage0_6[64], stage0_6[65]},
      {stage1_8[10],stage1_7[10],stage1_6[11],stage1_5[29],stage1_4[52]}
   );
   gpc606_5 gpc53 (
      {stage0_4[72], stage0_4[73], stage0_4[74], stage0_4[75], stage0_4[76], stage0_4[77]},
      {stage0_6[66], stage0_6[67], stage0_6[68], stage0_6[69], stage0_6[70], stage0_6[71]},
      {stage1_8[11],stage1_7[11],stage1_6[12],stage1_5[30],stage1_4[53]}
   );
   gpc606_5 gpc54 (
      {stage0_4[78], stage0_4[79], stage0_4[80], stage0_4[81], stage0_4[82], stage0_4[83]},
      {stage0_6[72], stage0_6[73], stage0_6[74], stage0_6[75], stage0_6[76], stage0_6[77]},
      {stage1_8[12],stage1_7[12],stage1_6[13],stage1_5[31],stage1_4[54]}
   );
   gpc606_5 gpc55 (
      {stage0_4[84], stage0_4[85], stage0_4[86], stage0_4[87], stage0_4[88], stage0_4[89]},
      {stage0_6[78], stage0_6[79], stage0_6[80], stage0_6[81], stage0_6[82], stage0_6[83]},
      {stage1_8[13],stage1_7[13],stage1_6[14],stage1_5[32],stage1_4[55]}
   );
   gpc606_5 gpc56 (
      {stage0_4[90], stage0_4[91], stage0_4[92], stage0_4[93], stage0_4[94], stage0_4[95]},
      {stage0_6[84], stage0_6[85], stage0_6[86], stage0_6[87], stage0_6[88], stage0_6[89]},
      {stage1_8[14],stage1_7[14],stage1_6[15],stage1_5[33],stage1_4[56]}
   );
   gpc606_5 gpc57 (
      {stage0_4[96], stage0_4[97], stage0_4[98], stage0_4[99], stage0_4[100], stage0_4[101]},
      {stage0_6[90], stage0_6[91], stage0_6[92], stage0_6[93], stage0_6[94], stage0_6[95]},
      {stage1_8[15],stage1_7[15],stage1_6[16],stage1_5[34],stage1_4[57]}
   );
   gpc606_5 gpc58 (
      {stage0_4[102], stage0_4[103], stage0_4[104], stage0_4[105], stage0_4[106], stage0_4[107]},
      {stage0_6[96], stage0_6[97], stage0_6[98], stage0_6[99], stage0_6[100], stage0_6[101]},
      {stage1_8[16],stage1_7[16],stage1_6[17],stage1_5[35],stage1_4[58]}
   );
   gpc606_5 gpc59 (
      {stage0_4[108], stage0_4[109], stage0_4[110], stage0_4[111], stage0_4[112], stage0_4[113]},
      {stage0_6[102], stage0_6[103], stage0_6[104], stage0_6[105], stage0_6[106], stage0_6[107]},
      {stage1_8[17],stage1_7[17],stage1_6[18],stage1_5[36],stage1_4[59]}
   );
   gpc606_5 gpc60 (
      {stage0_4[114], stage0_4[115], stage0_4[116], stage0_4[117], stage0_4[118], stage0_4[119]},
      {stage0_6[108], stage0_6[109], stage0_6[110], stage0_6[111], stage0_6[112], stage0_6[113]},
      {stage1_8[18],stage1_7[18],stage1_6[19],stage1_5[37],stage1_4[60]}
   );
   gpc606_5 gpc61 (
      {stage0_4[120], stage0_4[121], stage0_4[122], stage0_4[123], stage0_4[124], stage0_4[125]},
      {stage0_6[114], stage0_6[115], stage0_6[116], stage0_6[117], stage0_6[118], stage0_6[119]},
      {stage1_8[19],stage1_7[19],stage1_6[20],stage1_5[38],stage1_4[61]}
   );
   gpc606_5 gpc62 (
      {stage0_5[0], stage0_5[1], stage0_5[2], stage0_5[3], stage0_5[4], stage0_5[5]},
      {stage0_7[0], stage0_7[1], stage0_7[2], stage0_7[3], stage0_7[4], stage0_7[5]},
      {stage1_9[0],stage1_8[20],stage1_7[20],stage1_6[21],stage1_5[39]}
   );
   gpc606_5 gpc63 (
      {stage0_5[6], stage0_5[7], stage0_5[8], stage0_5[9], stage0_5[10], stage0_5[11]},
      {stage0_7[6], stage0_7[7], stage0_7[8], stage0_7[9], stage0_7[10], stage0_7[11]},
      {stage1_9[1],stage1_8[21],stage1_7[21],stage1_6[22],stage1_5[40]}
   );
   gpc606_5 gpc64 (
      {stage0_5[12], stage0_5[13], stage0_5[14], stage0_5[15], stage0_5[16], stage0_5[17]},
      {stage0_7[12], stage0_7[13], stage0_7[14], stage0_7[15], stage0_7[16], stage0_7[17]},
      {stage1_9[2],stage1_8[22],stage1_7[22],stage1_6[23],stage1_5[41]}
   );
   gpc606_5 gpc65 (
      {stage0_5[18], stage0_5[19], stage0_5[20], stage0_5[21], stage0_5[22], stage0_5[23]},
      {stage0_7[18], stage0_7[19], stage0_7[20], stage0_7[21], stage0_7[22], stage0_7[23]},
      {stage1_9[3],stage1_8[23],stage1_7[23],stage1_6[24],stage1_5[42]}
   );
   gpc606_5 gpc66 (
      {stage0_5[24], stage0_5[25], stage0_5[26], stage0_5[27], stage0_5[28], stage0_5[29]},
      {stage0_7[24], stage0_7[25], stage0_7[26], stage0_7[27], stage0_7[28], stage0_7[29]},
      {stage1_9[4],stage1_8[24],stage1_7[24],stage1_6[25],stage1_5[43]}
   );
   gpc606_5 gpc67 (
      {stage0_5[30], stage0_5[31], stage0_5[32], stage0_5[33], stage0_5[34], stage0_5[35]},
      {stage0_7[30], stage0_7[31], stage0_7[32], stage0_7[33], stage0_7[34], stage0_7[35]},
      {stage1_9[5],stage1_8[25],stage1_7[25],stage1_6[26],stage1_5[44]}
   );
   gpc606_5 gpc68 (
      {stage0_5[36], stage0_5[37], stage0_5[38], stage0_5[39], stage0_5[40], stage0_5[41]},
      {stage0_7[36], stage0_7[37], stage0_7[38], stage0_7[39], stage0_7[40], stage0_7[41]},
      {stage1_9[6],stage1_8[26],stage1_7[26],stage1_6[27],stage1_5[45]}
   );
   gpc606_5 gpc69 (
      {stage0_5[42], stage0_5[43], stage0_5[44], stage0_5[45], stage0_5[46], stage0_5[47]},
      {stage0_7[42], stage0_7[43], stage0_7[44], stage0_7[45], stage0_7[46], stage0_7[47]},
      {stage1_9[7],stage1_8[27],stage1_7[27],stage1_6[28],stage1_5[46]}
   );
   gpc606_5 gpc70 (
      {stage0_5[48], stage0_5[49], stage0_5[50], stage0_5[51], stage0_5[52], stage0_5[53]},
      {stage0_7[48], stage0_7[49], stage0_7[50], stage0_7[51], stage0_7[52], stage0_7[53]},
      {stage1_9[8],stage1_8[28],stage1_7[28],stage1_6[29],stage1_5[47]}
   );
   gpc606_5 gpc71 (
      {stage0_5[54], stage0_5[55], stage0_5[56], stage0_5[57], stage0_5[58], stage0_5[59]},
      {stage0_7[54], stage0_7[55], stage0_7[56], stage0_7[57], stage0_7[58], stage0_7[59]},
      {stage1_9[9],stage1_8[29],stage1_7[29],stage1_6[30],stage1_5[48]}
   );
   gpc606_5 gpc72 (
      {stage0_5[60], stage0_5[61], stage0_5[62], stage0_5[63], stage0_5[64], stage0_5[65]},
      {stage0_7[60], stage0_7[61], stage0_7[62], stage0_7[63], stage0_7[64], stage0_7[65]},
      {stage1_9[10],stage1_8[30],stage1_7[30],stage1_6[31],stage1_5[49]}
   );
   gpc606_5 gpc73 (
      {stage0_5[66], stage0_5[67], stage0_5[68], stage0_5[69], stage0_5[70], stage0_5[71]},
      {stage0_7[66], stage0_7[67], stage0_7[68], stage0_7[69], stage0_7[70], stage0_7[71]},
      {stage1_9[11],stage1_8[31],stage1_7[31],stage1_6[32],stage1_5[50]}
   );
   gpc606_5 gpc74 (
      {stage0_5[72], stage0_5[73], stage0_5[74], stage0_5[75], stage0_5[76], stage0_5[77]},
      {stage0_7[72], stage0_7[73], stage0_7[74], stage0_7[75], stage0_7[76], stage0_7[77]},
      {stage1_9[12],stage1_8[32],stage1_7[32],stage1_6[33],stage1_5[51]}
   );
   gpc606_5 gpc75 (
      {stage0_5[78], stage0_5[79], stage0_5[80], stage0_5[81], stage0_5[82], stage0_5[83]},
      {stage0_7[78], stage0_7[79], stage0_7[80], stage0_7[81], stage0_7[82], stage0_7[83]},
      {stage1_9[13],stage1_8[33],stage1_7[33],stage1_6[34],stage1_5[52]}
   );
   gpc606_5 gpc76 (
      {stage0_5[84], stage0_5[85], stage0_5[86], stage0_5[87], stage0_5[88], stage0_5[89]},
      {stage0_7[84], stage0_7[85], stage0_7[86], stage0_7[87], stage0_7[88], stage0_7[89]},
      {stage1_9[14],stage1_8[34],stage1_7[34],stage1_6[35],stage1_5[53]}
   );
   gpc606_5 gpc77 (
      {stage0_5[90], stage0_5[91], stage0_5[92], stage0_5[93], stage0_5[94], stage0_5[95]},
      {stage0_7[90], stage0_7[91], stage0_7[92], stage0_7[93], stage0_7[94], stage0_7[95]},
      {stage1_9[15],stage1_8[35],stage1_7[35],stage1_6[36],stage1_5[54]}
   );
   gpc606_5 gpc78 (
      {stage0_5[96], stage0_5[97], stage0_5[98], stage0_5[99], stage0_5[100], stage0_5[101]},
      {stage0_7[96], stage0_7[97], stage0_7[98], stage0_7[99], stage0_7[100], stage0_7[101]},
      {stage1_9[16],stage1_8[36],stage1_7[36],stage1_6[37],stage1_5[55]}
   );
   gpc606_5 gpc79 (
      {stage0_5[102], stage0_5[103], stage0_5[104], stage0_5[105], stage0_5[106], stage0_5[107]},
      {stage0_7[102], stage0_7[103], stage0_7[104], stage0_7[105], stage0_7[106], stage0_7[107]},
      {stage1_9[17],stage1_8[37],stage1_7[37],stage1_6[38],stage1_5[56]}
   );
   gpc606_5 gpc80 (
      {stage0_5[108], stage0_5[109], stage0_5[110], stage0_5[111], stage0_5[112], stage0_5[113]},
      {stage0_7[108], stage0_7[109], stage0_7[110], stage0_7[111], stage0_7[112], stage0_7[113]},
      {stage1_9[18],stage1_8[38],stage1_7[38],stage1_6[39],stage1_5[57]}
   );
   gpc606_5 gpc81 (
      {stage0_5[114], stage0_5[115], stage0_5[116], stage0_5[117], stage0_5[118], stage0_5[119]},
      {stage0_7[114], stage0_7[115], stage0_7[116], stage0_7[117], stage0_7[118], stage0_7[119]},
      {stage1_9[19],stage1_8[39],stage1_7[39],stage1_6[40],stage1_5[58]}
   );
   gpc606_5 gpc82 (
      {stage0_5[120], stage0_5[121], stage0_5[122], stage0_5[123], stage0_5[124], stage0_5[125]},
      {stage0_7[120], stage0_7[121], stage0_7[122], stage0_7[123], stage0_7[124], stage0_7[125]},
      {stage1_9[20],stage1_8[40],stage1_7[40],stage1_6[41],stage1_5[59]}
   );
   gpc606_5 gpc83 (
      {stage0_6[120], stage0_6[121], stage0_6[122], stage0_6[123], stage0_6[124], stage0_6[125]},
      {stage0_8[0], stage0_8[1], stage0_8[2], stage0_8[3], stage0_8[4], stage0_8[5]},
      {stage1_10[0],stage1_9[21],stage1_8[41],stage1_7[41],stage1_6[42]}
   );
   gpc606_5 gpc84 (
      {stage0_8[6], stage0_8[7], stage0_8[8], stage0_8[9], stage0_8[10], stage0_8[11]},
      {stage0_10[0], stage0_10[1], stage0_10[2], stage0_10[3], stage0_10[4], stage0_10[5]},
      {stage1_12[0],stage1_11[0],stage1_10[1],stage1_9[22],stage1_8[42]}
   );
   gpc606_5 gpc85 (
      {stage0_8[12], stage0_8[13], stage0_8[14], stage0_8[15], stage0_8[16], stage0_8[17]},
      {stage0_10[6], stage0_10[7], stage0_10[8], stage0_10[9], stage0_10[10], stage0_10[11]},
      {stage1_12[1],stage1_11[1],stage1_10[2],stage1_9[23],stage1_8[43]}
   );
   gpc606_5 gpc86 (
      {stage0_8[18], stage0_8[19], stage0_8[20], stage0_8[21], stage0_8[22], stage0_8[23]},
      {stage0_10[12], stage0_10[13], stage0_10[14], stage0_10[15], stage0_10[16], stage0_10[17]},
      {stage1_12[2],stage1_11[2],stage1_10[3],stage1_9[24],stage1_8[44]}
   );
   gpc606_5 gpc87 (
      {stage0_8[24], stage0_8[25], stage0_8[26], stage0_8[27], stage0_8[28], stage0_8[29]},
      {stage0_10[18], stage0_10[19], stage0_10[20], stage0_10[21], stage0_10[22], stage0_10[23]},
      {stage1_12[3],stage1_11[3],stage1_10[4],stage1_9[25],stage1_8[45]}
   );
   gpc606_5 gpc88 (
      {stage0_8[30], stage0_8[31], stage0_8[32], stage0_8[33], stage0_8[34], stage0_8[35]},
      {stage0_10[24], stage0_10[25], stage0_10[26], stage0_10[27], stage0_10[28], stage0_10[29]},
      {stage1_12[4],stage1_11[4],stage1_10[5],stage1_9[26],stage1_8[46]}
   );
   gpc606_5 gpc89 (
      {stage0_8[36], stage0_8[37], stage0_8[38], stage0_8[39], stage0_8[40], stage0_8[41]},
      {stage0_10[30], stage0_10[31], stage0_10[32], stage0_10[33], stage0_10[34], stage0_10[35]},
      {stage1_12[5],stage1_11[5],stage1_10[6],stage1_9[27],stage1_8[47]}
   );
   gpc606_5 gpc90 (
      {stage0_8[42], stage0_8[43], stage0_8[44], stage0_8[45], stage0_8[46], stage0_8[47]},
      {stage0_10[36], stage0_10[37], stage0_10[38], stage0_10[39], stage0_10[40], stage0_10[41]},
      {stage1_12[6],stage1_11[6],stage1_10[7],stage1_9[28],stage1_8[48]}
   );
   gpc606_5 gpc91 (
      {stage0_8[48], stage0_8[49], stage0_8[50], stage0_8[51], stage0_8[52], stage0_8[53]},
      {stage0_10[42], stage0_10[43], stage0_10[44], stage0_10[45], stage0_10[46], stage0_10[47]},
      {stage1_12[7],stage1_11[7],stage1_10[8],stage1_9[29],stage1_8[49]}
   );
   gpc606_5 gpc92 (
      {stage0_8[54], stage0_8[55], stage0_8[56], stage0_8[57], stage0_8[58], stage0_8[59]},
      {stage0_10[48], stage0_10[49], stage0_10[50], stage0_10[51], stage0_10[52], stage0_10[53]},
      {stage1_12[8],stage1_11[8],stage1_10[9],stage1_9[30],stage1_8[50]}
   );
   gpc606_5 gpc93 (
      {stage0_8[60], stage0_8[61], stage0_8[62], stage0_8[63], stage0_8[64], stage0_8[65]},
      {stage0_10[54], stage0_10[55], stage0_10[56], stage0_10[57], stage0_10[58], stage0_10[59]},
      {stage1_12[9],stage1_11[9],stage1_10[10],stage1_9[31],stage1_8[51]}
   );
   gpc606_5 gpc94 (
      {stage0_8[66], stage0_8[67], stage0_8[68], stage0_8[69], stage0_8[70], stage0_8[71]},
      {stage0_10[60], stage0_10[61], stage0_10[62], stage0_10[63], stage0_10[64], stage0_10[65]},
      {stage1_12[10],stage1_11[10],stage1_10[11],stage1_9[32],stage1_8[52]}
   );
   gpc606_5 gpc95 (
      {stage0_8[72], stage0_8[73], stage0_8[74], stage0_8[75], stage0_8[76], stage0_8[77]},
      {stage0_10[66], stage0_10[67], stage0_10[68], stage0_10[69], stage0_10[70], stage0_10[71]},
      {stage1_12[11],stage1_11[11],stage1_10[12],stage1_9[33],stage1_8[53]}
   );
   gpc606_5 gpc96 (
      {stage0_8[78], stage0_8[79], stage0_8[80], stage0_8[81], stage0_8[82], stage0_8[83]},
      {stage0_10[72], stage0_10[73], stage0_10[74], stage0_10[75], stage0_10[76], stage0_10[77]},
      {stage1_12[12],stage1_11[12],stage1_10[13],stage1_9[34],stage1_8[54]}
   );
   gpc606_5 gpc97 (
      {stage0_8[84], stage0_8[85], stage0_8[86], stage0_8[87], stage0_8[88], stage0_8[89]},
      {stage0_10[78], stage0_10[79], stage0_10[80], stage0_10[81], stage0_10[82], stage0_10[83]},
      {stage1_12[13],stage1_11[13],stage1_10[14],stage1_9[35],stage1_8[55]}
   );
   gpc606_5 gpc98 (
      {stage0_8[90], stage0_8[91], stage0_8[92], stage0_8[93], stage0_8[94], stage0_8[95]},
      {stage0_10[84], stage0_10[85], stage0_10[86], stage0_10[87], stage0_10[88], stage0_10[89]},
      {stage1_12[14],stage1_11[14],stage1_10[15],stage1_9[36],stage1_8[56]}
   );
   gpc606_5 gpc99 (
      {stage0_8[96], stage0_8[97], stage0_8[98], stage0_8[99], stage0_8[100], stage0_8[101]},
      {stage0_10[90], stage0_10[91], stage0_10[92], stage0_10[93], stage0_10[94], stage0_10[95]},
      {stage1_12[15],stage1_11[15],stage1_10[16],stage1_9[37],stage1_8[57]}
   );
   gpc606_5 gpc100 (
      {stage0_8[102], stage0_8[103], stage0_8[104], stage0_8[105], stage0_8[106], stage0_8[107]},
      {stage0_10[96], stage0_10[97], stage0_10[98], stage0_10[99], stage0_10[100], stage0_10[101]},
      {stage1_12[16],stage1_11[16],stage1_10[17],stage1_9[38],stage1_8[58]}
   );
   gpc615_5 gpc101 (
      {stage0_8[108], stage0_8[109], stage0_8[110], stage0_8[111], stage0_8[112]},
      {stage0_9[0]},
      {stage0_10[102], stage0_10[103], stage0_10[104], stage0_10[105], stage0_10[106], stage0_10[107]},
      {stage1_12[17],stage1_11[17],stage1_10[18],stage1_9[39],stage1_8[59]}
   );
   gpc615_5 gpc102 (
      {stage0_8[113], stage0_8[114], stage0_8[115], stage0_8[116], stage0_8[117]},
      {stage0_9[1]},
      {stage0_10[108], stage0_10[109], stage0_10[110], stage0_10[111], stage0_10[112], stage0_10[113]},
      {stage1_12[18],stage1_11[18],stage1_10[19],stage1_9[40],stage1_8[60]}
   );
   gpc615_5 gpc103 (
      {stage0_8[118], stage0_8[119], stage0_8[120], stage0_8[121], stage0_8[122]},
      {stage0_9[2]},
      {stage0_10[114], stage0_10[115], stage0_10[116], stage0_10[117], stage0_10[118], stage0_10[119]},
      {stage1_12[19],stage1_11[19],stage1_10[20],stage1_9[41],stage1_8[61]}
   );
   gpc615_5 gpc104 (
      {stage0_8[123], stage0_8[124], stage0_8[125], stage0_8[126], stage0_8[127]},
      {stage0_9[3]},
      {stage0_10[120], stage0_10[121], stage0_10[122], stage0_10[123], stage0_10[124], stage0_10[125]},
      {stage1_12[20],stage1_11[20],stage1_10[21],stage1_9[42],stage1_8[62]}
   );
   gpc606_5 gpc105 (
      {stage0_9[4], stage0_9[5], stage0_9[6], stage0_9[7], stage0_9[8], stage0_9[9]},
      {stage0_11[0], stage0_11[1], stage0_11[2], stage0_11[3], stage0_11[4], stage0_11[5]},
      {stage1_13[0],stage1_12[21],stage1_11[21],stage1_10[22],stage1_9[43]}
   );
   gpc606_5 gpc106 (
      {stage0_9[10], stage0_9[11], stage0_9[12], stage0_9[13], stage0_9[14], stage0_9[15]},
      {stage0_11[6], stage0_11[7], stage0_11[8], stage0_11[9], stage0_11[10], stage0_11[11]},
      {stage1_13[1],stage1_12[22],stage1_11[22],stage1_10[23],stage1_9[44]}
   );
   gpc606_5 gpc107 (
      {stage0_9[16], stage0_9[17], stage0_9[18], stage0_9[19], stage0_9[20], stage0_9[21]},
      {stage0_11[12], stage0_11[13], stage0_11[14], stage0_11[15], stage0_11[16], stage0_11[17]},
      {stage1_13[2],stage1_12[23],stage1_11[23],stage1_10[24],stage1_9[45]}
   );
   gpc606_5 gpc108 (
      {stage0_9[22], stage0_9[23], stage0_9[24], stage0_9[25], stage0_9[26], stage0_9[27]},
      {stage0_11[18], stage0_11[19], stage0_11[20], stage0_11[21], stage0_11[22], stage0_11[23]},
      {stage1_13[3],stage1_12[24],stage1_11[24],stage1_10[25],stage1_9[46]}
   );
   gpc606_5 gpc109 (
      {stage0_9[28], stage0_9[29], stage0_9[30], stage0_9[31], stage0_9[32], stage0_9[33]},
      {stage0_11[24], stage0_11[25], stage0_11[26], stage0_11[27], stage0_11[28], stage0_11[29]},
      {stage1_13[4],stage1_12[25],stage1_11[25],stage1_10[26],stage1_9[47]}
   );
   gpc606_5 gpc110 (
      {stage0_9[34], stage0_9[35], stage0_9[36], stage0_9[37], stage0_9[38], stage0_9[39]},
      {stage0_11[30], stage0_11[31], stage0_11[32], stage0_11[33], stage0_11[34], stage0_11[35]},
      {stage1_13[5],stage1_12[26],stage1_11[26],stage1_10[27],stage1_9[48]}
   );
   gpc606_5 gpc111 (
      {stage0_9[40], stage0_9[41], stage0_9[42], stage0_9[43], stage0_9[44], stage0_9[45]},
      {stage0_11[36], stage0_11[37], stage0_11[38], stage0_11[39], stage0_11[40], stage0_11[41]},
      {stage1_13[6],stage1_12[27],stage1_11[27],stage1_10[28],stage1_9[49]}
   );
   gpc606_5 gpc112 (
      {stage0_9[46], stage0_9[47], stage0_9[48], stage0_9[49], stage0_9[50], stage0_9[51]},
      {stage0_11[42], stage0_11[43], stage0_11[44], stage0_11[45], stage0_11[46], stage0_11[47]},
      {stage1_13[7],stage1_12[28],stage1_11[28],stage1_10[29],stage1_9[50]}
   );
   gpc606_5 gpc113 (
      {stage0_9[52], stage0_9[53], stage0_9[54], stage0_9[55], stage0_9[56], stage0_9[57]},
      {stage0_11[48], stage0_11[49], stage0_11[50], stage0_11[51], stage0_11[52], stage0_11[53]},
      {stage1_13[8],stage1_12[29],stage1_11[29],stage1_10[30],stage1_9[51]}
   );
   gpc606_5 gpc114 (
      {stage0_9[58], stage0_9[59], stage0_9[60], stage0_9[61], stage0_9[62], stage0_9[63]},
      {stage0_11[54], stage0_11[55], stage0_11[56], stage0_11[57], stage0_11[58], stage0_11[59]},
      {stage1_13[9],stage1_12[30],stage1_11[30],stage1_10[31],stage1_9[52]}
   );
   gpc606_5 gpc115 (
      {stage0_9[64], stage0_9[65], stage0_9[66], stage0_9[67], stage0_9[68], stage0_9[69]},
      {stage0_11[60], stage0_11[61], stage0_11[62], stage0_11[63], stage0_11[64], stage0_11[65]},
      {stage1_13[10],stage1_12[31],stage1_11[31],stage1_10[32],stage1_9[53]}
   );
   gpc606_5 gpc116 (
      {stage0_9[70], stage0_9[71], stage0_9[72], stage0_9[73], stage0_9[74], stage0_9[75]},
      {stage0_11[66], stage0_11[67], stage0_11[68], stage0_11[69], stage0_11[70], stage0_11[71]},
      {stage1_13[11],stage1_12[32],stage1_11[32],stage1_10[33],stage1_9[54]}
   );
   gpc606_5 gpc117 (
      {stage0_9[76], stage0_9[77], stage0_9[78], stage0_9[79], stage0_9[80], stage0_9[81]},
      {stage0_11[72], stage0_11[73], stage0_11[74], stage0_11[75], stage0_11[76], stage0_11[77]},
      {stage1_13[12],stage1_12[33],stage1_11[33],stage1_10[34],stage1_9[55]}
   );
   gpc606_5 gpc118 (
      {stage0_9[82], stage0_9[83], stage0_9[84], stage0_9[85], stage0_9[86], stage0_9[87]},
      {stage0_11[78], stage0_11[79], stage0_11[80], stage0_11[81], stage0_11[82], stage0_11[83]},
      {stage1_13[13],stage1_12[34],stage1_11[34],stage1_10[35],stage1_9[56]}
   );
   gpc606_5 gpc119 (
      {stage0_9[88], stage0_9[89], stage0_9[90], stage0_9[91], stage0_9[92], stage0_9[93]},
      {stage0_11[84], stage0_11[85], stage0_11[86], stage0_11[87], stage0_11[88], stage0_11[89]},
      {stage1_13[14],stage1_12[35],stage1_11[35],stage1_10[36],stage1_9[57]}
   );
   gpc606_5 gpc120 (
      {stage0_9[94], stage0_9[95], stage0_9[96], stage0_9[97], stage0_9[98], stage0_9[99]},
      {stage0_11[90], stage0_11[91], stage0_11[92], stage0_11[93], stage0_11[94], stage0_11[95]},
      {stage1_13[15],stage1_12[36],stage1_11[36],stage1_10[37],stage1_9[58]}
   );
   gpc606_5 gpc121 (
      {stage0_9[100], stage0_9[101], stage0_9[102], stage0_9[103], stage0_9[104], stage0_9[105]},
      {stage0_11[96], stage0_11[97], stage0_11[98], stage0_11[99], stage0_11[100], stage0_11[101]},
      {stage1_13[16],stage1_12[37],stage1_11[37],stage1_10[38],stage1_9[59]}
   );
   gpc606_5 gpc122 (
      {stage0_9[106], stage0_9[107], stage0_9[108], stage0_9[109], stage0_9[110], stage0_9[111]},
      {stage0_11[102], stage0_11[103], stage0_11[104], stage0_11[105], stage0_11[106], stage0_11[107]},
      {stage1_13[17],stage1_12[38],stage1_11[38],stage1_10[39],stage1_9[60]}
   );
   gpc606_5 gpc123 (
      {stage0_9[112], stage0_9[113], stage0_9[114], stage0_9[115], stage0_9[116], stage0_9[117]},
      {stage0_11[108], stage0_11[109], stage0_11[110], stage0_11[111], stage0_11[112], stage0_11[113]},
      {stage1_13[18],stage1_12[39],stage1_11[39],stage1_10[40],stage1_9[61]}
   );
   gpc615_5 gpc124 (
      {stage0_9[118], stage0_9[119], stage0_9[120], stage0_9[121], stage0_9[122]},
      {stage0_10[126]},
      {stage0_11[114], stage0_11[115], stage0_11[116], stage0_11[117], stage0_11[118], stage0_11[119]},
      {stage1_13[19],stage1_12[40],stage1_11[40],stage1_10[41],stage1_9[62]}
   );
   gpc615_5 gpc125 (
      {stage0_9[123], stage0_9[124], stage0_9[125], stage0_9[126], stage0_9[127]},
      {stage0_10[127]},
      {stage0_11[120], stage0_11[121], stage0_11[122], stage0_11[123], stage0_11[124], stage0_11[125]},
      {stage1_13[20],stage1_12[41],stage1_11[41],stage1_10[42],stage1_9[63]}
   );
   gpc1_1 gpc126 (
      {stage0_0[127]},
      {stage1_0[23]}
   );
   gpc1_1 gpc127 (
      {stage0_3[112]},
      {stage1_3[42]}
   );
   gpc1_1 gpc128 (
      {stage0_3[113]},
      {stage1_3[43]}
   );
   gpc1_1 gpc129 (
      {stage0_3[114]},
      {stage1_3[44]}
   );
   gpc1_1 gpc130 (
      {stage0_3[115]},
      {stage1_3[45]}
   );
   gpc1_1 gpc131 (
      {stage0_3[116]},
      {stage1_3[46]}
   );
   gpc1_1 gpc132 (
      {stage0_3[117]},
      {stage1_3[47]}
   );
   gpc1_1 gpc133 (
      {stage0_3[118]},
      {stage1_3[48]}
   );
   gpc1_1 gpc134 (
      {stage0_3[119]},
      {stage1_3[49]}
   );
   gpc1_1 gpc135 (
      {stage0_3[120]},
      {stage1_3[50]}
   );
   gpc1_1 gpc136 (
      {stage0_3[121]},
      {stage1_3[51]}
   );
   gpc1_1 gpc137 (
      {stage0_3[122]},
      {stage1_3[52]}
   );
   gpc1_1 gpc138 (
      {stage0_3[123]},
      {stage1_3[53]}
   );
   gpc1_1 gpc139 (
      {stage0_3[124]},
      {stage1_3[54]}
   );
   gpc1_1 gpc140 (
      {stage0_3[125]},
      {stage1_3[55]}
   );
   gpc1_1 gpc141 (
      {stage0_3[126]},
      {stage1_3[56]}
   );
   gpc1_1 gpc142 (
      {stage0_3[127]},
      {stage1_3[57]}
   );
   gpc1_1 gpc143 (
      {stage0_4[126]},
      {stage1_4[62]}
   );
   gpc1_1 gpc144 (
      {stage0_4[127]},
      {stage1_4[63]}
   );
   gpc1_1 gpc145 (
      {stage0_5[126]},
      {stage1_5[60]}
   );
   gpc1_1 gpc146 (
      {stage0_5[127]},
      {stage1_5[61]}
   );
   gpc1_1 gpc147 (
      {stage0_6[126]},
      {stage1_6[43]}
   );
   gpc1_1 gpc148 (
      {stage0_6[127]},
      {stage1_6[44]}
   );
   gpc1_1 gpc149 (
      {stage0_7[126]},
      {stage1_7[42]}
   );
   gpc1_1 gpc150 (
      {stage0_7[127]},
      {stage1_7[43]}
   );
   gpc1_1 gpc151 (
      {stage0_11[126]},
      {stage1_11[42]}
   );
   gpc1_1 gpc152 (
      {stage0_11[127]},
      {stage1_11[43]}
   );
   gpc2135_5 gpc153 (
      {stage1_0[0], stage1_0[1], stage1_0[2], stage1_0[3], stage1_0[4]},
      {stage1_1[0], stage1_1[1], stage1_1[2]},
      {stage1_2[0]},
      {stage1_3[0], stage1_3[1]},
      {stage2_4[0],stage2_3[0],stage2_2[0],stage2_1[0],stage2_0[0]}
   );
   gpc1163_5 gpc154 (
      {stage1_0[5], stage1_0[6], stage1_0[7]},
      {stage1_1[3], stage1_1[4], stage1_1[5], stage1_1[6], stage1_1[7], stage1_1[8]},
      {stage1_2[1]},
      {stage1_3[2]},
      {stage2_4[1],stage2_3[1],stage2_2[1],stage2_1[1],stage2_0[1]}
   );
   gpc1163_5 gpc155 (
      {stage1_0[8], stage1_0[9], stage1_0[10]},
      {stage1_1[9], stage1_1[10], stage1_1[11], stage1_1[12], stage1_1[13], stage1_1[14]},
      {stage1_2[2]},
      {stage1_3[3]},
      {stage2_4[2],stage2_3[2],stage2_2[2],stage2_1[2],stage2_0[2]}
   );
   gpc1163_5 gpc156 (
      {stage1_0[11], stage1_0[12], stage1_0[13]},
      {stage1_1[15], stage1_1[16], stage1_1[17], stage1_1[18], stage1_1[19], stage1_1[20]},
      {stage1_2[3]},
      {stage1_3[4]},
      {stage2_4[3],stage2_3[3],stage2_2[3],stage2_1[3],stage2_0[3]}
   );
   gpc1163_5 gpc157 (
      {stage1_0[14], stage1_0[15], stage1_0[16]},
      {stage1_1[21], stage1_1[22], stage1_1[23], stage1_1[24], stage1_1[25], stage1_1[26]},
      {stage1_2[4]},
      {stage1_3[5]},
      {stage2_4[4],stage2_3[4],stage2_2[4],stage2_1[4],stage2_0[4]}
   );
   gpc606_5 gpc158 (
      {stage1_1[27], stage1_1[28], stage1_1[29], stage1_1[30], stage1_1[31], stage1_1[32]},
      {stage1_3[6], stage1_3[7], stage1_3[8], stage1_3[9], stage1_3[10], stage1_3[11]},
      {stage2_5[0],stage2_4[5],stage2_3[5],stage2_2[5],stage2_1[5]}
   );
   gpc606_5 gpc159 (
      {stage1_1[33], stage1_1[34], stage1_1[35], stage1_1[36], stage1_1[37], stage1_1[38]},
      {stage1_3[12], stage1_3[13], stage1_3[14], stage1_3[15], stage1_3[16], stage1_3[17]},
      {stage2_5[1],stage2_4[6],stage2_3[6],stage2_2[6],stage2_1[6]}
   );
   gpc606_5 gpc160 (
      {stage1_2[5], stage1_2[6], stage1_2[7], stage1_2[8], stage1_2[9], stage1_2[10]},
      {stage1_4[0], stage1_4[1], stage1_4[2], stage1_4[3], stage1_4[4], stage1_4[5]},
      {stage2_6[0],stage2_5[2],stage2_4[7],stage2_3[7],stage2_2[7]}
   );
   gpc606_5 gpc161 (
      {stage1_2[11], stage1_2[12], stage1_2[13], stage1_2[14], stage1_2[15], stage1_2[16]},
      {stage1_4[6], stage1_4[7], stage1_4[8], stage1_4[9], stage1_4[10], stage1_4[11]},
      {stage2_6[1],stage2_5[3],stage2_4[8],stage2_3[8],stage2_2[8]}
   );
   gpc615_5 gpc162 (
      {stage1_2[17], stage1_2[18], stage1_2[19], stage1_2[20], stage1_2[21]},
      {stage1_3[18]},
      {stage1_4[12], stage1_4[13], stage1_4[14], stage1_4[15], stage1_4[16], stage1_4[17]},
      {stage2_6[2],stage2_5[4],stage2_4[9],stage2_3[9],stage2_2[9]}
   );
   gpc615_5 gpc163 (
      {stage1_2[22], stage1_2[23], stage1_2[24], stage1_2[25], stage1_2[26]},
      {stage1_3[19]},
      {stage1_4[18], stage1_4[19], stage1_4[20], stage1_4[21], stage1_4[22], stage1_4[23]},
      {stage2_6[3],stage2_5[5],stage2_4[10],stage2_3[10],stage2_2[10]}
   );
   gpc615_5 gpc164 (
      {stage1_2[27], stage1_2[28], stage1_2[29], stage1_2[30], stage1_2[31]},
      {stage1_3[20]},
      {stage1_4[24], stage1_4[25], stage1_4[26], stage1_4[27], stage1_4[28], stage1_4[29]},
      {stage2_6[4],stage2_5[6],stage2_4[11],stage2_3[11],stage2_2[11]}
   );
   gpc615_5 gpc165 (
      {stage1_2[32], stage1_2[33], stage1_2[34], stage1_2[35], stage1_2[36]},
      {stage1_3[21]},
      {stage1_4[30], stage1_4[31], stage1_4[32], stage1_4[33], stage1_4[34], stage1_4[35]},
      {stage2_6[5],stage2_5[7],stage2_4[12],stage2_3[12],stage2_2[12]}
   );
   gpc615_5 gpc166 (
      {stage1_2[37], stage1_2[38], stage1_2[39], stage1_2[40], stage1_2[41]},
      {stage1_3[22]},
      {stage1_4[36], stage1_4[37], stage1_4[38], stage1_4[39], stage1_4[40], stage1_4[41]},
      {stage2_6[6],stage2_5[8],stage2_4[13],stage2_3[13],stage2_2[13]}
   );
   gpc615_5 gpc167 (
      {stage1_3[23], stage1_3[24], stage1_3[25], stage1_3[26], stage1_3[27]},
      {stage1_4[42]},
      {stage1_5[0], stage1_5[1], stage1_5[2], stage1_5[3], stage1_5[4], stage1_5[5]},
      {stage2_7[0],stage2_6[7],stage2_5[9],stage2_4[14],stage2_3[14]}
   );
   gpc615_5 gpc168 (
      {stage1_3[28], stage1_3[29], stage1_3[30], stage1_3[31], stage1_3[32]},
      {stage1_4[43]},
      {stage1_5[6], stage1_5[7], stage1_5[8], stage1_5[9], stage1_5[10], stage1_5[11]},
      {stage2_7[1],stage2_6[8],stage2_5[10],stage2_4[15],stage2_3[15]}
   );
   gpc615_5 gpc169 (
      {stage1_3[33], stage1_3[34], stage1_3[35], stage1_3[36], stage1_3[37]},
      {stage1_4[44]},
      {stage1_5[12], stage1_5[13], stage1_5[14], stage1_5[15], stage1_5[16], stage1_5[17]},
      {stage2_7[2],stage2_6[9],stage2_5[11],stage2_4[16],stage2_3[16]}
   );
   gpc615_5 gpc170 (
      {stage1_3[38], stage1_3[39], stage1_3[40], stage1_3[41], stage1_3[42]},
      {stage1_4[45]},
      {stage1_5[18], stage1_5[19], stage1_5[20], stage1_5[21], stage1_5[22], stage1_5[23]},
      {stage2_7[3],stage2_6[10],stage2_5[12],stage2_4[17],stage2_3[17]}
   );
   gpc615_5 gpc171 (
      {stage1_3[43], stage1_3[44], stage1_3[45], stage1_3[46], stage1_3[47]},
      {stage1_4[46]},
      {stage1_5[24], stage1_5[25], stage1_5[26], stage1_5[27], stage1_5[28], stage1_5[29]},
      {stage2_7[4],stage2_6[11],stage2_5[13],stage2_4[18],stage2_3[18]}
   );
   gpc615_5 gpc172 (
      {stage1_3[48], stage1_3[49], stage1_3[50], stage1_3[51], stage1_3[52]},
      {stage1_4[47]},
      {stage1_5[30], stage1_5[31], stage1_5[32], stage1_5[33], stage1_5[34], stage1_5[35]},
      {stage2_7[5],stage2_6[12],stage2_5[14],stage2_4[19],stage2_3[19]}
   );
   gpc615_5 gpc173 (
      {stage1_3[53], stage1_3[54], stage1_3[55], stage1_3[56], stage1_3[57]},
      {stage1_4[48]},
      {stage1_5[36], stage1_5[37], stage1_5[38], stage1_5[39], stage1_5[40], stage1_5[41]},
      {stage2_7[6],stage2_6[13],stage2_5[15],stage2_4[20],stage2_3[20]}
   );
   gpc606_5 gpc174 (
      {stage1_4[49], stage1_4[50], stage1_4[51], stage1_4[52], stage1_4[53], stage1_4[54]},
      {stage1_6[0], stage1_6[1], stage1_6[2], stage1_6[3], stage1_6[4], stage1_6[5]},
      {stage2_8[0],stage2_7[7],stage2_6[14],stage2_5[16],stage2_4[21]}
   );
   gpc606_5 gpc175 (
      {stage1_4[55], stage1_4[56], stage1_4[57], stage1_4[58], stage1_4[59], stage1_4[60]},
      {stage1_6[6], stage1_6[7], stage1_6[8], stage1_6[9], stage1_6[10], stage1_6[11]},
      {stage2_8[1],stage2_7[8],stage2_6[15],stage2_5[17],stage2_4[22]}
   );
   gpc606_5 gpc176 (
      {stage1_5[42], stage1_5[43], stage1_5[44], stage1_5[45], stage1_5[46], stage1_5[47]},
      {stage1_7[0], stage1_7[1], stage1_7[2], stage1_7[3], stage1_7[4], stage1_7[5]},
      {stage2_9[0],stage2_8[2],stage2_7[9],stage2_6[16],stage2_5[18]}
   );
   gpc606_5 gpc177 (
      {stage1_5[48], stage1_5[49], stage1_5[50], stage1_5[51], stage1_5[52], stage1_5[53]},
      {stage1_7[6], stage1_7[7], stage1_7[8], stage1_7[9], stage1_7[10], stage1_7[11]},
      {stage2_9[1],stage2_8[3],stage2_7[10],stage2_6[17],stage2_5[19]}
   );
   gpc606_5 gpc178 (
      {stage1_5[54], stage1_5[55], stage1_5[56], stage1_5[57], stage1_5[58], stage1_5[59]},
      {stage1_7[12], stage1_7[13], stage1_7[14], stage1_7[15], stage1_7[16], stage1_7[17]},
      {stage2_9[2],stage2_8[4],stage2_7[11],stage2_6[18],stage2_5[20]}
   );
   gpc615_5 gpc179 (
      {stage1_6[12], stage1_6[13], stage1_6[14], stage1_6[15], stage1_6[16]},
      {stage1_7[18]},
      {stage1_8[0], stage1_8[1], stage1_8[2], stage1_8[3], stage1_8[4], stage1_8[5]},
      {stage2_10[0],stage2_9[3],stage2_8[5],stage2_7[12],stage2_6[19]}
   );
   gpc615_5 gpc180 (
      {stage1_6[17], stage1_6[18], stage1_6[19], stage1_6[20], stage1_6[21]},
      {stage1_7[19]},
      {stage1_8[6], stage1_8[7], stage1_8[8], stage1_8[9], stage1_8[10], stage1_8[11]},
      {stage2_10[1],stage2_9[4],stage2_8[6],stage2_7[13],stage2_6[20]}
   );
   gpc615_5 gpc181 (
      {stage1_6[22], stage1_6[23], stage1_6[24], stage1_6[25], stage1_6[26]},
      {stage1_7[20]},
      {stage1_8[12], stage1_8[13], stage1_8[14], stage1_8[15], stage1_8[16], stage1_8[17]},
      {stage2_10[2],stage2_9[5],stage2_8[7],stage2_7[14],stage2_6[21]}
   );
   gpc615_5 gpc182 (
      {stage1_6[27], stage1_6[28], stage1_6[29], stage1_6[30], stage1_6[31]},
      {stage1_7[21]},
      {stage1_8[18], stage1_8[19], stage1_8[20], stage1_8[21], stage1_8[22], stage1_8[23]},
      {stage2_10[3],stage2_9[6],stage2_8[8],stage2_7[15],stage2_6[22]}
   );
   gpc615_5 gpc183 (
      {stage1_6[32], stage1_6[33], stage1_6[34], stage1_6[35], stage1_6[36]},
      {stage1_7[22]},
      {stage1_8[24], stage1_8[25], stage1_8[26], stage1_8[27], stage1_8[28], stage1_8[29]},
      {stage2_10[4],stage2_9[7],stage2_8[9],stage2_7[16],stage2_6[23]}
   );
   gpc615_5 gpc184 (
      {stage1_6[37], stage1_6[38], stage1_6[39], stage1_6[40], stage1_6[41]},
      {stage1_7[23]},
      {stage1_8[30], stage1_8[31], stage1_8[32], stage1_8[33], stage1_8[34], stage1_8[35]},
      {stage2_10[5],stage2_9[8],stage2_8[10],stage2_7[17],stage2_6[24]}
   );
   gpc615_5 gpc185 (
      {stage1_7[24], stage1_7[25], stage1_7[26], stage1_7[27], stage1_7[28]},
      {stage1_8[36]},
      {stage1_9[0], stage1_9[1], stage1_9[2], stage1_9[3], stage1_9[4], stage1_9[5]},
      {stage2_11[0],stage2_10[6],stage2_9[9],stage2_8[11],stage2_7[18]}
   );
   gpc615_5 gpc186 (
      {stage1_7[29], stage1_7[30], stage1_7[31], stage1_7[32], stage1_7[33]},
      {stage1_8[37]},
      {stage1_9[6], stage1_9[7], stage1_9[8], stage1_9[9], stage1_9[10], stage1_9[11]},
      {stage2_11[1],stage2_10[7],stage2_9[10],stage2_8[12],stage2_7[19]}
   );
   gpc615_5 gpc187 (
      {stage1_7[34], stage1_7[35], stage1_7[36], stage1_7[37], stage1_7[38]},
      {stage1_8[38]},
      {stage1_9[12], stage1_9[13], stage1_9[14], stage1_9[15], stage1_9[16], stage1_9[17]},
      {stage2_11[2],stage2_10[8],stage2_9[11],stage2_8[13],stage2_7[20]}
   );
   gpc615_5 gpc188 (
      {stage1_7[39], stage1_7[40], stage1_7[41], stage1_7[42], stage1_7[43]},
      {stage1_8[39]},
      {stage1_9[18], stage1_9[19], stage1_9[20], stage1_9[21], stage1_9[22], stage1_9[23]},
      {stage2_11[3],stage2_10[9],stage2_9[12],stage2_8[14],stage2_7[21]}
   );
   gpc1163_5 gpc189 (
      {stage1_8[40], stage1_8[41], stage1_8[42]},
      {stage1_9[24], stage1_9[25], stage1_9[26], stage1_9[27], stage1_9[28], stage1_9[29]},
      {stage1_10[0]},
      {stage1_11[0]},
      {stage2_12[0],stage2_11[4],stage2_10[10],stage2_9[13],stage2_8[15]}
   );
   gpc606_5 gpc190 (
      {stage1_8[43], stage1_8[44], stage1_8[45], stage1_8[46], stage1_8[47], stage1_8[48]},
      {stage1_10[1], stage1_10[2], stage1_10[3], stage1_10[4], stage1_10[5], stage1_10[6]},
      {stage2_12[1],stage2_11[5],stage2_10[11],stage2_9[14],stage2_8[16]}
   );
   gpc615_5 gpc191 (
      {stage1_8[49], stage1_8[50], stage1_8[51], stage1_8[52], stage1_8[53]},
      {stage1_9[30]},
      {stage1_10[7], stage1_10[8], stage1_10[9], stage1_10[10], stage1_10[11], stage1_10[12]},
      {stage2_12[2],stage2_11[6],stage2_10[12],stage2_9[15],stage2_8[17]}
   );
   gpc2135_5 gpc192 (
      {stage1_9[31], stage1_9[32], stage1_9[33], stage1_9[34], stage1_9[35]},
      {stage1_10[13], stage1_10[14], stage1_10[15]},
      {stage1_11[1]},
      {stage1_12[0], stage1_12[1]},
      {stage2_13[0],stage2_12[3],stage2_11[7],stage2_10[13],stage2_9[16]}
   );
   gpc606_5 gpc193 (
      {stage1_9[36], stage1_9[37], stage1_9[38], stage1_9[39], stage1_9[40], stage1_9[41]},
      {stage1_11[2], stage1_11[3], stage1_11[4], stage1_11[5], stage1_11[6], stage1_11[7]},
      {stage2_13[1],stage2_12[4],stage2_11[8],stage2_10[14],stage2_9[17]}
   );
   gpc606_5 gpc194 (
      {stage1_9[42], stage1_9[43], stage1_9[44], stage1_9[45], stage1_9[46], stage1_9[47]},
      {stage1_11[8], stage1_11[9], stage1_11[10], stage1_11[11], stage1_11[12], stage1_11[13]},
      {stage2_13[2],stage2_12[5],stage2_11[9],stage2_10[15],stage2_9[18]}
   );
   gpc606_5 gpc195 (
      {stage1_9[48], stage1_9[49], stage1_9[50], stage1_9[51], stage1_9[52], stage1_9[53]},
      {stage1_11[14], stage1_11[15], stage1_11[16], stage1_11[17], stage1_11[18], stage1_11[19]},
      {stage2_13[3],stage2_12[6],stage2_11[10],stage2_10[16],stage2_9[19]}
   );
   gpc606_5 gpc196 (
      {stage1_9[54], stage1_9[55], stage1_9[56], stage1_9[57], stage1_9[58], stage1_9[59]},
      {stage1_11[20], stage1_11[21], stage1_11[22], stage1_11[23], stage1_11[24], stage1_11[25]},
      {stage2_13[4],stage2_12[7],stage2_11[11],stage2_10[17],stage2_9[20]}
   );
   gpc606_5 gpc197 (
      {stage1_10[16], stage1_10[17], stage1_10[18], stage1_10[19], stage1_10[20], stage1_10[21]},
      {stage1_12[2], stage1_12[3], stage1_12[4], stage1_12[5], stage1_12[6], stage1_12[7]},
      {stage2_14[0],stage2_13[5],stage2_12[8],stage2_11[12],stage2_10[18]}
   );
   gpc615_5 gpc198 (
      {stage1_10[22], stage1_10[23], stage1_10[24], stage1_10[25], stage1_10[26]},
      {stage1_11[26]},
      {stage1_12[8], stage1_12[9], stage1_12[10], stage1_12[11], stage1_12[12], stage1_12[13]},
      {stage2_14[1],stage2_13[6],stage2_12[9],stage2_11[13],stage2_10[19]}
   );
   gpc615_5 gpc199 (
      {stage1_10[27], stage1_10[28], stage1_10[29], stage1_10[30], stage1_10[31]},
      {stage1_11[27]},
      {stage1_12[14], stage1_12[15], stage1_12[16], stage1_12[17], stage1_12[18], stage1_12[19]},
      {stage2_14[2],stage2_13[7],stage2_12[10],stage2_11[14],stage2_10[20]}
   );
   gpc615_5 gpc200 (
      {stage1_10[32], stage1_10[33], stage1_10[34], stage1_10[35], stage1_10[36]},
      {stage1_11[28]},
      {stage1_12[20], stage1_12[21], stage1_12[22], stage1_12[23], stage1_12[24], stage1_12[25]},
      {stage2_14[3],stage2_13[8],stage2_12[11],stage2_11[15],stage2_10[21]}
   );
   gpc615_5 gpc201 (
      {stage1_10[37], stage1_10[38], stage1_10[39], stage1_10[40], stage1_10[41]},
      {stage1_11[29]},
      {stage1_12[26], stage1_12[27], stage1_12[28], stage1_12[29], stage1_12[30], stage1_12[31]},
      {stage2_14[4],stage2_13[9],stage2_12[12],stage2_11[16],stage2_10[22]}
   );
   gpc615_5 gpc202 (
      {stage1_11[30], stage1_11[31], stage1_11[32], stage1_11[33], stage1_11[34]},
      {stage1_12[32]},
      {stage1_13[0], stage1_13[1], stage1_13[2], stage1_13[3], stage1_13[4], stage1_13[5]},
      {stage2_15[0],stage2_14[5],stage2_13[10],stage2_12[13],stage2_11[17]}
   );
   gpc615_5 gpc203 (
      {stage1_11[35], stage1_11[36], stage1_11[37], stage1_11[38], stage1_11[39]},
      {stage1_12[33]},
      {stage1_13[6], stage1_13[7], stage1_13[8], stage1_13[9], stage1_13[10], stage1_13[11]},
      {stage2_15[1],stage2_14[6],stage2_13[11],stage2_12[14],stage2_11[18]}
   );
   gpc615_5 gpc204 (
      {stage1_11[40], stage1_11[41], stage1_11[42], stage1_11[43], 1'b0},
      {stage1_12[34]},
      {stage1_13[12], stage1_13[13], stage1_13[14], stage1_13[15], stage1_13[16], stage1_13[17]},
      {stage2_15[2],stage2_14[7],stage2_13[12],stage2_12[15],stage2_11[19]}
   );
   gpc117_4 gpc205 (
      {stage1_12[35], stage1_12[36], stage1_12[37], stage1_12[38], stage1_12[39], stage1_12[40], stage1_12[41]},
      {stage1_13[18]},
      {1'b0},
      {stage2_15[3],stage2_14[8],stage2_13[13],stage2_12[16]}
   );
   gpc1_1 gpc206 (
      {stage1_0[17]},
      {stage2_0[5]}
   );
   gpc1_1 gpc207 (
      {stage1_0[18]},
      {stage2_0[6]}
   );
   gpc1_1 gpc208 (
      {stage1_0[19]},
      {stage2_0[7]}
   );
   gpc1_1 gpc209 (
      {stage1_0[20]},
      {stage2_0[8]}
   );
   gpc1_1 gpc210 (
      {stage1_0[21]},
      {stage2_0[9]}
   );
   gpc1_1 gpc211 (
      {stage1_0[22]},
      {stage2_0[10]}
   );
   gpc1_1 gpc212 (
      {stage1_0[23]},
      {stage2_0[11]}
   );
   gpc1_1 gpc213 (
      {stage1_1[39]},
      {stage2_1[7]}
   );
   gpc1_1 gpc214 (
      {stage1_1[40]},
      {stage2_1[8]}
   );
   gpc1_1 gpc215 (
      {stage1_4[61]},
      {stage2_4[23]}
   );
   gpc1_1 gpc216 (
      {stage1_4[62]},
      {stage2_4[24]}
   );
   gpc1_1 gpc217 (
      {stage1_4[63]},
      {stage2_4[25]}
   );
   gpc1_1 gpc218 (
      {stage1_5[60]},
      {stage2_5[21]}
   );
   gpc1_1 gpc219 (
      {stage1_5[61]},
      {stage2_5[22]}
   );
   gpc1_1 gpc220 (
      {stage1_6[42]},
      {stage2_6[25]}
   );
   gpc1_1 gpc221 (
      {stage1_6[43]},
      {stage2_6[26]}
   );
   gpc1_1 gpc222 (
      {stage1_6[44]},
      {stage2_6[27]}
   );
   gpc1_1 gpc223 (
      {stage1_8[54]},
      {stage2_8[18]}
   );
   gpc1_1 gpc224 (
      {stage1_8[55]},
      {stage2_8[19]}
   );
   gpc1_1 gpc225 (
      {stage1_8[56]},
      {stage2_8[20]}
   );
   gpc1_1 gpc226 (
      {stage1_8[57]},
      {stage2_8[21]}
   );
   gpc1_1 gpc227 (
      {stage1_8[58]},
      {stage2_8[22]}
   );
   gpc1_1 gpc228 (
      {stage1_8[59]},
      {stage2_8[23]}
   );
   gpc1_1 gpc229 (
      {stage1_8[60]},
      {stage2_8[24]}
   );
   gpc1_1 gpc230 (
      {stage1_8[61]},
      {stage2_8[25]}
   );
   gpc1_1 gpc231 (
      {stage1_8[62]},
      {stage2_8[26]}
   );
   gpc1_1 gpc232 (
      {stage1_9[60]},
      {stage2_9[21]}
   );
   gpc1_1 gpc233 (
      {stage1_9[61]},
      {stage2_9[22]}
   );
   gpc1_1 gpc234 (
      {stage1_9[62]},
      {stage2_9[23]}
   );
   gpc1_1 gpc235 (
      {stage1_9[63]},
      {stage2_9[24]}
   );
   gpc1_1 gpc236 (
      {stage1_10[42]},
      {stage2_10[23]}
   );
   gpc1_1 gpc237 (
      {stage1_13[19]},
      {stage2_13[14]}
   );
   gpc1_1 gpc238 (
      {stage1_13[20]},
      {stage2_13[15]}
   );
   gpc606_5 gpc239 (
      {stage2_0[0], stage2_0[1], stage2_0[2], stage2_0[3], stage2_0[4], stage2_0[5]},
      {stage2_2[0], stage2_2[1], stage2_2[2], stage2_2[3], stage2_2[4], stage2_2[5]},
      {stage3_4[0],stage3_3[0],stage3_2[0],stage3_1[0],stage3_0[0]}
   );
   gpc606_5 gpc240 (
      {stage2_1[0], stage2_1[1], stage2_1[2], stage2_1[3], stage2_1[4], stage2_1[5]},
      {stage2_3[0], stage2_3[1], stage2_3[2], stage2_3[3], stage2_3[4], stage2_3[5]},
      {stage3_5[0],stage3_4[1],stage3_3[1],stage3_2[1],stage3_1[1]}
   );
   gpc615_5 gpc241 (
      {stage2_2[6], stage2_2[7], stage2_2[8], stage2_2[9], stage2_2[10]},
      {stage2_3[6]},
      {stage2_4[0], stage2_4[1], stage2_4[2], stage2_4[3], stage2_4[4], stage2_4[5]},
      {stage3_6[0],stage3_5[1],stage3_4[2],stage3_3[2],stage3_2[2]}
   );
   gpc615_5 gpc242 (
      {stage2_3[7], stage2_3[8], stage2_3[9], stage2_3[10], stage2_3[11]},
      {stage2_4[6]},
      {stage2_5[0], stage2_5[1], stage2_5[2], stage2_5[3], stage2_5[4], stage2_5[5]},
      {stage3_7[0],stage3_6[1],stage3_5[2],stage3_4[3],stage3_3[3]}
   );
   gpc615_5 gpc243 (
      {stage2_3[12], stage2_3[13], stage2_3[14], stage2_3[15], stage2_3[16]},
      {stage2_4[7]},
      {stage2_5[6], stage2_5[7], stage2_5[8], stage2_5[9], stage2_5[10], stage2_5[11]},
      {stage3_7[1],stage3_6[2],stage3_5[3],stage3_4[4],stage3_3[4]}
   );
   gpc615_5 gpc244 (
      {stage2_3[17], stage2_3[18], stage2_3[19], stage2_3[20], 1'b0},
      {stage2_4[8]},
      {stage2_5[12], stage2_5[13], stage2_5[14], stage2_5[15], stage2_5[16], stage2_5[17]},
      {stage3_7[2],stage3_6[3],stage3_5[4],stage3_4[5],stage3_3[5]}
   );
   gpc606_5 gpc245 (
      {stage2_4[9], stage2_4[10], stage2_4[11], stage2_4[12], stage2_4[13], stage2_4[14]},
      {stage2_6[0], stage2_6[1], stage2_6[2], stage2_6[3], stage2_6[4], stage2_6[5]},
      {stage3_8[0],stage3_7[3],stage3_6[4],stage3_5[5],stage3_4[6]}
   );
   gpc606_5 gpc246 (
      {stage2_4[15], stage2_4[16], stage2_4[17], stage2_4[18], stage2_4[19], stage2_4[20]},
      {stage2_6[6], stage2_6[7], stage2_6[8], stage2_6[9], stage2_6[10], stage2_6[11]},
      {stage3_8[1],stage3_7[4],stage3_6[5],stage3_5[6],stage3_4[7]}
   );
   gpc615_5 gpc247 (
      {stage2_4[21], stage2_4[22], stage2_4[23], stage2_4[24], stage2_4[25]},
      {stage2_5[18]},
      {stage2_6[12], stage2_6[13], stage2_6[14], stage2_6[15], stage2_6[16], stage2_6[17]},
      {stage3_8[2],stage3_7[5],stage3_6[6],stage3_5[7],stage3_4[8]}
   );
   gpc615_5 gpc248 (
      {stage2_6[18], stage2_6[19], stage2_6[20], stage2_6[21], stage2_6[22]},
      {stage2_7[0]},
      {stage2_8[0], stage2_8[1], stage2_8[2], stage2_8[3], stage2_8[4], stage2_8[5]},
      {stage3_10[0],stage3_9[0],stage3_8[3],stage3_7[6],stage3_6[7]}
   );
   gpc615_5 gpc249 (
      {stage2_6[23], stage2_6[24], stage2_6[25], stage2_6[26], stage2_6[27]},
      {stage2_7[1]},
      {stage2_8[6], stage2_8[7], stage2_8[8], stage2_8[9], stage2_8[10], stage2_8[11]},
      {stage3_10[1],stage3_9[1],stage3_8[4],stage3_7[7],stage3_6[8]}
   );
   gpc615_5 gpc250 (
      {stage2_7[2], stage2_7[3], stage2_7[4], stage2_7[5], stage2_7[6]},
      {stage2_8[12]},
      {stage2_9[0], stage2_9[1], stage2_9[2], stage2_9[3], stage2_9[4], stage2_9[5]},
      {stage3_11[0],stage3_10[2],stage3_9[2],stage3_8[5],stage3_7[8]}
   );
   gpc615_5 gpc251 (
      {stage2_7[7], stage2_7[8], stage2_7[9], stage2_7[10], stage2_7[11]},
      {stage2_8[13]},
      {stage2_9[6], stage2_9[7], stage2_9[8], stage2_9[9], stage2_9[10], stage2_9[11]},
      {stage3_11[1],stage3_10[3],stage3_9[3],stage3_8[6],stage3_7[9]}
   );
   gpc615_5 gpc252 (
      {stage2_7[12], stage2_7[13], stage2_7[14], stage2_7[15], stage2_7[16]},
      {stage2_8[14]},
      {stage2_9[12], stage2_9[13], stage2_9[14], stage2_9[15], stage2_9[16], stage2_9[17]},
      {stage3_11[2],stage3_10[4],stage3_9[4],stage3_8[7],stage3_7[10]}
   );
   gpc615_5 gpc253 (
      {stage2_7[17], stage2_7[18], stage2_7[19], stage2_7[20], stage2_7[21]},
      {stage2_8[15]},
      {stage2_9[18], stage2_9[19], stage2_9[20], stage2_9[21], stage2_9[22], stage2_9[23]},
      {stage3_11[3],stage3_10[5],stage3_9[5],stage3_8[8],stage3_7[11]}
   );
   gpc606_5 gpc254 (
      {stage2_8[16], stage2_8[17], stage2_8[18], stage2_8[19], stage2_8[20], stage2_8[21]},
      {stage2_10[0], stage2_10[1], stage2_10[2], stage2_10[3], stage2_10[4], stage2_10[5]},
      {stage3_12[0],stage3_11[4],stage3_10[6],stage3_9[6],stage3_8[9]}
   );
   gpc615_5 gpc255 (
      {stage2_8[22], stage2_8[23], stage2_8[24], stage2_8[25], stage2_8[26]},
      {stage2_9[24]},
      {stage2_10[6], stage2_10[7], stage2_10[8], stage2_10[9], stage2_10[10], stage2_10[11]},
      {stage3_12[1],stage3_11[5],stage3_10[7],stage3_9[7],stage3_8[10]}
   );
   gpc615_5 gpc256 (
      {stage2_10[12], stage2_10[13], stage2_10[14], stage2_10[15], stage2_10[16]},
      {stage2_11[0]},
      {stage2_12[0], stage2_12[1], stage2_12[2], stage2_12[3], stage2_12[4], stage2_12[5]},
      {stage3_14[0],stage3_13[0],stage3_12[2],stage3_11[6],stage3_10[8]}
   );
   gpc615_5 gpc257 (
      {stage2_10[17], stage2_10[18], stage2_10[19], stage2_10[20], stage2_10[21]},
      {stage2_11[1]},
      {stage2_12[6], stage2_12[7], stage2_12[8], stage2_12[9], stage2_12[10], stage2_12[11]},
      {stage3_14[1],stage3_13[1],stage3_12[3],stage3_11[7],stage3_10[9]}
   );
   gpc606_5 gpc258 (
      {stage2_11[2], stage2_11[3], stage2_11[4], stage2_11[5], stage2_11[6], stage2_11[7]},
      {stage2_13[0], stage2_13[1], stage2_13[2], stage2_13[3], stage2_13[4], stage2_13[5]},
      {stage3_15[0],stage3_14[2],stage3_13[2],stage3_12[4],stage3_11[8]}
   );
   gpc606_5 gpc259 (
      {stage2_11[8], stage2_11[9], stage2_11[10], stage2_11[11], stage2_11[12], stage2_11[13]},
      {stage2_13[6], stage2_13[7], stage2_13[8], stage2_13[9], stage2_13[10], stage2_13[11]},
      {stage3_15[1],stage3_14[3],stage3_13[3],stage3_12[5],stage3_11[9]}
   );
   gpc606_5 gpc260 (
      {stage2_11[14], stage2_11[15], stage2_11[16], stage2_11[17], stage2_11[18], stage2_11[19]},
      {stage2_13[12], stage2_13[13], stage2_13[14], stage2_13[15], 1'b0, 1'b0},
      {stage3_15[2],stage3_14[4],stage3_13[4],stage3_12[6],stage3_11[10]}
   );
   gpc606_5 gpc261 (
      {stage2_12[12], stage2_12[13], stage2_12[14], stage2_12[15], stage2_12[16], 1'b0},
      {stage2_14[0], stage2_14[1], stage2_14[2], stage2_14[3], stage2_14[4], stage2_14[5]},
      {stage3_16[0],stage3_15[3],stage3_14[5],stage3_13[5],stage3_12[7]}
   );
   gpc1_1 gpc262 (
      {stage2_0[6]},
      {stage3_0[1]}
   );
   gpc1_1 gpc263 (
      {stage2_0[7]},
      {stage3_0[2]}
   );
   gpc1_1 gpc264 (
      {stage2_0[8]},
      {stage3_0[3]}
   );
   gpc1_1 gpc265 (
      {stage2_0[9]},
      {stage3_0[4]}
   );
   gpc1_1 gpc266 (
      {stage2_0[10]},
      {stage3_0[5]}
   );
   gpc1_1 gpc267 (
      {stage2_0[11]},
      {stage3_0[6]}
   );
   gpc1_1 gpc268 (
      {stage2_1[6]},
      {stage3_1[2]}
   );
   gpc1_1 gpc269 (
      {stage2_1[7]},
      {stage3_1[3]}
   );
   gpc1_1 gpc270 (
      {stage2_1[8]},
      {stage3_1[4]}
   );
   gpc1_1 gpc271 (
      {stage2_2[11]},
      {stage3_2[3]}
   );
   gpc1_1 gpc272 (
      {stage2_2[12]},
      {stage3_2[4]}
   );
   gpc1_1 gpc273 (
      {stage2_2[13]},
      {stage3_2[5]}
   );
   gpc1_1 gpc274 (
      {stage2_5[19]},
      {stage3_5[8]}
   );
   gpc1_1 gpc275 (
      {stage2_5[20]},
      {stage3_5[9]}
   );
   gpc1_1 gpc276 (
      {stage2_5[21]},
      {stage3_5[10]}
   );
   gpc1_1 gpc277 (
      {stage2_5[22]},
      {stage3_5[11]}
   );
   gpc1_1 gpc278 (
      {stage2_10[22]},
      {stage3_10[10]}
   );
   gpc1_1 gpc279 (
      {stage2_10[23]},
      {stage3_10[11]}
   );
   gpc1_1 gpc280 (
      {stage2_14[6]},
      {stage3_14[6]}
   );
   gpc1_1 gpc281 (
      {stage2_14[7]},
      {stage3_14[7]}
   );
   gpc1_1 gpc282 (
      {stage2_14[8]},
      {stage3_14[8]}
   );
   gpc1_1 gpc283 (
      {stage2_15[0]},
      {stage3_15[4]}
   );
   gpc1_1 gpc284 (
      {stage2_15[1]},
      {stage3_15[5]}
   );
   gpc1_1 gpc285 (
      {stage2_15[2]},
      {stage3_15[6]}
   );
   gpc1_1 gpc286 (
      {stage2_15[3]},
      {stage3_15[7]}
   );
   gpc606_5 gpc287 (
      {stage3_1[0], stage3_1[1], stage3_1[2], stage3_1[3], stage3_1[4], 1'b0},
      {stage3_3[0], stage3_3[1], stage3_3[2], stage3_3[3], stage3_3[4], stage3_3[5]},
      {stage4_5[0],stage4_4[0],stage4_3[0],stage4_2[0],stage4_1[0]}
   );
   gpc606_5 gpc288 (
      {stage3_4[0], stage3_4[1], stage3_4[2], stage3_4[3], stage3_4[4], stage3_4[5]},
      {stage3_6[0], stage3_6[1], stage3_6[2], stage3_6[3], stage3_6[4], stage3_6[5]},
      {stage4_8[0],stage4_7[0],stage4_6[0],stage4_5[1],stage4_4[1]}
   );
   gpc606_5 gpc289 (
      {stage3_5[0], stage3_5[1], stage3_5[2], stage3_5[3], stage3_5[4], stage3_5[5]},
      {stage3_7[0], stage3_7[1], stage3_7[2], stage3_7[3], stage3_7[4], stage3_7[5]},
      {stage4_9[0],stage4_8[1],stage4_7[1],stage4_6[1],stage4_5[2]}
   );
   gpc606_5 gpc290 (
      {stage3_5[6], stage3_5[7], stage3_5[8], stage3_5[9], stage3_5[10], stage3_5[11]},
      {stage3_7[6], stage3_7[7], stage3_7[8], stage3_7[9], stage3_7[10], stage3_7[11]},
      {stage4_9[1],stage4_8[2],stage4_7[2],stage4_6[2],stage4_5[3]}
   );
   gpc615_5 gpc291 (
      {stage3_8[0], stage3_8[1], stage3_8[2], stage3_8[3], stage3_8[4]},
      {stage3_9[0]},
      {stage3_10[0], stage3_10[1], stage3_10[2], stage3_10[3], stage3_10[4], stage3_10[5]},
      {stage4_12[0],stage4_11[0],stage4_10[0],stage4_9[2],stage4_8[3]}
   );
   gpc615_5 gpc292 (
      {stage3_8[5], stage3_8[6], stage3_8[7], stage3_8[8], stage3_8[9]},
      {stage3_9[1]},
      {stage3_10[6], stage3_10[7], stage3_10[8], stage3_10[9], stage3_10[10], stage3_10[11]},
      {stage4_12[1],stage4_11[1],stage4_10[1],stage4_9[3],stage4_8[4]}
   );
   gpc606_5 gpc293 (
      {stage3_9[2], stage3_9[3], stage3_9[4], stage3_9[5], stage3_9[6], stage3_9[7]},
      {stage3_11[0], stage3_11[1], stage3_11[2], stage3_11[3], stage3_11[4], stage3_11[5]},
      {stage4_13[0],stage4_12[2],stage4_11[2],stage4_10[2],stage4_9[4]}
   );
   gpc615_5 gpc294 (
      {stage3_11[6], stage3_11[7], stage3_11[8], stage3_11[9], stage3_11[10]},
      {stage3_12[0]},
      {stage3_13[0], stage3_13[1], stage3_13[2], stage3_13[3], stage3_13[4], stage3_13[5]},
      {stage4_15[0],stage4_14[0],stage4_13[1],stage4_12[3],stage4_11[3]}
   );
   gpc606_5 gpc295 (
      {stage3_12[1], stage3_12[2], stage3_12[3], stage3_12[4], stage3_12[5], stage3_12[6]},
      {stage3_14[0], stage3_14[1], stage3_14[2], stage3_14[3], stage3_14[4], stage3_14[5]},
      {stage4_16[0],stage4_15[1],stage4_14[1],stage4_13[2],stage4_12[4]}
   );
   gpc1163_5 gpc296 (
      {stage3_14[6], stage3_14[7], stage3_14[8]},
      {stage3_15[0], stage3_15[1], stage3_15[2], stage3_15[3], stage3_15[4], stage3_15[5]},
      {stage3_16[0]},
      {1'b0},
      {stage4_18[0],stage4_17[0],stage4_16[1],stage4_15[2],stage4_14[2]}
   );
   gpc1_1 gpc297 (
      {stage3_0[0]},
      {stage4_0[0]}
   );
   gpc1_1 gpc298 (
      {stage3_0[1]},
      {stage4_0[1]}
   );
   gpc1_1 gpc299 (
      {stage3_0[2]},
      {stage4_0[2]}
   );
   gpc1_1 gpc300 (
      {stage3_0[3]},
      {stage4_0[3]}
   );
   gpc1_1 gpc301 (
      {stage3_0[4]},
      {stage4_0[4]}
   );
   gpc1_1 gpc302 (
      {stage3_0[5]},
      {stage4_0[5]}
   );
   gpc1_1 gpc303 (
      {stage3_0[6]},
      {stage4_0[6]}
   );
   gpc1_1 gpc304 (
      {stage3_2[0]},
      {stage4_2[1]}
   );
   gpc1_1 gpc305 (
      {stage3_2[1]},
      {stage4_2[2]}
   );
   gpc1_1 gpc306 (
      {stage3_2[2]},
      {stage4_2[3]}
   );
   gpc1_1 gpc307 (
      {stage3_2[3]},
      {stage4_2[4]}
   );
   gpc1_1 gpc308 (
      {stage3_2[4]},
      {stage4_2[5]}
   );
   gpc1_1 gpc309 (
      {stage3_2[5]},
      {stage4_2[6]}
   );
   gpc1_1 gpc310 (
      {stage3_4[6]},
      {stage4_4[2]}
   );
   gpc1_1 gpc311 (
      {stage3_4[7]},
      {stage4_4[3]}
   );
   gpc1_1 gpc312 (
      {stage3_4[8]},
      {stage4_4[4]}
   );
   gpc1_1 gpc313 (
      {stage3_6[6]},
      {stage4_6[3]}
   );
   gpc1_1 gpc314 (
      {stage3_6[7]},
      {stage4_6[4]}
   );
   gpc1_1 gpc315 (
      {stage3_6[8]},
      {stage4_6[5]}
   );
   gpc1_1 gpc316 (
      {stage3_8[10]},
      {stage4_8[5]}
   );
   gpc1_1 gpc317 (
      {stage3_12[7]},
      {stage4_12[5]}
   );
   gpc1_1 gpc318 (
      {stage3_15[6]},
      {stage4_15[3]}
   );
   gpc1_1 gpc319 (
      {stage3_15[7]},
      {stage4_15[4]}
   );
   gpc606_5 gpc320 (
      {stage4_0[0], stage4_0[1], stage4_0[2], stage4_0[3], stage4_0[4], stage4_0[5]},
      {stage4_2[0], stage4_2[1], stage4_2[2], stage4_2[3], stage4_2[4], stage4_2[5]},
      {stage5_4[0],stage5_3[0],stage5_2[0],stage5_1[0],stage5_0[0]}
   );
   gpc2135_5 gpc321 (
      {stage4_4[0], stage4_4[1], stage4_4[2], stage4_4[3], stage4_4[4]},
      {stage4_5[0], stage4_5[1], stage4_5[2]},
      {stage4_6[0]},
      {stage4_7[0], stage4_7[1]},
      {stage5_8[0],stage5_7[0],stage5_6[0],stage5_5[0],stage5_4[1]}
   );
   gpc615_5 gpc322 (
      {stage4_6[1], stage4_6[2], stage4_6[3], stage4_6[4], stage4_6[5]},
      {stage4_7[2]},
      {stage4_8[0], stage4_8[1], stage4_8[2], stage4_8[3], stage4_8[4], stage4_8[5]},
      {stage5_10[0],stage5_9[0],stage5_8[1],stage5_7[1],stage5_6[1]}
   );
   gpc2135_5 gpc323 (
      {stage4_9[0], stage4_9[1], stage4_9[2], stage4_9[3], stage4_9[4]},
      {stage4_10[0], stage4_10[1], stage4_10[2]},
      {stage4_11[0]},
      {stage4_12[0], stage4_12[1]},
      {stage5_13[0],stage5_12[0],stage5_11[0],stage5_10[1],stage5_9[1]}
   );
   gpc1343_5 gpc324 (
      {stage4_11[1], stage4_11[2], stage4_11[3]},
      {stage4_12[2], stage4_12[3], stage4_12[4], stage4_12[5]},
      {stage4_13[0], stage4_13[1], stage4_13[2]},
      {stage4_14[0]},
      {stage5_15[0],stage5_14[0],stage5_13[1],stage5_12[1],stage5_11[1]}
   );
   gpc1163_5 gpc325 (
      {stage4_14[1], stage4_14[2], 1'b0},
      {stage4_15[0], stage4_15[1], stage4_15[2], stage4_15[3], stage4_15[4], 1'b0},
      {stage4_16[0]},
      {stage4_17[0]},
      {stage5_18[0],stage5_17[0],stage5_16[0],stage5_15[1],stage5_14[1]}
   );
   gpc1_1 gpc326 (
      {stage4_0[6]},
      {stage5_0[1]}
   );
   gpc1_1 gpc327 (
      {stage4_1[0]},
      {stage5_1[1]}
   );
   gpc1_1 gpc328 (
      {stage4_2[6]},
      {stage5_2[1]}
   );
   gpc1_1 gpc329 (
      {stage4_3[0]},
      {stage5_3[1]}
   );
   gpc1_1 gpc330 (
      {stage4_5[3]},
      {stage5_5[1]}
   );
   gpc1_1 gpc331 (
      {stage4_16[1]},
      {stage5_16[1]}
   );
   gpc1_1 gpc332 (
      {stage4_18[0]},
      {stage5_18[1]}
   );
endmodule
module rowadder2_1_19(input [18:0] src0, input [18:0] src1, output [19:0] dst0);
    wire [18:0] gene;
    wire [18:0] prop;
    wire [19:0] out;
    wire [19:0] carryout;
    LUT2 #(
        .INIT(4'h8)
    ) lut_0_gene (
        .I0(src0[0]),
        .I1(src1[0]),
        .O(gene[0])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_0_prop (
        .I0(src0[0]),
        .I1(src1[0]),
        .O(prop[0])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_1_gene (
        .I0(src0[1]),
        .I1(src1[1]),
        .O(gene[1])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_1_prop (
        .I0(src0[1]),
        .I1(src1[1]),
        .O(prop[1])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_2_gene (
        .I0(src0[2]),
        .I1(src1[2]),
        .O(gene[2])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_2_prop (
        .I0(src0[2]),
        .I1(src1[2]),
        .O(prop[2])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_3_gene (
        .I0(src0[3]),
        .I1(src1[3]),
        .O(gene[3])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_3_prop (
        .I0(src0[3]),
        .I1(src1[3]),
        .O(prop[3])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_4_gene (
        .I0(src0[4]),
        .I1(src1[4]),
        .O(gene[4])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_4_prop (
        .I0(src0[4]),
        .I1(src1[4]),
        .O(prop[4])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_5_gene (
        .I0(src0[5]),
        .I1(src1[5]),
        .O(gene[5])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_5_prop (
        .I0(src0[5]),
        .I1(src1[5]),
        .O(prop[5])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_6_gene (
        .I0(src0[6]),
        .I1(src1[6]),
        .O(gene[6])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_6_prop (
        .I0(src0[6]),
        .I1(src1[6]),
        .O(prop[6])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_7_gene (
        .I0(src0[7]),
        .I1(src1[7]),
        .O(gene[7])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_7_prop (
        .I0(src0[7]),
        .I1(src1[7]),
        .O(prop[7])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_8_gene (
        .I0(src0[8]),
        .I1(src1[8]),
        .O(gene[8])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_8_prop (
        .I0(src0[8]),
        .I1(src1[8]),
        .O(prop[8])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_9_gene (
        .I0(src0[9]),
        .I1(src1[9]),
        .O(gene[9])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_9_prop (
        .I0(src0[9]),
        .I1(src1[9]),
        .O(prop[9])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_10_gene (
        .I0(src0[10]),
        .I1(src1[10]),
        .O(gene[10])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_10_prop (
        .I0(src0[10]),
        .I1(src1[10]),
        .O(prop[10])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_11_gene (
        .I0(src0[11]),
        .I1(src1[11]),
        .O(gene[11])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_11_prop (
        .I0(src0[11]),
        .I1(src1[11]),
        .O(prop[11])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_12_gene (
        .I0(src0[12]),
        .I1(src1[12]),
        .O(gene[12])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_12_prop (
        .I0(src0[12]),
        .I1(src1[12]),
        .O(prop[12])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_13_gene (
        .I0(src0[13]),
        .I1(src1[13]),
        .O(gene[13])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_13_prop (
        .I0(src0[13]),
        .I1(src1[13]),
        .O(prop[13])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_14_gene (
        .I0(src0[14]),
        .I1(src1[14]),
        .O(gene[14])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_14_prop (
        .I0(src0[14]),
        .I1(src1[14]),
        .O(prop[14])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_15_gene (
        .I0(src0[15]),
        .I1(src1[15]),
        .O(gene[15])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_15_prop (
        .I0(src0[15]),
        .I1(src1[15]),
        .O(prop[15])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_16_gene (
        .I0(src0[16]),
        .I1(src1[16]),
        .O(gene[16])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_16_prop (
        .I0(src0[16]),
        .I1(src1[16]),
        .O(prop[16])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_17_gene (
        .I0(src0[17]),
        .I1(src1[17]),
        .O(gene[17])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_17_prop (
        .I0(src0[17]),
        .I1(src1[17]),
        .O(prop[17])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_18_gene (
        .I0(src0[18]),
        .I1(src1[18]),
        .O(gene[18])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_18_prop (
        .I0(src0[18]),
        .I1(src1[18]),
        .O(prop[18])
    );
    CARRY4 carry4_3_0 (
        .CO(carryout[3:0]),
        .O(out[3:0]),
        .CI(1'h0),
        .CYINIT(1'h0),
        .DI(gene[3:0]),
        .S(prop[3:0])
    );
    CARRY4 carry4_7_4 (
        .CO(carryout[7:4]),
        .O(out[7:4]),
        .CI(carryout[3]),
        .CYINIT(1'h0),
        .DI(gene[7:4]),
        .S(prop[7:4])
    );
    CARRY4 carry4_11_8 (
        .CO(carryout[11:8]),
        .O(out[11:8]),
        .CI(carryout[7]),
        .CYINIT(1'h0),
        .DI(gene[11:8]),
        .S(prop[11:8])
    );
    CARRY4 carry4_15_12 (
        .CO(carryout[15:12]),
        .O(out[15:12]),
        .CI(carryout[11]),
        .CYINIT(1'h0),
        .DI(gene[15:12]),
        .S(prop[15:12])
    );
    CARRY4 carry4_19_16 (
        .CO(carryout[19:16]),
        .O(out[19:16]),
        .CI(carryout[15]),
        .CYINIT(1'h0),
        .DI({1'h0, gene[18:16]}),
        .S({1'h0, prop[18:16]})
    );
    assign dst0 = {carryout[18], out[18:0]};
endmodule


module testbench();
    reg [127:0] src0;
    reg [127:0] src1;
    reg [127:0] src2;
    reg [127:0] src3;
    reg [127:0] src4;
    reg [127:0] src5;
    reg [127:0] src6;
    reg [127:0] src7;
    reg [127:0] src8;
    reg [127:0] src9;
    reg [127:0] src10;
    reg [127:0] src11;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [18:0] srcsum;
    wire [18:0] dstsum;
    wire test;
    compressor2_1_128_12 compressor2_1_128_12(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13] + src0[14] + src0[15] + src0[16] + src0[17] + src0[18] + src0[19] + src0[20] + src0[21] + src0[22] + src0[23] + src0[24] + src0[25] + src0[26] + src0[27] + src0[28] + src0[29] + src0[30] + src0[31] + src0[32] + src0[33] + src0[34] + src0[35] + src0[36] + src0[37] + src0[38] + src0[39] + src0[40] + src0[41] + src0[42] + src0[43] + src0[44] + src0[45] + src0[46] + src0[47] + src0[48] + src0[49] + src0[50] + src0[51] + src0[52] + src0[53] + src0[54] + src0[55] + src0[56] + src0[57] + src0[58] + src0[59] + src0[60] + src0[61] + src0[62] + src0[63] + src0[64] + src0[65] + src0[66] + src0[67] + src0[68] + src0[69] + src0[70] + src0[71] + src0[72] + src0[73] + src0[74] + src0[75] + src0[76] + src0[77] + src0[78] + src0[79] + src0[80] + src0[81] + src0[82] + src0[83] + src0[84] + src0[85] + src0[86] + src0[87] + src0[88] + src0[89] + src0[90] + src0[91] + src0[92] + src0[93] + src0[94] + src0[95] + src0[96] + src0[97] + src0[98] + src0[99] + src0[100] + src0[101] + src0[102] + src0[103] + src0[104] + src0[105] + src0[106] + src0[107] + src0[108] + src0[109] + src0[110] + src0[111] + src0[112] + src0[113] + src0[114] + src0[115] + src0[116] + src0[117] + src0[118] + src0[119] + src0[120] + src0[121] + src0[122] + src0[123] + src0[124] + src0[125] + src0[126] + src0[127])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13] + src1[14] + src1[15] + src1[16] + src1[17] + src1[18] + src1[19] + src1[20] + src1[21] + src1[22] + src1[23] + src1[24] + src1[25] + src1[26] + src1[27] + src1[28] + src1[29] + src1[30] + src1[31] + src1[32] + src1[33] + src1[34] + src1[35] + src1[36] + src1[37] + src1[38] + src1[39] + src1[40] + src1[41] + src1[42] + src1[43] + src1[44] + src1[45] + src1[46] + src1[47] + src1[48] + src1[49] + src1[50] + src1[51] + src1[52] + src1[53] + src1[54] + src1[55] + src1[56] + src1[57] + src1[58] + src1[59] + src1[60] + src1[61] + src1[62] + src1[63] + src1[64] + src1[65] + src1[66] + src1[67] + src1[68] + src1[69] + src1[70] + src1[71] + src1[72] + src1[73] + src1[74] + src1[75] + src1[76] + src1[77] + src1[78] + src1[79] + src1[80] + src1[81] + src1[82] + src1[83] + src1[84] + src1[85] + src1[86] + src1[87] + src1[88] + src1[89] + src1[90] + src1[91] + src1[92] + src1[93] + src1[94] + src1[95] + src1[96] + src1[97] + src1[98] + src1[99] + src1[100] + src1[101] + src1[102] + src1[103] + src1[104] + src1[105] + src1[106] + src1[107] + src1[108] + src1[109] + src1[110] + src1[111] + src1[112] + src1[113] + src1[114] + src1[115] + src1[116] + src1[117] + src1[118] + src1[119] + src1[120] + src1[121] + src1[122] + src1[123] + src1[124] + src1[125] + src1[126] + src1[127])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13] + src2[14] + src2[15] + src2[16] + src2[17] + src2[18] + src2[19] + src2[20] + src2[21] + src2[22] + src2[23] + src2[24] + src2[25] + src2[26] + src2[27] + src2[28] + src2[29] + src2[30] + src2[31] + src2[32] + src2[33] + src2[34] + src2[35] + src2[36] + src2[37] + src2[38] + src2[39] + src2[40] + src2[41] + src2[42] + src2[43] + src2[44] + src2[45] + src2[46] + src2[47] + src2[48] + src2[49] + src2[50] + src2[51] + src2[52] + src2[53] + src2[54] + src2[55] + src2[56] + src2[57] + src2[58] + src2[59] + src2[60] + src2[61] + src2[62] + src2[63] + src2[64] + src2[65] + src2[66] + src2[67] + src2[68] + src2[69] + src2[70] + src2[71] + src2[72] + src2[73] + src2[74] + src2[75] + src2[76] + src2[77] + src2[78] + src2[79] + src2[80] + src2[81] + src2[82] + src2[83] + src2[84] + src2[85] + src2[86] + src2[87] + src2[88] + src2[89] + src2[90] + src2[91] + src2[92] + src2[93] + src2[94] + src2[95] + src2[96] + src2[97] + src2[98] + src2[99] + src2[100] + src2[101] + src2[102] + src2[103] + src2[104] + src2[105] + src2[106] + src2[107] + src2[108] + src2[109] + src2[110] + src2[111] + src2[112] + src2[113] + src2[114] + src2[115] + src2[116] + src2[117] + src2[118] + src2[119] + src2[120] + src2[121] + src2[122] + src2[123] + src2[124] + src2[125] + src2[126] + src2[127])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13] + src3[14] + src3[15] + src3[16] + src3[17] + src3[18] + src3[19] + src3[20] + src3[21] + src3[22] + src3[23] + src3[24] + src3[25] + src3[26] + src3[27] + src3[28] + src3[29] + src3[30] + src3[31] + src3[32] + src3[33] + src3[34] + src3[35] + src3[36] + src3[37] + src3[38] + src3[39] + src3[40] + src3[41] + src3[42] + src3[43] + src3[44] + src3[45] + src3[46] + src3[47] + src3[48] + src3[49] + src3[50] + src3[51] + src3[52] + src3[53] + src3[54] + src3[55] + src3[56] + src3[57] + src3[58] + src3[59] + src3[60] + src3[61] + src3[62] + src3[63] + src3[64] + src3[65] + src3[66] + src3[67] + src3[68] + src3[69] + src3[70] + src3[71] + src3[72] + src3[73] + src3[74] + src3[75] + src3[76] + src3[77] + src3[78] + src3[79] + src3[80] + src3[81] + src3[82] + src3[83] + src3[84] + src3[85] + src3[86] + src3[87] + src3[88] + src3[89] + src3[90] + src3[91] + src3[92] + src3[93] + src3[94] + src3[95] + src3[96] + src3[97] + src3[98] + src3[99] + src3[100] + src3[101] + src3[102] + src3[103] + src3[104] + src3[105] + src3[106] + src3[107] + src3[108] + src3[109] + src3[110] + src3[111] + src3[112] + src3[113] + src3[114] + src3[115] + src3[116] + src3[117] + src3[118] + src3[119] + src3[120] + src3[121] + src3[122] + src3[123] + src3[124] + src3[125] + src3[126] + src3[127])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13] + src4[14] + src4[15] + src4[16] + src4[17] + src4[18] + src4[19] + src4[20] + src4[21] + src4[22] + src4[23] + src4[24] + src4[25] + src4[26] + src4[27] + src4[28] + src4[29] + src4[30] + src4[31] + src4[32] + src4[33] + src4[34] + src4[35] + src4[36] + src4[37] + src4[38] + src4[39] + src4[40] + src4[41] + src4[42] + src4[43] + src4[44] + src4[45] + src4[46] + src4[47] + src4[48] + src4[49] + src4[50] + src4[51] + src4[52] + src4[53] + src4[54] + src4[55] + src4[56] + src4[57] + src4[58] + src4[59] + src4[60] + src4[61] + src4[62] + src4[63] + src4[64] + src4[65] + src4[66] + src4[67] + src4[68] + src4[69] + src4[70] + src4[71] + src4[72] + src4[73] + src4[74] + src4[75] + src4[76] + src4[77] + src4[78] + src4[79] + src4[80] + src4[81] + src4[82] + src4[83] + src4[84] + src4[85] + src4[86] + src4[87] + src4[88] + src4[89] + src4[90] + src4[91] + src4[92] + src4[93] + src4[94] + src4[95] + src4[96] + src4[97] + src4[98] + src4[99] + src4[100] + src4[101] + src4[102] + src4[103] + src4[104] + src4[105] + src4[106] + src4[107] + src4[108] + src4[109] + src4[110] + src4[111] + src4[112] + src4[113] + src4[114] + src4[115] + src4[116] + src4[117] + src4[118] + src4[119] + src4[120] + src4[121] + src4[122] + src4[123] + src4[124] + src4[125] + src4[126] + src4[127])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13] + src5[14] + src5[15] + src5[16] + src5[17] + src5[18] + src5[19] + src5[20] + src5[21] + src5[22] + src5[23] + src5[24] + src5[25] + src5[26] + src5[27] + src5[28] + src5[29] + src5[30] + src5[31] + src5[32] + src5[33] + src5[34] + src5[35] + src5[36] + src5[37] + src5[38] + src5[39] + src5[40] + src5[41] + src5[42] + src5[43] + src5[44] + src5[45] + src5[46] + src5[47] + src5[48] + src5[49] + src5[50] + src5[51] + src5[52] + src5[53] + src5[54] + src5[55] + src5[56] + src5[57] + src5[58] + src5[59] + src5[60] + src5[61] + src5[62] + src5[63] + src5[64] + src5[65] + src5[66] + src5[67] + src5[68] + src5[69] + src5[70] + src5[71] + src5[72] + src5[73] + src5[74] + src5[75] + src5[76] + src5[77] + src5[78] + src5[79] + src5[80] + src5[81] + src5[82] + src5[83] + src5[84] + src5[85] + src5[86] + src5[87] + src5[88] + src5[89] + src5[90] + src5[91] + src5[92] + src5[93] + src5[94] + src5[95] + src5[96] + src5[97] + src5[98] + src5[99] + src5[100] + src5[101] + src5[102] + src5[103] + src5[104] + src5[105] + src5[106] + src5[107] + src5[108] + src5[109] + src5[110] + src5[111] + src5[112] + src5[113] + src5[114] + src5[115] + src5[116] + src5[117] + src5[118] + src5[119] + src5[120] + src5[121] + src5[122] + src5[123] + src5[124] + src5[125] + src5[126] + src5[127])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13] + src6[14] + src6[15] + src6[16] + src6[17] + src6[18] + src6[19] + src6[20] + src6[21] + src6[22] + src6[23] + src6[24] + src6[25] + src6[26] + src6[27] + src6[28] + src6[29] + src6[30] + src6[31] + src6[32] + src6[33] + src6[34] + src6[35] + src6[36] + src6[37] + src6[38] + src6[39] + src6[40] + src6[41] + src6[42] + src6[43] + src6[44] + src6[45] + src6[46] + src6[47] + src6[48] + src6[49] + src6[50] + src6[51] + src6[52] + src6[53] + src6[54] + src6[55] + src6[56] + src6[57] + src6[58] + src6[59] + src6[60] + src6[61] + src6[62] + src6[63] + src6[64] + src6[65] + src6[66] + src6[67] + src6[68] + src6[69] + src6[70] + src6[71] + src6[72] + src6[73] + src6[74] + src6[75] + src6[76] + src6[77] + src6[78] + src6[79] + src6[80] + src6[81] + src6[82] + src6[83] + src6[84] + src6[85] + src6[86] + src6[87] + src6[88] + src6[89] + src6[90] + src6[91] + src6[92] + src6[93] + src6[94] + src6[95] + src6[96] + src6[97] + src6[98] + src6[99] + src6[100] + src6[101] + src6[102] + src6[103] + src6[104] + src6[105] + src6[106] + src6[107] + src6[108] + src6[109] + src6[110] + src6[111] + src6[112] + src6[113] + src6[114] + src6[115] + src6[116] + src6[117] + src6[118] + src6[119] + src6[120] + src6[121] + src6[122] + src6[123] + src6[124] + src6[125] + src6[126] + src6[127])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13] + src7[14] + src7[15] + src7[16] + src7[17] + src7[18] + src7[19] + src7[20] + src7[21] + src7[22] + src7[23] + src7[24] + src7[25] + src7[26] + src7[27] + src7[28] + src7[29] + src7[30] + src7[31] + src7[32] + src7[33] + src7[34] + src7[35] + src7[36] + src7[37] + src7[38] + src7[39] + src7[40] + src7[41] + src7[42] + src7[43] + src7[44] + src7[45] + src7[46] + src7[47] + src7[48] + src7[49] + src7[50] + src7[51] + src7[52] + src7[53] + src7[54] + src7[55] + src7[56] + src7[57] + src7[58] + src7[59] + src7[60] + src7[61] + src7[62] + src7[63] + src7[64] + src7[65] + src7[66] + src7[67] + src7[68] + src7[69] + src7[70] + src7[71] + src7[72] + src7[73] + src7[74] + src7[75] + src7[76] + src7[77] + src7[78] + src7[79] + src7[80] + src7[81] + src7[82] + src7[83] + src7[84] + src7[85] + src7[86] + src7[87] + src7[88] + src7[89] + src7[90] + src7[91] + src7[92] + src7[93] + src7[94] + src7[95] + src7[96] + src7[97] + src7[98] + src7[99] + src7[100] + src7[101] + src7[102] + src7[103] + src7[104] + src7[105] + src7[106] + src7[107] + src7[108] + src7[109] + src7[110] + src7[111] + src7[112] + src7[113] + src7[114] + src7[115] + src7[116] + src7[117] + src7[118] + src7[119] + src7[120] + src7[121] + src7[122] + src7[123] + src7[124] + src7[125] + src7[126] + src7[127])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13] + src8[14] + src8[15] + src8[16] + src8[17] + src8[18] + src8[19] + src8[20] + src8[21] + src8[22] + src8[23] + src8[24] + src8[25] + src8[26] + src8[27] + src8[28] + src8[29] + src8[30] + src8[31] + src8[32] + src8[33] + src8[34] + src8[35] + src8[36] + src8[37] + src8[38] + src8[39] + src8[40] + src8[41] + src8[42] + src8[43] + src8[44] + src8[45] + src8[46] + src8[47] + src8[48] + src8[49] + src8[50] + src8[51] + src8[52] + src8[53] + src8[54] + src8[55] + src8[56] + src8[57] + src8[58] + src8[59] + src8[60] + src8[61] + src8[62] + src8[63] + src8[64] + src8[65] + src8[66] + src8[67] + src8[68] + src8[69] + src8[70] + src8[71] + src8[72] + src8[73] + src8[74] + src8[75] + src8[76] + src8[77] + src8[78] + src8[79] + src8[80] + src8[81] + src8[82] + src8[83] + src8[84] + src8[85] + src8[86] + src8[87] + src8[88] + src8[89] + src8[90] + src8[91] + src8[92] + src8[93] + src8[94] + src8[95] + src8[96] + src8[97] + src8[98] + src8[99] + src8[100] + src8[101] + src8[102] + src8[103] + src8[104] + src8[105] + src8[106] + src8[107] + src8[108] + src8[109] + src8[110] + src8[111] + src8[112] + src8[113] + src8[114] + src8[115] + src8[116] + src8[117] + src8[118] + src8[119] + src8[120] + src8[121] + src8[122] + src8[123] + src8[124] + src8[125] + src8[126] + src8[127])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13] + src9[14] + src9[15] + src9[16] + src9[17] + src9[18] + src9[19] + src9[20] + src9[21] + src9[22] + src9[23] + src9[24] + src9[25] + src9[26] + src9[27] + src9[28] + src9[29] + src9[30] + src9[31] + src9[32] + src9[33] + src9[34] + src9[35] + src9[36] + src9[37] + src9[38] + src9[39] + src9[40] + src9[41] + src9[42] + src9[43] + src9[44] + src9[45] + src9[46] + src9[47] + src9[48] + src9[49] + src9[50] + src9[51] + src9[52] + src9[53] + src9[54] + src9[55] + src9[56] + src9[57] + src9[58] + src9[59] + src9[60] + src9[61] + src9[62] + src9[63] + src9[64] + src9[65] + src9[66] + src9[67] + src9[68] + src9[69] + src9[70] + src9[71] + src9[72] + src9[73] + src9[74] + src9[75] + src9[76] + src9[77] + src9[78] + src9[79] + src9[80] + src9[81] + src9[82] + src9[83] + src9[84] + src9[85] + src9[86] + src9[87] + src9[88] + src9[89] + src9[90] + src9[91] + src9[92] + src9[93] + src9[94] + src9[95] + src9[96] + src9[97] + src9[98] + src9[99] + src9[100] + src9[101] + src9[102] + src9[103] + src9[104] + src9[105] + src9[106] + src9[107] + src9[108] + src9[109] + src9[110] + src9[111] + src9[112] + src9[113] + src9[114] + src9[115] + src9[116] + src9[117] + src9[118] + src9[119] + src9[120] + src9[121] + src9[122] + src9[123] + src9[124] + src9[125] + src9[126] + src9[127])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13] + src10[14] + src10[15] + src10[16] + src10[17] + src10[18] + src10[19] + src10[20] + src10[21] + src10[22] + src10[23] + src10[24] + src10[25] + src10[26] + src10[27] + src10[28] + src10[29] + src10[30] + src10[31] + src10[32] + src10[33] + src10[34] + src10[35] + src10[36] + src10[37] + src10[38] + src10[39] + src10[40] + src10[41] + src10[42] + src10[43] + src10[44] + src10[45] + src10[46] + src10[47] + src10[48] + src10[49] + src10[50] + src10[51] + src10[52] + src10[53] + src10[54] + src10[55] + src10[56] + src10[57] + src10[58] + src10[59] + src10[60] + src10[61] + src10[62] + src10[63] + src10[64] + src10[65] + src10[66] + src10[67] + src10[68] + src10[69] + src10[70] + src10[71] + src10[72] + src10[73] + src10[74] + src10[75] + src10[76] + src10[77] + src10[78] + src10[79] + src10[80] + src10[81] + src10[82] + src10[83] + src10[84] + src10[85] + src10[86] + src10[87] + src10[88] + src10[89] + src10[90] + src10[91] + src10[92] + src10[93] + src10[94] + src10[95] + src10[96] + src10[97] + src10[98] + src10[99] + src10[100] + src10[101] + src10[102] + src10[103] + src10[104] + src10[105] + src10[106] + src10[107] + src10[108] + src10[109] + src10[110] + src10[111] + src10[112] + src10[113] + src10[114] + src10[115] + src10[116] + src10[117] + src10[118] + src10[119] + src10[120] + src10[121] + src10[122] + src10[123] + src10[124] + src10[125] + src10[126] + src10[127])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13] + src11[14] + src11[15] + src11[16] + src11[17] + src11[18] + src11[19] + src11[20] + src11[21] + src11[22] + src11[23] + src11[24] + src11[25] + src11[26] + src11[27] + src11[28] + src11[29] + src11[30] + src11[31] + src11[32] + src11[33] + src11[34] + src11[35] + src11[36] + src11[37] + src11[38] + src11[39] + src11[40] + src11[41] + src11[42] + src11[43] + src11[44] + src11[45] + src11[46] + src11[47] + src11[48] + src11[49] + src11[50] + src11[51] + src11[52] + src11[53] + src11[54] + src11[55] + src11[56] + src11[57] + src11[58] + src11[59] + src11[60] + src11[61] + src11[62] + src11[63] + src11[64] + src11[65] + src11[66] + src11[67] + src11[68] + src11[69] + src11[70] + src11[71] + src11[72] + src11[73] + src11[74] + src11[75] + src11[76] + src11[77] + src11[78] + src11[79] + src11[80] + src11[81] + src11[82] + src11[83] + src11[84] + src11[85] + src11[86] + src11[87] + src11[88] + src11[89] + src11[90] + src11[91] + src11[92] + src11[93] + src11[94] + src11[95] + src11[96] + src11[97] + src11[98] + src11[99] + src11[100] + src11[101] + src11[102] + src11[103] + src11[104] + src11[105] + src11[106] + src11[107] + src11[108] + src11[109] + src11[110] + src11[111] + src11[112] + src11[113] + src11[114] + src11[115] + src11[116] + src11[117] + src11[118] + src11[119] + src11[120] + src11[121] + src11[122] + src11[123] + src11[124] + src11[125] + src11[126] + src11[127])<<11);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'h0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'h2482e11dcd1d4c8e512c70fd120401ae1501d5f611bc58f7b1b40474ed60d33dac9f0a9c9ecde4667788788056de7bfc128565634c49309f7e037e83ead89fc13b906679156d33b401d46c19fe9d9b92749534d7fa0b5c35fe5426bb00804fcc44e7aabb119a88099b1a37c818f09421bbf2e3f08904846333aa3c94f14bc0b28caf44f5ff4306690d853e976e068bb60d10bc3883e9ee3c346d6b29df31a49e1e1325e0d3433ef8c431e516b4f05b721b8b7b97df698296fe0f6ed0ed7b8aa2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'ha3906ddb8999c2a88ae1651286e34a585cac2799b243a4d46183eec7c0c9109271c6bcc3a19f1d6cbc8cb7e8ca55b5e409a30e835d0021539fe721fbd9ad58c90473f61f3a8d7321f701f21ece6066b8f228e7d790711d9d7afe1e94d52de4e82538d2c6b0c5134476930d976d8e62e5feca9d684f182cdd49f919fb6b7563f68e01a75218b6c49fa54241cbdf4f67e93443e179d6502f978244c36effeb749684fc0da42c0e8f7f5892ca7024f10124f7e166be00bb9843f236f2e3e3a56103;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'h7e592afd317131426a65f7f045246869dc2db88008e70df64e771b6865f10c962cc2bb8fb681426b082458fb79929b0802d18caf5f9351a06066bf22a699931203e30d932ce62841375ed41898040d853cd9e71ce5f654b6e81056a17386a0451cd86698bf5e6653f5c925b6f7e43ec4b9ac4b47380d0aa55b4b438941c900e73d37410e10ba730f1f6201e58415403e4b13c6eb66422cc118d4154e43746f31407635f557b76cea817151475f4f7ab2679aeff82ff96a6329c5bdcfb38d600f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'hdb20009bb8c9a4a598ec96e0a08f8e9d4a61d3cc7275a7a662078a9e9a6d25d9baa1d4aa77cc5d5689ec2fb621a74a4750b26040a51ca816d72e180b194a98067471725d703789d7f13a098c3ad27c3fe73e1a68625de23ea3e4f77f9c56cb7eb168d2b2fe41cac242b8245218dbc6d064d3b12a36f91d7fabddea3db01a80c79a364f6deda823b7e519e49ff054dcb16a7740febd132cfd7554af088c144fa54237bebae0c73e5c8068cc851c413bb3f91664b7defb36f8729c911f9e67a7cb;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'h6f573e1903a1ea0d284aed77845bd7f04d96b5cdadbc3418c32c076d45df9252d2906e85c6a3e58dca4ecfafb5ab82ccf252232de37515b381dc9e84c3b9c25a522842482c9db01beefeae4d5ed3d7a195fda5123ff7e467dacd3c8fcebb6f22009676cbb8b7c7287fa34b33c1148b82cc7c2f2c7c8d5ff879e6730e4bb30272f0e86e294b4ed10aceb27bb5baf7b066bf5b8c83d422245b79cb655f517dbd51867308df163035e95ea350506b93228e1fbeef46f50fadd4c458d2df135a3e58;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'h519eb4dd611b33c377c9e8f799304e5eae2f76e4d6bee36e9b6cf5eb3e1dddc66d38e31fbc20a319b5215003d0dd2c11c0de253e605581018b7ae04120c9447224df56c06c8f1cf7f93b8a92069e86364fe789ba1fba5f0a29e74be83eb5b964d57abec0274ca3cc7bdd3df803d8702110abe5c14aeb7a8b7bd8831e298d2c9b4ab66a9700b88d378028d8e58957f6351837af0aa6d18072fdf6082158f885ed6b42162325fddab36feac4726873cf38b1fc2ecd952a9bab43bd95c41936905a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'hde0c2c45cf58a576b604b243c3e974db2daaffc704ca87d9a36cd8546879c71645ba518b3b565554fb03d5151427683102e3d1108b83777d10fb59c8bf57ab949a5259d0d6f5f277b67f1de450c9dacc4e394678a3e02b669c4ac1d0bfb6d4b0045f06525f9ab0bf18674abba7aecd9b2dfbd73f5c48ae1d0896d1076ed2849532462f631dd3e12d55b14e11a5f38d59d336b3b1ebf31dc1e56e67b817247740575b45a2d704b7d10a323bc9c829105591ca3f8cdd373aeba2d6ece50314df4c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'ha12dfc0000d953e4a9638b6954ff408ea910345be7ab340dc27075c710f4d5492a2b961eed019beacbc236109986d9eb3f8c6f0d77ed8365f183cbf5f129ca3fbed081d2d88645763bb046361c19a9501a7eda4533dba29e4dbfa90ca922063c92d6943d869d5dcf24f830e9fec7d18d0e6949740547696b9e280f28953dab4525e1a81400b5949205d01990ab2d8047d28828bbd34df4151a3496b110596982de42cf045204b8e1d4b5a493b0c3309325dd7704b23fa69a51c82bbc17a5fd00;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'h23e49e93d4869aec20908697abd5b8ca4eab5ae395bf045addfa13ac4a92cb75bb4642ec1308cbcb41ff9d5c95bef3c77b536e0e204ee1b71e4eac4b1a7b395f19ca263907b854949c5dbb66a845305f1a1ab107451690d22a78f08acaea4263df88a84610abb8aef4375a69541f5df327bae6b66545ed9534aa10adaecc9bbfda04998a42b2fb091fdf02872e1d956314e124085004d714ad174829b16906dec29ddd6b90a977ff154000dfd1ddd2dd99aab6979340937b6d496d59cf2fc585;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'hd9ffe887fd9bae02506ca3ca30d31e3c43592a5d9019f04bef8d0315553b0a1027e991cee1370f18e25f2e48c228702c73c3cae708a5d7077fe198e2a1f2e1aac057ac063a1a7a18a8254cc7b6b4b831d23eab0d51702ce016c0474e5ab286b6c96ba4a7a56a8bad0bef9f0d726aed7cadcb2c797e29b4b7dce19fc382b32b77163ed4d81197bd05de2920c7652f65b6b418434f4a1e8a57e7b73278c2fc7da65f55acc9fc29c503a2c017d210d8ea756304c7845a23f168002d8f4107fe11;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'h6c719bbd020b60425d8fafd1877bfdc82d7a50dbe2bd88e39d1d9a9e93d2b26f09325bd09e77a5a62b18a1da3b2647b1d2fc413aab47a1fcb4fbd9ce6ff68f3928c84401c0b0b7b46c902eff8453a7e4517347fe38a3e3c91c2f65cd25232ba37be3d24f08ea6cb68a87f5c9f142767aef6e69f33d326f17175dfe7842c1506f60447deb4c9e528bb9eb98f2ff9c9030521f748855d71b3228e0db26a331b1178abde95cf70e4cf4a867ff7c8b4f25f6e327c59cd8a0d908adaa42243647fd3b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'h4de7fa271d6ae8e9e99f1c5ef548544ca235a8393d0dd4a8bafe57dcf1742cbe762ba19f70f0e009bb82795f5f1038973b9de9adf1cd8e5f9b3473134dbebe6b23a0a51b0ce7d687cc2105a6adea7e4cb003c1dcc9c72caa76792f6fa98e62e1cbb6cdcb39bd87b37d02145d130025913ad58f3b9189eb8692b6a6d99944029089342b2b2b0ac49557cceae1a5e29b4f65bdb0bd7900706ddc18ec776f815ae95e47fb82118b7d3c8fc4252e7a69abd467fa8103d02a4f2c342ec9ec20baf550;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'hea16071bbcffd8924c8a3c4f96ca3160d47e39f8d0277284fd3c8bcae17b742ccae6ba20740b30c88fa077c5da63a7d780064216eb05bfe08fb22f2a51fe444ac6cbcbea869bfb7ac2156146bd74e7772620c2a599666f198009736890ff3cb0477fbdb9b653ad988ba08cec4c18d886dc422dbf9b841db2b3902a9ae6f6e07fd9dce0490b650dda7c0f9b699c9878d662c9b3cae44033034feff69a2da9edd0123b4261660461fbba369f0b9197d3aacfa8690507c910c50295d96b9ed2f0ba;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'h223eb9d02e419cf2bf946162ebfbae7fe84eb8f8f9f69316d0252f37104877207360c6926d829012788c3de395bf1915be0916376273b0ea35a013f3789d1a8076df7661235ff72247e8635368a797a8aa377479f0fff5045232747dad8f02395185d7720c8cb41816666a9618b3eccc30e264833e2f28aa21da432505646640c587e45a2cfe16ee0a011139d7b8b123162d0fe01f333afd19dc36a0c7bad79e70fd18e02d27fc847d8c73192421b9f6e6dcef674f1d20d9ddcd75c36492fc9d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'h307abc6588d6b3806051666f0193eb9b80f1e99507ba67f567eea4d8e04e9b36f384304335c9824740da0d22a715f5d127c269db86a787e7c7a15dd0b692533556623eb384a93d5ea345d056ae838897963d9ca81c93852b53dfcf78a81197df43be91c31d097f4c37964bd5f260e35e2ef44b298e5ca787ad5e67454c5a406baa5d8d048f9bd29e55f9acd549392e5abaa1c3c5ff567a9706496029b7584897c05d37e6d913c7b27fcf35738d04918bfe3dd973fa59cc3d5c72d543106a99c0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'h8e17e9bf9a026bab3f99e5b3e3021bf3be963dfc3060944737fb9372f633fba3406397dcf5856d34ee8dea84b0ccc6ac6b690893bf62563aff7735d7bdc49b11ff708bfb049d95ee4138cd931f365989b88b3f40d9493817c878f93be631793a1719db3fcedaed711db073ed350dffae767df827e9d57d6dd7b4d2c80fa85919b2847c173620f657aa868026a603ad8cf4811a23adde2f43861994e994be2f1babc1f9b513fc00309e3510c37f4e794c6293c3bc9c31ad0ab4ac0bed865e9a29;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'h37c26257e6426e8898f27d9d3b7b71c73f895f9c4ec998f5aa68f0c651a99fef264b3bea5b8e0e9b4eff0252644a1a70153b4d0f42127523739861a514c0652236b8c1afed72b010aa6baac4e611b5af1cab40618f9cc7614000ae8b39547bb8684163f79003dec59cf998f3ae3b1a07c8348274ad769ccb4f9c62d8701604eeb15c5f8292ac22b2c3bbf5ccaf89561565a0beb4df011441252575672170e86b4177e358b6782665e0da90c44034e12d076cb71d17f6b8a535d4f1c6ad7915fb;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'h5f6570218e8de26a22a54b20cb1bb1655f13268790ef75dc3c4c38b82245bc09f5f4bad26f3c31ba96dd1350b57fd5992b7ec1dda46f1590236019f44a1446a9a8e886a38fa640879c6db083470f7d9d782dcab23ecb517f773ab5b72eca0388b1112e9bdc371d035890a786c5788c9720ce127267fa141b9163ec34ece5b2a71fccb91728315c00caed7648c88398586eefac9cb3f94a047e2274ee60cafda06e8f3714f2092c7eee1901a39767dc5211813aea487ef305ee64a7904d8b4e52;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'ha230a046dc166c7ab03957ff0860f7419b92ca6581b2d1aba6f00272514563535a43df0f4cfe77846fa3dc9aefa7beb68d4cadcbe7a68e47483bfcc62927bf73600d5dd1905badf8e940b6299c89f23161b808c00941915b9df46c58dbfdad5514740102af9af1a381f6ebc8b3bb035ade8bfdcb7ce9234e2e145323372073d5d7d143f8d2fbba15ff5db07b40705bc3042b0dc9e7eb94f04498ff42b594e41046f6234e9305a87ec2d9ed19a81fa27f2d52ab88c4739352c4b15eb68904736a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'h85113ae3103367ca45df75ac90e337f62c80b0c8ca37b6899b9bbdd659f7b064aef54d80161dc64e3e31ed944130a457e5ae478190e00901a0f73d69dbaa03fafd55504c8e7e9d61f8f3e1c37cf3f5f9e1c5c032e0531d7d4a507b7b41e7852c12cb23e191e88db733d27a53febb31d2a3c7604fced433562de33f73ecc695af6bf0691a5d87bb5567b09ac53bd3d4d4d6d80666ffe8c8b3c9faee3c253e74bbe43cc110edc4ffcacba157b24d5c4613452d87ccb5f0cfa9d9d0efeb64954fe3;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'h2188b579ff566fd1e90e6ebbe1b7c1fff637ab017fe28bd99ae34d5ca9cb0e31285120a7fd967153e6e1a4cd3169265fbc704272e067b04709b2c4df1dc0b839c5fd36e0584c3fd7603946af5e1c1867beec0d725647d4fd87501e50af1ced4bc57ff2b33634c0179924210e727db81feaa4fbf88a2cc3c7a543b5f6401ef180cd854e11f2e38189fafef1c01b62b134c48673a9656957ab37eb021eb1009dc94645eb3e58d9ad1deb000de4373260b29f8c1c95bfa4e62548bf8b1b3df920c4;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'hde3b9c86d519853edce7e40065a7690c609f37ae42df6bd1f0759f3ec139611dfc5e48e1e5a59251d270f25fbe6d1c1a53d8ea485a07a665199ad86762138f4e2a769c318caf0b990b786231e2c6cf6855c0558e9e07cd4653324aafd8ea8fde584069c4907c2392f6e74d42d832c38f05d24383def2259a6e8de6e839e063f2bc272f2686b07ffdd288a141597bfc9bd6c86050556398d9dcbd01f473f7f1551d1c7662436a6b46554e8f9087f3c97ceb923ecac78efaa73e3b1575b931ef5e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'h3beec458f009d7e36b77339ddf7002216a987bcb2f3a9968cf14506eb466f43487ed7c80375d5a4dccd64a5dbac12653de20fee460089dd233aa956b616c3ab19710a8dba6e4c33f2080a9c7c6efb5b82b42ae6c72617c0029e0ebb7cc6ea24412aa1f2536a72f3511cd1a967543cd77ec8e4b89c5b3e4abf764c925c3639f154db32cd0a1d314f136ade76c8a282a9c0f4c3bc8117189385e614c2acefc0378917d019a1cbfc93b5f679dc50dddae372c3210987d88e076857471dcd36b2883;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'h17a06c8442be4d421c1bd24fd5175dd128b67a8fe759ec29a9da90001f1952850e8b10bd049b6435596ed18623418b26f906e5dbea2eb21a3582dda56a09b5f8d7e7d41c01fc6efd38383a9aec52c56b4c10c8afc6b274bfe64b5bddc183f7344c9a49bcec85910e695074ae929432a9a37d615a74563e3b5ed854836dd849f4db7292208996d46a31e3a619db405c1c058b6ea5766dcd314b3f46e2059ba51a675196da8916c2bde341cb88c97d0f3b1cbffc46583aba803fd64986c7994fd;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'h7f78086f1e238b3786d515487b81092207c6c7a556d6ca00a361941a2d38627d0e75a4f2fbdf65600b95245c13d3e6ac5940294729b940bbd69752d0aa3955ec702214fe0249892f8bb16148b4ff9135d24683d6ad0a543f1dfa4abd7de42b47733915cbd833809ac3af135ddc395271f218723e13e859ab19fab72cbc78bec58e1c447cf3584035034ea50b2d75c70e9b7cb1d057db367984b076c354e9c6a0f7abb0d7fb2fa49f832feace98c31afe0305a521522e308e6b5e9ccf3e0d8a89;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'hb9d8e52cc1b0713072e10b7b078dacfb2be4fb3e4255cf359ffd83e7cc606f36776254b08af2b8adc39dcaa7b0a7d58838802fe21fbd8ea259057b057a0ce8e57c8f06f5932f0d5f5de595709c33f4b339fa493338cf229923ad0faf174fafc63b073a436feee2c58adc4d1801a5c422b6881699ad32f30dc22b06b53a45f7a3b30ec5c3d3a665a14d9a66ac9fbb34a8538eafb26d26754a30d8f9cebeafdd8e70fec1a95b0cb7e2c9afea8308adfcb557a068a925bb55e3a93a9a5a9b7c2897;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'h5afdbd6151c3fa32a51bfd1e2fc732ecfa3404a5ba295ce1fbe797efc932919cf58031513763a85ade406479205b77f0c282ed6228b8aec8c18bf7a42c7b1486db7a3de4028035f64a0a717695cc56bec3fd7daa58c4ecb2ce8619a84add4af7f8b51427c8618f54eaf534e8bd54a272e2af5250b2d7d0237a1231f7ed77ba455bd5a1e351a36e1f04328f10b5b2c699b67c556b12beb306f6584ee7491efedc5fd9d8c79d8775100ecb6455f064185787d80591326d9f5d8db18d4046e066ec;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'h835e552edb18034cf86bc479bf7c05aa119b83a8d46c268f765eb39f22dd02f9f00dee9081aba6c0dccc4c8c7e439161f227a44ee9acff74ec9c256f6dfb612dfcb1791394357972926f1d02ab62bd562184a48ebb6cc6b30fc5f962eafe6432ac45c2053cc9fb6d688bd024ff956c1b519383806471e38e939c4218ca2046aaeee94cef4194e162aabfa0dcff12a5d385873da3c5dda19feaff83f3c4372b1161383540ee3ec1ba30207800bdef647fcb783eaba6f761def47cfa769b150b66;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'h35a5cc8fe694f0a17aaf83d6fc85e7d89cf118174afb709f2fed26626a220b90d87534164bd2cc9a5fc474b4382ff6d7d184a6070d1afd66adcdbfecc29aa178302f694df6b6c2c1ce0226fc9d9f4feb8197adc9dbc628138c04a32ef7bdae8f2896100f65b17c96054121a9bdd240d856fa7c47679d959308ea5f7bf518cf4a7ccd84b8d159b1d183af35e27306a4967fea4baf458e5dd275d635913982e6d28aea1e8d7b2510f693b2c41bd9145509c5839cb3823cc6fc544d27354dbe5556;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'h84890cd2916120dca035e6f76b5b7b0c473bde62c68e9c1909515b14c8c407c70e63771d1750b088a46867f826b22c0d411181ffadb388d3592e244f37b1baaa5e39da9083ec88a67c153dfbcfef3ed72e617e2348f8505683c75f6427daacd427ef8fa0fc4bd64f2a6b6e1a7aca0afe117cae33208b5cffa8f2627bd2fbfce9ae70b44b69469e7c70d1b77ee95c2be796f7c695113b3b67d14c6e2f9e6c529eda15c421e638e2cdb406260315205a5c8f53cbc8e9d0f9a7833788dfb88f6b93;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'h7fa2feafdc31ce1fc78002b89ac19bfa403fe538a0254af85467f359152ec32184cfda1da6bd828495885f95dba5a73257cb8904ee52f6d2fb076671e9da2271aac2b83a5446469b22c2ec3cb65f33b94da9e0a015756e37cac3138ecf763607cca2233a661d626b18540776ad56e585c06b894a93b27c1b6542617e32c1333cb688af6408f2d963dc2ed4f62ccc1b0b2f82f337f836ef462e6abd537f9d79b94778254aff372e7ab2bbcfc37d78a266df4e6df3dc957569c913321be651593f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'haf7b26bb76690dc0ba11a6ebebd22276a0b79f01d3f35f41dc14afb91d2a206edb2c445f42c1f3486b29234d4a52b230d5f5a782022331804593215b3d82033999bb7547153601eb82cfdca5442a9b78ba977748a74b2cbea9532abfa8b6d36eee108b1deb7376d7e6876ce8fbd173d282b12ce2d08f55d4ef15f6f9a0c91a312fa1626f2e2ab0b271b620d9b056cc34a9f7b0e454cafb9a8bbb456a0046819f938931c1de92f3c0971d3663c2b07d32afe93b123408111f587fff2ced057c6e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'h599020ab59720321441c39b5ff06be9b61e9394ea6530fe979f547a06243cf5830e79cffca8c33d9ad9c50fdfce30779cdd9d918b8d13877e3eb8069c36f9f83fc945af5c791fc44a79e34ca3386a76b6acd2aaeb8a2b4f511148dc64e75cd6d1f0cd9ea1b78a16d12684a9c82503e59338e44ff35d2fe1c537b71435f7a2b52c5c58885841e9d1f1dbec703fb4c06c59c1d1129dbd00dd935459113cf7d69aa76de429ee95338223fb06ea3ab260d45ca0b50771e0a794b5dc14fe984f9016d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'hbd6d447c57972bfe005a29cdf019fe09f55d15558a5bbb2fb4c0b0d60fe810f5fa7f6f02a34163ee75a875c67112ce1904e16366a2b9f66be487b9231d4e6f9cc2912425bd75f4cd8ae0073de0f6768803dea15ef088022a4ab86dcd61b4783353e0095b2087bdc254241fe7f3d2976342520055779c598f63eb8ccb21dd7a21547b665f3d7264a6a85e32898e556a2a7899a7a757867061629ecbadc62e40ec6aa67047a8e6641bd09002e67bbbc8453a4fd9702ae540c1ec80d00217a76e2f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'h853e698517dd89e1c40bab7d6e2c424a2af2937f9f5b813f16a707f2b63e463c7139bca598455ff237d6a7431cb9b871d5d127a9a44f7111025d883b4224620f6ece16f2fd96940461ae6c0fb8f9c0d61c7b90354ece21cd85505000693ee57ee38798f5e17bd20ba69b96185ba1c93ae9c8de4a41ea5611ce247d1d38ef0d4aeedbf197ac974f9ee6fade8553b87304b63c0252bce415851a55aa979ed90dadcc2d7acab4fef65ec11deaa309e28da886e13af1f425632e41da82d8027e7064;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'hea1100a6196c306408a441102c16222a52369f911a27baa18aad8f387eaf57408f20ef87d7563d30430c3f62610b107fec21014540a5e6764ec66f123c511f2f01da2214e5533794d5cd0522dd59a4589efbb3ebc1ce0255ccf7774c51e098d44521ffdb8052e1217ccbf3c4c0fb5e7c610fff6d54b1c20e8ac183a9bf1ab5b299a27f5d74d582c35d7bc9a8025438623a409ef42c02cc3d0fba657e083784e87a397fb159e8018f7801fbd84615318d842ba76f7134e6bd4cef44449a73f0c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'haf496341daa6f9faadb79141224f4ea4e5db349a1bb39af73826613f5252414b5c5a9d47d0ad4f6027d36107805c64c4bab208239554f51ec49ee9ec0ede3c5de8eb7a10001599c8290eda7eaf62dc1063ab3bfcb95a66d7780d174d9be6b3731137dd7f154bd560eceb97deca2d5b3d5bd6300580f3e7c271d54ac65c1ee18e6d5bd845e12812084bef847fa82a330c644a27cd171cc2a8c90effaf0637c7a3faa83f0ff6a6010572baa2f482bd805c86266449d8ad78deb44cba879314c492;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'hc31ca76f8f63d929caba06d0307f510b40377eb42932afb90b20bbb4e495fed0092f5ac4bc0d3518930df0cdcbcf00b3d591bfb0164d933c23aa51fe8a29aa195adcc625437e48e0fb7dfef2228150b641aafa2d57d41c3bb2168f205304c023bef0da6d24bff7a5fc6726ceae38ad138888edff3763411fb4358ba842bfc211ab0a293fc5c8e689500876cf58f92e1c2ea05d3dca755843d90215159ee5c4c4bb8711e2dea9e462a38e741cac17687f4f620278060bebf37cf13d9d6c58f200;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'ha014c5e77eaa0e0d59b388c74fa0d641497f445e3878d530428b79ff652ffd07cd728420c1fc1a5797b7f183bbaf614282ba45b5862e7e024810c50ba04347defc27d9b45ba5ecc983802b4f96163119577db874ee7cd35fbf8f10e577f9f6ebc7c6d7336503fe9463f4d452e5e3d6b285ed255e74fa274ece91bcf9efc1d452566d5fc8587909ac59f123e6584d82c857183948b3cd57924727d12d5bc113260eeb47f7607984a018039e48223c6c7eb7e33e28f362c7054590aa97e6456b8;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'h7501757220a4201d86d20aa837909340040415873b1f85b633a368b5de6ccb182ecc29afc2168736e0825584388c1cbf1ee74e6842cad9f5764e729d859bfe482f7fa82931051f8754be2f58e190451cadf1afa7690d2fdb5c446a6c54f42ea94184ac8743d0aa58d2d73c1893ab695af711a32140d987c9b2086a09fcceb9d7f92d3bf6c41334000bd3f65f61508e8ce0b77ff0db46aff6f7759bbb8c10701ef02043a55f3d5a74701a0db848174d87c6d2df35a302356bb05c0427f2667d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'h2bafb28feab1da9962543f8ebea057daede7da9d11bf50a16006446fca1f11596ced5a66c2fa9f72634426acc5f4276235868f700bb4221fc70eaccb15e292cc73a4f3d0dbeffd3e90738e9e7fe517977c849460b78b2f0adef886b8768bdfa6065f0501cf086c6125574877cfdb12665c0c948151faf39308702355acd13a1897d27e3e7ecd022446b2ac582a027a3680314dc933719cf72f8078be2706c0d190b68e34b464498c06443f0d5d358d94edab7903a70063f83809117250f5cdb8;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'hdf96e603bf6ad644d22b5302a271973e23d73fb7fa8f22e2c9bd499e2f88e392080936ed905b64ce7aa0b5e206113388da0484e16e21d00ad24dddd8ff29cc7047a116f2c7fafe3ab323f3da8f55f5e23e2127cc6bda1e566f76e801fd57516727ce62f4c6844ce228ebbb11a1f71f31337b410927189de1865a10e53dec5f03817a3faa1312ddda24c826ade3f6b248115fa07dc891c63c0bfea0ff88269f04be2182258d3fe9933788ae214a67889146e09c54c2eaeb404eb412945cae57f5;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'he6caa15f83af116c163649804a86c6ad3e9e472e4fa363147ce0ee8071c6a863f45182ed662e34c9e9bab4054522b37281577e2ca32f1dc21b3cf88ba41c9688768dd54adbb4fbe3f896c142e27477acf6435413455b6dd9179ef920825d14a9551272709bc0235cfda2f486a08698ddc0a5a06910b8a184b7740fd90104da19b74881e6615715b7757533b955b2346c120b5d00fda783473836004d021d174a47a391c6fa96b8d2ef725538688ad5c4f6b0b28e58f250026f5812d7cb188e59;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'h57ba6eb2026903ecb2d8fd40c6243eee57f96b040f1f7b083cd118bfce2a2adfabc6e0dd949dc4fb17383afae1d1706b67e16c913a5b73ab7ebc84b8d08f292e688cf493528480cd1c5087e792d130fd4c7f8476a18039599b3f90ae49d452ec1ca700ae2f8f832b829468d7f9543024cc95404a16e07d5b8d8fa980b76f4555f29a540df3d4274365a69c7cfeb0f81d631a8f0d569d4a1430c9891d0db41f4b969164a9494d26ae7096a22067a0d2369e06ec0f54bb7353b0cb609bbd32fc19;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'h5e98599d28958125a164b3d4762ccded39c30b6cc2506d7a281c71c8418f4b6213171d4f89ee98e576ea4937ad98f7feb625649cbbf52db753deaaeb049d022b33520e4116d9dc2c7e1baa98319af6170a37a957d8ae206e66643c1490357feecca7a21ef8b2fd7f9db38ccc001d0411e241c3f8939d3fe218a9e85303853d24b9815d52f3eab758e8126985b986beedfe62ec9a854f27d5c0281907ea388c42cee657e01d714cf27a671ce589ec8b1d35d7aabdc7a5087cb3b840893052a3ad;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'ha4cb406dbd48df3c7c2798e6b789090d2f56c3b1e6ac15b4b7103c59126e9a77a4a28b35809ae94d3164b3e6c7be0368da052fa6e196366176a1506a312d461e706ffad99c5527b3bf5e7c8de31321755cc214016e04b32f0e043c8da4d89cca6b9cd45ed7b6309e607b245ae7609c49dac92cb4a00ce8c3735e2c5675c29ce42e713cdf1a3f0643e45b87b47cb3bf294e2d4fe30260a4d673e668dbdede5a4dff315289d605b5fcc94fff8a96a9b9cf625851d65c4a81a9876be99fa78072c4;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'h95c949ec7d87c9ec8d22331b8fe64ea0e2fe9e5aa80d04785621f83e92e3b2413625b75e5e7ed798263505b1a26d4c70fae2d72e85717321089dfcd3d6553250c03cd6f675f5af68a5efdd9599e605adeb819814fb740b8bf3e55b6e0f340b6e93dff52c2e4842f73260e310a817033fb9d9bab47bb7584b5adaf762a51062e528a371f0cf047d7c53726f816c2e72db5be7729dcb67b505d09cea79843f378d9452155ec1ab26363f9db16e603aa904024a0a6ac370d0056c8023063b5b8787;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'h522850b9929054ab0cbe6be76cb3fee310d31fe7c729670bbed535439c2f06727c4a68e22e0d785266895b2825ef79f549a6a0b6af4ca7fa2fa0bb479f747d00202180ab716c851614203d553833d8ff0684fa45132a9af7cf72163a19199f4f519004b592056561b57e6cbc2ec3e1b212dcce44863d2316628d9d626d10c58f6aa57ebe51bb339a9bfb82106ded384ff343fc930d083763261af1889b6731e85a166bf09f2e2958d0c40b280b9c4c15fb6d624f1c90e5ad171defce5d00bb9b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'h772cf5686100fa5cfad47a39167d5f630cca76a1bce73b7f0edeca47cbea86161f71a54df9593634b6875397cb3d7c42409a53c798a70f4a993733d26c8b72eb4815961ac27d2fdc33afba2eccb01c8cfd7a7a1e9c4f1d2784dd6620e4c0588de9783969471150215f18336775d8752308904c743a79a0a492504f88b2cf9689f0c8f9ff97e83c155693c0d1f96bd5effd16dead2060f46b0df68577a71c9b9ea894fd6b02631260ca62b3068979beb49662ea470b8c30d7c5db4bc19c7776dd;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'hfa545aaca4e649c47eab67473e67df93d4288e009f395725157bd0f5226ca88799a020853a923aa986e46cd2334a1c4ff891468dd0ec015a3e96ba4a90b6c50821c38667be108844d23342a54da306aa2dc1866e0803cdfd074908e65bad041c1baf5c3887e2f312a9190e67c1e3d842a09c43eb3429aedf91eff7390f6b6bb357b1f92cc1e490059758c68f53497a174fc8ac5f9ded2c631ca272618280b27e899c18e09b6b5c5afbda60d8e96f3fc04550c6bf7290afc8bdc23bfbce1f9fc1;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'hec502f1ab847aabda99c8dc4dbcdc1d245f2159054e74f85b96cd018746c7c2896351ebad50e023cf234e836e82aecc0756fe60c96ad888fef80df2f13028fd4e05758a37a99795044cd0ec573fab76efa40f629a9c75866d40c081fae1bf1dc7cb9200e8705883b26a3f6f92eba06742876de2cdcc297b050cc82bc43732f9ff4a1ca222a4bfc38e2dceccfb0204b64425aa1737215951842f2a0f67bfca17cd51070951bf2bbe13202ea667f425886ae4d9ef9c93fd1151a74c98b0280efa2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'hcea71df46045ac0eab8b3ee01eaf46ae24507dc01b765cf5c5344a24a35f717ef21b4fd453c4f33e40f8978a32a02eb52e3cbe70fb162047883282ad5591ab98fa4d38a73cccd3932956faab62a59a0c6e0b0ff5690935b2e6a5c650a32cb39c9a8d3486c7a1dafa5830bdde02df6c45674fd0a57fdcceba5c2db0af61abbe518e07b5488b0677c78d192f785e21f1034b86ab58141bd0b197f30a0f7e3d33162351b5f5ab414f467b06c8731b06d00f1a420e88439bee0efab0f5817966d311;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'hb0f97ca4c3c9edfa85b470859758c8b6a1a5072d392559a06fdced9c2935fe18481c1e2d07a9ad21cfa953a9197d1fd2fe8800dc185a1e880885f1c18c7229f908a1d541ccc63c5bc959f91ddeedd5194b0912bcb5dbee372c5edfd2646117308237fd70f524662b13569be052117a3119eac451744604ab5a1c1679f42cbe9cd7f82dc989b908a0dd7939709e204d5a5606c2228afe84ed6bb0d776a77374d3736b97c013ad56df83471684590a4cf8cde2d811e32ac2274298e74fea221f90;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'h43b880b38e549f73552de7dbef85cf6822300161a57a1b254d1e47c4f2d6d215aca05b8606d675214cac15aa3de8d7f942549ac429fb991f9e568b5320bbb5e92459d0519e8279e789943d3b8f08653a598f2527709149621fcc9575d08ef5d722ab3169fee4f025cb2f68041af40ade5b6d419df65dc2c30a0a621dee8b44ea41e23e526bf5a739a6fa5d27bb3c27638b74882ff30711aeb9c638e93d0a8a709bfdea2bb6eb18ef4d43a28693eb11ea83f399f5733c2f9d7e813ba4e3d79c3;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'h815c174958152fd026f6ce7bf3999f7355ccd3b89c55590c5126b09b9613c665d666fe3502397165d87fe8b85064d943a3c233d90331c287920cc032fac1312ee9536f330c24f9a2e1fdc3cc2adcf1cd4881ffd13f827c04d86b5259cae61e65c9b6a7ec812b9236afe47e0824aa8f064fe1762cf6bb9bc5b7d268824dbb412fd4db8914c44059e4f6dc521817bb1b425d15bcb17a80fba13b63d2eab9a19511365d49f9d6443c164692ba01e17c8e913c27053f75f566f4375da3b7b5c2ebfd;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'hdb0661ce29fd69d3fac2546313163b1b24eafbadb567f2491d5a869e8bd71da370c793b642846da2fc5aa0bf6dc11facb23d948ba0fd0e57cbcdf7f0dc93fba1a2d1f755dd75d29b822b4f948261620e87d6de0bf0eaa0efa1960aa0bd0993a333613ad2c2e064180854fd08ee3a2d443f5c99a331e09888dd82bcce10049d0219a5e01cc62d81d6aaa45f0f108fd899a14f4fe80831bf895a149a89355312eacce9a667184ccf73e6731ed3c0c7c785bc4d0d881153cfcd76d7705556c94fd1;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'h2d2fb42644481c0bfbae515d90b9a60fe0993a00e7106adc5cde4dc45996a93c0685ffc319329cd840deffc196d80f8191416762cefe813595f72b84bf777eba410cd152efa3a1d868ec25c14ac5a39c933a79fc32323278cb8d2a65c9939452944c900bc53e281e69976747a00ed7da854b19a89552aedf97edc56ef919aa7c35b0a3dc8368761a9792cfd1c971e1a388e51552b0f58f07b8be1ecef6f5bb4e78f9c7a69e5bb995f378eaff6ee8082263f063946302dccc02fd8ff7b870c327;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'hdaa37d2babb9171aa2486a8e69dee1ccccebf1b493f17e67d95972c3c85736e9602a6ab301355f215fde2340e7dcf4f41236c2b58980f556d86225951fc59906738b530e06bdaa1368d879bd84cfa740736d8908ba537faae5c51f89c5799f9e8f1211aad497a8b0862d1b21e6cf1f13c40a3a623dace7aa958641bc9b7beffd958a58759e239e22d044cbe2f941848ec129ea76d85aad5dde0fb53efd51dddf38859b300febdef8d4d5bed7935a56334cac53004d884d7f93d938148e28ccdb;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'h3b05fd7460962aab36bfe93562aaf0e0053bc2f565fb086d83e073fabf433c66deb08b701738c7efc8275e440d36060902621564f9de940e6ef2c7cc71b9c7f20df46830e1d9ea2d1b1f528384ea77350c3a101bf06b172b257c11fd6e2e0b31c9d4e84d0933b24a7186980a0f534d3f511ab2a41ddb6f36c6541ed751d91abe6f7af63e6501c9554d7da8d3d6b07d9912c1909da861c425dfb9c9f3e17a315aec3f5b51a85eb04de179f4cf8ab35514da6f679c9c627dd0f414d32c5aec77e8;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'h9f51406b95624e3d2db0fab739852f6d55de81cd1ae0524a1b3072bdf8669c684b281b976356c1413d145632fc0be5f57be93bc64067059fb8fc34fd9c47430f15fef3556797ffcc724670e8eeb60d169c81d75b066c621c05a703a585aa4d4c6214ffd00895b3df9608f7271b6e31034ecbefbc3970df439bf30323c54b0c083b4bece37267349d0fefb406805b591b7db5feb4310d6231ec1fc620463625250369a9f752a2da2424f6796f64193de6dee4576a86c60d53be7402ecbb0d69e6;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'h86cddd34a5a13e85c0a9ca53be1b2ee9b1619068755ea0a4a4d6d2f013436f9d9235e694e4708241710ff9398f4dc4f04010729648baa1d83d4812a9d0198fc676b441e6e2a8bcd0eee9724350b9dc73e3782d95044ae3741fc1a3615c1a0af3230332ad5f81cf2df3aaca2961acf83aa74418f08e02b86d3c0ac223e4027712da640da38ba7bd0ab3bd8fea7972e1a6acb3f595688df514f3e3fb037077185882cba0e56a660803a1d47b5203bc8e8769af1e3617c25d03271f7e0bec58d3c5;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'hac968579b27e566e1b1b5423d78871bb6e75826a1649b0645bf11287716294b41d0a42f84774f5638501f7b40d299c0bd7169eeb186abacb17d4258159265c78114136d6f423f514fa57fb8e1636afe27423e337d8709a0e182180485617634a103ce015c55c794e01cf3c9a86ddcda76be884e75f77df543aba9256763d659d6327ac155b0b8557173cd2fd2e5ae1b15ab38c10a8a25a39891bfed90c24fcf70af203ecee3f56f361f445e4885b11e1d21e14169f0c349e624ff50fb8d916c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'h1c8ddbff940804b01a41fe01d4df3e8a10ceec7417794c79df83b8556393082fb1d27bff08a028b283ce3fd5861c10f93167a418c069819ddcdf71d6742e58b6997de679a013a7adbaccccc51db3a94f1720b95f3405aea81f4840b5f862e50d6d88c41799baff7297bba9e5ebd02d7a3f0d8590f2a8642d124493a27f668c45daeaee8908c1d34583c8a48a65ec1f803a10cf164d4f9f6e29dff651b58e434a170406fd4c67ba9099cfb586f63ee80b0868e997558d253fb570c3e52c6370f0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'hd2ddba860a361ff966a708b6723871eb0a4a843332920801d74624afc903e0b702083679e1a3be489909416404e696a3d42965839fca239e19cf1d7926dd7eb55be7413c650e29502c22c3223104b6806e3a2dd2130bb8f953c7f54ddafd8a128a0f6e712a48f5f97ce413dd668fab4100404d69762aa131fcd4f5c237d6d6148e17ba8be744304376a1823a00be6ada00bf2a2656e12c6be384b35a9b8ece8ffe7e3cf0ef3cfb6dfe308665f5b4cf686e9771ea965eb4d445c35b8aa9fccc3f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'h8e52140dacba89fac94c7aad78e9534a78a207b9947735a48255ab0bea833780eb52229e72cdd0ad23213e28a5fefdbd656aa7546dbbdd6a406107b63535f196cdd8722e7e04c7df2bbd6ae9865c222d71f680a3ccd0329b396e7aa94be81a045efaf711b49ec56975dda40128a245c3eaf2ef30e03d6683eb1f8661d5f85297d6361d893e842982d2e80fde22d99e51d6999045f6d78bca0cea4ccd5d77d1825c335f315ba1ac258681f8c12e2ad27acd4d26a65d5b08096c008841634e6925;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'h2903a1760fe0eeb736acb53156d6283d36341b3a96b82457100124f6588b490ce68d62d76973e3d0e03b94af4ad40f78fa672a968772d96c605f2ef6750012d1d8a02a53ce0fb3ca0bedfffe894f83de904f9f3e751e1bd8a25f13d1b03724d65e6e76afa5ca06209b99dcf1822fcbbb99e3c3685988c8bd94b7d1f86ea048f8a847624152d0ec35a6754190a3446e118390544eab88560d683ff4a44b2b4828ff5219ea08f7dafe4a281762b241d9e195844b35571ede51b07f7254ff030665;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'h67d4b139ff1ce7850522973c7032996241b2dcb97847e990fe4a5749810a27c59fc2188fdad91ec520a7b2a4f8100ed8ad7dd3a11e2fbafd1bab807682335a1382570e3d6430b495e68787d80a5b4c9c5a8310da76ee6c8ec4acd22ab0e7d810ad2bf335dc963d3219a9d5bc55c21bd909ec6e0f6acfb5ff329b29725b5bfacdf79344598fa9d6f5c9cf8e6ec4baa495d5859999dd336798e1fc9e166c92b5ae9f62477eeb36134d9743e62e697b4e784fb500f830637b4aef9eb343ac878e1e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'h9a8770156575018e06c2988d9f66c4a1753ea48b6dd0ee617296f5797168e21876a7180f0dc975b86827ae9b6179ed7f4a605a0f11e0b5b0e9c7ad7cc8e32459e3c8dd548a894f6af22ddb524e679c9c55fd486ae04103d87103e861dbd7df05dbadb552efdfc9bff853916f2cb04ec74fe207a50aef72fd24e793f54710b853b406b9bcdaa63115f6aa7f96310341cd7206306a074e3fc972503367b4fc61fb123c274e0df930b15124426e8380065be857663ff01c0e889bd50bc7e4b0fad4;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'he32c29a37c56d3ec05b73c5bb7d44dbca2510550566bc115d572f8109071538833f62f7c79e2fa39d9e9279bd3dbbbbc402af24538cd963789463d742e04a55b562f1d361215874a51d8b018055acd943823cfc1a17a17ca3006493aaf4edb8986da8615c72a38ec9c827fbbd0c1605222a999e385dc6f51170a69b9ae53cadec9534b8cfa366ba8f4e457a27bbae23b7d85d7b3b8a1d6a01e846ffa3653de30ae06c389133fe9a5d82b7c44346ab4b9f548cab766d340ec07bf823984fc5dc5;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'hf0ec7d9aa49e2ad1cc40ec1a07fd2cf40a0a3b673d1f24e08b454d853c2a7359d509e632a47714f51b864df621e40fcd0b06d13092a7b7b3f7eab98a349c91a6364f8bcc836296d18e630acf0f4ef6d6ed30db65e6e664e15dace1e4e362f1c8a9fb06fa3ad0021f4e6aa42362aeb86dd8240e838b910ba01a0d77d1deb538c61d727353224ee7ff6c71d37a543761477e13e5fa82eb317d162a8dbfb379dc44a7a1ba42ee7cb28bb92792ec5dabcb5fb94958876b326b5139330de058c1b2f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'h62a2b6c5af0a354ef730dc8f0f283bcd7bfa70950c90a691860206f5c83a890d8a677ea5e32019fa6714052cf383866e47ca7232d3cf39c5695876a2dab6f6b4e2b65a616c51d5eb226e894380ea8f41c65722fe768a83c1c056c47a9ee05d1cfb177e1af38507f3f6a0a3c1fdabb3c414f8413134b892f336efd4dd3380233ce14862f4f7e755736690b29d2da1995e6551ce69c66c3e8eb1bdbbe2c39ce1ceaccdfdc4fa478b71aee50f11429e6179373195c30ecf0d6824822196e38f4150;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'h1158839dd004a4b99ab572609c26f3e42ff9dc543375e3852e6d22c013dcbfae99a237aaf762168e4409f45f9cf8fceaf365f1d7bf0a0f33043608d57a9cfa6cdb41c66652db387dc779f35f1a39920d3e2e7ec9847ee891f166aa34877c87eadbb46b41d983da03b6ba3f5e88e7dcf6dca011e05127daf332b6676fda0a6a9e6c34f5c173f0b9fbee67ba632654147ab902d4f6c996a4d110eebaea394d3caf4771027fcf086382564de49a7fa198c47b28669bf96ea5ff073fc66fcec35124;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'h195bb798ec69608fa64dfc015826ab49663875e2b6d66bf97d5957771c58332224647a689db505baf52eeaf6665345b6d854894e6e892e8afdc4b3695c63fb98cec8c75f135c57a577f6261d9d73dd4bb76446f798f965d57377dac4e5f89f26582761963ed7ca29ec74eda7255b14b617b04eb653c6ec55bb1f60b291b1a854823c106e3c1f9a77652736b83617bc470a060d7d47ae8a39905a19d2dfaeef810253ecd7f98227ee8b40960f7c9b3d234f967a67f271afd0068773b3020c8040;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'hcc9dcc757dcf94a07618e0e48117e4a0b342cb0f9fa1546d860cf92e2e2b899a5bc5e73882bc9be83ced76f101c4f6310ac059a2e71afb4ba6d33dd7e296cf96657d1784b66d18ca8cce1ab5e18dd99b6470e8e0f73e8241878121bbc327d74926737b38af0580bd1936deb5efd66479843855a8c243f7d2a8e80eb4f7ac020041f51ef87e816c9aca9ed3c2e419a7c092dbaeb1e3e8bda5f3f2d34aa5bc867909118a1d87c8c3d8af4738a870c739ea94b3f90960481134dbfd0767284bfbb9;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'h688368ba6d3a26f5b53864f90e5462e5dda3e2271df5409cfdde95e49cec94d3d289fae95caad79fea45dad30d45211349c9f918f84440d429efc98321320062108f82b2252ace5b94170c9d9cefd5077310187d3ca8f194114806c85677af0e6e19090c38adf4ba92fa4ceccf97b27ed73effb83e5d89579ce46d76a9919563ced3eeb0d11f23833bdb86ef0a012b99ed0e241ff477137a01fe57b076a179ed9321b1fb1ccf49faf3e922a12ec8b730d0240bd03bae727c8e5c083164d3daff;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'h15872ba2d4bca5f82846a5eb4a3dbaa0821a1758ca0fee870d98462d7edc38b82e73382d7aa937582689be2ea70867181baa0b24fda6be2a069c2379fd0cca594772f719464a79538fd47d1cb2a7b894a2e72035c79e4504e821bd4e234ce38863392d7e1e6efa3f38ca6f4c8ec217d3894c1a21f655f2e821ead938de094d157a084ed84e69bd925eea6f3275bbf5a9c499e09bd7f61e79d6a0f9a48833eb719716b381ae6d9562c7a00fa566d0919747f9a4314b44ad5b7fcb8dcd06c97a29;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'h68f4b64d1261b2aafe6df3b9f9f3e176bcdad6ec989e1fbd3f4cb41123269d097cb5d653bc9c2d4b6ded925b9fa80e5abd038316e66afbb1cfa2567723a3fd801036c01bb085c8c571211615983755889e770f92e73306567c375f2466efd66dbd068d439034be6cc2754b7f4cebb0c23b62fd80cd52eca9a86a71aaa32c89c3c9df4da13f8ef520e15eb79774468408f929b24f2d166fd01b8056871c27abe93b5ecd87ca2a3b8f1353cfa8528743488c89f466e73fb865c7577cbe50011ea8;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'h3e31720d0234b0532bd748e0e3f188fb56e21d4940f54592c251461c9cedd9c2cd3945f38d277c67cbc14fe2487576f2f06c117b6a71302740e437e652aac0e310e5f7baae472792ddec1f159df8cb137a31d9220664305da5a2d9b03636f5ae1b2fe1c8fa8a1633fc24f76168407fba757b1fdd99c98458e1f973f7c3af4fc01ae05563ba3c9dfb41866937ed4c5399e0aa78b50f1949a4d81127c94e271e93e23185736dfc6e26eba2e14c4bfa770e1e794c876a51fc6f9d612b4ef117399e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'hddb34d3c587c43fb4bf226bcc5e18927a81c95cf32ec72f4df502aefb3e3b2c4579a22473a57d9d91e855866b65bdf77c1f483d6f040f1bd52376d6bff4a1cf881a2e0d529c6e09b9e21695079d3717f0d463bdaa27785dd84b52b4b194821659640638897072c4b2fd721a2d29df2f2ad663b5a11b877806a63c72c0617c926f80065e26f7dfc509a4712aab48ea1eb9ac30c0eabdb01ad21d3ac0a56f2bbe6940e4d4c3b25bb0458469c0559ccf967c7c246bfa5aba5228e79d1a6457efeda;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'h11e3067b625431b0e33db2d25687d65c27f6c0cbdefe64884523366da663a2b3c4645908ed10d2fa957a1de8b5354b6095b4103c8b34772e20ce0f915b65403618d8aaebbdb6c897f0d532e5bd3b2c8c4f9ca8bc8585a5b1711166602bc51167f5ab435e1f98dcb938cf9d08ed7f66a3566941c766ed3674328db1eb0d6373f7943ac7fcb8b65044da13fb99c5455b33fb49487dbe86f1b57a8ca79ea23dfa5d7b9a5814d179a3b5163c9c4ccc5c0297a663a3ea21d21ca1865c95daf4aa05bb;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'h57ae2ea8a5eb28360b9dc14e47c1086c3a1849b7e7a5223040fbc4d0604199b81733f1adb54df08a207ae700f782807a9427f888f5a1fd211d1b353d57a9900dad16a38541fafcf77a4452bc69011d9c551cced33ae1ecb150d80ae5f63e03a20be610344f1ecc04c4faf41ac701f65c3b01ab8a1df8b98d8c77d14417928286917bd330a7385e76307caedeafad9ecebd0d045edac6ecfa5777d20a2d5aa3c779b244e13ac2912b44db37f90fae2bd4016952cf96c4c60e12b3ff730d4c0337;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'hada3017de63ce91bcd4014372e4f0d700f56aa567d9ee24cb098b44fb6b5c505154e9620cf9cda919c5288d4cbac78be617a855b7f40892038932efc456e22fe38a366c7a644c5afff298dae0d35e09f6b2fc575e145444094ecb92965ed94e6f99e95aaaf7d12c5c2a5d85ba379269577c15e951961a8e5fcdbffcc1d51f1a295d4e069f9296f4c99c84a809e05b4566e549836fe7504bbb3ce084f4795f77b099088105e720b02a6ae3d4886fd0fa62408e0fbb39ad82e280ea19ab2779e02;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'h415c591d0fb63317caab23963d21ee40cd92f3fc0ca4d53b264548c149b2c3985e535cd205bac073996ad34e5a7378e2868d1033ea1349d35c71df6abd636c21df2ab3e4eec84a3c80a2b87359394d0594c9bba507e280b7fb2ab49d63e52e18a7edbac22f65a2becaa00542a16f69d1c046da5ec9948d9134cf349777b04c00b9ddb280b970370f8b02dd015a463df59bf9bf734e1bcc2ef080e055a863a9eea29eb68beaa0cbc54333208eab8d8e49333c16386b4e5c37bec9439a9504ae93;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'hb50f515061523bb27a2e6d959ac30de1a66f597a84228247b30efa267bc94fbd4710b3be4e58a033595492ce4b627a4a52488ef18a9e1ba5f767dafc0f6fc768e1a553f578b063dbd596aee56b5194db0f0e23e77f6fcdbefb9a8a087843313e10cdf7615a195238e4f0cc6b160151a68f27565347560141a017caf873b65c2898047998ba375066c68b41819935a826e36c45b82977df4941f51884f3a8db6e39035d95b8235c7af5d5aaec0869f25e3de6b06069dc9824b8ed8d377e1be9f9;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'hfc4704f2762423694ad3b45766b6cdc4108b4ed943d3e9e7f5a9b6b1bfa9b3b35d450b254a3bc47e0682ebb3177d01dacfa626ada1980fdf407830338ae2aafee67eb0527cc29b290879b65d4491877c6baa8e3c58f1e64a17a8e07de497f0586424d442dc866ad938e5144fa997fa1544947684ae90d9aebdb6a57f087bb0766c67b859006c71b31dd2cfdcb661257548d119e2efb69c6d44a6f77cd5e4554bccd5f96e951d6cb2c337acb27fa87cfe301c13a23cb0ce4a7832e67084f322ed;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'h1781248b706051ea93f9c137d9e02749c0b12aa7e695b62297cc26048c1b21fa8d808ed5863e1249bb7e2b57d7f35502eeab5121b82c37d6ab7402232a3e6842464a0fd1151baf8774d7d712cd10abf5d1caa596e23746109e1e6f4b8b2da155c7a8d1692476f156ffe357c332b512f6721d7274d9a289054aee308cb3d593685eb761c572b1281eaca01b512ab19a2c142fd9fe172baa77db48e5a474c63690b1893f9744f23b66d723241e6e65ff39f34d1d6de1deaada5c02f9d2339350e4;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'h4234d3840f8fc862e382453c451675b91af35729c2cf9489c6dfda250eadde2c4bc1284f20cda2b8f184cae0aa2043d6efeb2cb55524fa8fd879d14efbedfb1249326d9d8b240e6e75e255109358c344cac17b9528a420073f255ee26be48ca024dd71cbecc672a25e7a39e22051bba47179a191e155ee755f484b6d7754f817b44aec9a97c83ef17a15ad81204bff2ae67fe48415dc4be2c5a3c1152c0cd0574ef0f534d6ff953d808154d151f08a3591ece75b2ed16b4638288d5549fc2627;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'h31c62a2f2f9da4b02221fecf6c7a085f0616dfe623918cc894d0fb2d1aee59ac7fa8c1b1511d3ed175838644e2c4d24e6d5927693be291cea59253c65b34660bbb84dbfee6c760ebb91a415933c82899c89970ba568ce884f5f53e2324496436591a5b4617dc680de52e10c89d3844b4a84a529a5d123a76f13ed616ed14f465b6e0f7b8ff8ab9401943b2862cde13ce68d576fed5de5b79978946b0354d0ea21117b904f4d9434f9d0a761c8ba77b7adea677fc1bce0a880baac3d8db53c4ca;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'h737b174c8e51b506621d7cf30750154c7c4dd2405764e69707cc0131c2e3826c40f1d9943edf34f920b287e03241be23bb3691e4fa8410477bdb1e8afd1d767252da30ecb9a150f6498ffa411392b4dc592918d8df3a0f9c7c9562a259210874bccf619b8d645379106fdf2d7378345289afe09dcf7c49cd859d815f4f1723ab7d910ccfa45d9856d24781fe8e0968b72949c8c5fd5afac3ac3e3fb4ea52ba4c3c17ac542596c3f6c256a7ed1ab336d666f21a0b72062dfdafc345bc771a3dd;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'h819a03d03442a72031c0ecd1bbfa21d979a98d6c675f4851c67260a713f7c53ad43978aa3f0ce1c32628bcfdc035e51e450cfc250f83ea89cbc8c3c40e49bca217d4b1441c29172caf1506936b04ba8ffb787d86c1ef455c6cdfa3a8d3e81e5b33c3782c2a845b88b667e1b20fa5550a2ed42d1bea52b89d3d9032b61e27def4b8fa0698ead41d3f7685710a50ca46e7cf1f413daf91a8a57fc38d33e91d119041ec46919ef92d80f1b47d13da8622bbf71af862fedbf37e381ee38c98895d3c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'hcc2be72559583bea96f0597ed82837a0c6c455bc45476f287ba478d29fcf47bac8ca9af639fe1cd34c50e9649f5b822592e2c8a5e3705799833e34ad19af8143a06fc87a8f635deb2f43191b0cdf3ebd2027f777288fe78b5eec16c8d1815446cc750d9dc97bfa91b5601a592033e0711b8fff8009d31392d9a31075ee322de18167dc068994c8e0009517e64f925595c3ddc6dc894a27ccde59090966283ed6f7a0803d1f310c943b399b6c1d7bc82910b46b56457ba6f04cb4e988062e0588;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'hf8982830d920403ceb31746d809c989fff22a698388934ed5a767f9448291851cf54066182ef8526c9e223cec1f7fd906ab858ce35ebc628d92f9f638eb5d80d7085b029d00185d0bf97b33e54179dd5fa7f4eeb944e2aa3256ef203d28e492491c8625f806ce91cf303243d9bdcd8b5c69a60c3a2ec247d2d3456a47649672262b32ee808d59369415ef377c7c946cee523c5da6a5d6bad5834c521b4f1306e30b72772d6217324010365d18c8a54cacf181fd00172474824de003be7c0c070;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'h20fc53785cbd30423f3e44e5fdce93c481f6a190daeb2deae3ab660b453f05f0ce1bc2118ff80547623f8cdd52747c4413434b31cacb6f9d351f70cbaabbe9ee05a9fd7729da2e67cca4c5c20660a3306c1b68422a81346bf6d6d48a3314368a3b4927a7301822758e8daf763d63fea3cccdcdeae488edb8608ea0172c01edc3a91256720da801fc8561d502191cee25415e84d741a0f7cf6420b21dab570c665959d2535a36a7ef6a9230de9966b5a190ba23cf0b291d12db695b0bc04e9610;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'hba64afb2886bd7d47b7fe35a5e09747c0a03e94b59ffa6b06b1947cee8cc27f325c89f1c3b2a713e0b426ca9be04b17d7f2aff76e11f7bcf4ca0c6c507fddf6b7d97e116acc90f8f11df46254afaf3ebfbbd697279dd3d8e77ed468dc0df353a8aa9769acd1a65cfd2f8f742003a95982f46d354a2c22c2feacd2f9f38f99cf66898cbf59a280af6d23ec9b2768ceb418995a235b75774f5eff0fa3fd954b75b42d9aa4d6501b9d345355e07ff38b3e31bef65e103442718efc00d862be76d2e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'hb4be5684f164bd3e9b476e041d80f6b548f2f1bc37039e65aa64fb266f77a72174d392b7e74a5db23e79ac20887f8e19b3bc8d848098805e5a5be54306370e46819491513a66c38195091d2fbe996251463335a01c42dd71fe070ca18410a68eb419c899e1ff49958db1c8cb19dae571d39a577718ca9462c3ee9b781ea61132338cf7e7097d365eb4e09911b1355d979e6c169c13d427251db53edcde307c46e61425ea38881a604e7abc7559645cf39354aa8822401f68af67071d8808955b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'h7993d8b5a4527e52fede2b1af1e8b91c3148aeb4d502c2cb50eaa1566953c21f1ffbd2155f258096fb37031c62357a11137cd3a12a9107c6cae014473e6b51b34c50110b9964ef1366d1109c4a252e047f82a63814bc02bb41343454e6dc2b3126efa681c725770989aa4e7e0a41f190f844b03a80062d65815343b9294ac84947f2d273761e82b457a84b7c23f7ff132c7f90c2ea2cc6ceb3f1f40f6200aee415ab45808e75952157b27b0ba9831dad3d4ea6c6b08e284bc45f0108fbd8492c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'hd2254be1cc796fcac39b5c3a04f58adb9274a5d0c06d7adee89563973709dce13d54ad18d7348f519ae3c1e998c0c50090fa73a902c4a831916ad0c1cc251066852d4e2e8ec05e2d67ded4f36d7b9175f9ec1df1d3fc1bcf447294ee635cfa3c0e0fb6494b209beeb8835386181e4963dec74bd21bc7c6bc564ced194e67437800e3da772d90d7308dcad0afaaf4b482c7a5e1322fcc6dea632db87f4bc7cf81b0952dd179a7cb211431e1f49c528484ba270bfa99c51e8f7bcce08d9636ed32;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'h6898120c28741a47d34eccafb2ebe8a3f5e68c3918374333f52dc5eb62a2b7433dcdf625e8bf31b84719152d476cde67d3dbf4b31da8a715d34e01222923927f10bda004fe2067c2ec9d9ff1a37104d60cbcd43e1d36962ad98f835ef7b88ec481dfaaed23a2e044897d285e6843cff1bffe3f046390561712b0c40293ed54fe38366d27f242e9460e7b809797b260eb790c63f3ea52c0f8382d981cc9cdebe01251dc698f0a03702628ca1eff7e1dde6c901d384d72f383e126aa0f4ac41801;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'hac0cc21a65d4a97a2711ef8350edd72ccc24e7e6e92829d323376ee5ac3d574fade8c3f6c4686b5e46053f2508bb047ea385f8b09854e733a3c41e844141c8145e03a566ce9320465df844adc4014f8399bafdda939c603f117e9547897c538a5464354b9073293b81d4498fe1f3524bab428c5038df68e09923b9f22a58d166a951f98fef7baa62e1bd61860bd5526da2354088b85c77852930afbbaba5ba982b4d262aa9b9c990877dfe67241f13e103aa066ee7e0c0256831069aded58631;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'hd642538b1344a437d25f9716f866b72d16c53836b6f2561b9b0bbacacaf540a0be8adb38af2bc70ea1a6966defca97be991d572c36f173c1e238f00414da1c174be8a7c8232e5a3839770747d6bc0876038bfd7559db3ecee00de5b84df57c5c48d18e8b6d790e125bcfc594736530d653cc8e691beae6a9284973c4edd79bf65a7d0a1d3bae91e6ed17372eab0b92ebab0913851e773ea7c908f55549c634265c05d23de26e6e8f1af44b6c5151cd627a7cb93c4143c6ae8ad5bcacb85c1a89;
        #1
        $finish();
    end
endmodule
