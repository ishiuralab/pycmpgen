module compressor2_1_54_12_shiftregister(input clk, input in_data0, input in_data1, input in_data2, input in_data3, input in_data4, input in_data5, input in_data6, input in_data7, input in_data8, input in_data9, input in_data10, input in_data11, input in_data12, input in_data13, input in_data14, input in_data15, input in_data16, input in_data17, input in_data18, input in_data19, input in_data20, input in_data21, input in_data22, input in_data23, input in_data24, input in_data25, input in_data26, input in_data27, input in_data28, input in_data29, input in_data30, input in_data31, input in_data32, input in_data33, input in_data34, input in_data35, input in_data36, input in_data37, input in_data38, input in_data39, input in_data40, input in_data41, input in_data42, input in_data43, input in_data44, input in_data45, input in_data46, input in_data47, input in_data48, input in_data49, input in_data50, input in_data51, input in_data52, input in_data53, output [17:0]dst);
    reg [11:0] src0;
    reg [11:0] src1;
    reg [11:0] src2;
    reg [11:0] src3;
    reg [11:0] src4;
    reg [11:0] src5;
    reg [11:0] src6;
    reg [11:0] src7;
    reg [11:0] src8;
    reg [11:0] src9;
    reg [11:0] src10;
    reg [11:0] src11;
    reg [11:0] src12;
    reg [11:0] src13;
    reg [11:0] src14;
    reg [11:0] src15;
    reg [11:0] src16;
    reg [11:0] src17;
    reg [11:0] src18;
    reg [11:0] src19;
    reg [11:0] src20;
    reg [11:0] src21;
    reg [11:0] src22;
    reg [11:0] src23;
    reg [11:0] src24;
    reg [11:0] src25;
    reg [11:0] src26;
    reg [11:0] src27;
    reg [11:0] src28;
    reg [11:0] src29;
    reg [11:0] src30;
    reg [11:0] src31;
    reg [11:0] src32;
    reg [11:0] src33;
    reg [11:0] src34;
    reg [11:0] src35;
    reg [11:0] src36;
    reg [11:0] src37;
    reg [11:0] src38;
    reg [11:0] src39;
    reg [11:0] src40;
    reg [11:0] src41;
    reg [11:0] src42;
    reg [11:0] src43;
    reg [11:0] src44;
    reg [11:0] src45;
    reg [11:0] src46;
    reg [11:0] src47;
    reg [11:0] src48;
    reg [11:0] src49;
    reg [11:0] src50;
    reg [11:0] src51;
    reg [11:0] src52;
    reg [11:0] src53;
    compressor2_1_54_12 compressor2_1_54_12(.src0(src0), .src1(src1), .src2(src2), .src3(src3), .src4(src4), .src5(src5), .src6(src6), .src7(src7), .src8(src8), .src9(src9), .src10(src10), .src11(src11), .src12(src12), .src13(src13), .src14(src14), .src15(src15), .src16(src16), .src17(src17), .src18(src18), .src19(src19), .src20(src20), .src21(src21), .src22(src22), .src23(src23), .src24(src24), .src25(src25), .src26(src26), .src27(src27), .src28(src28), .src29(src29), .src30(src30), .src31(src31), .src32(src32), .src33(src33), .src34(src34), .src35(src35), .src36(src36), .src37(src37), .src38(src38), .src39(src39), .src40(src40), .src41(src41), .src42(src42), .src43(src43), .src44(src44), .src45(src45), .src46(src46), .src47(src47), .src48(src48), .src49(src49), .src50(src50), .src51(src51), .src52(src52), .src53(src53), .dst(dst));
    initial begin
        src0 <= 0;
        src1 <= 0;
        src2 <= 0;
        src3 <= 0;
        src4 <= 0;
        src5 <= 0;
        src6 <= 0;
        src7 <= 0;
        src8 <= 0;
        src9 <= 0;
        src10 <= 0;
        src11 <= 0;
        src12 <= 0;
        src13 <= 0;
        src14 <= 0;
        src15 <= 0;
        src16 <= 0;
        src17 <= 0;
        src18 <= 0;
        src19 <= 0;
        src20 <= 0;
        src21 <= 0;
        src22 <= 0;
        src23 <= 0;
        src24 <= 0;
        src25 <= 0;
        src26 <= 0;
        src27 <= 0;
        src28 <= 0;
        src29 <= 0;
        src30 <= 0;
        src31 <= 0;
        src32 <= 0;
        src33 <= 0;
        src34 <= 0;
        src35 <= 0;
        src36 <= 0;
        src37 <= 0;
        src38 <= 0;
        src39 <= 0;
        src40 <= 0;
        src41 <= 0;
        src42 <= 0;
        src43 <= 0;
        src44 <= 0;
        src45 <= 0;
        src46 <= 0;
        src47 <= 0;
        src48 <= 0;
        src49 <= 0;
        src50 <= 0;
        src51 <= 0;
        src52 <= 0;
        src53 <= 0;
    end
    always @(posedge clk) begin
        src0 <= {src0[10:0], in_data0};
        src1 <= {src1[10:0], in_data1};
        src2 <= {src2[10:0], in_data2};
        src3 <= {src3[10:0], in_data3};
        src4 <= {src4[10:0], in_data4};
        src5 <= {src5[10:0], in_data5};
        src6 <= {src6[10:0], in_data6};
        src7 <= {src7[10:0], in_data7};
        src8 <= {src8[10:0], in_data8};
        src9 <= {src9[10:0], in_data9};
        src10 <= {src10[10:0], in_data10};
        src11 <= {src11[10:0], in_data11};
        src12 <= {src12[10:0], in_data12};
        src13 <= {src13[10:0], in_data13};
        src14 <= {src14[10:0], in_data14};
        src15 <= {src15[10:0], in_data15};
        src16 <= {src16[10:0], in_data16};
        src17 <= {src17[10:0], in_data17};
        src18 <= {src18[10:0], in_data18};
        src19 <= {src19[10:0], in_data19};
        src20 <= {src20[10:0], in_data20};
        src21 <= {src21[10:0], in_data21};
        src22 <= {src22[10:0], in_data22};
        src23 <= {src23[10:0], in_data23};
        src24 <= {src24[10:0], in_data24};
        src25 <= {src25[10:0], in_data25};
        src26 <= {src26[10:0], in_data26};
        src27 <= {src27[10:0], in_data27};
        src28 <= {src28[10:0], in_data28};
        src29 <= {src29[10:0], in_data29};
        src30 <= {src30[10:0], in_data30};
        src31 <= {src31[10:0], in_data31};
        src32 <= {src32[10:0], in_data32};
        src33 <= {src33[10:0], in_data33};
        src34 <= {src34[10:0], in_data34};
        src35 <= {src35[10:0], in_data35};
        src36 <= {src36[10:0], in_data36};
        src37 <= {src37[10:0], in_data37};
        src38 <= {src38[10:0], in_data38};
        src39 <= {src39[10:0], in_data39};
        src40 <= {src40[10:0], in_data40};
        src41 <= {src41[10:0], in_data41};
        src42 <= {src42[10:0], in_data42};
        src43 <= {src43[10:0], in_data43};
        src44 <= {src44[10:0], in_data44};
        src45 <= {src45[10:0], in_data45};
        src46 <= {src46[10:0], in_data46};
        src47 <= {src47[10:0], in_data47};
        src48 <= {src48[10:0], in_data48};
        src49 <= {src49[10:0], in_data49};
        src50 <= {src50[10:0], in_data50};
        src51 <= {src51[10:0], in_data51};
        src52 <= {src52[10:0], in_data52};
        src53 <= {src53[10:0], in_data53};
    end
endmodule

module compressor2_1_54_12(
    input [11:0]src0,
    input [11:0]src1,
    input [11:0]src2,
    input [11:0]src3,
    input [11:0]src4,
    input [11:0]src5,
    input [11:0]src6,
    input [11:0]src7,
    input [11:0]src8,
    input [11:0]src9,
    input [11:0]src10,
    input [11:0]src11,
    input [11:0]src12,
    input [11:0]src13,
    input [11:0]src14,
    input [11:0]src15,
    input [11:0]src16,
    input [11:0]src17,
    input [11:0]src18,
    input [11:0]src19,
    input [11:0]src20,
    input [11:0]src21,
    input [11:0]src22,
    input [11:0]src23,
    input [11:0]src24,
    input [11:0]src25,
    input [11:0]src26,
    input [11:0]src27,
    input [11:0]src28,
    input [11:0]src29,
    input [11:0]src30,
    input [11:0]src31,
    input [11:0]src32,
    input [11:0]src33,
    input [11:0]src34,
    input [11:0]src35,
    input [11:0]src36,
    input [11:0]src37,
    input [11:0]src38,
    input [11:0]src39,
    input [11:0]src40,
    input [11:0]src41,
    input [11:0]src42,
    input [11:0]src43,
    input [11:0]src44,
    input [11:0]src45,
    input [11:0]src46,
    input [11:0]src47,
    input [11:0]src48,
    input [11:0]src49,
    input [11:0]src50,
    input [11:0]src51,
    input [11:0]src52,
    input [11:0]src53,
    output [17:0]dst);

    wire [1:0] comp_out0;
    wire [1:0] comp_out1;
    wire [1:0] comp_out2;
    wire [1:0] comp_out3;
    wire [1:0] comp_out4;
    wire [1:0] comp_out5;
    wire [1:0] comp_out6;
    wire [1:0] comp_out7;
    wire [1:0] comp_out8;
    wire [1:0] comp_out9;
    wire [1:0] comp_out10;
    wire [1:0] comp_out11;
    wire [1:0] comp_out12;
    wire [1:0] comp_out13;
    wire [1:0] comp_out14;
    wire [1:0] comp_out15;
    wire [1:0] comp_out16;
    wire [17:0] out;
    compressor compressor_inst(
        .src0({src53[0], src52[0], src51[0], src50[0], src49[0], src48[0], src47[0], src46[0], src45[0], src44[0], src43[0], src42[0], src41[0], src40[0], src39[0], src38[0], src37[0], src36[0], src35[0], src34[0], src33[0], src32[0], src31[0], src30[0], src29[0], src28[0], src27[0], src26[0], src25[0], src24[0], src23[0], src22[0], src21[0], src20[0], src19[0], src18[0], src17[0], src16[0], src15[0], src14[0], src13[0], src12[0], src11[0], src10[0], src9[0], src8[0], src7[0], src6[0], src5[0], src4[0], src3[0], src2[0], src1[0], src0[0]}),
        .src1({src53[1], src52[1], src51[1], src50[1], src49[1], src48[1], src47[1], src46[1], src45[1], src44[1], src43[1], src42[1], src41[1], src40[1], src39[1], src38[1], src37[1], src36[1], src35[1], src34[1], src33[1], src32[1], src31[1], src30[1], src29[1], src28[1], src27[1], src26[1], src25[1], src24[1], src23[1], src22[1], src21[1], src20[1], src19[1], src18[1], src17[1], src16[1], src15[1], src14[1], src13[1], src12[1], src11[1], src10[1], src9[1], src8[1], src7[1], src6[1], src5[1], src4[1], src3[1], src2[1], src1[1], src0[1]}),
        .src2({src53[2], src52[2], src51[2], src50[2], src49[2], src48[2], src47[2], src46[2], src45[2], src44[2], src43[2], src42[2], src41[2], src40[2], src39[2], src38[2], src37[2], src36[2], src35[2], src34[2], src33[2], src32[2], src31[2], src30[2], src29[2], src28[2], src27[2], src26[2], src25[2], src24[2], src23[2], src22[2], src21[2], src20[2], src19[2], src18[2], src17[2], src16[2], src15[2], src14[2], src13[2], src12[2], src11[2], src10[2], src9[2], src8[2], src7[2], src6[2], src5[2], src4[2], src3[2], src2[2], src1[2], src0[2]}),
        .src3({src53[3], src52[3], src51[3], src50[3], src49[3], src48[3], src47[3], src46[3], src45[3], src44[3], src43[3], src42[3], src41[3], src40[3], src39[3], src38[3], src37[3], src36[3], src35[3], src34[3], src33[3], src32[3], src31[3], src30[3], src29[3], src28[3], src27[3], src26[3], src25[3], src24[3], src23[3], src22[3], src21[3], src20[3], src19[3], src18[3], src17[3], src16[3], src15[3], src14[3], src13[3], src12[3], src11[3], src10[3], src9[3], src8[3], src7[3], src6[3], src5[3], src4[3], src3[3], src2[3], src1[3], src0[3]}),
        .src4({src53[4], src52[4], src51[4], src50[4], src49[4], src48[4], src47[4], src46[4], src45[4], src44[4], src43[4], src42[4], src41[4], src40[4], src39[4], src38[4], src37[4], src36[4], src35[4], src34[4], src33[4], src32[4], src31[4], src30[4], src29[4], src28[4], src27[4], src26[4], src25[4], src24[4], src23[4], src22[4], src21[4], src20[4], src19[4], src18[4], src17[4], src16[4], src15[4], src14[4], src13[4], src12[4], src11[4], src10[4], src9[4], src8[4], src7[4], src6[4], src5[4], src4[4], src3[4], src2[4], src1[4], src0[4]}),
        .src5({src53[5], src52[5], src51[5], src50[5], src49[5], src48[5], src47[5], src46[5], src45[5], src44[5], src43[5], src42[5], src41[5], src40[5], src39[5], src38[5], src37[5], src36[5], src35[5], src34[5], src33[5], src32[5], src31[5], src30[5], src29[5], src28[5], src27[5], src26[5], src25[5], src24[5], src23[5], src22[5], src21[5], src20[5], src19[5], src18[5], src17[5], src16[5], src15[5], src14[5], src13[5], src12[5], src11[5], src10[5], src9[5], src8[5], src7[5], src6[5], src5[5], src4[5], src3[5], src2[5], src1[5], src0[5]}),
        .src6({src53[6], src52[6], src51[6], src50[6], src49[6], src48[6], src47[6], src46[6], src45[6], src44[6], src43[6], src42[6], src41[6], src40[6], src39[6], src38[6], src37[6], src36[6], src35[6], src34[6], src33[6], src32[6], src31[6], src30[6], src29[6], src28[6], src27[6], src26[6], src25[6], src24[6], src23[6], src22[6], src21[6], src20[6], src19[6], src18[6], src17[6], src16[6], src15[6], src14[6], src13[6], src12[6], src11[6], src10[6], src9[6], src8[6], src7[6], src6[6], src5[6], src4[6], src3[6], src2[6], src1[6], src0[6]}),
        .src7({src53[7], src52[7], src51[7], src50[7], src49[7], src48[7], src47[7], src46[7], src45[7], src44[7], src43[7], src42[7], src41[7], src40[7], src39[7], src38[7], src37[7], src36[7], src35[7], src34[7], src33[7], src32[7], src31[7], src30[7], src29[7], src28[7], src27[7], src26[7], src25[7], src24[7], src23[7], src22[7], src21[7], src20[7], src19[7], src18[7], src17[7], src16[7], src15[7], src14[7], src13[7], src12[7], src11[7], src10[7], src9[7], src8[7], src7[7], src6[7], src5[7], src4[7], src3[7], src2[7], src1[7], src0[7]}),
        .src8({src53[8], src52[8], src51[8], src50[8], src49[8], src48[8], src47[8], src46[8], src45[8], src44[8], src43[8], src42[8], src41[8], src40[8], src39[8], src38[8], src37[8], src36[8], src35[8], src34[8], src33[8], src32[8], src31[8], src30[8], src29[8], src28[8], src27[8], src26[8], src25[8], src24[8], src23[8], src22[8], src21[8], src20[8], src19[8], src18[8], src17[8], src16[8], src15[8], src14[8], src13[8], src12[8], src11[8], src10[8], src9[8], src8[8], src7[8], src6[8], src5[8], src4[8], src3[8], src2[8], src1[8], src0[8]}),
        .src9({src53[9], src52[9], src51[9], src50[9], src49[9], src48[9], src47[9], src46[9], src45[9], src44[9], src43[9], src42[9], src41[9], src40[9], src39[9], src38[9], src37[9], src36[9], src35[9], src34[9], src33[9], src32[9], src31[9], src30[9], src29[9], src28[9], src27[9], src26[9], src25[9], src24[9], src23[9], src22[9], src21[9], src20[9], src19[9], src18[9], src17[9], src16[9], src15[9], src14[9], src13[9], src12[9], src11[9], src10[9], src9[9], src8[9], src7[9], src6[9], src5[9], src4[9], src3[9], src2[9], src1[9], src0[9]}),
        .src10({src53[10], src52[10], src51[10], src50[10], src49[10], src48[10], src47[10], src46[10], src45[10], src44[10], src43[10], src42[10], src41[10], src40[10], src39[10], src38[10], src37[10], src36[10], src35[10], src34[10], src33[10], src32[10], src31[10], src30[10], src29[10], src28[10], src27[10], src26[10], src25[10], src24[10], src23[10], src22[10], src21[10], src20[10], src19[10], src18[10], src17[10], src16[10], src15[10], src14[10], src13[10], src12[10], src11[10], src10[10], src9[10], src8[10], src7[10], src6[10], src5[10], src4[10], src3[10], src2[10], src1[10], src0[10]}),
        .src11({src53[11], src52[11], src51[11], src50[11], src49[11], src48[11], src47[11], src46[11], src45[11], src44[11], src43[11], src42[11], src41[11], src40[11], src39[11], src38[11], src37[11], src36[11], src35[11], src34[11], src33[11], src32[11], src31[11], src30[11], src29[11], src28[11], src27[11], src26[11], src25[11], src24[11], src23[11], src22[11], src21[11], src20[11], src19[11], src18[11], src17[11], src16[11], src15[11], src14[11], src13[11], src12[11], src11[11], src10[11], src9[11], src8[11], src7[11], src6[11], src5[11], src4[11], src3[11], src2[11], src1[11], src0[11]}),
        .dst0(comp_out0),
        .dst1(comp_out1),
        .dst2(comp_out2),
        .dst3(comp_out3),
        .dst4(comp_out4),
        .dst5(comp_out5),
        .dst6(comp_out6),
        .dst7(comp_out7),
        .dst8(comp_out8),
        .dst9(comp_out9),
        .dst10(comp_out10),
        .dst11(comp_out11),
        .dst12(comp_out12),
        .dst13(comp_out13),
        .dst14(comp_out14),
        .dst15(comp_out15),
        .dst16(comp_out16)
    );
    rowadder2_1_17 rowadder2_1inst(
        .src0({comp_out16[0], comp_out15[0], comp_out14[0], comp_out13[0], comp_out12[0], comp_out11[0], comp_out10[0], comp_out9[0], comp_out8[0], comp_out7[0], comp_out6[0], comp_out5[0], comp_out4[0], comp_out3[0], comp_out2[0], comp_out1[0], comp_out0[0]}),
        .src1({comp_out16[1], comp_out15[1], comp_out14[1], comp_out13[1], comp_out12[1], comp_out11[1], comp_out10[1], comp_out9[1], comp_out8[1], comp_out7[1], comp_out6[1], comp_out5[1], comp_out4[1], comp_out3[1], comp_out2[1], comp_out1[1], comp_out0[1]}),
        .dst0(out)
    );
    assign dst = out[17:0];
endmodule
module compressor (
      input wire [53:0] src0,
      input wire [53:0] src1,
      input wire [53:0] src2,
      input wire [53:0] src3,
      input wire [53:0] src4,
      input wire [53:0] src5,
      input wire [53:0] src6,
      input wire [53:0] src7,
      input wire [53:0] src8,
      input wire [53:0] src9,
      input wire [53:0] src10,
      input wire [53:0] src11,
      output wire [1:0] dst0,
      output wire [1:0] dst1,
      output wire [1:0] dst2,
      output wire [1:0] dst3,
      output wire [1:0] dst4,
      output wire [1:0] dst5,
      output wire [1:0] dst6,
      output wire [1:0] dst7,
      output wire [1:0] dst8,
      output wire [1:0] dst9,
      output wire [1:0] dst10,
      output wire [1:0] dst11,
      output wire [1:0] dst12,
      output wire [1:0] dst13,
      output wire [1:0] dst14,
      output wire [1:0] dst15,
      output wire [1:0] dst16);

   wire [53:0] stage0_0;
   wire [53:0] stage0_1;
   wire [53:0] stage0_2;
   wire [53:0] stage0_3;
   wire [53:0] stage0_4;
   wire [53:0] stage0_5;
   wire [53:0] stage0_6;
   wire [53:0] stage0_7;
   wire [53:0] stage0_8;
   wire [53:0] stage0_9;
   wire [53:0] stage0_10;
   wire [53:0] stage0_11;
   wire [17:0] stage1_0;
   wire [17:0] stage1_1;
   wire [17:0] stage1_2;
   wire [17:0] stage1_3;
   wire [25:0] stage1_4;
   wire [29:0] stage1_5;
   wire [18:0] stage1_6;
   wire [17:0] stage1_7;
   wire [26:0] stage1_8;
   wire [25:0] stage1_9;
   wire [19:0] stage1_10;
   wire [24:0] stage1_11;
   wire [16:0] stage1_12;
   wire [6:0] stage1_13;
   wire [7:0] stage2_0;
   wire [8:0] stage2_1;
   wire [5:0] stage2_2;
   wire [7:0] stage2_3;
   wire [11:0] stage2_4;
   wire [7:0] stage2_5;
   wire [12:0] stage2_6;
   wire [10:0] stage2_7;
   wire [7:0] stage2_8;
   wire [11:0] stage2_9;
   wire [10:0] stage2_10;
   wire [7:0] stage2_11;
   wire [12:0] stage2_12;
   wire [6:0] stage2_13;
   wire [2:0] stage2_14;
   wire [0:0] stage2_15;
   wire [3:0] stage3_0;
   wire [6:0] stage3_1;
   wire [5:0] stage3_2;
   wire [1:0] stage3_3;
   wire [5:0] stage3_4;
   wire [2:0] stage3_5;
   wire [3:0] stage3_6;
   wire [5:0] stage3_7;
   wire [4:0] stage3_8;
   wire [2:0] stage3_9;
   wire [3:0] stage3_10;
   wire [5:0] stage3_11;
   wire [5:0] stage3_12;
   wire [2:0] stage3_13;
   wire [2:0] stage3_14;
   wire [1:0] stage3_15;
   wire [0:0] stage3_16;
   wire [1:0] stage4_0;
   wire [1:0] stage4_1;
   wire [1:0] stage4_2;
   wire [1:0] stage4_3;
   wire [1:0] stage4_4;
   wire [1:0] stage4_5;
   wire [1:0] stage4_6;
   wire [1:0] stage4_7;
   wire [1:0] stage4_8;
   wire [1:0] stage4_9;
   wire [1:0] stage4_10;
   wire [1:0] stage4_11;
   wire [1:0] stage4_12;
   wire [1:0] stage4_13;
   wire [1:0] stage4_14;
   wire [1:0] stage4_15;
   wire [1:0] stage4_16;

   assign stage0_0 = src0;
   assign stage0_1 = src1;
   assign stage0_2 = src2;
   assign stage0_3 = src3;
   assign stage0_4 = src4;
   assign stage0_5 = src5;
   assign stage0_6 = src6;
   assign stage0_7 = src7;
   assign stage0_8 = src8;
   assign stage0_9 = src9;
   assign stage0_10 = src10;
   assign stage0_11 = src11;
   assign dst0 = stage4_0;
   assign dst1 = stage4_1;
   assign dst2 = stage4_2;
   assign dst3 = stage4_3;
   assign dst4 = stage4_4;
   assign dst5 = stage4_5;
   assign dst6 = stage4_6;
   assign dst7 = stage4_7;
   assign dst8 = stage4_8;
   assign dst9 = stage4_9;
   assign dst10 = stage4_10;
   assign dst11 = stage4_11;
   assign dst12 = stage4_12;
   assign dst13 = stage4_13;
   assign dst14 = stage4_14;
   assign dst15 = stage4_15;
   assign dst16 = stage4_16;

   gpc606_5 gpc0 (
      {stage0_0[0], stage0_0[1], stage0_0[2], stage0_0[3], stage0_0[4], stage0_0[5]},
      {stage0_2[0], stage0_2[1], stage0_2[2], stage0_2[3], stage0_2[4], stage0_2[5]},
      {stage1_4[0],stage1_3[0],stage1_2[0],stage1_1[0],stage1_0[0]}
   );
   gpc606_5 gpc1 (
      {stage0_0[6], stage0_0[7], stage0_0[8], stage0_0[9], stage0_0[10], stage0_0[11]},
      {stage0_2[6], stage0_2[7], stage0_2[8], stage0_2[9], stage0_2[10], stage0_2[11]},
      {stage1_4[1],stage1_3[1],stage1_2[1],stage1_1[1],stage1_0[1]}
   );
   gpc606_5 gpc2 (
      {stage0_0[12], stage0_0[13], stage0_0[14], stage0_0[15], stage0_0[16], stage0_0[17]},
      {stage0_2[12], stage0_2[13], stage0_2[14], stage0_2[15], stage0_2[16], stage0_2[17]},
      {stage1_4[2],stage1_3[2],stage1_2[2],stage1_1[2],stage1_0[2]}
   );
   gpc606_5 gpc3 (
      {stage0_0[18], stage0_0[19], stage0_0[20], stage0_0[21], stage0_0[22], stage0_0[23]},
      {stage0_2[18], stage0_2[19], stage0_2[20], stage0_2[21], stage0_2[22], stage0_2[23]},
      {stage1_4[3],stage1_3[3],stage1_2[3],stage1_1[3],stage1_0[3]}
   );
   gpc615_5 gpc4 (
      {stage0_0[24], stage0_0[25], stage0_0[26], stage0_0[27], stage0_0[28]},
      {stage0_1[0]},
      {stage0_2[24], stage0_2[25], stage0_2[26], stage0_2[27], stage0_2[28], stage0_2[29]},
      {stage1_4[4],stage1_3[4],stage1_2[4],stage1_1[4],stage1_0[4]}
   );
   gpc615_5 gpc5 (
      {stage0_0[29], stage0_0[30], stage0_0[31], stage0_0[32], stage0_0[33]},
      {stage0_1[1]},
      {stage0_2[30], stage0_2[31], stage0_2[32], stage0_2[33], stage0_2[34], stage0_2[35]},
      {stage1_4[5],stage1_3[5],stage1_2[5],stage1_1[5],stage1_0[5]}
   );
   gpc615_5 gpc6 (
      {stage0_0[34], stage0_0[35], stage0_0[36], stage0_0[37], stage0_0[38]},
      {stage0_1[2]},
      {stage0_2[36], stage0_2[37], stage0_2[38], stage0_2[39], stage0_2[40], stage0_2[41]},
      {stage1_4[6],stage1_3[6],stage1_2[6],stage1_1[6],stage1_0[6]}
   );
   gpc615_5 gpc7 (
      {stage0_0[39], stage0_0[40], stage0_0[41], stage0_0[42], stage0_0[43]},
      {stage0_1[3]},
      {stage0_2[42], stage0_2[43], stage0_2[44], stage0_2[45], stage0_2[46], stage0_2[47]},
      {stage1_4[7],stage1_3[7],stage1_2[7],stage1_1[7],stage1_0[7]}
   );
   gpc606_5 gpc8 (
      {stage0_1[4], stage0_1[5], stage0_1[6], stage0_1[7], stage0_1[8], stage0_1[9]},
      {stage0_3[0], stage0_3[1], stage0_3[2], stage0_3[3], stage0_3[4], stage0_3[5]},
      {stage1_5[0],stage1_4[8],stage1_3[8],stage1_2[8],stage1_1[8]}
   );
   gpc606_5 gpc9 (
      {stage0_1[10], stage0_1[11], stage0_1[12], stage0_1[13], stage0_1[14], stage0_1[15]},
      {stage0_3[6], stage0_3[7], stage0_3[8], stage0_3[9], stage0_3[10], stage0_3[11]},
      {stage1_5[1],stage1_4[9],stage1_3[9],stage1_2[9],stage1_1[9]}
   );
   gpc606_5 gpc10 (
      {stage0_1[16], stage0_1[17], stage0_1[18], stage0_1[19], stage0_1[20], stage0_1[21]},
      {stage0_3[12], stage0_3[13], stage0_3[14], stage0_3[15], stage0_3[16], stage0_3[17]},
      {stage1_5[2],stage1_4[10],stage1_3[10],stage1_2[10],stage1_1[10]}
   );
   gpc606_5 gpc11 (
      {stage0_1[22], stage0_1[23], stage0_1[24], stage0_1[25], stage0_1[26], stage0_1[27]},
      {stage0_3[18], stage0_3[19], stage0_3[20], stage0_3[21], stage0_3[22], stage0_3[23]},
      {stage1_5[3],stage1_4[11],stage1_3[11],stage1_2[11],stage1_1[11]}
   );
   gpc606_5 gpc12 (
      {stage0_1[28], stage0_1[29], stage0_1[30], stage0_1[31], stage0_1[32], stage0_1[33]},
      {stage0_3[24], stage0_3[25], stage0_3[26], stage0_3[27], stage0_3[28], stage0_3[29]},
      {stage1_5[4],stage1_4[12],stage1_3[12],stage1_2[12],stage1_1[12]}
   );
   gpc606_5 gpc13 (
      {stage0_1[34], stage0_1[35], stage0_1[36], stage0_1[37], stage0_1[38], stage0_1[39]},
      {stage0_3[30], stage0_3[31], stage0_3[32], stage0_3[33], stage0_3[34], stage0_3[35]},
      {stage1_5[5],stage1_4[13],stage1_3[13],stage1_2[13],stage1_1[13]}
   );
   gpc606_5 gpc14 (
      {stage0_1[40], stage0_1[41], stage0_1[42], stage0_1[43], stage0_1[44], stage0_1[45]},
      {stage0_3[36], stage0_3[37], stage0_3[38], stage0_3[39], stage0_3[40], stage0_3[41]},
      {stage1_5[6],stage1_4[14],stage1_3[14],stage1_2[14],stage1_1[14]}
   );
   gpc606_5 gpc15 (
      {stage0_1[46], stage0_1[47], stage0_1[48], stage0_1[49], stage0_1[50], stage0_1[51]},
      {stage0_3[42], stage0_3[43], stage0_3[44], stage0_3[45], stage0_3[46], stage0_3[47]},
      {stage1_5[7],stage1_4[15],stage1_3[15],stage1_2[15],stage1_1[15]}
   );
   gpc615_5 gpc16 (
      {stage0_2[48], stage0_2[49], stage0_2[50], stage0_2[51], stage0_2[52]},
      {stage0_3[48]},
      {stage0_4[0], stage0_4[1], stage0_4[2], stage0_4[3], stage0_4[4], stage0_4[5]},
      {stage1_6[0],stage1_5[8],stage1_4[16],stage1_3[16],stage1_2[16]}
   );
   gpc615_5 gpc17 (
      {stage0_3[49], stage0_3[50], stage0_3[51], stage0_3[52], stage0_3[53]},
      {stage0_4[6]},
      {stage0_5[0], stage0_5[1], stage0_5[2], stage0_5[3], stage0_5[4], stage0_5[5]},
      {stage1_7[0],stage1_6[1],stage1_5[9],stage1_4[17],stage1_3[17]}
   );
   gpc606_5 gpc18 (
      {stage0_4[7], stage0_4[8], stage0_4[9], stage0_4[10], stage0_4[11], stage0_4[12]},
      {stage0_6[0], stage0_6[1], stage0_6[2], stage0_6[3], stage0_6[4], stage0_6[5]},
      {stage1_8[0],stage1_7[1],stage1_6[2],stage1_5[10],stage1_4[18]}
   );
   gpc606_5 gpc19 (
      {stage0_4[13], stage0_4[14], stage0_4[15], stage0_4[16], stage0_4[17], stage0_4[18]},
      {stage0_6[6], stage0_6[7], stage0_6[8], stage0_6[9], stage0_6[10], stage0_6[11]},
      {stage1_8[1],stage1_7[2],stage1_6[3],stage1_5[11],stage1_4[19]}
   );
   gpc606_5 gpc20 (
      {stage0_4[19], stage0_4[20], stage0_4[21], stage0_4[22], stage0_4[23], stage0_4[24]},
      {stage0_6[12], stage0_6[13], stage0_6[14], stage0_6[15], stage0_6[16], stage0_6[17]},
      {stage1_8[2],stage1_7[3],stage1_6[4],stage1_5[12],stage1_4[20]}
   );
   gpc606_5 gpc21 (
      {stage0_4[25], stage0_4[26], stage0_4[27], stage0_4[28], stage0_4[29], stage0_4[30]},
      {stage0_6[18], stage0_6[19], stage0_6[20], stage0_6[21], stage0_6[22], stage0_6[23]},
      {stage1_8[3],stage1_7[4],stage1_6[5],stage1_5[13],stage1_4[21]}
   );
   gpc606_5 gpc22 (
      {stage0_4[31], stage0_4[32], stage0_4[33], stage0_4[34], stage0_4[35], stage0_4[36]},
      {stage0_6[24], stage0_6[25], stage0_6[26], stage0_6[27], stage0_6[28], stage0_6[29]},
      {stage1_8[4],stage1_7[5],stage1_6[6],stage1_5[14],stage1_4[22]}
   );
   gpc606_5 gpc23 (
      {stage0_4[37], stage0_4[38], stage0_4[39], stage0_4[40], stage0_4[41], stage0_4[42]},
      {stage0_6[30], stage0_6[31], stage0_6[32], stage0_6[33], stage0_6[34], stage0_6[35]},
      {stage1_8[5],stage1_7[6],stage1_6[7],stage1_5[15],stage1_4[23]}
   );
   gpc606_5 gpc24 (
      {stage0_4[43], stage0_4[44], stage0_4[45], stage0_4[46], stage0_4[47], stage0_4[48]},
      {stage0_6[36], stage0_6[37], stage0_6[38], stage0_6[39], stage0_6[40], stage0_6[41]},
      {stage1_8[6],stage1_7[7],stage1_6[8],stage1_5[16],stage1_4[24]}
   );
   gpc615_5 gpc25 (
      {stage0_4[49], stage0_4[50], stage0_4[51], stage0_4[52], stage0_4[53]},
      {stage0_5[6]},
      {stage0_6[42], stage0_6[43], stage0_6[44], stage0_6[45], stage0_6[46], stage0_6[47]},
      {stage1_8[7],stage1_7[8],stage1_6[9],stage1_5[17],stage1_4[25]}
   );
   gpc606_5 gpc26 (
      {stage0_5[7], stage0_5[8], stage0_5[9], stage0_5[10], stage0_5[11], stage0_5[12]},
      {stage0_7[0], stage0_7[1], stage0_7[2], stage0_7[3], stage0_7[4], stage0_7[5]},
      {stage1_9[0],stage1_8[8],stage1_7[9],stage1_6[10],stage1_5[18]}
   );
   gpc606_5 gpc27 (
      {stage0_5[13], stage0_5[14], stage0_5[15], stage0_5[16], stage0_5[17], stage0_5[18]},
      {stage0_7[6], stage0_7[7], stage0_7[8], stage0_7[9], stage0_7[10], stage0_7[11]},
      {stage1_9[1],stage1_8[9],stage1_7[10],stage1_6[11],stage1_5[19]}
   );
   gpc606_5 gpc28 (
      {stage0_5[19], stage0_5[20], stage0_5[21], stage0_5[22], stage0_5[23], stage0_5[24]},
      {stage0_7[12], stage0_7[13], stage0_7[14], stage0_7[15], stage0_7[16], stage0_7[17]},
      {stage1_9[2],stage1_8[10],stage1_7[11],stage1_6[12],stage1_5[20]}
   );
   gpc615_5 gpc29 (
      {stage0_5[25], stage0_5[26], stage0_5[27], stage0_5[28], stage0_5[29]},
      {stage0_6[48]},
      {stage0_7[18], stage0_7[19], stage0_7[20], stage0_7[21], stage0_7[22], stage0_7[23]},
      {stage1_9[3],stage1_8[11],stage1_7[12],stage1_6[13],stage1_5[21]}
   );
   gpc615_5 gpc30 (
      {stage0_5[30], stage0_5[31], stage0_5[32], stage0_5[33], stage0_5[34]},
      {stage0_6[49]},
      {stage0_7[24], stage0_7[25], stage0_7[26], stage0_7[27], stage0_7[28], stage0_7[29]},
      {stage1_9[4],stage1_8[12],stage1_7[13],stage1_6[14],stage1_5[22]}
   );
   gpc615_5 gpc31 (
      {stage0_5[35], stage0_5[36], stage0_5[37], stage0_5[38], stage0_5[39]},
      {stage0_6[50]},
      {stage0_7[30], stage0_7[31], stage0_7[32], stage0_7[33], stage0_7[34], stage0_7[35]},
      {stage1_9[5],stage1_8[13],stage1_7[14],stage1_6[15],stage1_5[23]}
   );
   gpc615_5 gpc32 (
      {stage0_5[40], stage0_5[41], stage0_5[42], stage0_5[43], stage0_5[44]},
      {stage0_6[51]},
      {stage0_7[36], stage0_7[37], stage0_7[38], stage0_7[39], stage0_7[40], stage0_7[41]},
      {stage1_9[6],stage1_8[14],stage1_7[15],stage1_6[16],stage1_5[24]}
   );
   gpc615_5 gpc33 (
      {stage0_5[45], stage0_5[46], stage0_5[47], stage0_5[48], stage0_5[49]},
      {stage0_6[52]},
      {stage0_7[42], stage0_7[43], stage0_7[44], stage0_7[45], stage0_7[46], stage0_7[47]},
      {stage1_9[7],stage1_8[15],stage1_7[16],stage1_6[17],stage1_5[25]}
   );
   gpc606_5 gpc34 (
      {stage0_7[48], stage0_7[49], stage0_7[50], stage0_7[51], stage0_7[52], stage0_7[53]},
      {stage0_9[0], stage0_9[1], stage0_9[2], stage0_9[3], stage0_9[4], stage0_9[5]},
      {stage1_11[0],stage1_10[0],stage1_9[8],stage1_8[16],stage1_7[17]}
   );
   gpc2135_5 gpc35 (
      {stage0_8[0], stage0_8[1], stage0_8[2], stage0_8[3], stage0_8[4]},
      {stage0_9[6], stage0_9[7], stage0_9[8]},
      {stage0_10[0]},
      {stage0_11[0], stage0_11[1]},
      {stage1_12[0],stage1_11[1],stage1_10[1],stage1_9[9],stage1_8[17]}
   );
   gpc2135_5 gpc36 (
      {stage0_8[5], stage0_8[6], stage0_8[7], stage0_8[8], stage0_8[9]},
      {stage0_9[9], stage0_9[10], stage0_9[11]},
      {stage0_10[1]},
      {stage0_11[2], stage0_11[3]},
      {stage1_12[1],stage1_11[2],stage1_10[2],stage1_9[10],stage1_8[18]}
   );
   gpc1406_5 gpc37 (
      {stage0_8[10], stage0_8[11], stage0_8[12], stage0_8[13], stage0_8[14], stage0_8[15]},
      {stage0_10[2], stage0_10[3], stage0_10[4], stage0_10[5]},
      {stage0_11[4]},
      {stage1_12[2],stage1_11[3],stage1_10[3],stage1_9[11],stage1_8[19]}
   );
   gpc606_5 gpc38 (
      {stage0_8[16], stage0_8[17], stage0_8[18], stage0_8[19], stage0_8[20], stage0_8[21]},
      {stage0_10[6], stage0_10[7], stage0_10[8], stage0_10[9], stage0_10[10], stage0_10[11]},
      {stage1_12[3],stage1_11[4],stage1_10[4],stage1_9[12],stage1_8[20]}
   );
   gpc606_5 gpc39 (
      {stage0_8[22], stage0_8[23], stage0_8[24], stage0_8[25], stage0_8[26], stage0_8[27]},
      {stage0_10[12], stage0_10[13], stage0_10[14], stage0_10[15], stage0_10[16], stage0_10[17]},
      {stage1_12[4],stage1_11[5],stage1_10[5],stage1_9[13],stage1_8[21]}
   );
   gpc606_5 gpc40 (
      {stage0_8[28], stage0_8[29], stage0_8[30], stage0_8[31], stage0_8[32], stage0_8[33]},
      {stage0_10[18], stage0_10[19], stage0_10[20], stage0_10[21], stage0_10[22], stage0_10[23]},
      {stage1_12[5],stage1_11[6],stage1_10[6],stage1_9[14],stage1_8[22]}
   );
   gpc615_5 gpc41 (
      {stage0_8[34], stage0_8[35], stage0_8[36], stage0_8[37], stage0_8[38]},
      {stage0_9[12]},
      {stage0_10[24], stage0_10[25], stage0_10[26], stage0_10[27], stage0_10[28], stage0_10[29]},
      {stage1_12[6],stage1_11[7],stage1_10[7],stage1_9[15],stage1_8[23]}
   );
   gpc615_5 gpc42 (
      {stage0_8[39], stage0_8[40], stage0_8[41], stage0_8[42], stage0_8[43]},
      {stage0_9[13]},
      {stage0_10[30], stage0_10[31], stage0_10[32], stage0_10[33], stage0_10[34], stage0_10[35]},
      {stage1_12[7],stage1_11[8],stage1_10[8],stage1_9[16],stage1_8[24]}
   );
   gpc615_5 gpc43 (
      {stage0_8[44], stage0_8[45], stage0_8[46], stage0_8[47], stage0_8[48]},
      {stage0_9[14]},
      {stage0_10[36], stage0_10[37], stage0_10[38], stage0_10[39], stage0_10[40], stage0_10[41]},
      {stage1_12[8],stage1_11[9],stage1_10[9],stage1_9[17],stage1_8[25]}
   );
   gpc615_5 gpc44 (
      {stage0_8[49], stage0_8[50], stage0_8[51], stage0_8[52], stage0_8[53]},
      {stage0_9[15]},
      {stage0_10[42], stage0_10[43], stage0_10[44], stage0_10[45], stage0_10[46], stage0_10[47]},
      {stage1_12[9],stage1_11[10],stage1_10[10],stage1_9[18],stage1_8[26]}
   );
   gpc606_5 gpc45 (
      {stage0_9[16], stage0_9[17], stage0_9[18], stage0_9[19], stage0_9[20], stage0_9[21]},
      {stage0_11[5], stage0_11[6], stage0_11[7], stage0_11[8], stage0_11[9], stage0_11[10]},
      {stage1_13[0],stage1_12[10],stage1_11[11],stage1_10[11],stage1_9[19]}
   );
   gpc606_5 gpc46 (
      {stage0_9[22], stage0_9[23], stage0_9[24], stage0_9[25], stage0_9[26], stage0_9[27]},
      {stage0_11[11], stage0_11[12], stage0_11[13], stage0_11[14], stage0_11[15], stage0_11[16]},
      {stage1_13[1],stage1_12[11],stage1_11[12],stage1_10[12],stage1_9[20]}
   );
   gpc606_5 gpc47 (
      {stage0_9[28], stage0_9[29], stage0_9[30], stage0_9[31], stage0_9[32], stage0_9[33]},
      {stage0_11[17], stage0_11[18], stage0_11[19], stage0_11[20], stage0_11[21], stage0_11[22]},
      {stage1_13[2],stage1_12[12],stage1_11[13],stage1_10[13],stage1_9[21]}
   );
   gpc615_5 gpc48 (
      {stage0_9[34], stage0_9[35], stage0_9[36], stage0_9[37], stage0_9[38]},
      {stage0_10[48]},
      {stage0_11[23], stage0_11[24], stage0_11[25], stage0_11[26], stage0_11[27], stage0_11[28]},
      {stage1_13[3],stage1_12[13],stage1_11[14],stage1_10[14],stage1_9[22]}
   );
   gpc615_5 gpc49 (
      {stage0_9[39], stage0_9[40], stage0_9[41], stage0_9[42], stage0_9[43]},
      {stage0_10[49]},
      {stage0_11[29], stage0_11[30], stage0_11[31], stage0_11[32], stage0_11[33], stage0_11[34]},
      {stage1_13[4],stage1_12[14],stage1_11[15],stage1_10[15],stage1_9[23]}
   );
   gpc615_5 gpc50 (
      {stage0_9[44], stage0_9[45], stage0_9[46], stage0_9[47], stage0_9[48]},
      {stage0_10[50]},
      {stage0_11[35], stage0_11[36], stage0_11[37], stage0_11[38], stage0_11[39], stage0_11[40]},
      {stage1_13[5],stage1_12[15],stage1_11[16],stage1_10[16],stage1_9[24]}
   );
   gpc615_5 gpc51 (
      {stage0_9[49], stage0_9[50], stage0_9[51], stage0_9[52], stage0_9[53]},
      {stage0_10[51]},
      {stage0_11[41], stage0_11[42], stage0_11[43], stage0_11[44], stage0_11[45], stage0_11[46]},
      {stage1_13[6],stage1_12[16],stage1_11[17],stage1_10[17],stage1_9[25]}
   );
   gpc1_1 gpc52 (
      {stage0_0[44]},
      {stage1_0[8]}
   );
   gpc1_1 gpc53 (
      {stage0_0[45]},
      {stage1_0[9]}
   );
   gpc1_1 gpc54 (
      {stage0_0[46]},
      {stage1_0[10]}
   );
   gpc1_1 gpc55 (
      {stage0_0[47]},
      {stage1_0[11]}
   );
   gpc1_1 gpc56 (
      {stage0_0[48]},
      {stage1_0[12]}
   );
   gpc1_1 gpc57 (
      {stage0_0[49]},
      {stage1_0[13]}
   );
   gpc1_1 gpc58 (
      {stage0_0[50]},
      {stage1_0[14]}
   );
   gpc1_1 gpc59 (
      {stage0_0[51]},
      {stage1_0[15]}
   );
   gpc1_1 gpc60 (
      {stage0_0[52]},
      {stage1_0[16]}
   );
   gpc1_1 gpc61 (
      {stage0_0[53]},
      {stage1_0[17]}
   );
   gpc1_1 gpc62 (
      {stage0_1[52]},
      {stage1_1[16]}
   );
   gpc1_1 gpc63 (
      {stage0_1[53]},
      {stage1_1[17]}
   );
   gpc1_1 gpc64 (
      {stage0_2[53]},
      {stage1_2[17]}
   );
   gpc1_1 gpc65 (
      {stage0_5[50]},
      {stage1_5[26]}
   );
   gpc1_1 gpc66 (
      {stage0_5[51]},
      {stage1_5[27]}
   );
   gpc1_1 gpc67 (
      {stage0_5[52]},
      {stage1_5[28]}
   );
   gpc1_1 gpc68 (
      {stage0_5[53]},
      {stage1_5[29]}
   );
   gpc1_1 gpc69 (
      {stage0_6[53]},
      {stage1_6[18]}
   );
   gpc1_1 gpc70 (
      {stage0_10[52]},
      {stage1_10[18]}
   );
   gpc1_1 gpc71 (
      {stage0_10[53]},
      {stage1_10[19]}
   );
   gpc1_1 gpc72 (
      {stage0_11[47]},
      {stage1_11[18]}
   );
   gpc1_1 gpc73 (
      {stage0_11[48]},
      {stage1_11[19]}
   );
   gpc1_1 gpc74 (
      {stage0_11[49]},
      {stage1_11[20]}
   );
   gpc1_1 gpc75 (
      {stage0_11[50]},
      {stage1_11[21]}
   );
   gpc1_1 gpc76 (
      {stage0_11[51]},
      {stage1_11[22]}
   );
   gpc1_1 gpc77 (
      {stage0_11[52]},
      {stage1_11[23]}
   );
   gpc1_1 gpc78 (
      {stage0_11[53]},
      {stage1_11[24]}
   );
   gpc2135_5 gpc79 (
      {stage1_0[0], stage1_0[1], stage1_0[2], stage1_0[3], stage1_0[4]},
      {stage1_1[0], stage1_1[1], stage1_1[2]},
      {stage1_2[0]},
      {stage1_3[0], stage1_3[1]},
      {stage2_4[0],stage2_3[0],stage2_2[0],stage2_1[0],stage2_0[0]}
   );
   gpc2135_5 gpc80 (
      {stage1_0[5], stage1_0[6], stage1_0[7], stage1_0[8], stage1_0[9]},
      {stage1_1[3], stage1_1[4], stage1_1[5]},
      {stage1_2[1]},
      {stage1_3[2], stage1_3[3]},
      {stage2_4[1],stage2_3[1],stage2_2[1],stage2_1[1],stage2_0[1]}
   );
   gpc1163_5 gpc81 (
      {stage1_0[10], stage1_0[11], stage1_0[12]},
      {stage1_1[6], stage1_1[7], stage1_1[8], stage1_1[9], stage1_1[10], stage1_1[11]},
      {stage1_2[2]},
      {stage1_3[4]},
      {stage2_4[2],stage2_3[2],stage2_2[2],stage2_1[2],stage2_0[2]}
   );
   gpc615_5 gpc82 (
      {stage1_2[3], stage1_2[4], stage1_2[5], stage1_2[6], stage1_2[7]},
      {stage1_3[5]},
      {stage1_4[0], stage1_4[1], stage1_4[2], stage1_4[3], stage1_4[4], stage1_4[5]},
      {stage2_6[0],stage2_5[0],stage2_4[3],stage2_3[3],stage2_2[3]}
   );
   gpc615_5 gpc83 (
      {stage1_2[8], stage1_2[9], stage1_2[10], stage1_2[11], stage1_2[12]},
      {stage1_3[6]},
      {stage1_4[6], stage1_4[7], stage1_4[8], stage1_4[9], stage1_4[10], stage1_4[11]},
      {stage2_6[1],stage2_5[1],stage2_4[4],stage2_3[4],stage2_2[4]}
   );
   gpc615_5 gpc84 (
      {stage1_2[13], stage1_2[14], stage1_2[15], stage1_2[16], stage1_2[17]},
      {stage1_3[7]},
      {stage1_4[12], stage1_4[13], stage1_4[14], stage1_4[15], stage1_4[16], stage1_4[17]},
      {stage2_6[2],stage2_5[2],stage2_4[5],stage2_3[5],stage2_2[5]}
   );
   gpc615_5 gpc85 (
      {stage1_3[8], stage1_3[9], stage1_3[10], stage1_3[11], stage1_3[12]},
      {stage1_4[18]},
      {stage1_5[0], stage1_5[1], stage1_5[2], stage1_5[3], stage1_5[4], stage1_5[5]},
      {stage2_7[0],stage2_6[3],stage2_5[3],stage2_4[6],stage2_3[6]}
   );
   gpc615_5 gpc86 (
      {stage1_3[13], stage1_3[14], stage1_3[15], stage1_3[16], stage1_3[17]},
      {stage1_4[19]},
      {stage1_5[6], stage1_5[7], stage1_5[8], stage1_5[9], stage1_5[10], stage1_5[11]},
      {stage2_7[1],stage2_6[4],stage2_5[4],stage2_4[7],stage2_3[7]}
   );
   gpc1163_5 gpc87 (
      {stage1_4[20], stage1_4[21], stage1_4[22]},
      {stage1_5[12], stage1_5[13], stage1_5[14], stage1_5[15], stage1_5[16], stage1_5[17]},
      {stage1_6[0]},
      {stage1_7[0]},
      {stage2_8[0],stage2_7[2],stage2_6[5],stage2_5[5],stage2_4[8]}
   );
   gpc606_5 gpc88 (
      {stage1_5[18], stage1_5[19], stage1_5[20], stage1_5[21], stage1_5[22], stage1_5[23]},
      {stage1_7[1], stage1_7[2], stage1_7[3], stage1_7[4], stage1_7[5], stage1_7[6]},
      {stage2_9[0],stage2_8[1],stage2_7[3],stage2_6[6],stage2_5[6]}
   );
   gpc606_5 gpc89 (
      {stage1_5[24], stage1_5[25], stage1_5[26], stage1_5[27], stage1_5[28], stage1_5[29]},
      {stage1_7[7], stage1_7[8], stage1_7[9], stage1_7[10], stage1_7[11], stage1_7[12]},
      {stage2_9[1],stage2_8[2],stage2_7[4],stage2_6[7],stage2_5[7]}
   );
   gpc606_5 gpc90 (
      {stage1_6[1], stage1_6[2], stage1_6[3], stage1_6[4], stage1_6[5], stage1_6[6]},
      {stage1_8[0], stage1_8[1], stage1_8[2], stage1_8[3], stage1_8[4], stage1_8[5]},
      {stage2_10[0],stage2_9[2],stage2_8[3],stage2_7[5],stage2_6[8]}
   );
   gpc615_5 gpc91 (
      {stage1_6[7], stage1_6[8], stage1_6[9], stage1_6[10], stage1_6[11]},
      {stage1_7[13]},
      {stage1_8[6], stage1_8[7], stage1_8[8], stage1_8[9], stage1_8[10], stage1_8[11]},
      {stage2_10[1],stage2_9[3],stage2_8[4],stage2_7[6],stage2_6[9]}
   );
   gpc615_5 gpc92 (
      {stage1_6[12], stage1_6[13], stage1_6[14], stage1_6[15], stage1_6[16]},
      {stage1_7[14]},
      {stage1_8[12], stage1_8[13], stage1_8[14], stage1_8[15], stage1_8[16], stage1_8[17]},
      {stage2_10[2],stage2_9[4],stage2_8[5],stage2_7[7],stage2_6[10]}
   );
   gpc1163_5 gpc93 (
      {stage1_8[18], stage1_8[19], stage1_8[20]},
      {stage1_9[0], stage1_9[1], stage1_9[2], stage1_9[3], stage1_9[4], stage1_9[5]},
      {stage1_10[0]},
      {stage1_11[0]},
      {stage2_12[0],stage2_11[0],stage2_10[3],stage2_9[5],stage2_8[6]}
   );
   gpc606_5 gpc94 (
      {stage1_8[21], stage1_8[22], stage1_8[23], stage1_8[24], stage1_8[25], stage1_8[26]},
      {stage1_10[1], stage1_10[2], stage1_10[3], stage1_10[4], stage1_10[5], stage1_10[6]},
      {stage2_12[1],stage2_11[1],stage2_10[4],stage2_9[6],stage2_8[7]}
   );
   gpc606_5 gpc95 (
      {stage1_9[6], stage1_9[7], stage1_9[8], stage1_9[9], stage1_9[10], stage1_9[11]},
      {stage1_11[1], stage1_11[2], stage1_11[3], stage1_11[4], stage1_11[5], stage1_11[6]},
      {stage2_13[0],stage2_12[2],stage2_11[2],stage2_10[5],stage2_9[7]}
   );
   gpc606_5 gpc96 (
      {stage1_9[12], stage1_9[13], stage1_9[14], stage1_9[15], stage1_9[16], stage1_9[17]},
      {stage1_11[7], stage1_11[8], stage1_11[9], stage1_11[10], stage1_11[11], stage1_11[12]},
      {stage2_13[1],stage2_12[3],stage2_11[3],stage2_10[6],stage2_9[8]}
   );
   gpc606_5 gpc97 (
      {stage1_9[18], stage1_9[19], stage1_9[20], stage1_9[21], stage1_9[22], stage1_9[23]},
      {stage1_11[13], stage1_11[14], stage1_11[15], stage1_11[16], stage1_11[17], stage1_11[18]},
      {stage2_13[2],stage2_12[4],stage2_11[4],stage2_10[7],stage2_9[9]}
   );
   gpc606_5 gpc98 (
      {stage1_10[7], stage1_10[8], stage1_10[9], stage1_10[10], stage1_10[11], stage1_10[12]},
      {stage1_12[0], stage1_12[1], stage1_12[2], stage1_12[3], stage1_12[4], stage1_12[5]},
      {stage2_14[0],stage2_13[3],stage2_12[5],stage2_11[5],stage2_10[8]}
   );
   gpc606_5 gpc99 (
      {stage1_10[13], stage1_10[14], stage1_10[15], stage1_10[16], stage1_10[17], stage1_10[18]},
      {stage1_12[6], stage1_12[7], stage1_12[8], stage1_12[9], stage1_12[10], stage1_12[11]},
      {stage2_14[1],stage2_13[4],stage2_12[6],stage2_11[6],stage2_10[9]}
   );
   gpc606_5 gpc100 (
      {stage1_11[19], stage1_11[20], stage1_11[21], stage1_11[22], stage1_11[23], stage1_11[24]},
      {stage1_13[0], stage1_13[1], stage1_13[2], stage1_13[3], stage1_13[4], stage1_13[5]},
      {stage2_15[0],stage2_14[2],stage2_13[5],stage2_12[7],stage2_11[7]}
   );
   gpc1_1 gpc101 (
      {stage1_0[13]},
      {stage2_0[3]}
   );
   gpc1_1 gpc102 (
      {stage1_0[14]},
      {stage2_0[4]}
   );
   gpc1_1 gpc103 (
      {stage1_0[15]},
      {stage2_0[5]}
   );
   gpc1_1 gpc104 (
      {stage1_0[16]},
      {stage2_0[6]}
   );
   gpc1_1 gpc105 (
      {stage1_0[17]},
      {stage2_0[7]}
   );
   gpc1_1 gpc106 (
      {stage1_1[12]},
      {stage2_1[3]}
   );
   gpc1_1 gpc107 (
      {stage1_1[13]},
      {stage2_1[4]}
   );
   gpc1_1 gpc108 (
      {stage1_1[14]},
      {stage2_1[5]}
   );
   gpc1_1 gpc109 (
      {stage1_1[15]},
      {stage2_1[6]}
   );
   gpc1_1 gpc110 (
      {stage1_1[16]},
      {stage2_1[7]}
   );
   gpc1_1 gpc111 (
      {stage1_1[17]},
      {stage2_1[8]}
   );
   gpc1_1 gpc112 (
      {stage1_4[23]},
      {stage2_4[9]}
   );
   gpc1_1 gpc113 (
      {stage1_4[24]},
      {stage2_4[10]}
   );
   gpc1_1 gpc114 (
      {stage1_4[25]},
      {stage2_4[11]}
   );
   gpc1_1 gpc115 (
      {stage1_6[17]},
      {stage2_6[11]}
   );
   gpc1_1 gpc116 (
      {stage1_6[18]},
      {stage2_6[12]}
   );
   gpc1_1 gpc117 (
      {stage1_7[15]},
      {stage2_7[8]}
   );
   gpc1_1 gpc118 (
      {stage1_7[16]},
      {stage2_7[9]}
   );
   gpc1_1 gpc119 (
      {stage1_7[17]},
      {stage2_7[10]}
   );
   gpc1_1 gpc120 (
      {stage1_9[24]},
      {stage2_9[10]}
   );
   gpc1_1 gpc121 (
      {stage1_9[25]},
      {stage2_9[11]}
   );
   gpc1_1 gpc122 (
      {stage1_10[19]},
      {stage2_10[10]}
   );
   gpc1_1 gpc123 (
      {stage1_12[12]},
      {stage2_12[8]}
   );
   gpc1_1 gpc124 (
      {stage1_12[13]},
      {stage2_12[9]}
   );
   gpc1_1 gpc125 (
      {stage1_12[14]},
      {stage2_12[10]}
   );
   gpc1_1 gpc126 (
      {stage1_12[15]},
      {stage2_12[11]}
   );
   gpc1_1 gpc127 (
      {stage1_12[16]},
      {stage2_12[12]}
   );
   gpc1_1 gpc128 (
      {stage1_13[6]},
      {stage2_13[6]}
   );
   gpc2135_5 gpc129 (
      {stage2_0[0], stage2_0[1], stage2_0[2], stage2_0[3], stage2_0[4]},
      {stage2_1[0], stage2_1[1], stage2_1[2]},
      {stage2_2[0]},
      {stage2_3[0], stage2_3[1]},
      {stage3_4[0],stage3_3[0],stage3_2[0],stage3_1[0],stage3_0[0]}
   );
   gpc606_5 gpc130 (
      {stage2_3[2], stage2_3[3], stage2_3[4], stage2_3[5], stage2_3[6], stage2_3[7]},
      {stage2_5[0], stage2_5[1], stage2_5[2], stage2_5[3], stage2_5[4], stage2_5[5]},
      {stage3_7[0],stage3_6[0],stage3_5[0],stage3_4[1],stage3_3[1]}
   );
   gpc615_5 gpc131 (
      {stage2_4[0], stage2_4[1], stage2_4[2], stage2_4[3], stage2_4[4]},
      {stage2_5[6]},
      {stage2_6[0], stage2_6[1], stage2_6[2], stage2_6[3], stage2_6[4], stage2_6[5]},
      {stage3_8[0],stage3_7[1],stage3_6[1],stage3_5[1],stage3_4[2]}
   );
   gpc615_5 gpc132 (
      {stage2_4[5], stage2_4[6], stage2_4[7], stage2_4[8], stage2_4[9]},
      {stage2_5[7]},
      {stage2_6[6], stage2_6[7], stage2_6[8], stage2_6[9], stage2_6[10], stage2_6[11]},
      {stage3_8[1],stage3_7[2],stage3_6[2],stage3_5[2],stage3_4[3]}
   );
   gpc615_5 gpc133 (
      {stage2_7[0], stage2_7[1], stage2_7[2], stage2_7[3], stage2_7[4]},
      {stage2_8[0]},
      {stage2_9[0], stage2_9[1], stage2_9[2], stage2_9[3], stage2_9[4], stage2_9[5]},
      {stage3_11[0],stage3_10[0],stage3_9[0],stage3_8[2],stage3_7[3]}
   );
   gpc615_5 gpc134 (
      {stage2_7[5], stage2_7[6], stage2_7[7], stage2_7[8], stage2_7[9]},
      {stage2_8[1]},
      {stage2_9[6], stage2_9[7], stage2_9[8], stage2_9[9], stage2_9[10], stage2_9[11]},
      {stage3_11[1],stage3_10[1],stage3_9[1],stage3_8[3],stage3_7[4]}
   );
   gpc606_5 gpc135 (
      {stage2_8[2], stage2_8[3], stage2_8[4], stage2_8[5], stage2_8[6], stage2_8[7]},
      {stage2_10[0], stage2_10[1], stage2_10[2], stage2_10[3], stage2_10[4], stage2_10[5]},
      {stage3_12[0],stage3_11[2],stage3_10[2],stage3_9[2],stage3_8[4]}
   );
   gpc615_5 gpc136 (
      {stage2_10[6], stage2_10[7], stage2_10[8], stage2_10[9], stage2_10[10]},
      {stage2_11[0]},
      {stage2_12[0], stage2_12[1], stage2_12[2], stage2_12[3], stage2_12[4], stage2_12[5]},
      {stage3_14[0],stage3_13[0],stage3_12[1],stage3_11[3],stage3_10[3]}
   );
   gpc606_5 gpc137 (
      {stage2_11[1], stage2_11[2], stage2_11[3], stage2_11[4], stage2_11[5], stage2_11[6]},
      {stage2_13[0], stage2_13[1], stage2_13[2], stage2_13[3], stage2_13[4], stage2_13[5]},
      {stage3_15[0],stage3_14[1],stage3_13[1],stage3_12[2],stage3_11[4]}
   );
   gpc1325_5 gpc138 (
      {stage2_12[6], stage2_12[7], stage2_12[8], stage2_12[9], stage2_12[10]},
      {stage2_13[6], 1'b0},
      {stage2_14[0], stage2_14[1], stage2_14[2]},
      {stage2_15[0]},
      {stage3_16[0],stage3_15[1],stage3_14[2],stage3_13[2],stage3_12[3]}
   );
   gpc1_1 gpc139 (
      {stage2_0[5]},
      {stage3_0[1]}
   );
   gpc1_1 gpc140 (
      {stage2_0[6]},
      {stage3_0[2]}
   );
   gpc1_1 gpc141 (
      {stage2_0[7]},
      {stage3_0[3]}
   );
   gpc1_1 gpc142 (
      {stage2_1[3]},
      {stage3_1[1]}
   );
   gpc1_1 gpc143 (
      {stage2_1[4]},
      {stage3_1[2]}
   );
   gpc1_1 gpc144 (
      {stage2_1[5]},
      {stage3_1[3]}
   );
   gpc1_1 gpc145 (
      {stage2_1[6]},
      {stage3_1[4]}
   );
   gpc1_1 gpc146 (
      {stage2_1[7]},
      {stage3_1[5]}
   );
   gpc1_1 gpc147 (
      {stage2_1[8]},
      {stage3_1[6]}
   );
   gpc1_1 gpc148 (
      {stage2_2[1]},
      {stage3_2[1]}
   );
   gpc1_1 gpc149 (
      {stage2_2[2]},
      {stage3_2[2]}
   );
   gpc1_1 gpc150 (
      {stage2_2[3]},
      {stage3_2[3]}
   );
   gpc1_1 gpc151 (
      {stage2_2[4]},
      {stage3_2[4]}
   );
   gpc1_1 gpc152 (
      {stage2_2[5]},
      {stage3_2[5]}
   );
   gpc1_1 gpc153 (
      {stage2_4[10]},
      {stage3_4[4]}
   );
   gpc1_1 gpc154 (
      {stage2_4[11]},
      {stage3_4[5]}
   );
   gpc1_1 gpc155 (
      {stage2_6[12]},
      {stage3_6[3]}
   );
   gpc1_1 gpc156 (
      {stage2_7[10]},
      {stage3_7[5]}
   );
   gpc1_1 gpc157 (
      {stage2_11[7]},
      {stage3_11[5]}
   );
   gpc1_1 gpc158 (
      {stage2_12[11]},
      {stage3_12[4]}
   );
   gpc1_1 gpc159 (
      {stage2_12[12]},
      {stage3_12[5]}
   );
   gpc1163_5 gpc160 (
      {stage3_0[0], stage3_0[1], stage3_0[2]},
      {stage3_1[0], stage3_1[1], stage3_1[2], stage3_1[3], stage3_1[4], stage3_1[5]},
      {stage3_2[0]},
      {stage3_3[0]},
      {stage4_4[0],stage4_3[0],stage4_2[0],stage4_1[0],stage4_0[0]}
   );
   gpc615_5 gpc161 (
      {stage3_2[1], stage3_2[2], stage3_2[3], stage3_2[4], stage3_2[5]},
      {stage3_3[1]},
      {stage3_4[0], stage3_4[1], stage3_4[2], stage3_4[3], stage3_4[4], stage3_4[5]},
      {stage4_6[0],stage4_5[0],stage4_4[1],stage4_3[1],stage4_2[1]}
   );
   gpc1343_5 gpc162 (
      {stage3_5[0], stage3_5[1], stage3_5[2]},
      {stage3_6[0], stage3_6[1], stage3_6[2], stage3_6[3]},
      {stage3_7[0], stage3_7[1], stage3_7[2]},
      {stage3_8[0]},
      {stage4_9[0],stage4_8[0],stage4_7[0],stage4_6[1],stage4_5[1]}
   );
   gpc1343_5 gpc163 (
      {stage3_7[3], stage3_7[4], stage3_7[5]},
      {stage3_8[1], stage3_8[2], stage3_8[3], stage3_8[4]},
      {stage3_9[0], stage3_9[1], stage3_9[2]},
      {stage3_10[0]},
      {stage4_11[0],stage4_10[0],stage4_9[1],stage4_8[1],stage4_7[1]}
   );
   gpc1163_5 gpc164 (
      {stage3_10[1], stage3_10[2], stage3_10[3]},
      {stage3_11[0], stage3_11[1], stage3_11[2], stage3_11[3], stage3_11[4], stage3_11[5]},
      {stage3_12[0]},
      {stage3_13[0]},
      {stage4_14[0],stage4_13[0],stage4_12[0],stage4_11[1],stage4_10[1]}
   );
   gpc1325_5 gpc165 (
      {stage3_12[1], stage3_12[2], stage3_12[3], stage3_12[4], stage3_12[5]},
      {stage3_13[1], stage3_13[2]},
      {stage3_14[0], stage3_14[1], stage3_14[2]},
      {stage3_15[0]},
      {stage4_16[0],stage4_15[0],stage4_14[1],stage4_13[1],stage4_12[1]}
   );
   gpc1_1 gpc166 (
      {stage3_0[3]},
      {stage4_0[1]}
   );
   gpc1_1 gpc167 (
      {stage3_1[6]},
      {stage4_1[1]}
   );
   gpc1_1 gpc168 (
      {stage3_15[1]},
      {stage4_15[1]}
   );
   gpc1_1 gpc169 (
      {stage3_16[0]},
      {stage4_16[1]}
   );
endmodule
module rowadder2_1_17(input [16:0] src0, input [16:0] src1, output [17:0] dst0);
    wire [16:0] gene;
    wire [16:0] prop;
    wire [19:0] out;
    wire [19:0] carryout;
    LUT2 #(
        .INIT(4'h8)
    ) lut_0_gene (
        .I0(src0[0]),
        .I1(src1[0]),
        .O(gene[0])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_0_prop (
        .I0(src0[0]),
        .I1(src1[0]),
        .O(prop[0])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_1_gene (
        .I0(src0[1]),
        .I1(src1[1]),
        .O(gene[1])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_1_prop (
        .I0(src0[1]),
        .I1(src1[1]),
        .O(prop[1])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_2_gene (
        .I0(src0[2]),
        .I1(src1[2]),
        .O(gene[2])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_2_prop (
        .I0(src0[2]),
        .I1(src1[2]),
        .O(prop[2])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_3_gene (
        .I0(src0[3]),
        .I1(src1[3]),
        .O(gene[3])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_3_prop (
        .I0(src0[3]),
        .I1(src1[3]),
        .O(prop[3])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_4_gene (
        .I0(src0[4]),
        .I1(src1[4]),
        .O(gene[4])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_4_prop (
        .I0(src0[4]),
        .I1(src1[4]),
        .O(prop[4])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_5_gene (
        .I0(src0[5]),
        .I1(src1[5]),
        .O(gene[5])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_5_prop (
        .I0(src0[5]),
        .I1(src1[5]),
        .O(prop[5])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_6_gene (
        .I0(src0[6]),
        .I1(src1[6]),
        .O(gene[6])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_6_prop (
        .I0(src0[6]),
        .I1(src1[6]),
        .O(prop[6])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_7_gene (
        .I0(src0[7]),
        .I1(src1[7]),
        .O(gene[7])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_7_prop (
        .I0(src0[7]),
        .I1(src1[7]),
        .O(prop[7])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_8_gene (
        .I0(src0[8]),
        .I1(src1[8]),
        .O(gene[8])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_8_prop (
        .I0(src0[8]),
        .I1(src1[8]),
        .O(prop[8])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_9_gene (
        .I0(src0[9]),
        .I1(src1[9]),
        .O(gene[9])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_9_prop (
        .I0(src0[9]),
        .I1(src1[9]),
        .O(prop[9])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_10_gene (
        .I0(src0[10]),
        .I1(src1[10]),
        .O(gene[10])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_10_prop (
        .I0(src0[10]),
        .I1(src1[10]),
        .O(prop[10])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_11_gene (
        .I0(src0[11]),
        .I1(src1[11]),
        .O(gene[11])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_11_prop (
        .I0(src0[11]),
        .I1(src1[11]),
        .O(prop[11])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_12_gene (
        .I0(src0[12]),
        .I1(src1[12]),
        .O(gene[12])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_12_prop (
        .I0(src0[12]),
        .I1(src1[12]),
        .O(prop[12])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_13_gene (
        .I0(src0[13]),
        .I1(src1[13]),
        .O(gene[13])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_13_prop (
        .I0(src0[13]),
        .I1(src1[13]),
        .O(prop[13])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_14_gene (
        .I0(src0[14]),
        .I1(src1[14]),
        .O(gene[14])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_14_prop (
        .I0(src0[14]),
        .I1(src1[14]),
        .O(prop[14])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_15_gene (
        .I0(src0[15]),
        .I1(src1[15]),
        .O(gene[15])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_15_prop (
        .I0(src0[15]),
        .I1(src1[15]),
        .O(prop[15])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_16_gene (
        .I0(src0[16]),
        .I1(src1[16]),
        .O(gene[16])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_16_prop (
        .I0(src0[16]),
        .I1(src1[16]),
        .O(prop[16])
    );
    CARRY4 carry4_3_0 (
        .CO(carryout[3:0]),
        .O(out[3:0]),
        .CI(1'h0),
        .CYINIT(1'h0),
        .DI(gene[3:0]),
        .S(prop[3:0])
    );
    CARRY4 carry4_7_4 (
        .CO(carryout[7:4]),
        .O(out[7:4]),
        .CI(carryout[3]),
        .CYINIT(1'h0),
        .DI(gene[7:4]),
        .S(prop[7:4])
    );
    CARRY4 carry4_11_8 (
        .CO(carryout[11:8]),
        .O(out[11:8]),
        .CI(carryout[7]),
        .CYINIT(1'h0),
        .DI(gene[11:8]),
        .S(prop[11:8])
    );
    CARRY4 carry4_15_12 (
        .CO(carryout[15:12]),
        .O(out[15:12]),
        .CI(carryout[11]),
        .CYINIT(1'h0),
        .DI(gene[15:12]),
        .S(prop[15:12])
    );
    CARRY4 carry4_19_16 (
        .CO(carryout[19:16]),
        .O(out[19:16]),
        .CI(carryout[15]),
        .CYINIT(1'h0),
        .DI({3'h0, gene[16:16]}),
        .S({3'h0, prop[16:16]})
    );
    assign dst0 = {carryout[16], out[16:0]};
endmodule


module comp2_1test_54_12();
    reg [11:0] src0;
    reg [11:0] src1;
    reg [11:0] src2;
    reg [11:0] src3;
    reg [11:0] src4;
    reg [11:0] src5;
    reg [11:0] src6;
    reg [11:0] src7;
    reg [11:0] src8;
    reg [11:0] src9;
    reg [11:0] src10;
    reg [11:0] src11;
    reg [11:0] src12;
    reg [11:0] src13;
    reg [11:0] src14;
    reg [11:0] src15;
    reg [11:0] src16;
    reg [11:0] src17;
    reg [11:0] src18;
    reg [11:0] src19;
    reg [11:0] src20;
    reg [11:0] src21;
    reg [11:0] src22;
    reg [11:0] src23;
    reg [11:0] src24;
    reg [11:0] src25;
    reg [11:0] src26;
    reg [11:0] src27;
    reg [11:0] src28;
    reg [11:0] src29;
    reg [11:0] src30;
    reg [11:0] src31;
    reg [11:0] src32;
    reg [11:0] src33;
    reg [11:0] src34;
    reg [11:0] src35;
    reg [11:0] src36;
    reg [11:0] src37;
    reg [11:0] src38;
    reg [11:0] src39;
    reg [11:0] src40;
    reg [11:0] src41;
    reg [11:0] src42;
    reg [11:0] src43;
    reg [11:0] src44;
    reg [11:0] src45;
    reg [11:0] src46;
    reg [11:0] src47;
    reg [11:0] src48;
    reg [11:0] src49;
    reg [11:0] src50;
    reg [11:0] src51;
    reg [11:0] src52;
    reg [11:0] src53;
    reg [17:0] exp;
    wire [17:0] dst;
    assign test = dst == exp;
    compressor2_1_54_12 compressor2_1_54_12_inst(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .src31(src31),
        .src32(src32),
        .src33(src33),
        .src34(src34),
        .src35(src35),
        .src36(src36),
        .src37(src37),
        .src38(src38),
        .src39(src39),
        .src40(src40),
        .src41(src41),
        .src42(src42),
        .src43(src43),
        .src44(src44),
        .src45(src45),
        .src46(src46),
        .src47(src47),
        .src48(src48),
        .src49(src49),
        .src50(src50),
        .src51(src51),
        .src52(src52),
        .src53(src53),
        .dst(dst)
    );
    initial begin
        $monitor("0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x %x", src0, src1, src2, src3, src4, src5, src6, src7, src8, src9, src10, src11, src12, src13, src14, src15, src16, src17, src18, src19, src20, src21, src22, src23, src24, src25, src26, src27, src28, src29, src30, src31, src32, src33, src34, src35, src36, src37, src38, src39, src40, src41, src42, src43, src44, src45, src46, src47, src48, src49, src50, src51, src52, src53, dst, exp, test);
        src0 <= 12'h254;
        src1 <= 12'hdb7;
        src2 <= 12'h5bf;
        src3 <= 12'h401;
        src4 <= 12'h1d4;
        src5 <= 12'h3c2;
        src6 <= 12'h678;
        src7 <= 12'hdf0;
        src8 <= 12'h6e0;
        src9 <= 12'h4e4;
        src10 <= 12'h2ff;
        src11 <= 12'h39f;
        src12 <= 12'h3cc;
        src13 <= 12'h9cc;
        src14 <= 12'h2c5;
        src15 <= 12'hd3e;
        src16 <= 12'h96f;
        src17 <= 12'h608;
        src18 <= 12'ha9e;
        src19 <= 12'h681;
        src20 <= 12'hab;
        src21 <= 12'h6ba;
        src22 <= 12'hd7d;
        src23 <= 12'h418;
        src24 <= 12'hb4e;
        src25 <= 12'hd64;
        src26 <= 12'h907;
        src27 <= 12'h596;
        src28 <= 12'h55e;
        src29 <= 12'ha55;
        src30 <= 12'h9fe;
        src31 <= 12'h9c4;
        src32 <= 12'h43;
        src33 <= 12'h928;
        src34 <= 12'hae2;
        src35 <= 12'hc20;
        src36 <= 12'h97c;
        src37 <= 12'he41;
        src38 <= 12'hd63;
        src39 <= 12'he18;
        src40 <= 12'h12d;
        src41 <= 12'hf22;
        src42 <= 12'h47;
        src43 <= 12'hdb1;
        src44 <= 12'h4b4;
        src45 <= 12'h145;
        src46 <= 12'hed6;
        src47 <= 12'hf1;
        src48 <= 12'hee3;
        src49 <= 12'hc11;
        src50 <= 12'hb15;
        src51 <= 12'h40a;
        src52 <= 12'h1f1;
        src53 <= 12'h921;
        exp <= 18'h1a4eb;
        #1
        src0 <= 12'h2c0;
        src1 <= 12'h8e0;
        src2 <= 12'h148;
        src3 <= 12'haeb;
        src4 <= 12'h4d1;
        src5 <= 12'h6aa;
        src6 <= 12'hd19;
        src7 <= 12'h4bf;
        src8 <= 12'hbb6;
        src9 <= 12'h537;
        src10 <= 12'h826;
        src11 <= 12'h9bc;
        src12 <= 12'h65a;
        src13 <= 12'h6b8;
        src14 <= 12'h63c;
        src15 <= 12'h81c;
        src16 <= 12'h264;
        src17 <= 12'h216;
        src18 <= 12'h1cc;
        src19 <= 12'h991;
        src20 <= 12'h56a;
        src21 <= 12'hf76;
        src22 <= 12'hd11;
        src23 <= 12'ha55;
        src24 <= 12'hc19;
        src25 <= 12'h7b7;
        src26 <= 12'h51c;
        src27 <= 12'hbd1;
        src28 <= 12'h2a3;
        src29 <= 12'hbdf;
        src30 <= 12'h528;
        src31 <= 12'hbf;
        src32 <= 12'h5ae;
        src33 <= 12'h4f7;
        src34 <= 12'h5e0;
        src35 <= 12'ha5a;
        src36 <= 12'hbcd;
        src37 <= 12'h689;
        src38 <= 12'hdb0;
        src39 <= 12'h89e;
        src40 <= 12'h6b3;
        src41 <= 12'hb77;
        src42 <= 12'hd8f;
        src43 <= 12'hbb1;
        src44 <= 12'ha78;
        src45 <= 12'hfb;
        src46 <= 12'he1f;
        src47 <= 12'h30;
        src48 <= 12'hf3a;
        src49 <= 12'hbfb;
        src50 <= 12'h59b;
        src51 <= 12'hae1;
        src52 <= 12'h119;
        src53 <= 12'h321;
        exp <= 18'h1a13c;
        #1
        src0 <= 12'h7de;
        src1 <= 12'he94;
        src2 <= 12'h780;
        src3 <= 12'h7b0;
        src4 <= 12'h42f;
        src5 <= 12'ha7;
        src6 <= 12'h947;
        src7 <= 12'h348;
        src8 <= 12'h5c0;
        src9 <= 12'hdd2;
        src10 <= 12'h2dc;
        src11 <= 12'hd22;
        src12 <= 12'hcbb;
        src13 <= 12'hb3d;
        src14 <= 12'h14c;
        src15 <= 12'ha5;
        src16 <= 12'h477;
        src17 <= 12'h113;
        src18 <= 12'h575;
        src19 <= 12'h2df;
        src20 <= 12'h3d2;
        src21 <= 12'h718;
        src22 <= 12'hd0b;
        src23 <= 12'h122;
        src24 <= 12'hf02;
        src25 <= 12'hbe3;
        src26 <= 12'h266;
        src27 <= 12'h29a;
        src28 <= 12'hdc6;
        src29 <= 12'h808;
        src30 <= 12'h88a;
        src31 <= 12'hfa4;
        src32 <= 12'h96d;
        src33 <= 12'hd20;
        src34 <= 12'h362;
        src35 <= 12'h252;
        src36 <= 12'h625;
        src37 <= 12'h6;
        src38 <= 12'h721;
        src39 <= 12'hb35;
        src40 <= 12'h123;
        src41 <= 12'h9bd;
        src42 <= 12'h4f1;
        src43 <= 12'he90;
        src44 <= 12'h1dd;
        src45 <= 12'h2d3;
        src46 <= 12'hbd8;
        src47 <= 12'h4b6;
        src48 <= 12'h9f3;
        src49 <= 12'h4fb;
        src50 <= 12'h9c9;
        src51 <= 12'h82;
        src52 <= 12'h47b;
        src53 <= 12'h46;
        exp <= 18'h16fb1;
        #1
        src0 <= 12'h853;
        src1 <= 12'hb0c;
        src2 <= 12'hd05;
        src3 <= 12'h451;
        src4 <= 12'h8e7;
        src5 <= 12'h82a;
        src6 <= 12'h384;
        src7 <= 12'h134;
        src8 <= 12'h7e4;
        src9 <= 12'he18;
        src10 <= 12'h1d3;
        src11 <= 12'h1f0;
        src12 <= 12'h2a7;
        src13 <= 12'h3fe;
        src14 <= 12'h7ce;
        src15 <= 12'hf47;
        src16 <= 12'h5b0;
        src17 <= 12'heed;
        src18 <= 12'hd08;
        src19 <= 12'h6a7;
        src20 <= 12'h832;
        src21 <= 12'h200;
        src22 <= 12'h17c;
        src23 <= 12'h983;
        src24 <= 12'h905;
        src25 <= 12'hbc0;
        src26 <= 12'h963;
        src27 <= 12'hd6c;
        src28 <= 12'he63;
        src29 <= 12'h6db;
        src30 <= 12'hc7f;
        src31 <= 12'h140;
        src32 <= 12'had4;
        src33 <= 12'hb25;
        src34 <= 12'h7f6;
        src35 <= 12'h3b5;
        src36 <= 12'he89;
        src37 <= 12'h61d;
        src38 <= 12'h11a;
        src39 <= 12'h90b;
        src40 <= 12'h1ac;
        src41 <= 12'h4ed;
        src42 <= 12'h981;
        src43 <= 12'h51e;
        src44 <= 12'h4fa;
        src45 <= 12'h540;
        src46 <= 12'h31;
        src47 <= 12'h57;
        src48 <= 12'hfe2;
        src49 <= 12'h6f3;
        src50 <= 12'h23d;
        src51 <= 12'h42e;
        src52 <= 12'h46b;
        src53 <= 12'h1bb;
        exp <= 18'h181d4;
        #1
        src0 <= 12'haab;
        src1 <= 12'h5eb;
        src2 <= 12'h9cb;
        src3 <= 12'hbda;
        src4 <= 12'h48f;
        src5 <= 12'h554;
        src6 <= 12'h166;
        src7 <= 12'h158;
        src8 <= 12'hb0;
        src9 <= 12'hd8;
        src10 <= 12'hf13;
        src11 <= 12'h896;
        src12 <= 12'hed;
        src13 <= 12'h4d8;
        src14 <= 12'h62b;
        src15 <= 12'hf1a;
        src16 <= 12'hfe5;
        src17 <= 12'h7f;
        src18 <= 12'hcc9;
        src19 <= 12'h70a;
        src20 <= 12'h875;
        src21 <= 12'h52;
        src22 <= 12'hf6a;
        src23 <= 12'he26;
        src24 <= 12'hcc6;
        src25 <= 12'h9d7;
        src26 <= 12'hfbf;
        src27 <= 12'h695;
        src28 <= 12'h205;
        src29 <= 12'habe;
        src30 <= 12'hbb;
        src31 <= 12'h248;
        src32 <= 12'hda5;
        src33 <= 12'hb3;
        src34 <= 12'h6e6;
        src35 <= 12'hb50;
        src36 <= 12'hf5d;
        src37 <= 12'h971;
        src38 <= 12'h374;
        src39 <= 12'h5fd;
        src40 <= 12'h9d8;
        src41 <= 12'h825;
        src42 <= 12'h868;
        src43 <= 12'h64c;
        src44 <= 12'hc20;
        src45 <= 12'h56e;
        src46 <= 12'h5f9;
        src47 <= 12'h879;
        src48 <= 12'h2c0;
        src49 <= 12'ha69;
        src50 <= 12'h7ff;
        src51 <= 12'hc11;
        src52 <= 12'hcb9;
        src53 <= 12'h752;
        exp <= 18'h1a71e;
        #1
        src0 <= 12'h91;
        src1 <= 12'h6b5;
        src2 <= 12'hcac;
        src3 <= 12'ha3f;
        src4 <= 12'hc00;
        src5 <= 12'h3f5;
        src6 <= 12'h97;
        src7 <= 12'hb49;
        src8 <= 12'h87c;
        src9 <= 12'hd3d;
        src10 <= 12'h3e7;
        src11 <= 12'h330;
        src12 <= 12'he79;
        src13 <= 12'h462;
        src14 <= 12'h78d;
        src15 <= 12'h5b0;
        src16 <= 12'hb63;
        src17 <= 12'h9b6;
        src18 <= 12'h13e;
        src19 <= 12'h9a1;
        src20 <= 12'h19c;
        src21 <= 12'h540;
        src22 <= 12'hfaa;
        src23 <= 12'hb23;
        src24 <= 12'h37e;
        src25 <= 12'hfac;
        src26 <= 12'h88a;
        src27 <= 12'h425;
        src28 <= 12'h786;
        src29 <= 12'h3a7;
        src30 <= 12'h4ff;
        src31 <= 12'h8f6;
        src32 <= 12'hb84;
        src33 <= 12'h345;
        src34 <= 12'h822;
        src35 <= 12'h978;
        src36 <= 12'h4fe;
        src37 <= 12'hd15;
        src38 <= 12'h1fd;
        src39 <= 12'haa8;
        src40 <= 12'h2b6;
        src41 <= 12'h791;
        src42 <= 12'h903;
        src43 <= 12'h537;
        src44 <= 12'h4fc;
        src45 <= 12'h363;
        src46 <= 12'he55;
        src47 <= 12'h4a5;
        src48 <= 12'hb62;
        src49 <= 12'h7c0;
        src50 <= 12'haf1;
        src51 <= 12'h1a3;
        src52 <= 12'h6f5;
        src53 <= 12'hda;
        exp <= 18'h18c04;
        #1
        src0 <= 12'ha6;
        src1 <= 12'h90d;
        src2 <= 12'h2e9;
        src3 <= 12'h967;
        src4 <= 12'h659;
        src5 <= 12'he3;
        src6 <= 12'hd17;
        src7 <= 12'hc98;
        src8 <= 12'hd54;
        src9 <= 12'h383;
        src10 <= 12'hf03;
        src11 <= 12'hb2c;
        src12 <= 12'h446;
        src13 <= 12'h7fe;
        src14 <= 12'h1aa;
        src15 <= 12'hd5e;
        src16 <= 12'hf7c;
        src17 <= 12'h3b7;
        src18 <= 12'h5ee;
        src19 <= 12'haf1;
        src20 <= 12'h64a;
        src21 <= 12'h857;
        src22 <= 12'hd92;
        src23 <= 12'h7ce;
        src24 <= 12'h2c6;
        src25 <= 12'hf5c;
        src26 <= 12'hb56;
        src27 <= 12'h849;
        src28 <= 12'hb97;
        src29 <= 12'h46d;
        src30 <= 12'h895;
        src31 <= 12'ha85;
        src32 <= 12'h22;
        src33 <= 12'h37b;
        src34 <= 12'he21;
        src35 <= 12'h571;
        src36 <= 12'hb03;
        src37 <= 12'h7e3;
        src38 <= 12'h6c0;
        src39 <= 12'hba;
        src40 <= 12'h985;
        src41 <= 12'hec5;
        src42 <= 12'h624;
        src43 <= 12'h6f5;
        src44 <= 12'hff3;
        src45 <= 12'hcd9;
        src46 <= 12'hef6;
        src47 <= 12'h759;
        src48 <= 12'h5ce;
        src49 <= 12'h210;
        src50 <= 12'h68b;
        src51 <= 12'h82;
        src52 <= 12'h1d7;
        src53 <= 12'haa;
        exp <= 18'h1a9ab;
        #1
        src0 <= 12'hf83;
        src1 <= 12'hc70;
        src2 <= 12'h11a;
        src3 <= 12'h633;
        src4 <= 12'hf04;
        src5 <= 12'hee1;
        src6 <= 12'hf96;
        src7 <= 12'hf55;
        src8 <= 12'h8d8;
        src9 <= 12'hf8b;
        src10 <= 12'ha66;
        src11 <= 12'h703;
        src12 <= 12'h46d;
        src13 <= 12'h972;
        src14 <= 12'h602;
        src15 <= 12'h88d;
        src16 <= 12'hd64;
        src17 <= 12'h719;
        src18 <= 12'h949;
        src19 <= 12'h3b1;
        src20 <= 12'h538;
        src21 <= 12'hda7;
        src22 <= 12'h714;
        src23 <= 12'h8a0;
        src24 <= 12'h466;
        src25 <= 12'hea9;
        src26 <= 12'h11c;
        src27 <= 12'hb69;
        src28 <= 12'h361;
        src29 <= 12'hf5c;
        src30 <= 12'h5b8;
        src31 <= 12'hf5c;
        src32 <= 12'hbb;
        src33 <= 12'ha0b;
        src34 <= 12'h144;
        src35 <= 12'hac8;
        src36 <= 12'hc31;
        src37 <= 12'h422;
        src38 <= 12'h6e;
        src39 <= 12'h78e;
        src40 <= 12'h9c5;
        src41 <= 12'hb8a;
        src42 <= 12'h2ca;
        src43 <= 12'hc73;
        src44 <= 12'hbea;
        src45 <= 12'heee;
        src46 <= 12'h656;
        src47 <= 12'h31b;
        src48 <= 12'h78;
        src49 <= 12'he06;
        src50 <= 12'h28e;
        src51 <= 12'ha2c;
        src52 <= 12'h98;
        src53 <= 12'h7d0;
        exp <= 18'h1cd4f;
        #1
        src0 <= 12'h385;
        src1 <= 12'h226;
        src2 <= 12'hd4a;
        src3 <= 12'h82;
        src4 <= 12'h4f1;
        src5 <= 12'hf7a;
        src6 <= 12'h676;
        src7 <= 12'hae8;
        src8 <= 12'h63;
        src9 <= 12'h72d;
        src10 <= 12'h1b2;
        src11 <= 12'h17b;
        src12 <= 12'hb3a;
        src13 <= 12'hc77;
        src14 <= 12'h8f7;
        src15 <= 12'hfc4;
        src16 <= 12'ha95;
        src17 <= 12'h934;
        src18 <= 12'h88c;
        src19 <= 12'h890;
        src20 <= 12'h589;
        src21 <= 12'h52c;
        src22 <= 12'h7c9;
        src23 <= 12'hf15;
        src24 <= 12'h25c;
        src25 <= 12'h293;
        src26 <= 12'hfaa;
        src27 <= 12'hc9;
        src28 <= 12'h959;
        src29 <= 12'h275;
        src30 <= 12'hd9c;
        src31 <= 12'h57e;
        src32 <= 12'h98;
        src33 <= 12'h834;
        src34 <= 12'h557;
        src35 <= 12'h996;
        src36 <= 12'h555;
        src37 <= 12'ha9e;
        src38 <= 12'h735;
        src39 <= 12'h8f6;
        src40 <= 12'h1da;
        src41 <= 12'h1f6;
        src42 <= 12'he49;
        src43 <= 12'h5c6;
        src44 <= 12'h43d;
        src45 <= 12'h77c;
        src46 <= 12'he83;
        src47 <= 12'hf44;
        src48 <= 12'h5eb;
        src49 <= 12'hb79;
        src50 <= 12'hc90;
        src51 <= 12'h1e7;
        src52 <= 12'h799;
        src53 <= 12'h59f;
        exp <= 18'h19574;
        #1
        src0 <= 12'h53a;
        src1 <= 12'h8dd;
        src2 <= 12'h70a;
        src3 <= 12'h785;
        src4 <= 12'h9fe;
        src5 <= 12'h97a;
        src6 <= 12'h21c;
        src7 <= 12'h562;
        src8 <= 12'h66;
        src9 <= 12'h723;
        src10 <= 12'h50;
        src11 <= 12'h419;
        src12 <= 12'hca2;
        src13 <= 12'h9dc;
        src14 <= 12'h905;
        src15 <= 12'h1fc;
        src16 <= 12'h94f;
        src17 <= 12'h6f5;
        src18 <= 12'h702;
        src19 <= 12'h31;
        src20 <= 12'hf09;
        src21 <= 12'h609;
        src22 <= 12'he9d;
        src23 <= 12'h2c0;
        src24 <= 12'hd77;
        src25 <= 12'hd2b;
        src26 <= 12'h1af;
        src27 <= 12'he02;
        src28 <= 12'h2ea;
        src29 <= 12'h31c;
        src30 <= 12'he8f;
        src31 <= 12'hacc;
        src32 <= 12'h6fd;
        src33 <= 12'hd52;
        src34 <= 12'h2b2;
        src35 <= 12'h59b;
        src36 <= 12'h824;
        src37 <= 12'hb87;
        src38 <= 12'h160;
        src39 <= 12'h8a2;
        src40 <= 12'h108;
        src41 <= 12'h785;
        src42 <= 12'h547;
        src43 <= 12'h323;
        src44 <= 12'h59;
        src45 <= 12'hd19;
        src46 <= 12'h322;
        src47 <= 12'h760;
        src48 <= 12'h256;
        src49 <= 12'ha65;
        src50 <= 12'hed2;
        src51 <= 12'hf1;
        src52 <= 12'hf71;
        src53 <= 12'h720;
        exp <= 18'h182ea;
        #1
        src0 <= 12'h57d;
        src1 <= 12'h5a6;
        src2 <= 12'h641;
        src3 <= 12'h7d4;
        src4 <= 12'hac2;
        src5 <= 12'h6bf;
        src6 <= 12'hca9;
        src7 <= 12'h27a;
        src8 <= 12'hc6e;
        src9 <= 12'h32d;
        src10 <= 12'hc25;
        src11 <= 12'h7f5;
        src12 <= 12'ha82;
        src13 <= 12'he43;
        src14 <= 12'h382;
        src15 <= 12'h6a;
        src16 <= 12'h17a;
        src17 <= 12'h17b;
        src18 <= 12'ha1d;
        src19 <= 12'h6eb;
        src20 <= 12'h921;
        src21 <= 12'h34a;
        src22 <= 12'hf31;
        src23 <= 12'hbe3;
        src24 <= 12'h5e8;
        src25 <= 12'h9c1;
        src26 <= 12'h7de;
        src27 <= 12'h3b2;
        src28 <= 12'h82b;
        src29 <= 12'h778;
        src30 <= 12'h325;
        src31 <= 12'h3f9;
        src32 <= 12'h5dc;
        src33 <= 12'h5a3;
        src34 <= 12'h32c;
        src35 <= 12'h38e;
        src36 <= 12'h8ca;
        src37 <= 12'h1c2;
        src38 <= 12'h6ad;
        src39 <= 12'hc14;
        src40 <= 12'h42f;
        src41 <= 12'hdc4;
        src42 <= 12'h4c0;
        src43 <= 12'h9b2;
        src44 <= 12'h2cb;
        src45 <= 12'hb89;
        src46 <= 12'h9f9;
        src47 <= 12'h34f;
        src48 <= 12'hafa;
        src49 <= 12'h332;
        src50 <= 12'h670;
        src51 <= 12'h8cf;
        src52 <= 12'hb7;
        src53 <= 12'hdaa;
        exp <= 18'h17f0b;
        #1
        src0 <= 12'he0;
        src1 <= 12'hffa;
        src2 <= 12'h98e;
        src3 <= 12'hf61;
        src4 <= 12'h1e;
        src5 <= 12'hd52;
        src6 <= 12'hcbf;
        src7 <= 12'h700;
        src8 <= 12'h623;
        src9 <= 12'h215;
        src10 <= 12'he52;
        src11 <= 12'hdfe;
        src12 <= 12'hb67;
        src13 <= 12'ha5b;
        src14 <= 12'hecf;
        src15 <= 12'h570;
        src16 <= 12'h22a;
        src17 <= 12'h88f;
        src18 <= 12'h692;
        src19 <= 12'h87a;
        src20 <= 12'h2a3;
        src21 <= 12'h58e;
        src22 <= 12'he7a;
        src23 <= 12'hf57;
        src24 <= 12'h74a;
        src25 <= 12'he8d;
        src26 <= 12'h6cc;
        src27 <= 12'hd48;
        src28 <= 12'hf00;
        src29 <= 12'h3c;
        src30 <= 12'h28;
        src31 <= 12'he8d;
        src32 <= 12'h7f2;
        src33 <= 12'h361;
        src34 <= 12'hdcd;
        src35 <= 12'h98e;
        src36 <= 12'h8b5;
        src37 <= 12'h5f3;
        src38 <= 12'h999;
        src39 <= 12'hd93;
        src40 <= 12'hc83;
        src41 <= 12'hb39;
        src42 <= 12'hdb5;
        src43 <= 12'h14f;
        src44 <= 12'ha8f;
        src45 <= 12'ha98;
        src46 <= 12'h67f;
        src47 <= 12'hc60;
        src48 <= 12'h670;
        src49 <= 12'h12a;
        src50 <= 12'hcde;
        src51 <= 12'h7e4;
        src52 <= 12'ha12;
        src53 <= 12'h9aa;
        exp <= 18'h1e884;
        #1
        src0 <= 12'hc24;
        src1 <= 12'h635;
        src2 <= 12'hb0c;
        src3 <= 12'h6a4;
        src4 <= 12'h5ef;
        src5 <= 12'hba2;
        src6 <= 12'h11c;
        src7 <= 12'h4fc;
        src8 <= 12'h4ba;
        src9 <= 12'h39;
        src10 <= 12'h649;
        src11 <= 12'heae;
        src12 <= 12'hfd6;
        src13 <= 12'h4b3;
        src14 <= 12'h688;
        src15 <= 12'h238;
        src16 <= 12'h908;
        src17 <= 12'he9b;
        src18 <= 12'h9f1;
        src19 <= 12'h3f3;
        src20 <= 12'hc2b;
        src21 <= 12'hfc0;
        src22 <= 12'hfbe;
        src23 <= 12'h247;
        src24 <= 12'h1fa;
        src25 <= 12'h7f2;
        src26 <= 12'h7c3;
        src27 <= 12'h945;
        src28 <= 12'h2b5;
        src29 <= 12'he56;
        src30 <= 12'h57e;
        src31 <= 12'h36a;
        src32 <= 12'h27b;
        src33 <= 12'he02;
        src34 <= 12'h268;
        src35 <= 12'h57c;
        src36 <= 12'h627;
        src37 <= 12'hd91;
        src38 <= 12'hcd8;
        src39 <= 12'h749;
        src40 <= 12'h765;
        src41 <= 12'hca0;
        src42 <= 12'h123;
        src43 <= 12'haaa;
        src44 <= 12'hd29;
        src45 <= 12'hcc0;
        src46 <= 12'h680;
        src47 <= 12'hb88;
        src48 <= 12'h6e;
        src49 <= 12'hcef;
        src50 <= 12'h6af;
        src51 <= 12'h57e;
        src52 <= 12'h85;
        src53 <= 12'hb85;
        exp <= 18'h1acd4;
        #1
        src0 <= 12'h438;
        src1 <= 12'hfe3;
        src2 <= 12'h16f;
        src3 <= 12'hcf7;
        src4 <= 12'h72;
        src5 <= 12'h408;
        src6 <= 12'h40f;
        src7 <= 12'h6c;
        src8 <= 12'h22d;
        src9 <= 12'hd78;
        src10 <= 12'h97f;
        src11 <= 12'hf03;
        src12 <= 12'h76b;
        src13 <= 12'hadc;
        src14 <= 12'hec4;
        src15 <= 12'hfb0;
        src16 <= 12'h84b;
        src17 <= 12'ha50;
        src18 <= 12'h2b3;
        src19 <= 12'h1c4;
        src20 <= 12'hb19;
        src21 <= 12'h9fb;
        src22 <= 12'h79d;
        src23 <= 12'hb1f;
        src24 <= 12'h7c4;
        src25 <= 12'hbe4;
        src26 <= 12'h505;
        src27 <= 12'h507;
        src28 <= 12'h8ec;
        src29 <= 12'h47e;
        src30 <= 12'h2c4;
        src31 <= 12'hd7c;
        src32 <= 12'h562;
        src33 <= 12'h4dc;
        src34 <= 12'hd2e;
        src35 <= 12'haf5;
        src36 <= 12'ha9;
        src37 <= 12'h502;
        src38 <= 12'hfe;
        src39 <= 12'hae5;
        src40 <= 12'h32a;
        src41 <= 12'hea8;
        src42 <= 12'h998;
        src43 <= 12'h1d7;
        src44 <= 12'hda7;
        src45 <= 12'hcfe;
        src46 <= 12'h5be;
        src47 <= 12'h6d0;
        src48 <= 12'hf1c;
        src49 <= 12'hbf9;
        src50 <= 12'h8c1;
        src51 <= 12'h21e;
        src52 <= 12'ha9a;
        src53 <= 12'h71;
        exp <= 18'h1a7fa;
        #1
        src0 <= 12'h415;
        src1 <= 12'h5d3;
        src2 <= 12'hd2a;
        src3 <= 12'ha1;
        src4 <= 12'he02;
        src5 <= 12'hc91;
        src6 <= 12'h36c;
        src7 <= 12'h951;
        src8 <= 12'h513;
        src9 <= 12'h552;
        src10 <= 12'h4ad;
        src11 <= 12'h434;
        src12 <= 12'hc66;
        src13 <= 12'h292;
        src14 <= 12'h7d1;
        src15 <= 12'h37d;
        src16 <= 12'h28f;
        src17 <= 12'h1ad;
        src18 <= 12'h752;
        src19 <= 12'hd05;
        src20 <= 12'hc6;
        src21 <= 12'h53e;
        src22 <= 12'h6fd;
        src23 <= 12'hb78;
        src24 <= 12'h41a;
        src25 <= 12'hf8d;
        src26 <= 12'he57;
        src27 <= 12'h1b5;
        src28 <= 12'h91a;
        src29 <= 12'h61f;
        src30 <= 12'hd97;
        src31 <= 12'h241;
        src32 <= 12'h979;
        src33 <= 12'h9a8;
        src34 <= 12'hfaf;
        src35 <= 12'h4a3;
        src36 <= 12'hc5c;
        src37 <= 12'h6d;
        src38 <= 12'h7aa;
        src39 <= 12'hd1;
        src40 <= 12'hb49;
        src41 <= 12'h103;
        src42 <= 12'h774;
        src43 <= 12'hb30;
        src44 <= 12'ha27;
        src45 <= 12'h38b;
        src46 <= 12'h495;
        src47 <= 12'h384;
        src48 <= 12'hfcb;
        src49 <= 12'h12c;
        src50 <= 12'hf9f;
        src51 <= 12'hd95;
        src52 <= 12'h383;
        src53 <= 12'hd3a;
        exp <= 18'h190b9;
        #1
        src0 <= 12'he5;
        src1 <= 12'h86f;
        src2 <= 12'h683;
        src3 <= 12'ha40;
        src4 <= 12'h7b2;
        src5 <= 12'h35a;
        src6 <= 12'he3d;
        src7 <= 12'hdd7;
        src8 <= 12'h141;
        src9 <= 12'h1dd;
        src10 <= 12'h600;
        src11 <= 12'h2a7;
        src12 <= 12'hbfc;
        src13 <= 12'h188;
        src14 <= 12'h130;
        src15 <= 12'h32f;
        src16 <= 12'hb3a;
        src17 <= 12'h569;
        src18 <= 12'hd4;
        src19 <= 12'hf91;
        src20 <= 12'h447;
        src21 <= 12'hc4;
        src22 <= 12'ha03;
        src23 <= 12'hf83;
        src24 <= 12'h948;
        src25 <= 12'h317;
        src26 <= 12'h896;
        src27 <= 12'hd5f;
        src28 <= 12'hb5c;
        src29 <= 12'h575;
        src30 <= 12'h5c4;
        src31 <= 12'hdac;
        src32 <= 12'ha6;
        src33 <= 12'h284;
        src34 <= 12'hf79;
        src35 <= 12'h118;
        src36 <= 12'hf56;
        src37 <= 12'hb6d;
        src38 <= 12'hd19;
        src39 <= 12'h873;
        src40 <= 12'he92;
        src41 <= 12'hd9a;
        src42 <= 12'h1ca;
        src43 <= 12'hf46;
        src44 <= 12'h367;
        src45 <= 12'h4da;
        src46 <= 12'h968;
        src47 <= 12'hb85;
        src48 <= 12'h356;
        src49 <= 12'h170;
        src50 <= 12'h184;
        src51 <= 12'h4b7;
        src52 <= 12'h311;
        src53 <= 12'he4a;
        exp <= 18'h18fdd;
        #1
        src0 <= 12'hc7f;
        src1 <= 12'h32b;
        src2 <= 12'hd0d;
        src3 <= 12'h34c;
        src4 <= 12'h2ef;
        src5 <= 12'h6d;
        src6 <= 12'h178;
        src7 <= 12'h979;
        src8 <= 12'hf94;
        src9 <= 12'h3ca;
        src10 <= 12'h5b3;
        src11 <= 12'hbdc;
        src12 <= 12'h1bb;
        src13 <= 12'h85b;
        src14 <= 12'h7c8;
        src15 <= 12'hc15;
        src16 <= 12'h765;
        src17 <= 12'h654;
        src18 <= 12'hce0;
        src19 <= 12'h7a5;
        src20 <= 12'h89c;
        src21 <= 12'h23b;
        src22 <= 12'hb81;
        src23 <= 12'h5cd;
        src24 <= 12'h7f1;
        src25 <= 12'h851;
        src26 <= 12'h109;
        src27 <= 12'hc91;
        src28 <= 12'hbdd;
        src29 <= 12'h379;
        src30 <= 12'hea3;
        src31 <= 12'h83d;
        src32 <= 12'h7a8;
        src33 <= 12'hdca;
        src34 <= 12'h57f;
        src35 <= 12'h98a;
        src36 <= 12'h48c;
        src37 <= 12'h6b5;
        src38 <= 12'h72b;
        src39 <= 12'hae;
        src40 <= 12'h1c5;
        src41 <= 12'h473;
        src42 <= 12'h32b;
        src43 <= 12'h3a;
        src44 <= 12'h15;
        src45 <= 12'h549;
        src46 <= 12'h738;
        src47 <= 12'h7de;
        src48 <= 12'h504;
        src49 <= 12'h48;
        src50 <= 12'h1c5;
        src51 <= 12'h504;
        src52 <= 12'h73e;
        src53 <= 12'h22a;
        exp <= 18'h15ec8;
        #1
        src0 <= 12'h4d8;
        src1 <= 12'hbfc;
        src2 <= 12'h5e9;
        src3 <= 12'h50a;
        src4 <= 12'hc4;
        src5 <= 12'h466;
        src6 <= 12'he14;
        src7 <= 12'h321;
        src8 <= 12'he49;
        src9 <= 12'h4f5;
        src10 <= 12'h595;
        src11 <= 12'h8b8;
        src12 <= 12'hed2;
        src13 <= 12'h781;
        src14 <= 12'h4d;
        src15 <= 12'h747;
        src16 <= 12'ha26;
        src17 <= 12'hb4f;
        src18 <= 12'h6a7;
        src19 <= 12'hf3f;
        src20 <= 12'h7ab;
        src21 <= 12'h59a;
        src22 <= 12'h6f4;
        src23 <= 12'ha28;
        src24 <= 12'h44e;
        src25 <= 12'h615;
        src26 <= 12'h30c;
        src27 <= 12'hda1;
        src28 <= 12'h307;
        src29 <= 12'h9c6;
        src30 <= 12'h363;
        src31 <= 12'hfed;
        src32 <= 12'hbd3;
        src33 <= 12'h407;
        src34 <= 12'h4eb;
        src35 <= 12'hafa;
        src36 <= 12'h2bc;
        src37 <= 12'h347;
        src38 <= 12'he56;
        src39 <= 12'hb70;
        src40 <= 12'h9e7;
        src41 <= 12'h80;
        src42 <= 12'h786;
        src43 <= 12'hb59;
        src44 <= 12'hf38;
        src45 <= 12'hfb1;
        src46 <= 12'he7;
        src47 <= 12'h24f;
        src48 <= 12'hdb1;
        src49 <= 12'hf3c;
        src50 <= 12'h8d;
        src51 <= 12'h242;
        src52 <= 12'h7a4;
        src53 <= 12'hb0b;
        exp <= 18'h1a7d9;
        #1
        src0 <= 12'h613;
        src1 <= 12'hc2b;
        src2 <= 12'h27d;
        src3 <= 12'h740;
        src4 <= 12'h866;
        src5 <= 12'h65d;
        src6 <= 12'h947;
        src7 <= 12'hd1e;
        src8 <= 12'h8e3;
        src9 <= 12'hc31;
        src10 <= 12'h513;
        src11 <= 12'hd12;
        src12 <= 12'h4e6;
        src13 <= 12'h58b;
        src14 <= 12'h779;
        src15 <= 12'hbe2;
        src16 <= 12'h87a;
        src17 <= 12'h608;
        src18 <= 12'h8d4;
        src19 <= 12'hc4;
        src20 <= 12'h49;
        src21 <= 12'h3ed;
        src22 <= 12'h66f;
        src23 <= 12'h418;
        src24 <= 12'he00;
        src25 <= 12'h6f4;
        src26 <= 12'h676;
        src27 <= 12'h639;
        src28 <= 12'hc9d;
        src29 <= 12'h12f;
        src30 <= 12'h110;
        src31 <= 12'ha38;
        src32 <= 12'h6a3;
        src33 <= 12'h73a;
        src34 <= 12'h1a2;
        src35 <= 12'hfc0;
        src36 <= 12'h4ba;
        src37 <= 12'h303;
        src38 <= 12'h6ff;
        src39 <= 12'h461;
        src40 <= 12'h2cb;
        src41 <= 12'hc13;
        src42 <= 12'ha3d;
        src43 <= 12'h30b;
        src44 <= 12'h97;
        src45 <= 12'hd3f;
        src46 <= 12'h1e6;
        src47 <= 12'h452;
        src48 <= 12'hf8a;
        src49 <= 12'h1f6;
        src50 <= 12'hf01;
        src51 <= 12'h22a;
        src52 <= 12'h5e4;
        src53 <= 12'h738;
        exp <= 18'h17a0d;
        #1
        src0 <= 12'hbd;
        src1 <= 12'h7d9;
        src2 <= 12'hcaa;
        src3 <= 12'h40e;
        src4 <= 12'h1ec;
        src5 <= 12'h37d;
        src6 <= 12'h389;
        src7 <= 12'h412;
        src8 <= 12'h5dd;
        src9 <= 12'h2ee;
        src10 <= 12'h3c6;
        src11 <= 12'h91f;
        src12 <= 12'hba5;
        src13 <= 12'h5be;
        src14 <= 12'h68b;
        src15 <= 12'h33d;
        src16 <= 12'h648;
        src17 <= 12'h6a3;
        src18 <= 12'h7a6;
        src19 <= 12'hec8;
        src20 <= 12'h796;
        src21 <= 12'h335;
        src22 <= 12'hd29;
        src23 <= 12'h6e7;
        src24 <= 12'hf95;
        src25 <= 12'h72a;
        src26 <= 12'h918;
        src27 <= 12'hd5f;
        src28 <= 12'he5e;
        src29 <= 12'haa9;
        src30 <= 12'h603;
        src31 <= 12'hd3c;
        src32 <= 12'hfe6;
        src33 <= 12'hd07;
        src34 <= 12'h89d;
        src35 <= 12'h8df;
        src36 <= 12'h79c;
        src37 <= 12'h75d;
        src38 <= 12'h554;
        src39 <= 12'hfce;
        src40 <= 12'hb7e;
        src41 <= 12'he05;
        src42 <= 12'he62;
        src43 <= 12'h79d;
        src44 <= 12'h12a;
        src45 <= 12'h36b;
        src46 <= 12'h234;
        src47 <= 12'h7e9;
        src48 <= 12'h6b;
        src49 <= 12'h223;
        src50 <= 12'h24d;
        src51 <= 12'ha2d;
        src52 <= 12'h56a;
        src53 <= 12'hf44;
        exp <= 18'h1a74b;
        #1
        src0 <= 12'hf71;
        src1 <= 12'hd1;
        src2 <= 12'h70e;
        src3 <= 12'h717;
        src4 <= 12'h367;
        src5 <= 12'hab2;
        src6 <= 12'hbed;
        src7 <= 12'h6db;
        src8 <= 12'hff3;
        src9 <= 12'hf3d;
        src10 <= 12'haeb;
        src11 <= 12'h94c;
        src12 <= 12'hcdc;
        src13 <= 12'hee3;
        src14 <= 12'h6b7;
        src15 <= 12'h92a;
        src16 <= 12'hafc;
        src17 <= 12'h4aa;
        src18 <= 12'h53f;
        src19 <= 12'h2f1;
        src20 <= 12'h891;
        src21 <= 12'hf6f;
        src22 <= 12'h1fe;
        src23 <= 12'h95b;
        src24 <= 12'hfe9;
        src25 <= 12'h793;
        src26 <= 12'hb40;
        src27 <= 12'h994;
        src28 <= 12'hfbf;
        src29 <= 12'h9c2;
        src30 <= 12'ha76;
        src31 <= 12'he26;
        src32 <= 12'h401;
        src33 <= 12'h231;
        src34 <= 12'hebf;
        src35 <= 12'ha1f;
        src36 <= 12'hc8e;
        src37 <= 12'hb7;
        src38 <= 12'he1c;
        src39 <= 12'hc4c;
        src40 <= 12'h28f;
        src41 <= 12'h2ed;
        src42 <= 12'h27c;
        src43 <= 12'h7d7;
        src44 <= 12'h30f;
        src45 <= 12'h21d;
        src46 <= 12'h52e;
        src47 <= 12'h488;
        src48 <= 12'h6d5;
        src49 <= 12'hbcc;
        src50 <= 12'h286;
        src51 <= 12'h8a2;
        src52 <= 12'ha97;
        src53 <= 12'h16;
        exp <= 18'h1c5cf;
        #1
        src0 <= 12'hbf8;
        src1 <= 12'h467;
        src2 <= 12'hd79;
        src3 <= 12'h113;
        src4 <= 12'hf7e;
        src5 <= 12'hb3a;
        src6 <= 12'h19d;
        src7 <= 12'h49c;
        src8 <= 12'h13b;
        src9 <= 12'h31d;
        src10 <= 12'h654;
        src11 <= 12'h31c;
        src12 <= 12'h10f;
        src13 <= 12'h759;
        src14 <= 12'hb44;
        src15 <= 12'hb33;
        src16 <= 12'h821;
        src17 <= 12'h5a6;
        src18 <= 12'h59e;
        src19 <= 12'hbe2;
        src20 <= 12'h1d1;
        src21 <= 12'h1dd;
        src22 <= 12'h512;
        src23 <= 12'h41e;
        src24 <= 12'hf97;
        src25 <= 12'h949;
        src26 <= 12'h6f7;
        src27 <= 12'ha60;
        src28 <= 12'hab3;
        src29 <= 12'h571;
        src30 <= 12'h531;
        src31 <= 12'h780;
        src32 <= 12'h5d7;
        src33 <= 12'hbc5;
        src34 <= 12'h487;
        src35 <= 12'hb8d;
        src36 <= 12'h317;
        src37 <= 12'hb50;
        src38 <= 12'hc32;
        src39 <= 12'hc59;
        src40 <= 12'h3de;
        src41 <= 12'h94b;
        src42 <= 12'h5e0;
        src43 <= 12'h83a;
        src44 <= 12'h3e5;
        src45 <= 12'h30d;
        src46 <= 12'hf2e;
        src47 <= 12'h2e3;
        src48 <= 12'heca;
        src49 <= 12'hd45;
        src50 <= 12'ha8;
        src51 <= 12'h4ae;
        src52 <= 12'h37;
        src53 <= 12'h15f;
        exp <= 18'h17f97;
        #1
        src0 <= 12'ha7a;
        src1 <= 12'ha4b;
        src2 <= 12'h834;
        src3 <= 12'h415;
        src4 <= 12'h35c;
        src5 <= 12'h63c;
        src6 <= 12'h62f;
        src7 <= 12'hb2d;
        src8 <= 12'h155;
        src9 <= 12'h515;
        src10 <= 12'h78c;
        src11 <= 12'hbb0;
        src12 <= 12'h7e1;
        src13 <= 12'hb47;
        src14 <= 12'h2c2;
        src15 <= 12'hac8;
        src16 <= 12'h18;
        src17 <= 12'hc4f;
        src18 <= 12'h405;
        src19 <= 12'h755;
        src20 <= 12'h2f8;
        src21 <= 12'h5f3;
        src22 <= 12'h1fa;
        src23 <= 12'h204;
        src24 <= 12'h397;
        src25 <= 12'hc09;
        src26 <= 12'h96a;
        src27 <= 12'h2a6;
        src28 <= 12'h90a;
        src29 <= 12'hd02;
        src30 <= 12'h5fa;
        src31 <= 12'h8a0;
        src32 <= 12'h1bd;
        src33 <= 12'h1cb;
        src34 <= 12'hb35;
        src35 <= 12'h697;
        src36 <= 12'h702;
        src37 <= 12'h8a2;
        src38 <= 12'h391;
        src39 <= 12'h5b;
        src40 <= 12'had2;
        src41 <= 12'hf7c;
        src42 <= 12'h3c6;
        src43 <= 12'h1bb;
        src44 <= 12'h54b;
        src45 <= 12'h30f;
        src46 <= 12'h3f1;
        src47 <= 12'hcb4;
        src48 <= 12'hbe5;
        src49 <= 12'hbac;
        src50 <= 12'hbf6;
        src51 <= 12'h97b;
        src52 <= 12'haeb;
        src53 <= 12'h3e9;
        exp <= 18'h178e2;
        #1
        src0 <= 12'h44e;
        src1 <= 12'hcb3;
        src2 <= 12'h2d5;
        src3 <= 12'hb1;
        src4 <= 12'h849;
        src5 <= 12'hb7e;
        src6 <= 12'h1fd;
        src7 <= 12'hace;
        src8 <= 12'ha88;
        src9 <= 12'h5f8;
        src10 <= 12'h39b;
        src11 <= 12'h6ff;
        src12 <= 12'h6a1;
        src13 <= 12'hef7;
        src14 <= 12'had2;
        src15 <= 12'hdfc;
        src16 <= 12'he9a;
        src17 <= 12'h1ee;
        src18 <= 12'h4c5;
        src19 <= 12'hacb;
        src20 <= 12'h482;
        src21 <= 12'h600;
        src22 <= 12'hd34;
        src23 <= 12'h38b;
        src24 <= 12'h82f;
        src25 <= 12'h1a7;
        src26 <= 12'hb8b;
        src27 <= 12'hfce;
        src28 <= 12'h671;
        src29 <= 12'ha04;
        src30 <= 12'h7f;
        src31 <= 12'h199;
        src32 <= 12'hf2;
        src33 <= 12'h24c;
        src34 <= 12'h9ee;
        src35 <= 12'h3bd;
        src36 <= 12'h87d;
        src37 <= 12'h47a;
        src38 <= 12'h1e0;
        src39 <= 12'h2cb;
        src40 <= 12'h1a1;
        src41 <= 12'hb4c;
        src42 <= 12'h1ed;
        src43 <= 12'h734;
        src44 <= 12'h854;
        src45 <= 12'hd99;
        src46 <= 12'he67;
        src47 <= 12'h84;
        src48 <= 12'h4b2;
        src49 <= 12'hf2a;
        src50 <= 12'h33;
        src51 <= 12'h3f2;
        src52 <= 12'hcad;
        src53 <= 12'h17d;
        exp <= 18'h1754a;
        #1
        src0 <= 12'h6da;
        src1 <= 12'h1c7;
        src2 <= 12'h963;
        src3 <= 12'h248;
        src4 <= 12'hb8;
        src5 <= 12'h621;
        src6 <= 12'he10;
        src7 <= 12'hbbe;
        src8 <= 12'h7ca;
        src9 <= 12'h554;
        src10 <= 12'h255;
        src11 <= 12'hc60;
        src12 <= 12'h921;
        src13 <= 12'h63e;
        src14 <= 12'h9f9;
        src15 <= 12'h7cf;
        src16 <= 12'h1a0;
        src17 <= 12'h6e9;
        src18 <= 12'h4ff;
        src19 <= 12'hc1;
        src20 <= 12'h8a3;
        src21 <= 12'hb2f;
        src22 <= 12'h8b0;
        src23 <= 12'h415;
        src24 <= 12'h96e;
        src25 <= 12'h1c6;
        src26 <= 12'h163;
        src27 <= 12'h15b;
        src28 <= 12'hd38;
        src29 <= 12'h78f;
        src30 <= 12'hb3a;
        src31 <= 12'h3c4;
        src32 <= 12'h573;
        src33 <= 12'h280;
        src34 <= 12'hd1e;
        src35 <= 12'h37f;
        src36 <= 12'hf78;
        src37 <= 12'hd35;
        src38 <= 12'h894;
        src39 <= 12'h246;
        src40 <= 12'h3ac;
        src41 <= 12'h148;
        src42 <= 12'h135;
        src43 <= 12'h70a;
        src44 <= 12'h2eb;
        src45 <= 12'hb85;
        src46 <= 12'h29b;
        src47 <= 12'hbb6;
        src48 <= 12'h7f3;
        src49 <= 12'h994;
        src50 <= 12'hb9c;
        src51 <= 12'h712;
        src52 <= 12'h596;
        src53 <= 12'h8c4;
        exp <= 18'h16f1e;
        #1
        src0 <= 12'hb73;
        src1 <= 12'hf60;
        src2 <= 12'h3b8;
        src3 <= 12'h32e;
        src4 <= 12'hb38;
        src5 <= 12'h5ac;
        src6 <= 12'h31b;
        src7 <= 12'hbe6;
        src8 <= 12'h4a1;
        src9 <= 12'h548;
        src10 <= 12'hd52;
        src11 <= 12'h227;
        src12 <= 12'h140;
        src13 <= 12'h202;
        src14 <= 12'heaf;
        src15 <= 12'hed9;
        src16 <= 12'h9cb;
        src17 <= 12'he0a;
        src18 <= 12'hc6f;
        src19 <= 12'h8d9;
        src20 <= 12'hd90;
        src21 <= 12'h6ba;
        src22 <= 12'h711;
        src23 <= 12'h1dc;
        src24 <= 12'h16f;
        src25 <= 12'h19c;
        src26 <= 12'ha73;
        src27 <= 12'h9b8;
        src28 <= 12'h620;
        src29 <= 12'h737;
        src30 <= 12'h250;
        src31 <= 12'hb12;
        src32 <= 12'hefc;
        src33 <= 12'ha94;
        src34 <= 12'h132;
        src35 <= 12'h6ac;
        src36 <= 12'h289;
        src37 <= 12'h35e;
        src38 <= 12'hd2f;
        src39 <= 12'hf03;
        src40 <= 12'h273;
        src41 <= 12'h268;
        src42 <= 12'h8c0;
        src43 <= 12'h3eb;
        src44 <= 12'hecc;
        src45 <= 12'h708;
        src46 <= 12'h96b;
        src47 <= 12'hbb6;
        src48 <= 12'hd25;
        src49 <= 12'hbbb;
        src50 <= 12'hac3;
        src51 <= 12'h3d;
        src52 <= 12'h689;
        src53 <= 12'hc06;
        exp <= 18'h1ae7e;
        #1
        src0 <= 12'h34;
        src1 <= 12'h7fc;
        src2 <= 12'he3b;
        src3 <= 12'hcbf;
        src4 <= 12'h68e;
        src5 <= 12'h12b;
        src6 <= 12'h838;
        src7 <= 12'h126;
        src8 <= 12'h5fd;
        src9 <= 12'hdcd;
        src10 <= 12'hff3;
        src11 <= 12'h60e;
        src12 <= 12'h2b3;
        src13 <= 12'hb6d;
        src14 <= 12'hcac;
        src15 <= 12'ha97;
        src16 <= 12'h2c3;
        src17 <= 12'hd0b;
        src18 <= 12'h63f;
        src19 <= 12'hea5;
        src20 <= 12'hff0;
        src21 <= 12'hb88;
        src22 <= 12'h77b;
        src23 <= 12'h41e;
        src24 <= 12'h3db;
        src25 <= 12'hcb6;
        src26 <= 12'h22f;
        src27 <= 12'h8f;
        src28 <= 12'h8b8;
        src29 <= 12'h304;
        src30 <= 12'hbb8;
        src31 <= 12'h725;
        src32 <= 12'hc35;
        src33 <= 12'h25b;
        src34 <= 12'h67;
        src35 <= 12'hab8;
        src36 <= 12'hab5;
        src37 <= 12'hfb5;
        src38 <= 12'hdb1;
        src39 <= 12'hd7b;
        src40 <= 12'hc9c;
        src41 <= 12'h166;
        src42 <= 12'h387;
        src43 <= 12'h8b;
        src44 <= 12'h129;
        src45 <= 12'h43b;
        src46 <= 12'hfb5;
        src47 <= 12'h192;
        src48 <= 12'h90b;
        src49 <= 12'h9f3;
        src50 <= 12'h153;
        src51 <= 12'hb6f;
        src52 <= 12'h8ce;
        src53 <= 12'haa0;
        exp <= 18'h1ac4c;
        #1
        src0 <= 12'h5c5;
        src1 <= 12'he09;
        src2 <= 12'h56e;
        src3 <= 12'h14e;
        src4 <= 12'h8cc;
        src5 <= 12'hf5d;
        src6 <= 12'h704;
        src7 <= 12'hd6c;
        src8 <= 12'h162;
        src9 <= 12'h13b;
        src10 <= 12'h87a;
        src11 <= 12'h5ec;
        src12 <= 12'hf56;
        src13 <= 12'h2d1;
        src14 <= 12'hba0;
        src15 <= 12'he1f;
        src16 <= 12'h823;
        src17 <= 12'hfd1;
        src18 <= 12'hc34;
        src19 <= 12'h295;
        src20 <= 12'h71c;
        src21 <= 12'hd5f;
        src22 <= 12'had4;
        src23 <= 12'ha5f;
        src24 <= 12'hd79;
        src25 <= 12'h428;
        src26 <= 12'he49;
        src27 <= 12'hb39;
        src28 <= 12'h577;
        src29 <= 12'hea3;
        src30 <= 12'hd28;
        src31 <= 12'h155;
        src32 <= 12'h9e2;
        src33 <= 12'h948;
        src34 <= 12'h67f;
        src35 <= 12'had2;
        src36 <= 12'h336;
        src37 <= 12'h251;
        src38 <= 12'hdb4;
        src39 <= 12'ha38;
        src40 <= 12'h17b;
        src41 <= 12'hbd9;
        src42 <= 12'ha9d;
        src43 <= 12'he79;
        src44 <= 12'h164;
        src45 <= 12'h992;
        src46 <= 12'hedf;
        src47 <= 12'h1ad;
        src48 <= 12'h655;
        src49 <= 12'h1db;
        src50 <= 12'hd86;
        src51 <= 12'hd63;
        src52 <= 12'hd1d;
        src53 <= 12'h6d0;
        exp <= 18'h1dd11;
        #1
        src0 <= 12'h1e;
        src1 <= 12'h752;
        src2 <= 12'h52a;
        src3 <= 12'h253;
        src4 <= 12'h2ea;
        src5 <= 12'h3bf;
        src6 <= 12'hacf;
        src7 <= 12'hb5c;
        src8 <= 12'hd4f;
        src9 <= 12'hd33;
        src10 <= 12'h826;
        src11 <= 12'h50b;
        src12 <= 12'hcc;
        src13 <= 12'h80e;
        src14 <= 12'h45e;
        src15 <= 12'h18e;
        src16 <= 12'h6dd;
        src17 <= 12'h5a;
        src18 <= 12'hd17;
        src19 <= 12'hf3;
        src20 <= 12'hcd5;
        src21 <= 12'hc40;
        src22 <= 12'ha52;
        src23 <= 12'h190;
        src24 <= 12'h1bd;
        src25 <= 12'h9d1;
        src26 <= 12'h3ef;
        src27 <= 12'h400;
        src28 <= 12'h3d6;
        src29 <= 12'h453;
        src30 <= 12'hc66;
        src31 <= 12'h27;
        src32 <= 12'h632;
        src33 <= 12'h806;
        src34 <= 12'h123;
        src35 <= 12'h1c0;
        src36 <= 12'h79b;
        src37 <= 12'hc0e;
        src38 <= 12'h197;
        src39 <= 12'hb9a;
        src40 <= 12'h94e;
        src41 <= 12'h91a;
        src42 <= 12'h676;
        src43 <= 12'h56d;
        src44 <= 12'h681;
        src45 <= 12'h9d6;
        src46 <= 12'h158;
        src47 <= 12'h705;
        src48 <= 12'h82;
        src49 <= 12'h29a;
        src50 <= 12'hfbf;
        src51 <= 12'h79b;
        src52 <= 12'h202;
        src53 <= 12'h10b;
        exp <= 18'h14b1c;
        #1
        src0 <= 12'hb3a;
        src1 <= 12'h86c;
        src2 <= 12'hf3a;
        src3 <= 12'hb8e;
        src4 <= 12'hece;
        src5 <= 12'h9a6;
        src6 <= 12'h36b;
        src7 <= 12'hec8;
        src8 <= 12'h39c;
        src9 <= 12'h2b4;
        src10 <= 12'h394;
        src11 <= 12'hc6b;
        src12 <= 12'h9b1;
        src13 <= 12'hcaf;
        src14 <= 12'h4d;
        src15 <= 12'ha2e;
        src16 <= 12'hdb4;
        src17 <= 12'h863;
        src18 <= 12'h6d5;
        src19 <= 12'h124;
        src20 <= 12'h582;
        src21 <= 12'ha78;
        src22 <= 12'h4d9;
        src23 <= 12'h223;
        src24 <= 12'h89d;
        src25 <= 12'h77f;
        src26 <= 12'hf91;
        src27 <= 12'h5f9;
        src28 <= 12'hd4e;
        src29 <= 12'hae3;
        src30 <= 12'hc2;
        src31 <= 12'h493;
        src32 <= 12'h9e3;
        src33 <= 12'hdb6;
        src34 <= 12'h833;
        src35 <= 12'ha33;
        src36 <= 12'hb6e;
        src37 <= 12'hc70;
        src38 <= 12'h67b;
        src39 <= 12'h9fc;
        src40 <= 12'h29c;
        src41 <= 12'h4f2;
        src42 <= 12'h936;
        src43 <= 12'h5b6;
        src44 <= 12'he7f;
        src45 <= 12'hb68;
        src46 <= 12'h3cc;
        src47 <= 12'hb63;
        src48 <= 12'h7cb;
        src49 <= 12'hfe4;
        src50 <= 12'h3ef;
        src51 <= 12'h7f1;
        src52 <= 12'h17b;
        src53 <= 12'h383;
        exp <= 18'h1c2e2;
        #1
        src0 <= 12'ha23;
        src1 <= 12'h456;
        src2 <= 12'h472;
        src3 <= 12'hcc2;
        src4 <= 12'h7dc;
        src5 <= 12'h9ce;
        src6 <= 12'h95a;
        src7 <= 12'he87;
        src8 <= 12'h73d;
        src9 <= 12'h31d;
        src10 <= 12'h19c;
        src11 <= 12'h67d;
        src12 <= 12'hcb1;
        src13 <= 12'h5a7;
        src14 <= 12'hdd5;
        src15 <= 12'hc62;
        src16 <= 12'ha10;
        src17 <= 12'ha01;
        src18 <= 12'h399;
        src19 <= 12'hd35;
        src20 <= 12'hba8;
        src21 <= 12'hc10;
        src22 <= 12'h140;
        src23 <= 12'h681;
        src24 <= 12'h117;
        src25 <= 12'hffd;
        src26 <= 12'h8e6;
        src27 <= 12'hd40;
        src28 <= 12'hf02;
        src29 <= 12'h22f;
        src30 <= 12'h8ca;
        src31 <= 12'hf7b;
        src32 <= 12'hc1e;
        src33 <= 12'hae9;
        src34 <= 12'h55;
        src35 <= 12'hde0;
        src36 <= 12'hc5f;
        src37 <= 12'hf7;
        src38 <= 12'h83a;
        src39 <= 12'h472;
        src40 <= 12'ha8d;
        src41 <= 12'h602;
        src42 <= 12'hcc5;
        src43 <= 12'h969;
        src44 <= 12'h804;
        src45 <= 12'hc84;
        src46 <= 12'haaa;
        src47 <= 12'h391;
        src48 <= 12'h92b;
        src49 <= 12'hdbc;
        src50 <= 12'hc7f;
        src51 <= 12'h3b;
        src52 <= 12'h6e4;
        src53 <= 12'h1fe;
        exp <= 18'h1d283;
        #1
        src0 <= 12'h94a;
        src1 <= 12'hfb7;
        src2 <= 12'h7c0;
        src3 <= 12'hedc;
        src4 <= 12'h127;
        src5 <= 12'h135;
        src6 <= 12'h2ce;
        src7 <= 12'hc4f;
        src8 <= 12'ha0e;
        src9 <= 12'hcd3;
        src10 <= 12'h64a;
        src11 <= 12'h588;
        src12 <= 12'h9c1;
        src13 <= 12'haa6;
        src14 <= 12'h236;
        src15 <= 12'hec7;
        src16 <= 12'h34c;
        src17 <= 12'h45b;
        src18 <= 12'hd3a;
        src19 <= 12'h37a;
        src20 <= 12'ha83;
        src21 <= 12'h317;
        src22 <= 12'h346;
        src23 <= 12'hbf8;
        src24 <= 12'h26f;
        src25 <= 12'h8a3;
        src26 <= 12'h438;
        src27 <= 12'h244;
        src28 <= 12'he2f;
        src29 <= 12'h992;
        src30 <= 12'h2b9;
        src31 <= 12'he3f;
        src32 <= 12'h77d;
        src33 <= 12'hced;
        src34 <= 12'h507;
        src35 <= 12'h8ec;
        src36 <= 12'h4c2;
        src37 <= 12'hce2;
        src38 <= 12'h6d8;
        src39 <= 12'h94c;
        src40 <= 12'h699;
        src41 <= 12'h901;
        src42 <= 12'ha73;
        src43 <= 12'h3d0;
        src44 <= 12'he3c;
        src45 <= 12'h45f;
        src46 <= 12'hada;
        src47 <= 12'hf3;
        src48 <= 12'h353;
        src49 <= 12'h1c7;
        src50 <= 12'h4b1;
        src51 <= 12'h962;
        src52 <= 12'h878;
        src53 <= 12'hbb2;
        exp <= 18'h1a068;
        #1
        src0 <= 12'h83b;
        src1 <= 12'h197;
        src2 <= 12'hae2;
        src3 <= 12'hd74;
        src4 <= 12'h313;
        src5 <= 12'h37e;
        src6 <= 12'h590;
        src7 <= 12'hcb8;
        src8 <= 12'h5e8;
        src9 <= 12'hedc;
        src10 <= 12'h93a;
        src11 <= 12'h21b;
        src12 <= 12'h20a;
        src13 <= 12'h3dc;
        src14 <= 12'h9f0;
        src15 <= 12'h34f;
        src16 <= 12'hfbe;
        src17 <= 12'h4a9;
        src18 <= 12'h48d;
        src19 <= 12'h651;
        src20 <= 12'h78d;
        src21 <= 12'hf22;
        src22 <= 12'he40;
        src23 <= 12'h5c1;
        src24 <= 12'h880;
        src25 <= 12'h6be;
        src26 <= 12'h82e;
        src27 <= 12'hdcd;
        src28 <= 12'h70c;
        src29 <= 12'h169;
        src30 <= 12'h1ed;
        src31 <= 12'h598;
        src32 <= 12'h50;
        src33 <= 12'h3f2;
        src34 <= 12'h996;
        src35 <= 12'h58a;
        src36 <= 12'h210;
        src37 <= 12'h606;
        src38 <= 12'h47d;
        src39 <= 12'h3b;
        src40 <= 12'h5c4;
        src41 <= 12'h52;
        src42 <= 12'h99d;
        src43 <= 12'h671;
        src44 <= 12'hc06;
        src45 <= 12'heef;
        src46 <= 12'h31;
        src47 <= 12'h556;
        src48 <= 12'h70f;
        src49 <= 12'he6d;
        src50 <= 12'hcdc;
        src51 <= 12'hc15;
        src52 <= 12'h9be;
        src53 <= 12'h302;
        exp <= 18'h17f64;
        #1
        src0 <= 12'h4e9;
        src1 <= 12'hcc8;
        src2 <= 12'he24;
        src3 <= 12'hd9a;
        src4 <= 12'h1e9;
        src5 <= 12'hd3;
        src6 <= 12'h74f;
        src7 <= 12'hdf8;
        src8 <= 12'h9c5;
        src9 <= 12'h673;
        src10 <= 12'hdac;
        src11 <= 12'h542;
        src12 <= 12'h3b0;
        src13 <= 12'h3c1;
        src14 <= 12'he78;
        src15 <= 12'h573;
        src16 <= 12'h3a4;
        src17 <= 12'hf6b;
        src18 <= 12'h222;
        src19 <= 12'h33b;
        src20 <= 12'hbf9;
        src21 <= 12'h34b;
        src22 <= 12'h514;
        src23 <= 12'hcd2;
        src24 <= 12'h569;
        src25 <= 12'h8ac;
        src26 <= 12'h5e0;
        src27 <= 12'h209;
        src28 <= 12'h25a;
        src29 <= 12'h181;
        src30 <= 12'hfd8;
        src31 <= 12'h27a;
        src32 <= 12'h3e5;
        src33 <= 12'hdda;
        src34 <= 12'h3b5;
        src35 <= 12'hecd;
        src36 <= 12'hfe0;
        src37 <= 12'hf44;
        src38 <= 12'h3ac;
        src39 <= 12'h461;
        src40 <= 12'h91c;
        src41 <= 12'h335;
        src42 <= 12'h1db;
        src43 <= 12'he86;
        src44 <= 12'hece;
        src45 <= 12'h98;
        src46 <= 12'h35a;
        src47 <= 12'h61;
        src48 <= 12'h3ad;
        src49 <= 12'hd02;
        src50 <= 12'hdb6;
        src51 <= 12'h8f8;
        src52 <= 12'hf2;
        src53 <= 12'h550;
        exp <= 18'h19299;
        #1
        src0 <= 12'h1ec;
        src1 <= 12'hbaf;
        src2 <= 12'h489;
        src3 <= 12'hd28;
        src4 <= 12'hd6e;
        src5 <= 12'h245;
        src6 <= 12'h132;
        src7 <= 12'hb18;
        src8 <= 12'hcaf;
        src9 <= 12'h2c4;
        src10 <= 12'h294;
        src11 <= 12'he49;
        src12 <= 12'ha25;
        src13 <= 12'h60c;
        src14 <= 12'h249;
        src15 <= 12'hdd0;
        src16 <= 12'hc0a;
        src17 <= 12'h6b5;
        src18 <= 12'h1e4;
        src19 <= 12'h4a8;
        src20 <= 12'hbd4;
        src21 <= 12'hee6;
        src22 <= 12'h100;
        src23 <= 12'hf99;
        src24 <= 12'hda;
        src25 <= 12'h53e;
        src26 <= 12'hb30;
        src27 <= 12'h584;
        src28 <= 12'h225;
        src29 <= 12'hbcd;
        src30 <= 12'hb3c;
        src31 <= 12'h953;
        src32 <= 12'hfb3;
        src33 <= 12'h971;
        src34 <= 12'heb1;
        src35 <= 12'hfdf;
        src36 <= 12'hf9d;
        src37 <= 12'h180;
        src38 <= 12'h3da;
        src39 <= 12'hf1c;
        src40 <= 12'h688;
        src41 <= 12'hdec;
        src42 <= 12'hdb;
        src43 <= 12'h42e;
        src44 <= 12'ha0e;
        src45 <= 12'hf0d;
        src46 <= 12'h293;
        src47 <= 12'h147;
        src48 <= 12'hf2d;
        src49 <= 12'h790;
        src50 <= 12'h5f5;
        src51 <= 12'h4b1;
        src52 <= 12'hd5;
        src53 <= 12'h141;
        exp <= 18'h1af80;
        #1
        src0 <= 12'hed2;
        src1 <= 12'h465;
        src2 <= 12'h896;
        src3 <= 12'he0f;
        src4 <= 12'h916;
        src5 <= 12'h891;
        src6 <= 12'h51d;
        src7 <= 12'h164;
        src8 <= 12'h551;
        src9 <= 12'h9eb;
        src10 <= 12'h20d;
        src11 <= 12'hc49;
        src12 <= 12'hb20;
        src13 <= 12'h37d;
        src14 <= 12'hd43;
        src15 <= 12'haad;
        src16 <= 12'h568;
        src17 <= 12'h7ce;
        src18 <= 12'hc36;
        src19 <= 12'h578;
        src20 <= 12'hcce;
        src21 <= 12'h260;
        src22 <= 12'h58;
        src23 <= 12'h6ac;
        src24 <= 12'h53;
        src25 <= 12'h70;
        src26 <= 12'h735;
        src27 <= 12'h3a2;
        src28 <= 12'h1be;
        src29 <= 12'h56f;
        src30 <= 12'h1b9;
        src31 <= 12'h800;
        src32 <= 12'hb0;
        src33 <= 12'h8b6;
        src34 <= 12'h1e8;
        src35 <= 12'hc07;
        src36 <= 12'hb66;
        src37 <= 12'hb42;
        src38 <= 12'hac6;
        src39 <= 12'h65b;
        src40 <= 12'h8c7;
        src41 <= 12'h5de;
        src42 <= 12'h964;
        src43 <= 12'hff2;
        src44 <= 12'hb2d;
        src45 <= 12'hf83;
        src46 <= 12'h980;
        src47 <= 12'hb26;
        src48 <= 12'h994;
        src49 <= 12'h1f5;
        src50 <= 12'hd77;
        src51 <= 12'h86;
        src52 <= 12'h679;
        src53 <= 12'h911;
        exp <= 18'h19738;
        #1
        src0 <= 12'h173;
        src1 <= 12'hb8e;
        src2 <= 12'h3a9;
        src3 <= 12'h3e0;
        src4 <= 12'hc2a;
        src5 <= 12'h280;
        src6 <= 12'hefa;
        src7 <= 12'h709;
        src8 <= 12'hf17;
        src9 <= 12'h77d;
        src10 <= 12'h488;
        src11 <= 12'h5be;
        src12 <= 12'h7af;
        src13 <= 12'h8e7;
        src14 <= 12'h3e8;
        src15 <= 12'hb26;
        src16 <= 12'hb15;
        src17 <= 12'h72d;
        src18 <= 12'h572;
        src19 <= 12'hda3;
        src20 <= 12'h5ba;
        src21 <= 12'h33f;
        src22 <= 12'h8b7;
        src23 <= 12'h4d6;
        src24 <= 12'hb87;
        src25 <= 12'h78e;
        src26 <= 12'hf41;
        src27 <= 12'h663;
        src28 <= 12'h9cb;
        src29 <= 12'h8fa;
        src30 <= 12'h208;
        src31 <= 12'hae4;
        src32 <= 12'ha6b;
        src33 <= 12'hd96;
        src34 <= 12'h365;
        src35 <= 12'h763;
        src36 <= 12'h63d;
        src37 <= 12'h49a;
        src38 <= 12'h57f;
        src39 <= 12'h560;
        src40 <= 12'hf41;
        src41 <= 12'h30a;
        src42 <= 12'h8f0;
        src43 <= 12'h1c5;
        src44 <= 12'he96;
        src45 <= 12'h94f;
        src46 <= 12'h541;
        src47 <= 12'h97d;
        src48 <= 12'h5cb;
        src49 <= 12'h6b4;
        src50 <= 12'hb1;
        src51 <= 12'h5be;
        src52 <= 12'he39;
        src53 <= 12'hac6;
        exp <= 18'h1a60b;
        #1
        src0 <= 12'ha7b;
        src1 <= 12'hf4c;
        src2 <= 12'h7a4;
        src3 <= 12'hd05;
        src4 <= 12'h113;
        src5 <= 12'hbd0;
        src6 <= 12'h93a;
        src7 <= 12'h7b6;
        src8 <= 12'hf88;
        src9 <= 12'h7c5;
        src10 <= 12'haa;
        src11 <= 12'h24e;
        src12 <= 12'h7f8;
        src13 <= 12'hd39;
        src14 <= 12'hb7e;
        src15 <= 12'haf1;
        src16 <= 12'h613;
        src17 <= 12'h66d;
        src18 <= 12'h38;
        src19 <= 12'h175;
        src20 <= 12'hef7;
        src21 <= 12'h508;
        src22 <= 12'h4a9;
        src23 <= 12'h9ef;
        src24 <= 12'he5b;
        src25 <= 12'hb4a;
        src26 <= 12'h189;
        src27 <= 12'h1db;
        src28 <= 12'h1f7;
        src29 <= 12'haaf;
        src30 <= 12'h3f5;
        src31 <= 12'h868;
        src32 <= 12'hd06;
        src33 <= 12'h2c8;
        src34 <= 12'h822;
        src35 <= 12'had1;
        src36 <= 12'hf23;
        src37 <= 12'hbe9;
        src38 <= 12'h603;
        src39 <= 12'hbff;
        src40 <= 12'hc16;
        src41 <= 12'he1a;
        src42 <= 12'h692;
        src43 <= 12'h769;
        src44 <= 12'h612;
        src45 <= 12'h2ac;
        src46 <= 12'h6c6;
        src47 <= 12'h3d5;
        src48 <= 12'h50b;
        src49 <= 12'hc50;
        src50 <= 12'h9b1;
        src51 <= 12'hef6;
        src52 <= 12'h9ae;
        src53 <= 12'h3f;
        exp <= 18'h1b83a;
        #1
        src0 <= 12'h485;
        src1 <= 12'h62e;
        src2 <= 12'h537;
        src3 <= 12'hbfb;
        src4 <= 12'ha16;
        src5 <= 12'h71;
        src6 <= 12'h1b3;
        src7 <= 12'hc57;
        src8 <= 12'h94;
        src9 <= 12'hc08;
        src10 <= 12'h20c;
        src11 <= 12'hc4b;
        src12 <= 12'hd27;
        src13 <= 12'he1c;
        src14 <= 12'h379;
        src15 <= 12'h9ed;
        src16 <= 12'ha01;
        src17 <= 12'hfcb;
        src18 <= 12'hde8;
        src19 <= 12'had9;
        src20 <= 12'h936;
        src21 <= 12'h995;
        src22 <= 12'h6e8;
        src23 <= 12'h77f;
        src24 <= 12'h877;
        src25 <= 12'h1c4;
        src26 <= 12'h271;
        src27 <= 12'h3d3;
        src28 <= 12'hcce;
        src29 <= 12'h7e6;
        src30 <= 12'hf67;
        src31 <= 12'ha5c;
        src32 <= 12'ha95;
        src33 <= 12'h591;
        src34 <= 12'h2ee;
        src35 <= 12'h4f8;
        src36 <= 12'hb76;
        src37 <= 12'h7e9;
        src38 <= 12'h1a6;
        src39 <= 12'heae;
        src40 <= 12'h3d9;
        src41 <= 12'hd4e;
        src42 <= 12'hf29;
        src43 <= 12'h353;
        src44 <= 12'h32f;
        src45 <= 12'hdb;
        src46 <= 12'h770;
        src47 <= 12'he0d;
        src48 <= 12'h38f;
        src49 <= 12'h42a;
        src50 <= 12'hb;
        src51 <= 12'h7dd;
        src52 <= 12'hdc7;
        src53 <= 12'h837;
        exp <= 18'h1a94f;
        #1
        src0 <= 12'he09;
        src1 <= 12'h6dd;
        src2 <= 12'h5e;
        src3 <= 12'ha1a;
        src4 <= 12'h4f3;
        src5 <= 12'h777;
        src6 <= 12'hcb5;
        src7 <= 12'hf75;
        src8 <= 12'h222;
        src9 <= 12'h674;
        src10 <= 12'heaf;
        src11 <= 12'h1b0;
        src12 <= 12'hb72;
        src13 <= 12'h7fd;
        src14 <= 12'he09;
        src15 <= 12'habf;
        src16 <= 12'hc4f;
        src17 <= 12'h76e;
        src18 <= 12'h9ba;
        src19 <= 12'h7d7;
        src20 <= 12'hed8;
        src21 <= 12'hbee;
        src22 <= 12'h262;
        src23 <= 12'hce5;
        src24 <= 12'hfab;
        src25 <= 12'hdb4;
        src26 <= 12'h108;
        src27 <= 12'h6c7;
        src28 <= 12'h8d4;
        src29 <= 12'h596;
        src30 <= 12'haf4;
        src31 <= 12'h322;
        src32 <= 12'h926;
        src33 <= 12'h420;
        src34 <= 12'hb7b;
        src35 <= 12'h83f;
        src36 <= 12'h952;
        src37 <= 12'hc23;
        src38 <= 12'hbfd;
        src39 <= 12'h717;
        src40 <= 12'h1d9;
        src41 <= 12'h83d;
        src42 <= 12'h8aa;
        src43 <= 12'h1e5;
        src44 <= 12'ha93;
        src45 <= 12'h906;
        src46 <= 12'h3aa;
        src47 <= 12'h7cc;
        src48 <= 12'h189;
        src49 <= 12'h8b;
        src50 <= 12'hdaa;
        src51 <= 12'hab0;
        src52 <= 12'h69;
        src53 <= 12'h877;
        exp <= 18'h1beb2;
        #1
        src0 <= 12'h1f;
        src1 <= 12'ha31;
        src2 <= 12'h4a5;
        src3 <= 12'h1b9;
        src4 <= 12'h699;
        src5 <= 12'haf7;
        src6 <= 12'h9c0;
        src7 <= 12'h7db;
        src8 <= 12'h544;
        src9 <= 12'hf6;
        src10 <= 12'hb64;
        src11 <= 12'h6d3;
        src12 <= 12'h5dc;
        src13 <= 12'ha13;
        src14 <= 12'he23;
        src15 <= 12'hf8c;
        src16 <= 12'h966;
        src17 <= 12'h54a;
        src18 <= 12'ha54;
        src19 <= 12'h302;
        src20 <= 12'h4d6;
        src21 <= 12'h219;
        src22 <= 12'h8bc;
        src23 <= 12'h943;
        src24 <= 12'h250;
        src25 <= 12'h49f;
        src26 <= 12'h50;
        src27 <= 12'hc95;
        src28 <= 12'h60f;
        src29 <= 12'h2d3;
        src30 <= 12'h2d1;
        src31 <= 12'h720;
        src32 <= 12'h79d;
        src33 <= 12'h350;
        src34 <= 12'h468;
        src35 <= 12'h719;
        src36 <= 12'h745;
        src37 <= 12'h67a;
        src38 <= 12'h7b8;
        src39 <= 12'h1f4;
        src40 <= 12'h86f;
        src41 <= 12'hd95;
        src42 <= 12'h76f;
        src43 <= 12'ha35;
        src44 <= 12'hcc2;
        src45 <= 12'hcb2;
        src46 <= 12'hee3;
        src47 <= 12'hd2a;
        src48 <= 12'hb17;
        src49 <= 12'haf0;
        src50 <= 12'ha33;
        src51 <= 12'h97f;
        src52 <= 12'h36c;
        src53 <= 12'h59c;
        exp <= 18'h19346;
        #1
        src0 <= 12'h738;
        src1 <= 12'hc97;
        src2 <= 12'h287;
        src3 <= 12'hd55;
        src4 <= 12'hf83;
        src5 <= 12'he9d;
        src6 <= 12'h99d;
        src7 <= 12'hd9;
        src8 <= 12'he61;
        src9 <= 12'h3cc;
        src10 <= 12'h4f3;
        src11 <= 12'hd00;
        src12 <= 12'hdd9;
        src13 <= 12'haea;
        src14 <= 12'h3ce;
        src15 <= 12'hb3d;
        src16 <= 12'he86;
        src17 <= 12'h371;
        src18 <= 12'h107;
        src19 <= 12'hd97;
        src20 <= 12'he32;
        src21 <= 12'h952;
        src22 <= 12'hd6d;
        src23 <= 12'h4d4;
        src24 <= 12'h20c;
        src25 <= 12'h374;
        src26 <= 12'h491;
        src27 <= 12'hd3b;
        src28 <= 12'h54b;
        src29 <= 12'heda;
        src30 <= 12'hf43;
        src31 <= 12'he53;
        src32 <= 12'hd3d;
        src33 <= 12'h1bb;
        src34 <= 12'he9c;
        src35 <= 12'h9f7;
        src36 <= 12'hf77;
        src37 <= 12'h801;
        src38 <= 12'h25a;
        src39 <= 12'h1ae;
        src40 <= 12'h76b;
        src41 <= 12'h305;
        src42 <= 12'h356;
        src43 <= 12'hc6a;
        src44 <= 12'h270;
        src45 <= 12'h947;
        src46 <= 12'hef9;
        src47 <= 12'h178;
        src48 <= 12'h385;
        src49 <= 12'h259;
        src50 <= 12'hb56;
        src51 <= 12'ha40;
        src52 <= 12'h1b4;
        src53 <= 12'h819;
        exp <= 18'h1ca34;
        #1
        src0 <= 12'he29;
        src1 <= 12'ha65;
        src2 <= 12'he01;
        src3 <= 12'h1a;
        src4 <= 12'h7c5;
        src5 <= 12'h4c1;
        src6 <= 12'h73f;
        src7 <= 12'h44d;
        src8 <= 12'hc90;
        src9 <= 12'h69c;
        src10 <= 12'hd59;
        src11 <= 12'h8c5;
        src12 <= 12'h575;
        src13 <= 12'h8e5;
        src14 <= 12'hd48;
        src15 <= 12'hfbe;
        src16 <= 12'h532;
        src17 <= 12'ha0d;
        src18 <= 12'h5ab;
        src19 <= 12'h400;
        src20 <= 12'h9b4;
        src21 <= 12'h373;
        src22 <= 12'h656;
        src23 <= 12'h1c;
        src24 <= 12'h6ed;
        src25 <= 12'heb1;
        src26 <= 12'h418;
        src27 <= 12'hb5b;
        src28 <= 12'hbc8;
        src29 <= 12'hebf;
        src30 <= 12'h1a6;
        src31 <= 12'hf6d;
        src32 <= 12'ha3d;
        src33 <= 12'h53f;
        src34 <= 12'h163;
        src35 <= 12'hca7;
        src36 <= 12'h499;
        src37 <= 12'hf8a;
        src38 <= 12'h99b;
        src39 <= 12'h14d;
        src40 <= 12'h59a;
        src41 <= 12'hebd;
        src42 <= 12'hb2e;
        src43 <= 12'hd04;
        src44 <= 12'h2e0;
        src45 <= 12'he8a;
        src46 <= 12'h939;
        src47 <= 12'h7f;
        src48 <= 12'h101;
        src49 <= 12'h63;
        src50 <= 12'h722;
        src51 <= 12'h15e;
        src52 <= 12'h776;
        src53 <= 12'haeb;
        exp <= 18'h1b114;
        #1
        src0 <= 12'h9f1;
        src1 <= 12'h45f;
        src2 <= 12'h7c9;
        src3 <= 12'hb49;
        src4 <= 12'h370;
        src5 <= 12'ha3c;
        src6 <= 12'hde1;
        src7 <= 12'hc26;
        src8 <= 12'h722;
        src9 <= 12'hc6f;
        src10 <= 12'ha3e;
        src11 <= 12'heba;
        src12 <= 12'h9d6;
        src13 <= 12'h281;
        src14 <= 12'hd62;
        src15 <= 12'hf04;
        src16 <= 12'h11b;
        src17 <= 12'h7b4;
        src18 <= 12'hf;
        src19 <= 12'h7ee;
        src20 <= 12'h23b;
        src21 <= 12'h873;
        src22 <= 12'h119;
        src23 <= 12'hd80;
        src24 <= 12'h2b5;
        src25 <= 12'h1df;
        src26 <= 12'hf3;
        src27 <= 12'ha6e;
        src28 <= 12'hf79;
        src29 <= 12'h10;
        src30 <= 12'h270;
        src31 <= 12'h505;
        src32 <= 12'h7bf;
        src33 <= 12'h359;
        src34 <= 12'h8be;
        src35 <= 12'h54f;
        src36 <= 12'hbcb;
        src37 <= 12'h44d;
        src38 <= 12'h512;
        src39 <= 12'heb7;
        src40 <= 12'h402;
        src41 <= 12'h92b;
        src42 <= 12'hdcc;
        src43 <= 12'h1a;
        src44 <= 12'hf83;
        src45 <= 12'ha38;
        src46 <= 12'hff0;
        src47 <= 12'h922;
        src48 <= 12'h8c9;
        src49 <= 12'h2f2;
        src50 <= 12'h744;
        src51 <= 12'hde8;
        src52 <= 12'hd6e;
        src53 <= 12'he60;
        exp <= 18'h1b6fc;
        #1
        src0 <= 12'hf56;
        src1 <= 12'h6ed;
        src2 <= 12'h2dd;
        src3 <= 12'hc81;
        src4 <= 12'h23e;
        src5 <= 12'hf42;
        src6 <= 12'h377;
        src7 <= 12'hb53;
        src8 <= 12'hef7;
        src9 <= 12'hc20;
        src10 <= 12'h2e;
        src11 <= 12'hf13;
        src12 <= 12'h521;
        src13 <= 12'h391;
        src14 <= 12'h69e;
        src15 <= 12'h87a;
        src16 <= 12'h1a;
        src17 <= 12'ha09;
        src18 <= 12'he2d;
        src19 <= 12'he83;
        src20 <= 12'h4a;
        src21 <= 12'hf25;
        src22 <= 12'hb07;
        src23 <= 12'h506;
        src24 <= 12'h538;
        src25 <= 12'he;
        src26 <= 12'h8d4;
        src27 <= 12'hc2d;
        src28 <= 12'h2ec;
        src29 <= 12'h6cc;
        src30 <= 12'h4ae;
        src31 <= 12'h127;
        src32 <= 12'h2f2;
        src33 <= 12'h687;
        src34 <= 12'h1e6;
        src35 <= 12'hd54;
        src36 <= 12'h766;
        src37 <= 12'hf21;
        src38 <= 12'hcbf;
        src39 <= 12'h3fa;
        src40 <= 12'he80;
        src41 <= 12'h70e;
        src42 <= 12'hcc;
        src43 <= 12'hdf0;
        src44 <= 12'h97f;
        src45 <= 12'hb4e;
        src46 <= 12'hc14;
        src47 <= 12'hb28;
        src48 <= 12'hbf8;
        src49 <= 12'hac4;
        src50 <= 12'h1ee;
        src51 <= 12'he;
        src52 <= 12'hc65;
        src53 <= 12'h743;
        exp <= 18'h1b4d6;
        #1
        src0 <= 12'h528;
        src1 <= 12'ha6b;
        src2 <= 12'h21a;
        src3 <= 12'hd82;
        src4 <= 12'hb0f;
        src5 <= 12'h84;
        src6 <= 12'hcba;
        src7 <= 12'h8d0;
        src8 <= 12'h5fe;
        src9 <= 12'he1b;
        src10 <= 12'hd4d;
        src11 <= 12'hea0;
        src12 <= 12'h39a;
        src13 <= 12'hc55;
        src14 <= 12'hbb5;
        src15 <= 12'h86a;
        src16 <= 12'ha0f;
        src17 <= 12'h98e;
        src18 <= 12'hbd6;
        src19 <= 12'h94b;
        src20 <= 12'h9a9;
        src21 <= 12'h37b;
        src22 <= 12'h441;
        src23 <= 12'h10e;
        src24 <= 12'hc8;
        src25 <= 12'h2ee;
        src26 <= 12'hc66;
        src27 <= 12'h48d;
        src28 <= 12'ha6;
        src29 <= 12'h733;
        src30 <= 12'hb2f;
        src31 <= 12'h810;
        src32 <= 12'h213;
        src33 <= 12'h571;
        src34 <= 12'h585;
        src35 <= 12'h573;
        src36 <= 12'hc0f;
        src37 <= 12'h8f1;
        src38 <= 12'h384;
        src39 <= 12'h10c;
        src40 <= 12'h13c;
        src41 <= 12'h95f;
        src42 <= 12'hfe0;
        src43 <= 12'h5a;
        src44 <= 12'h9b3;
        src45 <= 12'h21f;
        src46 <= 12'hc6e;
        src47 <= 12'hca8;
        src48 <= 12'he53;
        src49 <= 12'h3fd;
        src50 <= 12'h1fb;
        src51 <= 12'hb36;
        src52 <= 12'hc59;
        src53 <= 12'hdf7;
        exp <= 18'h1a4ec;
        #1
        src0 <= 12'hcee;
        src1 <= 12'h6fb;
        src2 <= 12'hf25;
        src3 <= 12'hf10;
        src4 <= 12'hf65;
        src5 <= 12'h26;
        src6 <= 12'h3e8;
        src7 <= 12'hc3b;
        src8 <= 12'h26;
        src9 <= 12'hd47;
        src10 <= 12'h18f;
        src11 <= 12'h60f;
        src12 <= 12'h35b;
        src13 <= 12'h35b;
        src14 <= 12'h32d;
        src15 <= 12'h192;
        src16 <= 12'h8ac;
        src17 <= 12'h50e;
        src18 <= 12'h17d;
        src19 <= 12'h249;
        src20 <= 12'h622;
        src21 <= 12'h8cd;
        src22 <= 12'h6b5;
        src23 <= 12'h602;
        src24 <= 12'h824;
        src25 <= 12'hd8d;
        src26 <= 12'h8b6;
        src27 <= 12'h437;
        src28 <= 12'h242;
        src29 <= 12'hb9d;
        src30 <= 12'h3a1;
        src31 <= 12'h324;
        src32 <= 12'he09;
        src33 <= 12'he27;
        src34 <= 12'h8a7;
        src35 <= 12'hed7;
        src36 <= 12'h8cb;
        src37 <= 12'hbd7;
        src38 <= 12'hd87;
        src39 <= 12'h33c;
        src40 <= 12'h48;
        src41 <= 12'hbe8;
        src42 <= 12'hd9d;
        src43 <= 12'h9a9;
        src44 <= 12'hb14;
        src45 <= 12'h274;
        src46 <= 12'hd2a;
        src47 <= 12'h9ab;
        src48 <= 12'hbaa;
        src49 <= 12'h17d;
        src50 <= 12'ha4;
        src51 <= 12'ha1a;
        src52 <= 12'h1ca;
        src53 <= 12'heb4;
        exp <= 18'h19ffd;
        #1
        src0 <= 12'h9ec;
        src1 <= 12'h16f;
        src2 <= 12'hfbb;
        src3 <= 12'h18c;
        src4 <= 12'h137;
        src5 <= 12'h783;
        src6 <= 12'he95;
        src7 <= 12'h80d;
        src8 <= 12'hf78;
        src9 <= 12'hc2;
        src10 <= 12'hdcd;
        src11 <= 12'h8be;
        src12 <= 12'hed3;
        src13 <= 12'h2e3;
        src14 <= 12'h577;
        src15 <= 12'h46f;
        src16 <= 12'h3bf;
        src17 <= 12'h286;
        src18 <= 12'h7d5;
        src19 <= 12'h9c1;
        src20 <= 12'hed8;
        src21 <= 12'hfdf;
        src22 <= 12'h5d7;
        src23 <= 12'hb1e;
        src24 <= 12'hdea;
        src25 <= 12'h240;
        src26 <= 12'h529;
        src27 <= 12'h576;
        src28 <= 12'h752;
        src29 <= 12'h238;
        src30 <= 12'h308;
        src31 <= 12'h183;
        src32 <= 12'h4d6;
        src33 <= 12'h886;
        src34 <= 12'h5e7;
        src35 <= 12'h476;
        src36 <= 12'h2ac;
        src37 <= 12'hc25;
        src38 <= 12'h7a7;
        src39 <= 12'hd8c;
        src40 <= 12'hfb3;
        src41 <= 12'hea7;
        src42 <= 12'h807;
        src43 <= 12'h26d;
        src44 <= 12'h218;
        src45 <= 12'hc89;
        src46 <= 12'h4e3;
        src47 <= 12'h88;
        src48 <= 12'h481;
        src49 <= 12'he3c;
        src50 <= 12'hc5f;
        src51 <= 12'h77a;
        src52 <= 12'h6cb;
        src53 <= 12'hb17;
        exp <= 18'h19fd3;
        #1
        src0 <= 12'hec0;
        src1 <= 12'ha49;
        src2 <= 12'hbbd;
        src3 <= 12'h4cb;
        src4 <= 12'had4;
        src5 <= 12'h92f;
        src6 <= 12'ha7f;
        src7 <= 12'h6af;
        src8 <= 12'h3c;
        src9 <= 12'hb41;
        src10 <= 12'h391;
        src11 <= 12'h6ba;
        src12 <= 12'head;
        src13 <= 12'h2d7;
        src14 <= 12'h8d9;
        src15 <= 12'hc15;
        src16 <= 12'h463;
        src17 <= 12'hcb5;
        src18 <= 12'ha4b;
        src19 <= 12'h48c;
        src20 <= 12'hddf;
        src21 <= 12'hde9;
        src22 <= 12'h2a;
        src23 <= 12'h1d1;
        src24 <= 12'h889;
        src25 <= 12'hcf7;
        src26 <= 12'h55f;
        src27 <= 12'h708;
        src28 <= 12'h404;
        src29 <= 12'h870;
        src30 <= 12'h8ca;
        src31 <= 12'h915;
        src32 <= 12'h937;
        src33 <= 12'h33;
        src34 <= 12'h70a;
        src35 <= 12'h853;
        src36 <= 12'h6a1;
        src37 <= 12'hc96;
        src38 <= 12'hd2e;
        src39 <= 12'h392;
        src40 <= 12'ha6e;
        src41 <= 12'h59b;
        src42 <= 12'h8a1;
        src43 <= 12'h2c7;
        src44 <= 12'h2c;
        src45 <= 12'h389;
        src46 <= 12'he64;
        src47 <= 12'h5cd;
        src48 <= 12'hb26;
        src49 <= 12'h918;
        src50 <= 12'he90;
        src51 <= 12'h9e2;
        src52 <= 12'h2f0;
        src53 <= 12'haf3;
        exp <= 18'h1b390;
        #1
        src0 <= 12'h6ad;
        src1 <= 12'h245;
        src2 <= 12'h1c8;
        src3 <= 12'hdfe;
        src4 <= 12'h692;
        src5 <= 12'hf75;
        src6 <= 12'h372;
        src7 <= 12'h7c4;
        src8 <= 12'hb6e;
        src9 <= 12'h33f;
        src10 <= 12'hfd4;
        src11 <= 12'h847;
        src12 <= 12'h4ad;
        src13 <= 12'hc1d;
        src14 <= 12'hc4f;
        src15 <= 12'h705;
        src16 <= 12'h381;
        src17 <= 12'he83;
        src18 <= 12'h734;
        src19 <= 12'hc33;
        src20 <= 12'h522;
        src21 <= 12'h82b;
        src22 <= 12'he64;
        src23 <= 12'hdb3;
        src24 <= 12'h99c;
        src25 <= 12'hd4a;
        src26 <= 12'hf1b;
        src27 <= 12'hf9c;
        src28 <= 12'h204;
        src29 <= 12'h283;
        src30 <= 12'h716;
        src31 <= 12'he98;
        src32 <= 12'h31a;
        src33 <= 12'hb7f;
        src34 <= 12'h78e;
        src35 <= 12'h9e7;
        src36 <= 12'hbcc;
        src37 <= 12'hbfd;
        src38 <= 12'h5e2;
        src39 <= 12'h195;
        src40 <= 12'h83e;
        src41 <= 12'h87a;
        src42 <= 12'hbe5;
        src43 <= 12'hc90;
        src44 <= 12'h6ee;
        src45 <= 12'h993;
        src46 <= 12'hf68;
        src47 <= 12'h1cf;
        src48 <= 12'hd6a;
        src49 <= 12'h55;
        src50 <= 12'h886;
        src51 <= 12'he9d;
        src52 <= 12'h8ff;
        src53 <= 12'hd8b;
        exp <= 18'h1e91b;
        #1
        src0 <= 12'h40b;
        src1 <= 12'h2ad;
        src2 <= 12'hbd4;
        src3 <= 12'hd95;
        src4 <= 12'h931;
        src5 <= 12'hd85;
        src6 <= 12'h86a;
        src7 <= 12'h1c1;
        src8 <= 12'h26f;
        src9 <= 12'h3e3;
        src10 <= 12'hd76;
        src11 <= 12'h383;
        src12 <= 12'hf2e;
        src13 <= 12'hf7c;
        src14 <= 12'h908;
        src15 <= 12'h4b5;
        src16 <= 12'h48c;
        src17 <= 12'h583;
        src18 <= 12'hecb;
        src19 <= 12'h118;
        src20 <= 12'h5be;
        src21 <= 12'h688;
        src22 <= 12'hb98;
        src23 <= 12'h2cc;
        src24 <= 12'h6c7;
        src25 <= 12'h205;
        src26 <= 12'h520;
        src27 <= 12'h519;
        src28 <= 12'h6e9;
        src29 <= 12'hb65;
        src30 <= 12'hccc;
        src31 <= 12'h7f1;
        src32 <= 12'h4b5;
        src33 <= 12'hdc5;
        src34 <= 12'hb90;
        src35 <= 12'h769;
        src36 <= 12'h7bb;
        src37 <= 12'h935;
        src38 <= 12'h496;
        src39 <= 12'hea6;
        src40 <= 12'h333;
        src41 <= 12'h488;
        src42 <= 12'h8f5;
        src43 <= 12'h36e;
        src44 <= 12'habe;
        src45 <= 12'hc12;
        src46 <= 12'h3b3;
        src47 <= 12'hd4e;
        src48 <= 12'hdb4;
        src49 <= 12'h356;
        src50 <= 12'h96e;
        src51 <= 12'h4fb;
        src52 <= 12'h50a;
        src53 <= 12'h25c;
        exp <= 18'h19fc7;
        #1
        src0 <= 12'h4e1;
        src1 <= 12'hedb;
        src2 <= 12'h62;
        src3 <= 12'h760;
        src4 <= 12'h931;
        src5 <= 12'hcdb;
        src6 <= 12'hac5;
        src7 <= 12'h35e;
        src8 <= 12'h782;
        src9 <= 12'h2bb;
        src10 <= 12'h1cc;
        src11 <= 12'he94;
        src12 <= 12'hc79;
        src13 <= 12'h110;
        src14 <= 12'h725;
        src15 <= 12'h7ed;
        src16 <= 12'h104;
        src17 <= 12'h675;
        src18 <= 12'h696;
        src19 <= 12'ha1b;
        src20 <= 12'h272;
        src21 <= 12'h1b6;
        src22 <= 12'h8cd;
        src23 <= 12'h63c;
        src24 <= 12'haa8;
        src25 <= 12'h865;
        src26 <= 12'h250;
        src27 <= 12'haa4;
        src28 <= 12'ha36;
        src29 <= 12'h8a0;
        src30 <= 12'h92e;
        src31 <= 12'h26f;
        src32 <= 12'haf6;
        src33 <= 12'hf6c;
        src34 <= 12'hd5f;
        src35 <= 12'h9b9;
        src36 <= 12'hfb3;
        src37 <= 12'hc4f;
        src38 <= 12'h381;
        src39 <= 12'h125;
        src40 <= 12'hdcc;
        src41 <= 12'hf27;
        src42 <= 12'hcc4;
        src43 <= 12'hfcf;
        src44 <= 12'hb39;
        src45 <= 12'hc76;
        src46 <= 12'h2b;
        src47 <= 12'hbce;
        src48 <= 12'hf8b;
        src49 <= 12'h31d;
        src50 <= 12'hee3;
        src51 <= 12'h362;
        src52 <= 12'h26e;
        src53 <= 12'hde9;
        exp <= 18'h1c548;
        #1
        src0 <= 12'he44;
        src1 <= 12'h65f;
        src2 <= 12'h5fb;
        src3 <= 12'h354;
        src4 <= 12'h547;
        src5 <= 12'hb0b;
        src6 <= 12'hb62;
        src7 <= 12'h7cf;
        src8 <= 12'hf2f;
        src9 <= 12'hf83;
        src10 <= 12'h959;
        src11 <= 12'h724;
        src12 <= 12'h3b1;
        src13 <= 12'h9e8;
        src14 <= 12'h8d9;
        src15 <= 12'h97c;
        src16 <= 12'hc34;
        src17 <= 12'hc88;
        src18 <= 12'h499;
        src19 <= 12'hf60;
        src20 <= 12'h176;
        src21 <= 12'ha33;
        src22 <= 12'h536;
        src23 <= 12'he7;
        src24 <= 12'hcbb;
        src25 <= 12'h73;
        src26 <= 12'h316;
        src27 <= 12'h4ef;
        src28 <= 12'h33e;
        src29 <= 12'h136;
        src30 <= 12'hbef;
        src31 <= 12'h5ea;
        src32 <= 12'h1b1;
        src33 <= 12'hab6;
        src34 <= 12'h691;
        src35 <= 12'h275;
        src36 <= 12'hbcb;
        src37 <= 12'hedb;
        src38 <= 12'h77f;
        src39 <= 12'h60f;
        src40 <= 12'ha49;
        src41 <= 12'h613;
        src42 <= 12'h0;
        src43 <= 12'h3fe;
        src44 <= 12'h528;
        src45 <= 12'hf50;
        src46 <= 12'hf12;
        src47 <= 12'haba;
        src48 <= 12'hd74;
        src49 <= 12'h6fd;
        src50 <= 12'h6d9;
        src51 <= 12'h26f;
        src52 <= 12'h72d;
        src53 <= 12'h76a;
        exp <= 18'h1a71c;
        #1
        src0 <= 12'h4fd;
        src1 <= 12'h510;
        src2 <= 12'hf91;
        src3 <= 12'h6f3;
        src4 <= 12'he5d;
        src5 <= 12'h4f1;
        src6 <= 12'he78;
        src7 <= 12'hcb9;
        src8 <= 12'h6f5;
        src9 <= 12'h42a;
        src10 <= 12'h605;
        src11 <= 12'he47;
        src12 <= 12'h1dc;
        src13 <= 12'he37;
        src14 <= 12'h31c;
        src15 <= 12'h868;
        src16 <= 12'h523;
        src17 <= 12'hb63;
        src18 <= 12'h4f3;
        src19 <= 12'h4c6;
        src20 <= 12'h610;
        src21 <= 12'h589;
        src22 <= 12'h981;
        src23 <= 12'h6a3;
        src24 <= 12'he27;
        src25 <= 12'h357;
        src26 <= 12'h413;
        src27 <= 12'h9ed;
        src28 <= 12'he28;
        src29 <= 12'h722;
        src30 <= 12'h5e2;
        src31 <= 12'ha05;
        src32 <= 12'h9c7;
        src33 <= 12'h85c;
        src34 <= 12'h6bc;
        src35 <= 12'h6;
        src36 <= 12'he1;
        src37 <= 12'ha39;
        src38 <= 12'h13a;
        src39 <= 12'h3fa;
        src40 <= 12'h4cb;
        src41 <= 12'h7f5;
        src42 <= 12'hf46;
        src43 <= 12'h4ac;
        src44 <= 12'h2ef;
        src45 <= 12'hd9b;
        src46 <= 12'h874;
        src47 <= 12'hf13;
        src48 <= 12'hf72;
        src49 <= 12'hd08;
        src50 <= 12'h610;
        src51 <= 12'h2f8;
        src52 <= 12'h903;
        src53 <= 12'hc9e;
        exp <= 18'h1b1d6;
        #1
        src0 <= 12'h9b7;
        src1 <= 12'h9b4;
        src2 <= 12'hcbd;
        src3 <= 12'h8f;
        src4 <= 12'he1f;
        src5 <= 12'h4f5;
        src6 <= 12'h49d;
        src7 <= 12'he0f;
        src8 <= 12'hd1d;
        src9 <= 12'hd0f;
        src10 <= 12'hd62;
        src11 <= 12'hfc9;
        src12 <= 12'h303;
        src13 <= 12'h778;
        src14 <= 12'hc02;
        src15 <= 12'h257;
        src16 <= 12'h4c4;
        src17 <= 12'hb76;
        src18 <= 12'h583;
        src19 <= 12'h45f;
        src20 <= 12'h97b;
        src21 <= 12'h9b1;
        src22 <= 12'h8cd;
        src23 <= 12'h729;
        src24 <= 12'hf2e;
        src25 <= 12'h576;
        src26 <= 12'h8f8;
        src27 <= 12'h510;
        src28 <= 12'h9a4;
        src29 <= 12'ha94;
        src30 <= 12'h59;
        src31 <= 12'h8a0;
        src32 <= 12'h2be;
        src33 <= 12'h613;
        src34 <= 12'h973;
        src35 <= 12'h4d3;
        src36 <= 12'h8cc;
        src37 <= 12'h431;
        src38 <= 12'h759;
        src39 <= 12'h80c;
        src40 <= 12'h2e2;
        src41 <= 12'he7c;
        src42 <= 12'hb54;
        src43 <= 12'hf6b;
        src44 <= 12'heff;
        src45 <= 12'haa5;
        src46 <= 12'h515;
        src47 <= 12'hd5;
        src48 <= 12'h557;
        src49 <= 12'hf96;
        src50 <= 12'hcd3;
        src51 <= 12'hc47;
        src52 <= 12'ha55;
        src53 <= 12'h52;
        exp <= 18'h1cb8f;
        #1
        src0 <= 12'h900;
        src1 <= 12'h475;
        src2 <= 12'hed2;
        src3 <= 12'h9bd;
        src4 <= 12'h7c4;
        src5 <= 12'h4f8;
        src6 <= 12'h6d7;
        src7 <= 12'h1ca;
        src8 <= 12'h467;
        src9 <= 12'hab2;
        src10 <= 12'h946;
        src11 <= 12'haaf;
        src12 <= 12'heeb;
        src13 <= 12'ha94;
        src14 <= 12'ha6c;
        src15 <= 12'h4cb;
        src16 <= 12'h9b6;
        src17 <= 12'h9d4;
        src18 <= 12'h153;
        src19 <= 12'h79;
        src20 <= 12'h361;
        src21 <= 12'h1fd;
        src22 <= 12'hf54;
        src23 <= 12'h9a8;
        src24 <= 12'hd95;
        src25 <= 12'ha45;
        src26 <= 12'h6cb;
        src27 <= 12'he22;
        src28 <= 12'hf1c;
        src29 <= 12'hd03;
        src30 <= 12'h6ff;
        src31 <= 12'h5ed;
        src32 <= 12'h581;
        src33 <= 12'h68a;
        src34 <= 12'hb19;
        src35 <= 12'h7fe;
        src36 <= 12'hdf6;
        src37 <= 12'h19f;
        src38 <= 12'h74f;
        src39 <= 12'h659;
        src40 <= 12'h155;
        src41 <= 12'h1b6;
        src42 <= 12'h8e8;
        src43 <= 12'h2fc;
        src44 <= 12'hc0;
        src45 <= 12'h34a;
        src46 <= 12'he01;
        src47 <= 12'h5f0;
        src48 <= 12'he6a;
        src49 <= 12'h885;
        src50 <= 12'hdbe;
        src51 <= 12'h305;
        src52 <= 12'hd4d;
        src53 <= 12'hd39;
        exp <= 18'h1b628;
        #1
        src0 <= 12'h4b3;
        src1 <= 12'h221;
        src2 <= 12'h3b1;
        src3 <= 12'ha7f;
        src4 <= 12'h2a;
        src5 <= 12'hc18;
        src6 <= 12'h563;
        src7 <= 12'h3ab;
        src8 <= 12'hac2;
        src9 <= 12'h69;
        src10 <= 12'h4e;
        src11 <= 12'hba8;
        src12 <= 12'h179;
        src13 <= 12'he44;
        src14 <= 12'hb0;
        src15 <= 12'h6d2;
        src16 <= 12'h8b8;
        src17 <= 12'h452;
        src18 <= 12'h6e7;
        src19 <= 12'h8a9;
        src20 <= 12'hb14;
        src21 <= 12'h91;
        src22 <= 12'h62a;
        src23 <= 12'h80a;
        src24 <= 12'h447;
        src25 <= 12'h44d;
        src26 <= 12'h8dd;
        src27 <= 12'h484;
        src28 <= 12'h9ee;
        src29 <= 12'h2d1;
        src30 <= 12'hf28;
        src31 <= 12'h8fd;
        src32 <= 12'h671;
        src33 <= 12'h601;
        src34 <= 12'haff;
        src35 <= 12'h9bc;
        src36 <= 12'hd17;
        src37 <= 12'h7a9;
        src38 <= 12'h1c2;
        src39 <= 12'h92;
        src40 <= 12'h9bc;
        src41 <= 12'hc15;
        src42 <= 12'hde0;
        src43 <= 12'h7c0;
        src44 <= 12'he95;
        src45 <= 12'hc65;
        src46 <= 12'h7c3;
        src47 <= 12'h9d1;
        src48 <= 12'h9e3;
        src49 <= 12'h60f;
        src50 <= 12'h67;
        src51 <= 12'h2d9;
        src52 <= 12'hac4;
        src53 <= 12'h60b;
        exp <= 18'h17e41;
        #1
        src0 <= 12'h7bc;
        src1 <= 12'h30e;
        src2 <= 12'h772;
        src3 <= 12'hc10;
        src4 <= 12'hef5;
        src5 <= 12'h9fb;
        src6 <= 12'h561;
        src7 <= 12'hafb;
        src8 <= 12'h4b3;
        src9 <= 12'h734;
        src10 <= 12'h2fb;
        src11 <= 12'h243;
        src12 <= 12'h846;
        src13 <= 12'he0;
        src14 <= 12'h3c2;
        src15 <= 12'h75d;
        src16 <= 12'h814;
        src17 <= 12'h66a;
        src18 <= 12'h1fa;
        src19 <= 12'hcfd;
        src20 <= 12'h923;
        src21 <= 12'h700;
        src22 <= 12'h1da;
        src23 <= 12'h7d;
        src24 <= 12'h9a6;
        src25 <= 12'h49d;
        src26 <= 12'h78f;
        src27 <= 12'hafc;
        src28 <= 12'h237;
        src29 <= 12'hdd9;
        src30 <= 12'hda1;
        src31 <= 12'h9c0;
        src32 <= 12'hfe;
        src33 <= 12'h594;
        src34 <= 12'he21;
        src35 <= 12'h6b3;
        src36 <= 12'hc90;
        src37 <= 12'hb10;
        src38 <= 12'h4a5;
        src39 <= 12'hecd;
        src40 <= 12'haef;
        src41 <= 12'hcab;
        src42 <= 12'h2c0;
        src43 <= 12'hdab;
        src44 <= 12'he68;
        src45 <= 12'h7c9;
        src46 <= 12'h1e5;
        src47 <= 12'hb3c;
        src48 <= 12'h8f2;
        src49 <= 12'ha9b;
        src50 <= 12'h8a5;
        src51 <= 12'h2e4;
        src52 <= 12'h98f;
        src53 <= 12'ha0d;
        exp <= 18'h1a9b1;
        #1
        src0 <= 12'h974;
        src1 <= 12'h9d;
        src2 <= 12'ha33;
        src3 <= 12'ha41;
        src4 <= 12'h73a;
        src5 <= 12'hc65;
        src6 <= 12'hc7e;
        src7 <= 12'h126;
        src8 <= 12'h62c;
        src9 <= 12'h24;
        src10 <= 12'h675;
        src11 <= 12'hfc4;
        src12 <= 12'hd3e;
        src13 <= 12'h629;
        src14 <= 12'h35;
        src15 <= 12'h4d5;
        src16 <= 12'h311;
        src17 <= 12'he63;
        src18 <= 12'hf66;
        src19 <= 12'hb0e;
        src20 <= 12'h534;
        src21 <= 12'h60d;
        src22 <= 12'hfb8;
        src23 <= 12'hace;
        src24 <= 12'h150;
        src25 <= 12'hc0f;
        src26 <= 12'h2f3;
        src27 <= 12'h822;
        src28 <= 12'h99a;
        src29 <= 12'h38e;
        src30 <= 12'h3ee;
        src31 <= 12'h257;
        src32 <= 12'h9d2;
        src33 <= 12'ha6b;
        src34 <= 12'h53c;
        src35 <= 12'h2f0;
        src36 <= 12'h86d;
        src37 <= 12'h69b;
        src38 <= 12'h425;
        src39 <= 12'h75;
        src40 <= 12'hf52;
        src41 <= 12'ha44;
        src42 <= 12'h750;
        src43 <= 12'hfc9;
        src44 <= 12'h324;
        src45 <= 12'hccd;
        src46 <= 12'h90d;
        src47 <= 12'hd5d;
        src48 <= 12'hf68;
        src49 <= 12'h59b;
        src50 <= 12'heeb;
        src51 <= 12'hec8;
        src52 <= 12'h3d;
        src53 <= 12'h4bc;
        exp <= 18'h1b116;
        #1
        src0 <= 12'h9f5;
        src1 <= 12'h711;
        src2 <= 12'h86f;
        src3 <= 12'heb0;
        src4 <= 12'h994;
        src5 <= 12'h7a8;
        src6 <= 12'h8e5;
        src7 <= 12'h75b;
        src8 <= 12'h3ae;
        src9 <= 12'hd12;
        src10 <= 12'h625;
        src11 <= 12'h52a;
        src12 <= 12'he99;
        src13 <= 12'h575;
        src14 <= 12'h57e;
        src15 <= 12'h964;
        src16 <= 12'h1db;
        src17 <= 12'h32;
        src18 <= 12'h5e2;
        src19 <= 12'he3d;
        src20 <= 12'h3db;
        src21 <= 12'hae2;
        src22 <= 12'h356;
        src23 <= 12'h51a;
        src24 <= 12'h4c6;
        src25 <= 12'h90b;
        src26 <= 12'h27d;
        src27 <= 12'hdf5;
        src28 <= 12'hc39;
        src29 <= 12'hc5e;
        src30 <= 12'h874;
        src31 <= 12'h5d6;
        src32 <= 12'ha3d;
        src33 <= 12'h4c4;
        src34 <= 12'h21;
        src35 <= 12'h1cf;
        src36 <= 12'h617;
        src37 <= 12'h75d;
        src38 <= 12'h85e;
        src39 <= 12'h73a;
        src40 <= 12'h57a;
        src41 <= 12'h624;
        src42 <= 12'h24a;
        src43 <= 12'haad;
        src44 <= 12'hd81;
        src45 <= 12'h72c;
        src46 <= 12'hbf7;
        src47 <= 12'hc16;
        src48 <= 12'hfbc;
        src49 <= 12'hee7;
        src50 <= 12'ha60;
        src51 <= 12'hbcb;
        src52 <= 12'h94;
        src53 <= 12'h9e2;
        exp <= 18'h1adad;
        #1
        src0 <= 12'h289;
        src1 <= 12'h9dd;
        src2 <= 12'h2c1;
        src3 <= 12'hc0a;
        src4 <= 12'h1e6;
        src5 <= 12'h528;
        src6 <= 12'h1c5;
        src7 <= 12'hc59;
        src8 <= 12'he86;
        src9 <= 12'h69d;
        src10 <= 12'hac9;
        src11 <= 12'hf15;
        src12 <= 12'h718;
        src13 <= 12'hd35;
        src14 <= 12'ha28;
        src15 <= 12'h1af;
        src16 <= 12'h70a;
        src17 <= 12'hfd5;
        src18 <= 12'h838;
        src19 <= 12'hf9a;
        src20 <= 12'hedc;
        src21 <= 12'h356;
        src22 <= 12'h6fa;
        src23 <= 12'he65;
        src24 <= 12'hc21;
        src25 <= 12'h71c;
        src26 <= 12'h5f7;
        src27 <= 12'hf58;
        src28 <= 12'h818;
        src29 <= 12'h579;
        src30 <= 12'h50a;
        src31 <= 12'h58e;
        src32 <= 12'h48;
        src33 <= 12'had;
        src34 <= 12'h4c9;
        src35 <= 12'h64a;
        src36 <= 12'h968;
        src37 <= 12'h6a6;
        src38 <= 12'hc4c;
        src39 <= 12'h633;
        src40 <= 12'had5;
        src41 <= 12'h89c;
        src42 <= 12'hd89;
        src43 <= 12'h14e;
        src44 <= 12'h54d;
        src45 <= 12'hd4c;
        src46 <= 12'h69f;
        src47 <= 12'h20b;
        src48 <= 12'h114;
        src49 <= 12'h6bc;
        src50 <= 12'h49b;
        src51 <= 12'he31;
        src52 <= 12'h3ac;
        src53 <= 12'h23f;
        exp <= 18'h1a320;
        #1
        src0 <= 12'h4a4;
        src1 <= 12'h51d;
        src2 <= 12'hf5a;
        src3 <= 12'hb92;
        src4 <= 12'h79c;
        src5 <= 12'h321;
        src6 <= 12'ha7a;
        src7 <= 12'h491;
        src8 <= 12'h4ad;
        src9 <= 12'hcf7;
        src10 <= 12'hd89;
        src11 <= 12'h5cc;
        src12 <= 12'h25d;
        src13 <= 12'hc62;
        src14 <= 12'h8bb;
        src15 <= 12'h87e;
        src16 <= 12'h75e;
        src17 <= 12'h5d1;
        src18 <= 12'hc3d;
        src19 <= 12'h5e9;
        src20 <= 12'hb8e;
        src21 <= 12'hc51;
        src22 <= 12'h134;
        src23 <= 12'h35;
        src24 <= 12'h3b9;
        src25 <= 12'h43b;
        src26 <= 12'h7ff;
        src27 <= 12'he62;
        src28 <= 12'hbc6;
        src29 <= 12'h92b;
        src30 <= 12'hde3;
        src31 <= 12'hcf2;
        src32 <= 12'h48d;
        src33 <= 12'h29a;
        src34 <= 12'h196;
        src35 <= 12'h8d8;
        src36 <= 12'h872;
        src37 <= 12'h55f;
        src38 <= 12'hfe1;
        src39 <= 12'h888;
        src40 <= 12'ha82;
        src41 <= 12'had3;
        src42 <= 12'ha20;
        src43 <= 12'hbec;
        src44 <= 12'ha1b;
        src45 <= 12'h32c;
        src46 <= 12'h7e5;
        src47 <= 12'h89d;
        src48 <= 12'hfdb;
        src49 <= 12'h83e;
        src50 <= 12'hf9e;
        src51 <= 12'hc47;
        src52 <= 12'h10c;
        src53 <= 12'h358;
        exp <= 18'h1c379;
        #1
        src0 <= 12'h742;
        src1 <= 12'h851;
        src2 <= 12'h9c3;
        src3 <= 12'h809;
        src4 <= 12'h2fa;
        src5 <= 12'ha66;
        src6 <= 12'h31c;
        src7 <= 12'hcf7;
        src8 <= 12'h890;
        src9 <= 12'h6de;
        src10 <= 12'hd85;
        src11 <= 12'h948;
        src12 <= 12'h577;
        src13 <= 12'hd17;
        src14 <= 12'hb11;
        src15 <= 12'h197;
        src16 <= 12'h807;
        src17 <= 12'h7ae;
        src18 <= 12'h9a5;
        src19 <= 12'h396;
        src20 <= 12'h608;
        src21 <= 12'h58d;
        src22 <= 12'hb36;
        src23 <= 12'h5ed;
        src24 <= 12'h356;
        src25 <= 12'h2cc;
        src26 <= 12'h3b8;
        src27 <= 12'h9cb;
        src28 <= 12'h3e;
        src29 <= 12'h2ae;
        src30 <= 12'h5d1;
        src31 <= 12'h841;
        src32 <= 12'hd55;
        src33 <= 12'hc11;
        src34 <= 12'h354;
        src35 <= 12'haf6;
        src36 <= 12'h4b;
        src37 <= 12'ha50;
        src38 <= 12'h384;
        src39 <= 12'h394;
        src40 <= 12'h38;
        src41 <= 12'h3c;
        src42 <= 12'h278;
        src43 <= 12'h72c;
        src44 <= 12'he65;
        src45 <= 12'hb1;
        src46 <= 12'ha84;
        src47 <= 12'h2c;
        src48 <= 12'ha78;
        src49 <= 12'hd50;
        src50 <= 12'h69;
        src51 <= 12'h844;
        src52 <= 12'h69c;
        src53 <= 12'h8de;
        exp <= 18'h16fbe;
        #1
        src0 <= 12'hc3d;
        src1 <= 12'h6b6;
        src2 <= 12'ha86;
        src3 <= 12'hf63;
        src4 <= 12'h4;
        src5 <= 12'h38a;
        src6 <= 12'h9d3;
        src7 <= 12'h6f2;
        src8 <= 12'h3a7;
        src9 <= 12'h188;
        src10 <= 12'h8b4;
        src11 <= 12'hd6e;
        src12 <= 12'haa9;
        src13 <= 12'h9d7;
        src14 <= 12'hc0a;
        src15 <= 12'h6a0;
        src16 <= 12'hc34;
        src17 <= 12'h38e;
        src18 <= 12'h47f;
        src19 <= 12'h3b4;
        src20 <= 12'h468;
        src21 <= 12'hb63;
        src22 <= 12'h799;
        src23 <= 12'hbdb;
        src24 <= 12'h115;
        src25 <= 12'h25b;
        src26 <= 12'h813;
        src27 <= 12'hbdb;
        src28 <= 12'h665;
        src29 <= 12'hd4c;
        src30 <= 12'hd0d;
        src31 <= 12'h217;
        src32 <= 12'h6f3;
        src33 <= 12'h167;
        src34 <= 12'hd81;
        src35 <= 12'hd1f;
        src36 <= 12'h584;
        src37 <= 12'hc2e;
        src38 <= 12'hea8;
        src39 <= 12'h958;
        src40 <= 12'hb35;
        src41 <= 12'h3fa;
        src42 <= 12'hef8;
        src43 <= 12'h143;
        src44 <= 12'h97;
        src45 <= 12'hfb4;
        src46 <= 12'h2e9;
        src47 <= 12'h315;
        src48 <= 12'h397;
        src49 <= 12'h390;
        src50 <= 12'h168;
        src51 <= 12'hd17;
        src52 <= 12'he91;
        src53 <= 12'hd20;
        exp <= 18'h1acc7;
        #1
        src0 <= 12'heb7;
        src1 <= 12'h6e;
        src2 <= 12'h2b3;
        src3 <= 12'h7f3;
        src4 <= 12'hc9;
        src5 <= 12'hb7e;
        src6 <= 12'h32c;
        src7 <= 12'hdef;
        src8 <= 12'hb31;
        src9 <= 12'hbd0;
        src10 <= 12'h5cb;
        src11 <= 12'h9f9;
        src12 <= 12'h3bf;
        src13 <= 12'h336;
        src14 <= 12'h4cd;
        src15 <= 12'h9f0;
        src16 <= 12'h128;
        src17 <= 12'hdd9;
        src18 <= 12'h88;
        src19 <= 12'h9b1;
        src20 <= 12'h1e0;
        src21 <= 12'h45e;
        src22 <= 12'h1b8;
        src23 <= 12'h3d4;
        src24 <= 12'h64e;
        src25 <= 12'h493;
        src26 <= 12'h6c9;
        src27 <= 12'hd08;
        src28 <= 12'h5e3;
        src29 <= 12'hcd6;
        src30 <= 12'h775;
        src31 <= 12'hd2f;
        src32 <= 12'hbd7;
        src33 <= 12'heb6;
        src34 <= 12'h867;
        src35 <= 12'h782;
        src36 <= 12'h919;
        src37 <= 12'h869;
        src38 <= 12'hc1e;
        src39 <= 12'hf9d;
        src40 <= 12'hf8c;
        src41 <= 12'h2bc;
        src42 <= 12'h819;
        src43 <= 12'h6a0;
        src44 <= 12'he50;
        src45 <= 12'hc94;
        src46 <= 12'hc19;
        src47 <= 12'h26c;
        src48 <= 12'h4e;
        src49 <= 12'hbd7;
        src50 <= 12'h173;
        src51 <= 12'h578;
        src52 <= 12'h48;
        src53 <= 12'h54c;
        exp <= 18'h19978;
        #1
        src0 <= 12'hdd9;
        src1 <= 12'h199;
        src2 <= 12'h9cf;
        src3 <= 12'h60b;
        src4 <= 12'hdfd;
        src5 <= 12'h5b5;
        src6 <= 12'haf7;
        src7 <= 12'h362;
        src8 <= 12'h9f;
        src9 <= 12'h9d9;
        src10 <= 12'hb90;
        src11 <= 12'hd20;
        src12 <= 12'hbf8;
        src13 <= 12'h963;
        src14 <= 12'hf58;
        src15 <= 12'h8c4;
        src16 <= 12'h7ed;
        src17 <= 12'h13d;
        src18 <= 12'hf3e;
        src19 <= 12'hc25;
        src20 <= 12'h183;
        src21 <= 12'hdf6;
        src22 <= 12'h609;
        src23 <= 12'h649;
        src24 <= 12'h2f4;
        src25 <= 12'h5a8;
        src26 <= 12'h227;
        src27 <= 12'h781;
        src28 <= 12'hfa1;
        src29 <= 12'h967;
        src30 <= 12'h8e8;
        src31 <= 12'h216;
        src32 <= 12'hc62;
        src33 <= 12'h2e2;
        src34 <= 12'h35;
        src35 <= 12'h1de;
        src36 <= 12'he1a;
        src37 <= 12'h91;
        src38 <= 12'h349;
        src39 <= 12'h734;
        src40 <= 12'h522;
        src41 <= 12'hc1;
        src42 <= 12'hb72;
        src43 <= 12'h242;
        src44 <= 12'h710;
        src45 <= 12'hea3;
        src46 <= 12'h758;
        src47 <= 12'h73b;
        src48 <= 12'h7e0;
        src49 <= 12'hf3c;
        src50 <= 12'h5b5;
        src51 <= 12'h887;
        src52 <= 12'h90c;
        src53 <= 12'hb5d;
        exp <= 18'h1a4b5;
        #1
        src0 <= 12'h41d;
        src1 <= 12'hd0;
        src2 <= 12'h298;
        src3 <= 12'ha11;
        src4 <= 12'h8b8;
        src5 <= 12'h81b;
        src6 <= 12'hd9d;
        src7 <= 12'hec1;
        src8 <= 12'hbae;
        src9 <= 12'hbd6;
        src10 <= 12'h691;
        src11 <= 12'h642;
        src12 <= 12'hc2d;
        src13 <= 12'h126;
        src14 <= 12'h179;
        src15 <= 12'hcd3;
        src16 <= 12'hee6;
        src17 <= 12'hb3e;
        src18 <= 12'h821;
        src19 <= 12'h3;
        src20 <= 12'h225;
        src21 <= 12'h28b;
        src22 <= 12'h454;
        src23 <= 12'h555;
        src24 <= 12'hb25;
        src25 <= 12'hb70;
        src26 <= 12'h44f;
        src27 <= 12'hdfd;
        src28 <= 12'h17;
        src29 <= 12'hc35;
        src30 <= 12'heb3;
        src31 <= 12'h57b;
        src32 <= 12'hac5;
        src33 <= 12'h25e;
        src34 <= 12'h69e;
        src35 <= 12'h7c4;
        src36 <= 12'h1b6;
        src37 <= 12'hbbb;
        src38 <= 12'ha9e;
        src39 <= 12'h478;
        src40 <= 12'hc6e;
        src41 <= 12'h770;
        src42 <= 12'h4ea;
        src43 <= 12'hf34;
        src44 <= 12'h33e;
        src45 <= 12'h1ff;
        src46 <= 12'h3c4;
        src47 <= 12'hf81;
        src48 <= 12'hee;
        src49 <= 12'hd67;
        src50 <= 12'h358;
        src51 <= 12'h37e;
        src52 <= 12'h1fb;
        src53 <= 12'h93e;
        exp <= 18'h191a7;
        #1
        src0 <= 12'h95d;
        src1 <= 12'he9c;
        src2 <= 12'hefa;
        src3 <= 12'h56;
        src4 <= 12'h25d;
        src5 <= 12'hf1b;
        src6 <= 12'hbcb;
        src7 <= 12'he76;
        src8 <= 12'hc55;
        src9 <= 12'h980;
        src10 <= 12'h23;
        src11 <= 12'h74a;
        src12 <= 12'h11a;
        src13 <= 12'h824;
        src14 <= 12'he1d;
        src15 <= 12'h44a;
        src16 <= 12'hdfd;
        src17 <= 12'heff;
        src18 <= 12'hadb;
        src19 <= 12'h8e6;
        src20 <= 12'he78;
        src21 <= 12'hbc3;
        src22 <= 12'h26e;
        src23 <= 12'h225;
        src24 <= 12'he58;
        src25 <= 12'hde1;
        src26 <= 12'hd5e;
        src27 <= 12'hf05;
        src28 <= 12'hf72;
        src29 <= 12'h115;
        src30 <= 12'hee2;
        src31 <= 12'hb88;
        src32 <= 12'haf5;
        src33 <= 12'he92;
        src34 <= 12'hfe5;
        src35 <= 12'h9ba;
        src36 <= 12'he4b;
        src37 <= 12'ha20;
        src38 <= 12'hef;
        src39 <= 12'hab9;
        src40 <= 12'h6b7;
        src41 <= 12'hb77;
        src42 <= 12'h8af;
        src43 <= 12'hfff;
        src44 <= 12'he37;
        src45 <= 12'h637;
        src46 <= 12'hba9;
        src47 <= 12'hf4a;
        src48 <= 12'hf2b;
        src49 <= 12'h584;
        src50 <= 12'h3;
        src51 <= 12'hf5;
        src52 <= 12'h11;
        src53 <= 12'h835;
        exp <= 18'h20e64;
        #1
        src0 <= 12'h8b8;
        src1 <= 12'he4c;
        src2 <= 12'h9e8;
        src3 <= 12'h170;
        src4 <= 12'h244;
        src5 <= 12'h985;
        src6 <= 12'h7f4;
        src7 <= 12'hffa;
        src8 <= 12'h431;
        src9 <= 12'hae4;
        src10 <= 12'h26b;
        src11 <= 12'h83;
        src12 <= 12'hc38;
        src13 <= 12'h8bd;
        src14 <= 12'h3b7;
        src15 <= 12'h3e9;
        src16 <= 12'h8c7;
        src17 <= 12'h3af;
        src18 <= 12'h9de;
        src19 <= 12'h326;
        src20 <= 12'h469;
        src21 <= 12'hdfb;
        src22 <= 12'h9d5;
        src23 <= 12'hd59;
        src24 <= 12'hb0f;
        src25 <= 12'h8d0;
        src26 <= 12'haf6;
        src27 <= 12'hd0;
        src28 <= 12'hb17;
        src29 <= 12'h22c;
        src30 <= 12'h59c;
        src31 <= 12'hffd;
        src32 <= 12'h2b3;
        src33 <= 12'hfdc;
        src34 <= 12'h9c7;
        src35 <= 12'he21;
        src36 <= 12'h528;
        src37 <= 12'hdb6;
        src38 <= 12'h60d;
        src39 <= 12'h987;
        src40 <= 12'hd0d;
        src41 <= 12'h351;
        src42 <= 12'h223;
        src43 <= 12'h41d;
        src44 <= 12'hc7c;
        src45 <= 12'hf84;
        src46 <= 12'hbad;
        src47 <= 12'h726;
        src48 <= 12'h814;
        src49 <= 12'hfec;
        src50 <= 12'hdaa;
        src51 <= 12'hf5d;
        src52 <= 12'h678;
        src53 <= 12'ha83;
        exp <= 18'h1d294;
        #1
        src0 <= 12'h55b;
        src1 <= 12'ha97;
        src2 <= 12'h27d;
        src3 <= 12'h50;
        src4 <= 12'hba4;
        src5 <= 12'hb87;
        src6 <= 12'hda7;
        src7 <= 12'h89b;
        src8 <= 12'hf7f;
        src9 <= 12'hf7;
        src10 <= 12'ha5e;
        src11 <= 12'hc17;
        src12 <= 12'hef1;
        src13 <= 12'h95d;
        src14 <= 12'h40;
        src15 <= 12'hbc1;
        src16 <= 12'h4f5;
        src17 <= 12'h120;
        src18 <= 12'h64b;
        src19 <= 12'hf0;
        src20 <= 12'h17e;
        src21 <= 12'hb58;
        src22 <= 12'he90;
        src23 <= 12'he54;
        src24 <= 12'hef5;
        src25 <= 12'h7bd;
        src26 <= 12'hb6b;
        src27 <= 12'h35f;
        src28 <= 12'hefd;
        src29 <= 12'haba;
        src30 <= 12'he24;
        src31 <= 12'h829;
        src32 <= 12'h510;
        src33 <= 12'h542;
        src34 <= 12'h6f0;
        src35 <= 12'hc03;
        src36 <= 12'h675;
        src37 <= 12'h32a;
        src38 <= 12'h512;
        src39 <= 12'h271;
        src40 <= 12'h7b0;
        src41 <= 12'heb6;
        src42 <= 12'h7d7;
        src43 <= 12'hb0f;
        src44 <= 12'h56b;
        src45 <= 12'hfa2;
        src46 <= 12'h141;
        src47 <= 12'h439;
        src48 <= 12'hee;
        src49 <= 12'h529;
        src50 <= 12'h1e0;
        src51 <= 12'ha2c;
        src52 <= 12'h679;
        src53 <= 12'h7bc;
        exp <= 18'h1aa82;
        #1
        src0 <= 12'hcf8;
        src1 <= 12'hb88;
        src2 <= 12'h46e;
        src3 <= 12'hd5a;
        src4 <= 12'ha3d;
        src5 <= 12'h507;
        src6 <= 12'hb67;
        src7 <= 12'h3e4;
        src8 <= 12'h896;
        src9 <= 12'ha85;
        src10 <= 12'h756;
        src11 <= 12'h33f;
        src12 <= 12'hc4e;
        src13 <= 12'hc80;
        src14 <= 12'he6b;
        src15 <= 12'h2a;
        src16 <= 12'h8b2;
        src17 <= 12'haa3;
        src18 <= 12'h2c1;
        src19 <= 12'h7ae;
        src20 <= 12'h176;
        src21 <= 12'hb23;
        src22 <= 12'h993;
        src23 <= 12'h8f0;
        src24 <= 12'h8fd;
        src25 <= 12'hbbf;
        src26 <= 12'h6c3;
        src27 <= 12'hb3c;
        src28 <= 12'hf73;
        src29 <= 12'hdf9;
        src30 <= 12'h33f;
        src31 <= 12'h157;
        src32 <= 12'h17c;
        src33 <= 12'h24c;
        src34 <= 12'h4a0;
        src35 <= 12'h1f9;
        src36 <= 12'h267;
        src37 <= 12'h24a;
        src38 <= 12'hce3;
        src39 <= 12'h450;
        src40 <= 12'hac9;
        src41 <= 12'haae;
        src42 <= 12'hc5;
        src43 <= 12'h2d0;
        src44 <= 12'h62b;
        src45 <= 12'h53e;
        src46 <= 12'h511;
        src47 <= 12'h7a7;
        src48 <= 12'h3ba;
        src49 <= 12'h63f;
        src50 <= 12'h7f9;
        src51 <= 12'hb7c;
        src52 <= 12'h8e1;
        src53 <= 12'h830;
        exp <= 18'h19378;
        #1
        src0 <= 12'h182;
        src1 <= 12'h9e5;
        src2 <= 12'h3f7;
        src3 <= 12'hf62;
        src4 <= 12'hf99;
        src5 <= 12'hedf;
        src6 <= 12'h83f;
        src7 <= 12'h20f;
        src8 <= 12'h1c;
        src9 <= 12'hb5c;
        src10 <= 12'h4c2;
        src11 <= 12'hf8;
        src12 <= 12'ha13;
        src13 <= 12'h800;
        src14 <= 12'hfa8;
        src15 <= 12'h431;
        src16 <= 12'hd34;
        src17 <= 12'h8cc;
        src18 <= 12'h6a0;
        src19 <= 12'hdab;
        src20 <= 12'h8a0;
        src21 <= 12'h58c;
        src22 <= 12'h8a7;
        src23 <= 12'hd3c;
        src24 <= 12'hc33;
        src25 <= 12'hf8a;
        src26 <= 12'h135;
        src27 <= 12'h524;
        src28 <= 12'hec7;
        src29 <= 12'h424;
        src30 <= 12'ha0a;
        src31 <= 12'ha02;
        src32 <= 12'hbde;
        src33 <= 12'hc86;
        src34 <= 12'hc50;
        src35 <= 12'he5f;
        src36 <= 12'h243;
        src37 <= 12'h753;
        src38 <= 12'h7e3;
        src39 <= 12'h8e4;
        src40 <= 12'hb8f;
        src41 <= 12'h6c7;
        src42 <= 12'h6f5;
        src43 <= 12'h3d8;
        src44 <= 12'h93c;
        src45 <= 12'h706;
        src46 <= 12'he;
        src47 <= 12'h610;
        src48 <= 12'h4ee;
        src49 <= 12'hdfd;
        src50 <= 12'ha52;
        src51 <= 12'h2a3;
        src52 <= 12'hfeb;
        src53 <= 12'h435;
        exp <= 18'h1cafe;
        #1
        src0 <= 12'h3a4;
        src1 <= 12'hf7a;
        src2 <= 12'h738;
        src3 <= 12'ha63;
        src4 <= 12'hf84;
        src5 <= 12'hdaa;
        src6 <= 12'h249;
        src7 <= 12'hec1;
        src8 <= 12'hd01;
        src9 <= 12'h28;
        src10 <= 12'h68e;
        src11 <= 12'h807;
        src12 <= 12'heba;
        src13 <= 12'h20;
        src14 <= 12'h1e4;
        src15 <= 12'h808;
        src16 <= 12'h82e;
        src17 <= 12'hdcb;
        src18 <= 12'hc41;
        src19 <= 12'hc92;
        src20 <= 12'h4cc;
        src21 <= 12'he7a;
        src22 <= 12'he23;
        src23 <= 12'hcaf;
        src24 <= 12'hf57;
        src25 <= 12'ha1f;
        src26 <= 12'hfd;
        src27 <= 12'h859;
        src28 <= 12'h6d6;
        src29 <= 12'hdc2;
        src30 <= 12'he29;
        src31 <= 12'h4f9;
        src32 <= 12'hc;
        src33 <= 12'ha49;
        src34 <= 12'hf2d;
        src35 <= 12'h8aa;
        src36 <= 12'he79;
        src37 <= 12'he2;
        src38 <= 12'hbcd;
        src39 <= 12'h53c;
        src40 <= 12'h4f1;
        src41 <= 12'hc6b;
        src42 <= 12'hd98;
        src43 <= 12'h437;
        src44 <= 12'hc02;
        src45 <= 12'h6da;
        src46 <= 12'hefd;
        src47 <= 12'h676;
        src48 <= 12'hc9f;
        src49 <= 12'h212;
        src50 <= 12'h1dd;
        src51 <= 12'h83f;
        src52 <= 12'hb0d;
        src53 <= 12'hd30;
        exp <= 18'h1edf3;
        #1
        src0 <= 12'h407;
        src1 <= 12'haf9;
        src2 <= 12'hbad;
        src3 <= 12'h24d;
        src4 <= 12'hedc;
        src5 <= 12'h539;
        src6 <= 12'h601;
        src7 <= 12'h3f7;
        src8 <= 12'h485;
        src9 <= 12'h978;
        src10 <= 12'h3b9;
        src11 <= 12'hfed;
        src12 <= 12'h34f;
        src13 <= 12'h834;
        src14 <= 12'hd61;
        src15 <= 12'h8cb;
        src16 <= 12'h186;
        src17 <= 12'hf9f;
        src18 <= 12'he4a;
        src19 <= 12'h64a;
        src20 <= 12'h922;
        src21 <= 12'hcfc;
        src22 <= 12'h894;
        src23 <= 12'h8eb;
        src24 <= 12'h1d8;
        src25 <= 12'h68d;
        src26 <= 12'h81d;
        src27 <= 12'h14e;
        src28 <= 12'ha70;
        src29 <= 12'h21a;
        src30 <= 12'hdc5;
        src31 <= 12'hc44;
        src32 <= 12'habf;
        src33 <= 12'hc30;
        src34 <= 12'hf47;
        src35 <= 12'h6a3;
        src36 <= 12'h1b9;
        src37 <= 12'h9c;
        src38 <= 12'h4ba;
        src39 <= 12'he55;
        src40 <= 12'h608;
        src41 <= 12'h144;
        src42 <= 12'h6ef;
        src43 <= 12'h238;
        src44 <= 12'hac8;
        src45 <= 12'hf20;
        src46 <= 12'h56d;
        src47 <= 12'hb7a;
        src48 <= 12'h987;
        src49 <= 12'h72b;
        src50 <= 12'h286;
        src51 <= 12'he51;
        src52 <= 12'hc5d;
        src53 <= 12'h88f;
        exp <= 18'h1b806;
        #1
        src0 <= 12'heaf;
        src1 <= 12'h2e6;
        src2 <= 12'h767;
        src3 <= 12'he4;
        src4 <= 12'hc69;
        src5 <= 12'he8c;
        src6 <= 12'hcf8;
        src7 <= 12'h93c;
        src8 <= 12'h2f8;
        src9 <= 12'hb6e;
        src10 <= 12'h2d1;
        src11 <= 12'he9;
        src12 <= 12'h52;
        src13 <= 12'hd7e;
        src14 <= 12'h32c;
        src15 <= 12'hc1;
        src16 <= 12'hd97;
        src17 <= 12'h18b;
        src18 <= 12'h35c;
        src19 <= 12'ha02;
        src20 <= 12'h81d;
        src21 <= 12'h3fa;
        src22 <= 12'h905;
        src23 <= 12'h286;
        src24 <= 12'ha50;
        src25 <= 12'h88a;
        src26 <= 12'hea9;
        src27 <= 12'h221;
        src28 <= 12'h247;
        src29 <= 12'hbef;
        src30 <= 12'h5ea;
        src31 <= 12'h1c7;
        src32 <= 12'h856;
        src33 <= 12'ha8;
        src34 <= 12'hfde;
        src35 <= 12'he7;
        src36 <= 12'h7d2;
        src37 <= 12'h1c0;
        src38 <= 12'hf93;
        src39 <= 12'h7ad;
        src40 <= 12'h847;
        src41 <= 12'h82e;
        src42 <= 12'h143;
        src43 <= 12'h203;
        src44 <= 12'h7c4;
        src45 <= 12'h8f9;
        src46 <= 12'hd05;
        src47 <= 12'h862;
        src48 <= 12'h80;
        src49 <= 12'h167;
        src50 <= 12'h8a1;
        src51 <= 12'h5bb;
        src52 <= 12'h784;
        src53 <= 12'hd9;
        exp <= 18'h169a7;
        #1
        src0 <= 12'hdb8;
        src1 <= 12'hdfc;
        src2 <= 12'h36c;
        src3 <= 12'h16a;
        src4 <= 12'h30b;
        src5 <= 12'h7ba;
        src6 <= 12'h285;
        src7 <= 12'hf1f;
        src8 <= 12'h6e1;
        src9 <= 12'hd44;
        src10 <= 12'h6fd;
        src11 <= 12'ha20;
        src12 <= 12'ha17;
        src13 <= 12'h955;
        src14 <= 12'ha7;
        src15 <= 12'hadb;
        src16 <= 12'h8ac;
        src17 <= 12'ha45;
        src18 <= 12'h28b;
        src19 <= 12'hd5;
        src20 <= 12'he2a;
        src21 <= 12'h6c7;
        src22 <= 12'hc90;
        src23 <= 12'h695;
        src24 <= 12'h565;
        src25 <= 12'hb84;
        src26 <= 12'hd4f;
        src27 <= 12'hece;
        src28 <= 12'h4dc;
        src29 <= 12'hf91;
        src30 <= 12'hbb5;
        src31 <= 12'he45;
        src32 <= 12'he8e;
        src33 <= 12'hafb;
        src34 <= 12'ha8;
        src35 <= 12'h61d;
        src36 <= 12'hf9a;
        src37 <= 12'h84f;
        src38 <= 12'h9a;
        src39 <= 12'hd12;
        src40 <= 12'hf1;
        src41 <= 12'h5e4;
        src42 <= 12'hcb8;
        src43 <= 12'hf32;
        src44 <= 12'hbe0;
        src45 <= 12'h309;
        src46 <= 12'h205;
        src47 <= 12'h4ae;
        src48 <= 12'h29c;
        src49 <= 12'he1c;
        src50 <= 12'hc3e;
        src51 <= 12'hf41;
        src52 <= 12'hb7b;
        src53 <= 12'h877;
        exp <= 18'h1d95e;
        #1
        src0 <= 12'haa0;
        src1 <= 12'h4fa;
        src2 <= 12'h54d;
        src3 <= 12'h202;
        src4 <= 12'h886;
        src5 <= 12'h6d6;
        src6 <= 12'h82b;
        src7 <= 12'h661;
        src8 <= 12'h5c1;
        src9 <= 12'hed9;
        src10 <= 12'h200;
        src11 <= 12'he53;
        src12 <= 12'h6c5;
        src13 <= 12'h596;
        src14 <= 12'h742;
        src15 <= 12'hfb9;
        src16 <= 12'h68f;
        src17 <= 12'habb;
        src18 <= 12'he60;
        src19 <= 12'hdf8;
        src20 <= 12'h638;
        src21 <= 12'h11c;
        src22 <= 12'h495;
        src23 <= 12'hd6d;
        src24 <= 12'h89a;
        src25 <= 12'h308;
        src26 <= 12'h54f;
        src27 <= 12'h80a;
        src28 <= 12'h49f;
        src29 <= 12'h4fd;
        src30 <= 12'hb7c;
        src31 <= 12'h936;
        src32 <= 12'hfcf;
        src33 <= 12'h735;
        src34 <= 12'h466;
        src35 <= 12'hcf5;
        src36 <= 12'h471;
        src37 <= 12'h90f;
        src38 <= 12'h65f;
        src39 <= 12'h8d4;
        src40 <= 12'hff6;
        src41 <= 12'h6ac;
        src42 <= 12'h23a;
        src43 <= 12'h1d;
        src44 <= 12'hfcf;
        src45 <= 12'h445;
        src46 <= 12'h6e6;
        src47 <= 12'h154;
        src48 <= 12'h95f;
        src49 <= 12'h963;
        src50 <= 12'hfcd;
        src51 <= 12'he00;
        src52 <= 12'h502;
        src53 <= 12'he09;
        exp <= 18'h1b948;
        #1
        src0 <= 12'h329;
        src1 <= 12'h5d2;
        src2 <= 12'h6f6;
        src3 <= 12'hc17;
        src4 <= 12'h39a;
        src5 <= 12'hc1d;
        src6 <= 12'h236;
        src7 <= 12'h26f;
        src8 <= 12'hfa4;
        src9 <= 12'h78c;
        src10 <= 12'hb17;
        src11 <= 12'hd98;
        src12 <= 12'h193;
        src13 <= 12'h271;
        src14 <= 12'h957;
        src15 <= 12'h112;
        src16 <= 12'h9f5;
        src17 <= 12'hefe;
        src18 <= 12'h62c;
        src19 <= 12'hd91;
        src20 <= 12'h613;
        src21 <= 12'hf6;
        src22 <= 12'h89e;
        src23 <= 12'hd42;
        src24 <= 12'h49c;
        src25 <= 12'h489;
        src26 <= 12'hbab;
        src27 <= 12'hc28;
        src28 <= 12'h465;
        src29 <= 12'h922;
        src30 <= 12'hb5e;
        src31 <= 12'h7e2;
        src32 <= 12'hfd;
        src33 <= 12'hcab;
        src34 <= 12'h596;
        src35 <= 12'h9ef;
        src36 <= 12'h4e9;
        src37 <= 12'h78d;
        src38 <= 12'h531;
        src39 <= 12'h20b;
        src40 <= 12'haad;
        src41 <= 12'h75e;
        src42 <= 12'h8b7;
        src43 <= 12'h319;
        src44 <= 12'h623;
        src45 <= 12'h50c;
        src46 <= 12'hcaa;
        src47 <= 12'h75;
        src48 <= 12'hb59;
        src49 <= 12'h42a;
        src50 <= 12'h95f;
        src51 <= 12'h17b;
        src52 <= 12'h75d;
        src53 <= 12'hc6e;
        exp <= 18'h18f38;
        #1
        src0 <= 12'hfb7;
        src1 <= 12'h27a;
        src2 <= 12'h5f6;
        src3 <= 12'hc67;
        src4 <= 12'hb7a;
        src5 <= 12'hab9;
        src6 <= 12'h877;
        src7 <= 12'h328;
        src8 <= 12'h3ec;
        src9 <= 12'hbdd;
        src10 <= 12'h9ce;
        src11 <= 12'h7d4;
        src12 <= 12'h9ca;
        src13 <= 12'h936;
        src14 <= 12'h441;
        src15 <= 12'h99;
        src16 <= 12'hf0b;
        src17 <= 12'ha7e;
        src18 <= 12'hec;
        src19 <= 12'h42a;
        src20 <= 12'h5b4;
        src21 <= 12'habd;
        src22 <= 12'hb27;
        src23 <= 12'hca1;
        src24 <= 12'h355;
        src25 <= 12'h162;
        src26 <= 12'hb13;
        src27 <= 12'hb86;
        src28 <= 12'h210;
        src29 <= 12'ha06;
        src30 <= 12'h53a;
        src31 <= 12'h8a9;
        src32 <= 12'he4b;
        src33 <= 12'hb00;
        src34 <= 12'h890;
        src35 <= 12'h8e7;
        src36 <= 12'h804;
        src37 <= 12'h302;
        src38 <= 12'h3d9;
        src39 <= 12'h427;
        src40 <= 12'hf05;
        src41 <= 12'h56d;
        src42 <= 12'hc12;
        src43 <= 12'h663;
        src44 <= 12'hfcd;
        src45 <= 12'h6e3;
        src46 <= 12'ha1f;
        src47 <= 12'hd22;
        src48 <= 12'hfe3;
        src49 <= 12'h813;
        src50 <= 12'hf5f;
        src51 <= 12'hbf1;
        src52 <= 12'h10e;
        src53 <= 12'h56e;
        exp <= 18'h1c828;
        #1
        src0 <= 12'h795;
        src1 <= 12'h92b;
        src2 <= 12'h476;
        src3 <= 12'hbc6;
        src4 <= 12'hcab;
        src5 <= 12'h228;
        src6 <= 12'h666;
        src7 <= 12'hdae;
        src8 <= 12'h23c;
        src9 <= 12'hcbc;
        src10 <= 12'h1eb;
        src11 <= 12'hb34;
        src12 <= 12'h3a;
        src13 <= 12'hd1a;
        src14 <= 12'h8;
        src15 <= 12'h33;
        src16 <= 12'hcd1;
        src17 <= 12'habe;
        src18 <= 12'hafd;
        src19 <= 12'h981;
        src20 <= 12'h949;
        src21 <= 12'hbfe;
        src22 <= 12'h1ad;
        src23 <= 12'he67;
        src24 <= 12'h46d;
        src25 <= 12'h83b;
        src26 <= 12'h25d;
        src27 <= 12'h606;
        src28 <= 12'h7ac;
        src29 <= 12'h6dd;
        src30 <= 12'hc01;
        src31 <= 12'hadb;
        src32 <= 12'h46f;
        src33 <= 12'h52b;
        src34 <= 12'h7c9;
        src35 <= 12'hff7;
        src36 <= 12'hf60;
        src37 <= 12'h649;
        src38 <= 12'h6;
        src39 <= 12'h2eb;
        src40 <= 12'h91d;
        src41 <= 12'h22a;
        src42 <= 12'ha11;
        src43 <= 12'hcc4;
        src44 <= 12'hfe2;
        src45 <= 12'hb00;
        src46 <= 12'ha39;
        src47 <= 12'h5ce;
        src48 <= 12'h48c;
        src49 <= 12'h7e7;
        src50 <= 12'hd9b;
        src51 <= 12'h21e;
        src52 <= 12'h39b;
        src53 <= 12'h3bc;
        exp <= 18'h1a3dd;
        #1
        src0 <= 12'h753;
        src1 <= 12'h51a;
        src2 <= 12'h8c1;
        src3 <= 12'h86e;
        src4 <= 12'h96a;
        src5 <= 12'h334;
        src6 <= 12'hfe6;
        src7 <= 12'h21c;
        src8 <= 12'hdca;
        src9 <= 12'h38f;
        src10 <= 12'hf2a;
        src11 <= 12'h41f;
        src12 <= 12'hebe;
        src13 <= 12'h87f;
        src14 <= 12'h6fd;
        src15 <= 12'ha55;
        src16 <= 12'ha9e;
        src17 <= 12'h491;
        src18 <= 12'h67c;
        src19 <= 12'hd7b;
        src20 <= 12'hcc7;
        src21 <= 12'hfe0;
        src22 <= 12'hcca;
        src23 <= 12'h2b3;
        src24 <= 12'h3d3;
        src25 <= 12'h4ae;
        src26 <= 12'hfee;
        src27 <= 12'hf3a;
        src28 <= 12'h156;
        src29 <= 12'h45d;
        src30 <= 12'h21d;
        src31 <= 12'hea6;
        src32 <= 12'h6b3;
        src33 <= 12'h32b;
        src34 <= 12'h336;
        src35 <= 12'hcec;
        src36 <= 12'hcb8;
        src37 <= 12'hb7;
        src38 <= 12'h690;
        src39 <= 12'h62f;
        src40 <= 12'h46f;
        src41 <= 12'h3ba;
        src42 <= 12'h67e;
        src43 <= 12'h8e0;
        src44 <= 12'h85e;
        src45 <= 12'ha7b;
        src46 <= 12'h749;
        src47 <= 12'h9b8;
        src48 <= 12'h8bd;
        src49 <= 12'h7b4;
        src50 <= 12'hc6a;
        src51 <= 12'h7fb;
        src52 <= 12'he94;
        src53 <= 12'hb10;
        exp <= 18'h1c4df;
        #1
        src0 <= 12'ha1e;
        src1 <= 12'h378;
        src2 <= 12'h40d;
        src3 <= 12'h676;
        src4 <= 12'heaf;
        src5 <= 12'hfd6;
        src6 <= 12'hcab;
        src7 <= 12'h8bc;
        src8 <= 12'he2d;
        src9 <= 12'hf62;
        src10 <= 12'h7b2;
        src11 <= 12'h918;
        src12 <= 12'he92;
        src13 <= 12'ha44;
        src14 <= 12'h685;
        src15 <= 12'hc4d;
        src16 <= 12'h18d;
        src17 <= 12'h4d1;
        src18 <= 12'h4e9;
        src19 <= 12'hd08;
        src20 <= 12'h97;
        src21 <= 12'h5ee;
        src22 <= 12'he5;
        src23 <= 12'hb71;
        src24 <= 12'h486;
        src25 <= 12'hd4c;
        src26 <= 12'hf83;
        src27 <= 12'h6e1;
        src28 <= 12'h522;
        src29 <= 12'h243;
        src30 <= 12'hb4e;
        src31 <= 12'h1d9;
        src32 <= 12'h30d;
        src33 <= 12'h269;
        src34 <= 12'h820;
        src35 <= 12'h6b9;
        src36 <= 12'h224;
        src37 <= 12'hd27;
        src38 <= 12'h475;
        src39 <= 12'hbea;
        src40 <= 12'h988;
        src41 <= 12'hdce;
        src42 <= 12'hfb4;
        src43 <= 12'h7c;
        src44 <= 12'hf0e;
        src45 <= 12'h325;
        src46 <= 12'hb1d;
        src47 <= 12'h8c7;
        src48 <= 12'h98e;
        src49 <= 12'hb9c;
        src50 <= 12'h8a5;
        src51 <= 12'h74f;
        src52 <= 12'h658;
        src53 <= 12'ha8b;
        exp <= 18'h1c589;
        #1
        src0 <= 12'hc40;
        src1 <= 12'h72e;
        src2 <= 12'hc5d;
        src3 <= 12'h9fe;
        src4 <= 12'h346;
        src5 <= 12'ha73;
        src6 <= 12'hacf;
        src7 <= 12'h643;
        src8 <= 12'h57e;
        src9 <= 12'h81b;
        src10 <= 12'h638;
        src11 <= 12'h6c3;
        src12 <= 12'h956;
        src13 <= 12'hf40;
        src14 <= 12'h77a;
        src15 <= 12'h69f;
        src16 <= 12'h66b;
        src17 <= 12'h5a7;
        src18 <= 12'h277;
        src19 <= 12'hedb;
        src20 <= 12'hb5a;
        src21 <= 12'h95d;
        src22 <= 12'h3b1;
        src23 <= 12'h68b;
        src24 <= 12'hec8;
        src25 <= 12'h168;
        src26 <= 12'h37a;
        src27 <= 12'h77a;
        src28 <= 12'h2ca;
        src29 <= 12'hec3;
        src30 <= 12'h6d7;
        src31 <= 12'hd43;
        src32 <= 12'ha2d;
        src33 <= 12'had1;
        src34 <= 12'hb03;
        src35 <= 12'h7ca;
        src36 <= 12'h6fd;
        src37 <= 12'he86;
        src38 <= 12'h8e;
        src39 <= 12'h7dd;
        src40 <= 12'hb0a;
        src41 <= 12'h9ee;
        src42 <= 12'h648;
        src43 <= 12'ha63;
        src44 <= 12'h1a6;
        src45 <= 12'h69c;
        src46 <= 12'h78e;
        src47 <= 12'h66f;
        src48 <= 12'hc3e;
        src49 <= 12'h41e;
        src50 <= 12'hfa;
        src51 <= 12'hae3;
        src52 <= 12'h47d;
        src53 <= 12'h3fd;
        exp <= 18'h1ad47;
        #1
        src0 <= 12'h2b3;
        src1 <= 12'he77;
        src2 <= 12'h6ab;
        src3 <= 12'h317;
        src4 <= 12'hf70;
        src5 <= 12'h620;
        src6 <= 12'h2f4;
        src7 <= 12'h9ce;
        src8 <= 12'ha15;
        src9 <= 12'h243;
        src10 <= 12'h96;
        src11 <= 12'hc63;
        src12 <= 12'h5;
        src13 <= 12'h59;
        src14 <= 12'h903;
        src15 <= 12'h9e6;
        src16 <= 12'h490;
        src17 <= 12'h262;
        src18 <= 12'hd34;
        src19 <= 12'ha5b;
        src20 <= 12'he0a;
        src21 <= 12'h247;
        src22 <= 12'h577;
        src23 <= 12'h2f7;
        src24 <= 12'h10b;
        src25 <= 12'h2f2;
        src26 <= 12'h7b4;
        src27 <= 12'h43c;
        src28 <= 12'h531;
        src29 <= 12'h43f;
        src30 <= 12'he9c;
        src31 <= 12'ha8b;
        src32 <= 12'he7c;
        src33 <= 12'h664;
        src34 <= 12'h3bd;
        src35 <= 12'hae7;
        src36 <= 12'h6e3;
        src37 <= 12'hd46;
        src38 <= 12'h58c;
        src39 <= 12'h7ec;
        src40 <= 12'h1c7;
        src41 <= 12'h458;
        src42 <= 12'hfa6;
        src43 <= 12'h480;
        src44 <= 12'h8be;
        src45 <= 12'h1fe;
        src46 <= 12'hc5b;
        src47 <= 12'hd1;
        src48 <= 12'hc4d;
        src49 <= 12'h245;
        src50 <= 12'h10;
        src51 <= 12'hb2f;
        src52 <= 12'hedb;
        src53 <= 12'h492;
        exp <= 18'h1782a;
        #1
        src0 <= 12'hd5e;
        src1 <= 12'h64e;
        src2 <= 12'h67a;
        src3 <= 12'h8f;
        src4 <= 12'h45d;
        src5 <= 12'h2d7;
        src6 <= 12'h57c;
        src7 <= 12'h8db;
        src8 <= 12'h3be;
        src9 <= 12'hebe;
        src10 <= 12'hb98;
        src11 <= 12'hf93;
        src12 <= 12'h358;
        src13 <= 12'hc69;
        src14 <= 12'hf5b;
        src15 <= 12'h5a9;
        src16 <= 12'hd16;
        src17 <= 12'h527;
        src18 <= 12'h43;
        src19 <= 12'hef8;
        src20 <= 12'h9b1;
        src21 <= 12'h73e;
        src22 <= 12'h37e;
        src23 <= 12'h4de;
        src24 <= 12'h4dc;
        src25 <= 12'heb8;
        src26 <= 12'h6db;
        src27 <= 12'h174;
        src28 <= 12'h73d;
        src29 <= 12'hb7b;
        src30 <= 12'hae7;
        src31 <= 12'h416;
        src32 <= 12'hdef;
        src33 <= 12'h15f;
        src34 <= 12'h5ef;
        src35 <= 12'hf05;
        src36 <= 12'hfe3;
        src37 <= 12'hd63;
        src38 <= 12'h811;
        src39 <= 12'h668;
        src40 <= 12'he02;
        src41 <= 12'he14;
        src42 <= 12'he61;
        src43 <= 12'hbb9;
        src44 <= 12'h1b2;
        src45 <= 12'hda3;
        src46 <= 12'hd4a;
        src47 <= 12'h8de;
        src48 <= 12'hc6f;
        src49 <= 12'h208;
        src50 <= 12'he5b;
        src51 <= 12'h235;
        src52 <= 12'h1a3;
        src53 <= 12'ha4b;
        exp <= 18'h1d1aa;
        #1
        src0 <= 12'h50a;
        src1 <= 12'h5b0;
        src2 <= 12'he9e;
        src3 <= 12'h4e2;
        src4 <= 12'h1d1;
        src5 <= 12'hbb5;
        src6 <= 12'h72f;
        src7 <= 12'h9e0;
        src8 <= 12'hc65;
        src9 <= 12'h628;
        src10 <= 12'hbd4;
        src11 <= 12'ha34;
        src12 <= 12'h837;
        src13 <= 12'hca3;
        src14 <= 12'hf1a;
        src15 <= 12'h379;
        src16 <= 12'h2a3;
        src17 <= 12'hf0;
        src18 <= 12'hc4a;
        src19 <= 12'hd31;
        src20 <= 12'h69;
        src21 <= 12'h84c;
        src22 <= 12'h704;
        src23 <= 12'h3f2;
        src24 <= 12'h17f;
        src25 <= 12'h65b;
        src26 <= 12'hf08;
        src27 <= 12'h3d4;
        src28 <= 12'hcae;
        src29 <= 12'hbae;
        src30 <= 12'h934;
        src31 <= 12'hf0f;
        src32 <= 12'h8b2;
        src33 <= 12'hfda;
        src34 <= 12'hcb2;
        src35 <= 12'h4f1;
        src36 <= 12'hf9;
        src37 <= 12'h4f1;
        src38 <= 12'h9d7;
        src39 <= 12'h982;
        src40 <= 12'h3e9;
        src41 <= 12'h1f3;
        src42 <= 12'hd81;
        src43 <= 12'h7fb;
        src44 <= 12'hb3d;
        src45 <= 12'hb7d;
        src46 <= 12'h1b;
        src47 <= 12'h25f;
        src48 <= 12'h810;
        src49 <= 12'hb8f;
        src50 <= 12'h931;
        src51 <= 12'h115;
        src52 <= 12'h9ef;
        src53 <= 12'h8e9;
        exp <= 18'h1b19a;
        #1
        src0 <= 12'h544;
        src1 <= 12'hbbf;
        src2 <= 12'h48b;
        src3 <= 12'haae;
        src4 <= 12'h385;
        src5 <= 12'hf2a;
        src6 <= 12'h95a;
        src7 <= 12'hf5b;
        src8 <= 12'hf99;
        src9 <= 12'ha8e;
        src10 <= 12'h65b;
        src11 <= 12'h724;
        src12 <= 12'hab6;
        src13 <= 12'hd0d;
        src14 <= 12'h61a;
        src15 <= 12'h49e;
        src16 <= 12'hcc8;
        src17 <= 12'h6bd;
        src18 <= 12'h83;
        src19 <= 12'ha96;
        src20 <= 12'hc8e;
        src21 <= 12'h481;
        src22 <= 12'h930;
        src23 <= 12'h17a;
        src24 <= 12'h2a;
        src25 <= 12'hd5b;
        src26 <= 12'hcf9;
        src27 <= 12'hace;
        src28 <= 12'h5a7;
        src29 <= 12'h120;
        src30 <= 12'h99f;
        src31 <= 12'h79b;
        src32 <= 12'hc87;
        src33 <= 12'h748;
        src34 <= 12'h659;
        src35 <= 12'h184;
        src36 <= 12'h78e;
        src37 <= 12'hdee;
        src38 <= 12'hf0;
        src39 <= 12'hc17;
        src40 <= 12'h7b;
        src41 <= 12'h92;
        src42 <= 12'hdee;
        src43 <= 12'h248;
        src44 <= 12'h57f;
        src45 <= 12'hb00;
        src46 <= 12'he9a;
        src47 <= 12'h8b8;
        src48 <= 12'hfaf;
        src49 <= 12'hfd8;
        src50 <= 12'h7e3;
        src51 <= 12'h941;
        src52 <= 12'ha60;
        src53 <= 12'hdbf;
        exp <= 18'h1cd72;
        #1
        src0 <= 12'he2c;
        src1 <= 12'h70d;
        src2 <= 12'hd7;
        src3 <= 12'h395;
        src4 <= 12'h5ee;
        src5 <= 12'hc48;
        src6 <= 12'h99;
        src7 <= 12'hbc2;
        src8 <= 12'h74d;
        src9 <= 12'ha3;
        src10 <= 12'h112;
        src11 <= 12'h76;
        src12 <= 12'hd8e;
        src13 <= 12'h430;
        src14 <= 12'haa5;
        src15 <= 12'h799;
        src16 <= 12'h242;
        src17 <= 12'h539;
        src18 <= 12'h3d9;
        src19 <= 12'h873;
        src20 <= 12'ha97;
        src21 <= 12'hdf6;
        src22 <= 12'hbaf;
        src23 <= 12'hc1;
        src24 <= 12'hcc0;
        src25 <= 12'had9;
        src26 <= 12'hf85;
        src27 <= 12'h8ac;
        src28 <= 12'h6c2;
        src29 <= 12'h9c8;
        src30 <= 12'he49;
        src31 <= 12'h15b;
        src32 <= 12'h5a8;
        src33 <= 12'h847;
        src34 <= 12'hd70;
        src35 <= 12'hc7c;
        src36 <= 12'h8a2;
        src37 <= 12'he5c;
        src38 <= 12'hde1;
        src39 <= 12'h41;
        src40 <= 12'h4da;
        src41 <= 12'hc21;
        src42 <= 12'h92c;
        src43 <= 12'h1b8;
        src44 <= 12'h643;
        src45 <= 12'h317;
        src46 <= 12'h264;
        src47 <= 12'h493;
        src48 <= 12'hafa;
        src49 <= 12'hd28;
        src50 <= 12'hab5;
        src51 <= 12'h9b7;
        src52 <= 12'hc0;
        src53 <= 12'hf6d;
        exp <= 18'h1a44c;
        #1
        src0 <= 12'h4d1;
        src1 <= 12'h94b;
        src2 <= 12'h5ab;
        src3 <= 12'he36;
        src4 <= 12'ha74;
        src5 <= 12'h791;
        src6 <= 12'h213;
        src7 <= 12'h22a;
        src8 <= 12'h2cd;
        src9 <= 12'h3ef;
        src10 <= 12'hb4c;
        src11 <= 12'h5f5;
        src12 <= 12'hbe7;
        src13 <= 12'h6e4;
        src14 <= 12'h3db;
        src15 <= 12'h4d6;
        src16 <= 12'hcd;
        src17 <= 12'ha4f;
        src18 <= 12'hf81;
        src19 <= 12'h575;
        src20 <= 12'hf0b;
        src21 <= 12'hc58;
        src22 <= 12'h1a7;
        src23 <= 12'h38b;
        src24 <= 12'h354;
        src25 <= 12'hc8c;
        src26 <= 12'hdfc;
        src27 <= 12'hfda;
        src28 <= 12'h20b;
        src29 <= 12'hd93;
        src30 <= 12'h36c;
        src31 <= 12'h93;
        src32 <= 12'he47;
        src33 <= 12'h8d1;
        src34 <= 12'h9e8;
        src35 <= 12'hafa;
        src36 <= 12'h14;
        src37 <= 12'hbc2;
        src38 <= 12'h5c2;
        src39 <= 12'h716;
        src40 <= 12'hed5;
        src41 <= 12'h468;
        src42 <= 12'h8c4;
        src43 <= 12'h47e;
        src44 <= 12'hdd3;
        src45 <= 12'h32;
        src46 <= 12'h9c4;
        src47 <= 12'hcd3;
        src48 <= 12'h3cf;
        src49 <= 12'he84;
        src50 <= 12'h5e5;
        src51 <= 12'h68d;
        src52 <= 12'hbb9;
        src53 <= 12'hc37;
        exp <= 18'h1ae2a;
        #1
        src0 <= 12'hb63;
        src1 <= 12'h557;
        src2 <= 12'h1aa;
        src3 <= 12'h344;
        src4 <= 12'hea;
        src5 <= 12'hafe;
        src6 <= 12'h665;
        src7 <= 12'h4b;
        src8 <= 12'hc5c;
        src9 <= 12'hacf;
        src10 <= 12'h62e;
        src11 <= 12'hf55;
        src12 <= 12'hfdd;
        src13 <= 12'he56;
        src14 <= 12'ha83;
        src15 <= 12'hc00;
        src16 <= 12'h77b;
        src17 <= 12'h9f4;
        src18 <= 12'h5af;
        src19 <= 12'hcfc;
        src20 <= 12'h985;
        src21 <= 12'haea;
        src22 <= 12'h69;
        src23 <= 12'h79a;
        src24 <= 12'hc58;
        src25 <= 12'h4a0;
        src26 <= 12'h6cc;
        src27 <= 12'h3d6;
        src28 <= 12'hb72;
        src29 <= 12'h9ec;
        src30 <= 12'hdb5;
        src31 <= 12'hb16;
        src32 <= 12'h258;
        src33 <= 12'h8e0;
        src34 <= 12'h6e3;
        src35 <= 12'hd5f;
        src36 <= 12'h94c;
        src37 <= 12'hc1a;
        src38 <= 12'h828;
        src39 <= 12'h71b;
        src40 <= 12'h3d7;
        src41 <= 12'h11;
        src42 <= 12'h41f;
        src43 <= 12'h50;
        src44 <= 12'hbae;
        src45 <= 12'h78e;
        src46 <= 12'he8;
        src47 <= 12'h16c;
        src48 <= 12'haa9;
        src49 <= 12'h812;
        src50 <= 12'hf22;
        src51 <= 12'hc0b;
        src52 <= 12'hefb;
        src53 <= 12'h60b;
        exp <= 18'h1b8eb;
        #1
        src0 <= 12'h465;
        src1 <= 12'hafa;
        src2 <= 12'h157;
        src3 <= 12'hda6;
        src4 <= 12'h6bf;
        src5 <= 12'h5ea;
        src6 <= 12'h7f2;
        src7 <= 12'ha20;
        src8 <= 12'h586;
        src9 <= 12'hfd5;
        src10 <= 12'h883;
        src11 <= 12'h6f0;
        src12 <= 12'hb4e;
        src13 <= 12'h98e;
        src14 <= 12'h7b2;
        src15 <= 12'hbb0;
        src16 <= 12'h94b;
        src17 <= 12'h379;
        src18 <= 12'haaf;
        src19 <= 12'h8d5;
        src20 <= 12'h742;
        src21 <= 12'h78b;
        src22 <= 12'h4f7;
        src23 <= 12'h4d2;
        src24 <= 12'h286;
        src25 <= 12'h99;
        src26 <= 12'hdd3;
        src27 <= 12'h4;
        src28 <= 12'hea9;
        src29 <= 12'hbf7;
        src30 <= 12'h5c6;
        src31 <= 12'heb9;
        src32 <= 12'h2c6;
        src33 <= 12'he0d;
        src34 <= 12'hc73;
        src35 <= 12'h869;
        src36 <= 12'h229;
        src37 <= 12'hb59;
        src38 <= 12'h81d;
        src39 <= 12'hf17;
        src40 <= 12'h8b1;
        src41 <= 12'h8ae;
        src42 <= 12'h9c6;
        src43 <= 12'hf75;
        src44 <= 12'he65;
        src45 <= 12'h440;
        src46 <= 12'hb65;
        src47 <= 12'h9bd;
        src48 <= 12'h9e8;
        src49 <= 12'hf95;
        src50 <= 12'hafc;
        src51 <= 12'hcaf;
        src52 <= 12'h374;
        src53 <= 12'h5a0;
        exp <= 18'h1da18;
        #1
        src0 <= 12'h3f9;
        src1 <= 12'h187;
        src2 <= 12'h94d;
        src3 <= 12'hd11;
        src4 <= 12'h28;
        src5 <= 12'h906;
        src6 <= 12'h24d;
        src7 <= 12'h8ea;
        src8 <= 12'hcdf;
        src9 <= 12'hd6;
        src10 <= 12'h674;
        src11 <= 12'hac0;
        src12 <= 12'h40d;
        src13 <= 12'hf4f;
        src14 <= 12'hb11;
        src15 <= 12'h64b;
        src16 <= 12'hdf;
        src17 <= 12'h5ee;
        src18 <= 12'h66a;
        src19 <= 12'h1f7;
        src20 <= 12'h107;
        src21 <= 12'h80b;
        src22 <= 12'hda6;
        src23 <= 12'h97d;
        src24 <= 12'h301;
        src25 <= 12'h325;
        src26 <= 12'ha10;
        src27 <= 12'h793;
        src28 <= 12'h478;
        src29 <= 12'h9e7;
        src30 <= 12'hc40;
        src31 <= 12'h480;
        src32 <= 12'h94c;
        src33 <= 12'h464;
        src34 <= 12'h2e;
        src35 <= 12'h3bc;
        src36 <= 12'h91c;
        src37 <= 12'h6a1;
        src38 <= 12'hc3b;
        src39 <= 12'hb82;
        src40 <= 12'h4a7;
        src41 <= 12'hb1a;
        src42 <= 12'heeb;
        src43 <= 12'he16;
        src44 <= 12'hbb8;
        src45 <= 12'h710;
        src46 <= 12'h507;
        src47 <= 12'ha7c;
        src48 <= 12'h192;
        src49 <= 12'h64;
        src50 <= 12'h904;
        src51 <= 12'hf25;
        src52 <= 12'hf6;
        src53 <= 12'h5ec;
        exp <= 18'h18351;
        #1
        src0 <= 12'h2fe;
        src1 <= 12'he70;
        src2 <= 12'hac5;
        src3 <= 12'h88e;
        src4 <= 12'hdf2;
        src5 <= 12'h4f0;
        src6 <= 12'h800;
        src7 <= 12'h385;
        src8 <= 12'h141;
        src9 <= 12'hd90;
        src10 <= 12'h467;
        src11 <= 12'h465;
        src12 <= 12'h613;
        src13 <= 12'h440;
        src14 <= 12'ha50;
        src15 <= 12'h589;
        src16 <= 12'h7c0;
        src17 <= 12'h93b;
        src18 <= 12'hfbc;
        src19 <= 12'h40b;
        src20 <= 12'h9e5;
        src21 <= 12'h7df;
        src22 <= 12'h72;
        src23 <= 12'h974;
        src24 <= 12'h487;
        src25 <= 12'h46b;
        src26 <= 12'h671;
        src27 <= 12'h241;
        src28 <= 12'h1f3;
        src29 <= 12'h63;
        src30 <= 12'h1a1;
        src31 <= 12'h404;
        src32 <= 12'h90;
        src33 <= 12'h798;
        src34 <= 12'h9c1;
        src35 <= 12'h83a;
        src36 <= 12'h168;
        src37 <= 12'h59b;
        src38 <= 12'hc4f;
        src39 <= 12'h7c9;
        src40 <= 12'hea1;
        src41 <= 12'h81b;
        src42 <= 12'hd2f;
        src43 <= 12'hc4c;
        src44 <= 12'hc9b;
        src45 <= 12'heab;
        src46 <= 12'h811;
        src47 <= 12'hac0;
        src48 <= 12'h212;
        src49 <= 12'hbe4;
        src50 <= 12'h844;
        src51 <= 12'h7b2;
        src52 <= 12'h269;
        src53 <= 12'hb61;
        exp <= 18'h18e3e;
        #1
        src0 <= 12'h810;
        src1 <= 12'hc39;
        src2 <= 12'h76d;
        src3 <= 12'ha99;
        src4 <= 12'hda0;
        src5 <= 12'hf9d;
        src6 <= 12'h7fc;
        src7 <= 12'he09;
        src8 <= 12'hdd2;
        src9 <= 12'hfcd;
        src10 <= 12'h623;
        src11 <= 12'h2d6;
        src12 <= 12'h830;
        src13 <= 12'ha4c;
        src14 <= 12'hd24;
        src15 <= 12'hb44;
        src16 <= 12'hdb1;
        src17 <= 12'hc43;
        src18 <= 12'h917;
        src19 <= 12'hbbf;
        src20 <= 12'hdf;
        src21 <= 12'hfca;
        src22 <= 12'hc6e;
        src23 <= 12'h2aa;
        src24 <= 12'ha9b;
        src25 <= 12'hb7f;
        src26 <= 12'h52b;
        src27 <= 12'heba;
        src28 <= 12'h1ab;
        src29 <= 12'h5c0;
        src30 <= 12'h2af;
        src31 <= 12'h9f0;
        src32 <= 12'h800;
        src33 <= 12'ha9;
        src34 <= 12'h359;
        src35 <= 12'hbcc;
        src36 <= 12'h3a4;
        src37 <= 12'h934;
        src38 <= 12'h2fd;
        src39 <= 12'h2ee;
        src40 <= 12'hd2e;
        src41 <= 12'h258;
        src42 <= 12'hc88;
        src43 <= 12'he23;
        src44 <= 12'hf13;
        src45 <= 12'hbf8;
        src46 <= 12'h6b5;
        src47 <= 12'h519;
        src48 <= 12'h57b;
        src49 <= 12'hf02;
        src50 <= 12'h3d;
        src51 <= 12'hfa0;
        src52 <= 12'hafd;
        src53 <= 12'h80;
        exp <= 18'h1e313;
        #1
        src0 <= 12'h7c7;
        src1 <= 12'h141;
        src2 <= 12'hc94;
        src3 <= 12'hd8c;
        src4 <= 12'h5ea;
        src5 <= 12'h362;
        src6 <= 12'hc75;
        src7 <= 12'h905;
        src8 <= 12'he0f;
        src9 <= 12'h832;
        src10 <= 12'h9cf;
        src11 <= 12'ha18;
        src12 <= 12'h478;
        src13 <= 12'hbea;
        src14 <= 12'h825;
        src15 <= 12'h6f6;
        src16 <= 12'he29;
        src17 <= 12'ha99;
        src18 <= 12'h6c1;
        src19 <= 12'h928;
        src20 <= 12'h884;
        src21 <= 12'h524;
        src22 <= 12'had9;
        src23 <= 12'he54;
        src24 <= 12'hb19;
        src25 <= 12'hb4c;
        src26 <= 12'hfcc;
        src27 <= 12'h802;
        src28 <= 12'ha68;
        src29 <= 12'h154;
        src30 <= 12'h76c;
        src31 <= 12'hd0b;
        src32 <= 12'h6e0;
        src33 <= 12'hac4;
        src34 <= 12'hb0b;
        src35 <= 12'h11d;
        src36 <= 12'h839;
        src37 <= 12'h184;
        src38 <= 12'h72b;
        src39 <= 12'hcff;
        src40 <= 12'h7f7;
        src41 <= 12'h2c5;
        src42 <= 12'h70f;
        src43 <= 12'h6b2;
        src44 <= 12'h86b;
        src45 <= 12'h9fd;
        src46 <= 12'hbd7;
        src47 <= 12'he2d;
        src48 <= 12'h8d2;
        src49 <= 12'h927;
        src50 <= 12'h23b;
        src51 <= 12'h6dd;
        src52 <= 12'h882;
        src53 <= 12'h9c9;
        exp <= 18'h1d771;
        #1
        src0 <= 12'h10f;
        src1 <= 12'hc36;
        src2 <= 12'he1d;
        src3 <= 12'h5a1;
        src4 <= 12'h6ac;
        src5 <= 12'hdf3;
        src6 <= 12'hd6f;
        src7 <= 12'heaa;
        src8 <= 12'h1ff;
        src9 <= 12'h109;
        src10 <= 12'hc80;
        src11 <= 12'ha0e;
        src12 <= 12'h810;
        src13 <= 12'h6d6;
        src14 <= 12'h180;
        src15 <= 12'hc4d;
        src16 <= 12'hb9e;
        src17 <= 12'h551;
        src18 <= 12'h7e1;
        src19 <= 12'he7e;
        src20 <= 12'h758;
        src21 <= 12'h80;
        src22 <= 12'hbd4;
        src23 <= 12'h531;
        src24 <= 12'ha41;
        src25 <= 12'h975;
        src26 <= 12'he3c;
        src27 <= 12'h6dc;
        src28 <= 12'hb1a;
        src29 <= 12'he6f;
        src30 <= 12'h972;
        src31 <= 12'h952;
        src32 <= 12'hc0e;
        src33 <= 12'h673;
        src34 <= 12'hcc6;
        src35 <= 12'h7d3;
        src36 <= 12'hb51;
        src37 <= 12'h4f;
        src38 <= 12'haf0;
        src39 <= 12'h49e;
        src40 <= 12'hcfa;
        src41 <= 12'h45a;
        src42 <= 12'hc8b;
        src43 <= 12'h999;
        src44 <= 12'h177;
        src45 <= 12'h125;
        src46 <= 12'h95a;
        src47 <= 12'hd27;
        src48 <= 12'h97c;
        src49 <= 12'h1be;
        src50 <= 12'hf7e;
        src51 <= 12'h7af;
        src52 <= 12'hf31;
        src53 <= 12'hdd3;
        exp <= 18'h1df92;
        #1
        src0 <= 12'h2f0;
        src1 <= 12'ha3d;
        src2 <= 12'h4b4;
        src3 <= 12'he53;
        src4 <= 12'hd21;
        src5 <= 12'h375;
        src6 <= 12'hfb3;
        src7 <= 12'h6e8;
        src8 <= 12'h2fd;
        src9 <= 12'hd6f;
        src10 <= 12'h375;
        src11 <= 12'h813;
        src12 <= 12'hdbf;
        src13 <= 12'h702;
        src14 <= 12'h3b5;
        src15 <= 12'hec2;
        src16 <= 12'h2d6;
        src17 <= 12'h269;
        src18 <= 12'haf8;
        src19 <= 12'hae0;
        src20 <= 12'hff3;
        src21 <= 12'h218;
        src22 <= 12'h29c;
        src23 <= 12'ha7d;
        src24 <= 12'h1d2;
        src25 <= 12'h9c3;
        src26 <= 12'hb6d;
        src27 <= 12'h166;
        src28 <= 12'ha9d;
        src29 <= 12'haf;
        src30 <= 12'hbbc;
        src31 <= 12'h624;
        src32 <= 12'hb6f;
        src33 <= 12'h325;
        src34 <= 12'h635;
        src35 <= 12'hab3;
        src36 <= 12'h5a9;
        src37 <= 12'h409;
        src38 <= 12'h6ac;
        src39 <= 12'ha5a;
        src40 <= 12'h2ab;
        src41 <= 12'hda0;
        src42 <= 12'hec3;
        src43 <= 12'h62a;
        src44 <= 12'h45c;
        src45 <= 12'hf34;
        src46 <= 12'h6d9;
        src47 <= 12'h243;
        src48 <= 12'h44c;
        src49 <= 12'h10d;
        src50 <= 12'h201;
        src51 <= 12'h5b2;
        src52 <= 12'h368;
        src53 <= 12'h25;
        exp <= 18'h18711;
        #1
        src0 <= 12'h11d;
        src1 <= 12'h568;
        src2 <= 12'h113;
        src3 <= 12'hf73;
        src4 <= 12'hbec;
        src5 <= 12'h886;
        src6 <= 12'hdce;
        src7 <= 12'h139;
        src8 <= 12'h178;
        src9 <= 12'h709;
        src10 <= 12'h104;
        src11 <= 12'hec3;
        src12 <= 12'hf93;
        src13 <= 12'h2d8;
        src14 <= 12'h8c1;
        src15 <= 12'h880;
        src16 <= 12'h2ef;
        src17 <= 12'h732;
        src18 <= 12'h855;
        src19 <= 12'ha1b;
        src20 <= 12'h85e;
        src21 <= 12'h158;
        src22 <= 12'hdf9;
        src23 <= 12'h6e8;
        src24 <= 12'h30c;
        src25 <= 12'h11c;
        src26 <= 12'h1ad;
        src27 <= 12'hb5f;
        src28 <= 12'haa3;
        src29 <= 12'hb1b;
        src30 <= 12'h749;
        src31 <= 12'h2f2;
        src32 <= 12'hc60;
        src33 <= 12'h791;
        src34 <= 12'ha25;
        src35 <= 12'h7c2;
        src36 <= 12'ha56;
        src37 <= 12'h975;
        src38 <= 12'hc05;
        src39 <= 12'hb05;
        src40 <= 12'hd93;
        src41 <= 12'hc3;
        src42 <= 12'h742;
        src43 <= 12'h6f;
        src44 <= 12'h70d;
        src45 <= 12'heb9;
        src46 <= 12'hd8e;
        src47 <= 12'h6f8;
        src48 <= 12'ha72;
        src49 <= 12'h192;
        src50 <= 12'h9b8;
        src51 <= 12'h579;
        src52 <= 12'h83c;
        src53 <= 12'hc25;
        exp <= 18'h1a363;
        #1
        src0 <= 12'h646;
        src1 <= 12'ha2e;
        src2 <= 12'h5a0;
        src3 <= 12'h669;
        src4 <= 12'h817;
        src5 <= 12'hae4;
        src6 <= 12'h226;
        src7 <= 12'hdd6;
        src8 <= 12'h5f4;
        src9 <= 12'he11;
        src10 <= 12'hea1;
        src11 <= 12'hc2f;
        src12 <= 12'h420;
        src13 <= 12'h78a;
        src14 <= 12'h6df;
        src15 <= 12'hcbe;
        src16 <= 12'h107;
        src17 <= 12'hb6;
        src18 <= 12'hccb;
        src19 <= 12'h979;
        src20 <= 12'hab;
        src21 <= 12'hbba;
        src22 <= 12'hc95;
        src23 <= 12'h770;
        src24 <= 12'h7d7;
        src25 <= 12'hd94;
        src26 <= 12'h721;
        src27 <= 12'hf90;
        src28 <= 12'h496;
        src29 <= 12'he88;
        src30 <= 12'hb4e;
        src31 <= 12'hfc4;
        src32 <= 12'h792;
        src33 <= 12'h785;
        src34 <= 12'h3c8;
        src35 <= 12'he4b;
        src36 <= 12'h175;
        src37 <= 12'hd49;
        src38 <= 12'h175;
        src39 <= 12'h797;
        src40 <= 12'h5a8;
        src41 <= 12'h533;
        src42 <= 12'hf5;
        src43 <= 12'h6f9;
        src44 <= 12'h553;
        src45 <= 12'hdd2;
        src46 <= 12'h531;
        src47 <= 12'h36a;
        src48 <= 12'h85a;
        src49 <= 12'h963;
        src50 <= 12'h487;
        src51 <= 12'h2bc;
        src52 <= 12'hab5;
        src53 <= 12'hbaa;
        exp <= 18'h1b723;
        #1
        src0 <= 12'he6b;
        src1 <= 12'h659;
        src2 <= 12'hb26;
        src3 <= 12'h93e;
        src4 <= 12'h98e;
        src5 <= 12'hcce;
        src6 <= 12'h269;
        src7 <= 12'h3d3;
        src8 <= 12'h1f9;
        src9 <= 12'h872;
        src10 <= 12'h83c;
        src11 <= 12'hc18;
        src12 <= 12'hfe;
        src13 <= 12'h429;
        src14 <= 12'hf2;
        src15 <= 12'h7ad;
        src16 <= 12'hd76;
        src17 <= 12'had5;
        src18 <= 12'h6b5;
        src19 <= 12'h89c;
        src20 <= 12'h53d;
        src21 <= 12'hcfe;
        src22 <= 12'hd3e;
        src23 <= 12'hb3;
        src24 <= 12'hcc4;
        src25 <= 12'h2fc;
        src26 <= 12'h373;
        src27 <= 12'h601;
        src28 <= 12'h801;
        src29 <= 12'hbc3;
        src30 <= 12'h9d4;
        src31 <= 12'h143;
        src32 <= 12'h9ee;
        src33 <= 12'h291;
        src34 <= 12'hc2f;
        src35 <= 12'hcf9;
        src36 <= 12'h7ff;
        src37 <= 12'hcf;
        src38 <= 12'he65;
        src39 <= 12'h4af;
        src40 <= 12'h754;
        src41 <= 12'ha0a;
        src42 <= 12'h8aa;
        src43 <= 12'h2ec;
        src44 <= 12'hf39;
        src45 <= 12'h8cf;
        src46 <= 12'h877;
        src47 <= 12'hb6b;
        src48 <= 12'h981;
        src49 <= 12'h6b4;
        src50 <= 12'h336;
        src51 <= 12'h6fb;
        src52 <= 12'h9c8;
        src53 <= 12'h63;
        exp <= 18'h1a114;
        #1
        $finish;
    end
endmodule

