module testbench();
    reg [28:0] src0;
    reg [28:0] src1;
    reg [28:0] src2;
    reg [28:0] src3;
    reg [28:0] src4;
    reg [28:0] src5;
    reg [28:0] src6;
    reg [28:0] src7;
    reg [28:0] src8;
    reg [28:0] src9;
    reg [28:0] src10;
    reg [28:0] src11;
    reg [28:0] src12;
    reg [28:0] src13;
    reg [28:0] src14;
    reg [28:0] src15;
    reg [28:0] src16;
    reg [28:0] src17;
    reg [28:0] src18;
    reg [28:0] src19;
    reg [28:0] src20;
    reg [28:0] src21;
    reg [28:0] src22;
    reg [28:0] src23;
    reg [28:0] src24;
    reg [28:0] src25;
    reg [28:0] src26;
    reg [28:0] src27;
    reg [28:0] src28;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [0:0] dst26;
    wire [0:0] dst27;
    wire [0:0] dst28;
    wire [0:0] dst29;
    wire [0:0] dst30;
    wire [0:0] dst31;
    wire [0:0] dst32;
    wire [0:0] dst33;
    wire [0:0] dst34;
    wire [33:0] srcsum;
    wire [33:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25),
        .dst26(dst26),
        .dst27(dst27),
        .dst28(dst28),
        .dst29(dst29),
        .dst30(dst30),
        .dst31(dst31),
        .dst32(dst32),
        .dst33(dst33),
        .dst34(dst34));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13] + src0[14] + src0[15] + src0[16] + src0[17] + src0[18] + src0[19] + src0[20] + src0[21] + src0[22] + src0[23] + src0[24] + src0[25] + src0[26] + src0[27] + src0[28])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13] + src1[14] + src1[15] + src1[16] + src1[17] + src1[18] + src1[19] + src1[20] + src1[21] + src1[22] + src1[23] + src1[24] + src1[25] + src1[26] + src1[27] + src1[28])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13] + src2[14] + src2[15] + src2[16] + src2[17] + src2[18] + src2[19] + src2[20] + src2[21] + src2[22] + src2[23] + src2[24] + src2[25] + src2[26] + src2[27] + src2[28])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13] + src3[14] + src3[15] + src3[16] + src3[17] + src3[18] + src3[19] + src3[20] + src3[21] + src3[22] + src3[23] + src3[24] + src3[25] + src3[26] + src3[27] + src3[28])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13] + src4[14] + src4[15] + src4[16] + src4[17] + src4[18] + src4[19] + src4[20] + src4[21] + src4[22] + src4[23] + src4[24] + src4[25] + src4[26] + src4[27] + src4[28])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13] + src5[14] + src5[15] + src5[16] + src5[17] + src5[18] + src5[19] + src5[20] + src5[21] + src5[22] + src5[23] + src5[24] + src5[25] + src5[26] + src5[27] + src5[28])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13] + src6[14] + src6[15] + src6[16] + src6[17] + src6[18] + src6[19] + src6[20] + src6[21] + src6[22] + src6[23] + src6[24] + src6[25] + src6[26] + src6[27] + src6[28])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13] + src7[14] + src7[15] + src7[16] + src7[17] + src7[18] + src7[19] + src7[20] + src7[21] + src7[22] + src7[23] + src7[24] + src7[25] + src7[26] + src7[27] + src7[28])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13] + src8[14] + src8[15] + src8[16] + src8[17] + src8[18] + src8[19] + src8[20] + src8[21] + src8[22] + src8[23] + src8[24] + src8[25] + src8[26] + src8[27] + src8[28])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13] + src9[14] + src9[15] + src9[16] + src9[17] + src9[18] + src9[19] + src9[20] + src9[21] + src9[22] + src9[23] + src9[24] + src9[25] + src9[26] + src9[27] + src9[28])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13] + src10[14] + src10[15] + src10[16] + src10[17] + src10[18] + src10[19] + src10[20] + src10[21] + src10[22] + src10[23] + src10[24] + src10[25] + src10[26] + src10[27] + src10[28])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13] + src11[14] + src11[15] + src11[16] + src11[17] + src11[18] + src11[19] + src11[20] + src11[21] + src11[22] + src11[23] + src11[24] + src11[25] + src11[26] + src11[27] + src11[28])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12] + src12[13] + src12[14] + src12[15] + src12[16] + src12[17] + src12[18] + src12[19] + src12[20] + src12[21] + src12[22] + src12[23] + src12[24] + src12[25] + src12[26] + src12[27] + src12[28])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13] + src13[14] + src13[15] + src13[16] + src13[17] + src13[18] + src13[19] + src13[20] + src13[21] + src13[22] + src13[23] + src13[24] + src13[25] + src13[26] + src13[27] + src13[28])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14] + src14[15] + src14[16] + src14[17] + src14[18] + src14[19] + src14[20] + src14[21] + src14[22] + src14[23] + src14[24] + src14[25] + src14[26] + src14[27] + src14[28])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15] + src15[16] + src15[17] + src15[18] + src15[19] + src15[20] + src15[21] + src15[22] + src15[23] + src15[24] + src15[25] + src15[26] + src15[27] + src15[28])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16] + src16[17] + src16[18] + src16[19] + src16[20] + src16[21] + src16[22] + src16[23] + src16[24] + src16[25] + src16[26] + src16[27] + src16[28])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17] + src17[18] + src17[19] + src17[20] + src17[21] + src17[22] + src17[23] + src17[24] + src17[25] + src17[26] + src17[27] + src17[28])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15] + src18[16] + src18[17] + src18[18] + src18[19] + src18[20] + src18[21] + src18[22] + src18[23] + src18[24] + src18[25] + src18[26] + src18[27] + src18[28])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13] + src19[14] + src19[15] + src19[16] + src19[17] + src19[18] + src19[19] + src19[20] + src19[21] + src19[22] + src19[23] + src19[24] + src19[25] + src19[26] + src19[27] + src19[28])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6] + src20[7] + src20[8] + src20[9] + src20[10] + src20[11] + src20[12] + src20[13] + src20[14] + src20[15] + src20[16] + src20[17] + src20[18] + src20[19] + src20[20] + src20[21] + src20[22] + src20[23] + src20[24] + src20[25] + src20[26] + src20[27] + src20[28])<<20) + ((src21[0] + src21[1] + src21[2] + src21[3] + src21[4] + src21[5] + src21[6] + src21[7] + src21[8] + src21[9] + src21[10] + src21[11] + src21[12] + src21[13] + src21[14] + src21[15] + src21[16] + src21[17] + src21[18] + src21[19] + src21[20] + src21[21] + src21[22] + src21[23] + src21[24] + src21[25] + src21[26] + src21[27] + src21[28])<<21) + ((src22[0] + src22[1] + src22[2] + src22[3] + src22[4] + src22[5] + src22[6] + src22[7] + src22[8] + src22[9] + src22[10] + src22[11] + src22[12] + src22[13] + src22[14] + src22[15] + src22[16] + src22[17] + src22[18] + src22[19] + src22[20] + src22[21] + src22[22] + src22[23] + src22[24] + src22[25] + src22[26] + src22[27] + src22[28])<<22) + ((src23[0] + src23[1] + src23[2] + src23[3] + src23[4] + src23[5] + src23[6] + src23[7] + src23[8] + src23[9] + src23[10] + src23[11] + src23[12] + src23[13] + src23[14] + src23[15] + src23[16] + src23[17] + src23[18] + src23[19] + src23[20] + src23[21] + src23[22] + src23[23] + src23[24] + src23[25] + src23[26] + src23[27] + src23[28])<<23) + ((src24[0] + src24[1] + src24[2] + src24[3] + src24[4] + src24[5] + src24[6] + src24[7] + src24[8] + src24[9] + src24[10] + src24[11] + src24[12] + src24[13] + src24[14] + src24[15] + src24[16] + src24[17] + src24[18] + src24[19] + src24[20] + src24[21] + src24[22] + src24[23] + src24[24] + src24[25] + src24[26] + src24[27] + src24[28])<<24) + ((src25[0] + src25[1] + src25[2] + src25[3] + src25[4] + src25[5] + src25[6] + src25[7] + src25[8] + src25[9] + src25[10] + src25[11] + src25[12] + src25[13] + src25[14] + src25[15] + src25[16] + src25[17] + src25[18] + src25[19] + src25[20] + src25[21] + src25[22] + src25[23] + src25[24] + src25[25] + src25[26] + src25[27] + src25[28])<<25) + ((src26[0] + src26[1] + src26[2] + src26[3] + src26[4] + src26[5] + src26[6] + src26[7] + src26[8] + src26[9] + src26[10] + src26[11] + src26[12] + src26[13] + src26[14] + src26[15] + src26[16] + src26[17] + src26[18] + src26[19] + src26[20] + src26[21] + src26[22] + src26[23] + src26[24] + src26[25] + src26[26] + src26[27] + src26[28])<<26) + ((src27[0] + src27[1] + src27[2] + src27[3] + src27[4] + src27[5] + src27[6] + src27[7] + src27[8] + src27[9] + src27[10] + src27[11] + src27[12] + src27[13] + src27[14] + src27[15] + src27[16] + src27[17] + src27[18] + src27[19] + src27[20] + src27[21] + src27[22] + src27[23] + src27[24] + src27[25] + src27[26] + src27[27] + src27[28])<<27) + ((src28[0] + src28[1] + src28[2] + src28[3] + src28[4] + src28[5] + src28[6] + src28[7] + src28[8] + src28[9] + src28[10] + src28[11] + src28[12] + src28[13] + src28[14] + src28[15] + src28[16] + src28[17] + src28[18] + src28[19] + src28[20] + src28[21] + src28[22] + src28[23] + src28[24] + src28[25] + src28[26] + src28[27] + src28[28])<<28);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25) + ((dst26[0])<<26) + ((dst27[0])<<27) + ((dst28[0])<<28) + ((dst29[0])<<29) + ((dst30[0])<<30) + ((dst31[0])<<31) + ((dst32[0])<<32) + ((dst33[0])<<33) + ((dst34[0])<<34);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h0;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h12a7b5a0e71b9f6be39122e49f82e9a7c40b55ffd0823f7468eb0f568f7a8dff1ae318d4349112550d554a1beebd99abb3017df7bad3fea18315082eb1ad7ce2be1b12717da14717efb6ae114989c1dae4c03397f5a2d07d731ef44b9f4a5bbec07ac22493ef9c78e9f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c69ccfecbff3c2726ef2dc8ab7ca1337175082888fdef6bef77e086273b5c4efd423ea3cbfa8f227fd8997d62fd46e389d2212d99ad0f2f2929b5ce7bd6355ef7847ad6394ff98f33c5e34a20c8743c2036c4c017fce9354de5c199c072000e14b805ab5098fdfc8f9;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hccd80b1b2bebde156e9877654e47593fb7d87489f64539f2fdd2fda54661fc49db0652a23f4244946881ed4acfc2d59f9db28311fe6768f92c26fa4f54469d3c4bb306ba330ae724a563c43b23c867592b5b634a4601893bda8801f86d2c8029be024afbd7a6a5ba0c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h112c537aed08e846e0868c6fc59c5f78b636600fa334649a228eabc10a1edaa50621cb3573fa36ed472001d60987f8f45ada08666a64d0a06b655419b25099623a99c040c8b14f33663a4a4fd356878abb956585584869178d7defe3c3be104f7e11099a0f74f6ddb6f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1aa7d5cbfa667375ca2b2287de7f686a976821261487c0342d5dc20c79baaf472d2e69b0eaee4898624787c00010d308ee511cc8f4c283bb40e17ef25b724e2d51fa7cf01c96965de7ca4f4af725d605a12befb1d7a54a5d33d48f8bbd4667a2d372f59603657988b67;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h14898372c958f9b41e88032b535edb4b636da1300be6a45ff9fc6dc5ddc0af43ad5dd136f46cbac5335b53ac856127ec9d7c124427f300864a82b304691d82b0ffc7df08567c1be75ff1a0d87a651da9ff43f87fb19300fd81f0df3bb7838e7e78ad9b9b2b394cb49c0;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf7c4709c56f066c8a947a1f01b2f77e38eb0368ef8bec2a1681aeac0bc5794d10e78772424780110074cd2d887df83324540997938f34e436c6e8d168a9be81212ca7a1e81411cb0c245a824bd27f82e53bfe07f75ed2eeae49cd70f94cf46e0786dc1c8b42e9f872c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h20296111b56670338d8a0d2b5db741ed92500ed4d8d72c5564a6d0d1e36322bba34dace88d47437906d43300b11c3f50d3a11d4bc3d359228aee03c385f2a51760c0a5e02fbd580e92191971a6f71192241febb8d4a5db075cec8ce65f48480dad2c078e64b23e2b55;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h13f38ceea3c9fa4633035ed935f97f899645ea32d21e5f50155522c60dbed1753599ab04507a773fc9af523103a7e836ddf76e25abe563b5bd2a2d8854ccc2775cefd80ab5c5e99d9c185225567b0495df42cdcb658fb839b4db4ad3719d501c198d959ff688bea4ebf;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h15436f3ff7ea0160319308b8ca4c771a2e43321eca9f565d51130a658d1368bee841d94fb41508eb6be011fb942bf2ac57ad942f2aed4e116dea4086ceb4d4ff4024a4955725a07599053b3a9a4f28b79fac8d817b85dde1d3e3094ad3d68c1034f51aa0dd22bd3bf1b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d0e074de28ed694e8549839dcd09cf1f5437ab9531ae1fc9d27381614062a012eb862d0e62c12cea2acf0962263d746af48ee07a484d165f650e2176d34ada1b665f2f4f62d3a58f7f54d90c9dc95bb6fa06085e6c6026326b00b8dfc785d005cb120e429c86cefc0e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h3730fdb4bab5c2c87d1e47150ba87feacc8a37721d7523f5a3a4cad0ccaa5f13146e3de6581b4cdb74a7f1f4533550a7e798c7c6a5644ac9d1c457eb941a2713da7824e00b28d787431598b1433ab549e1e26a8d4e4a5ea9ed8bb4725acd06409c990cd37922fa070;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha55b77dcb7469397b2b3893c8925c0198a2cc173014707aa138a1053b270560ea250f18fb9ff538ff02f1aaeb28f42e8d5339b325953733db42e2434b0f56836e92945d52750c64069416c1c4c2d07e53cbc4dccffd2e7caae7e33f0e77d199d1aa0900ee4606cbc64;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h2d86633036278218ed1296f8625db1b9e8456e1538cd4269e813baef23b4a39b7c467ecea98f3e218de2506b3c236b9f805552e0f4326a90e3e6f5fce4f34995614b138639030c9eb724b6da3905ebe649709db4ae46c63ea3e814fec95b18545aee6e3f96371c63f2;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a5dd74904bfacb038d9b436fb9ea102a67f7ca3ac07a5fcb798cef2100129bfbfcd00708f476943f5e7c9aa4ed9154739c5b9cf9ca0f2c2503f32af23f2684e959818102e8f40e8345669d68bee5a96488bc5f96c8c4391044193ace3b43399281f5acb924ef8b07fe;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf9fa515a5bc8fef5f2d0af3fcf8131835b2ff279f3db63a61144c8f68e9f9a64d466cac80dd618ababf90925cbfc7ae707d48764d3b784c897a30dfa721a8f2594cdcf91a4c4fc6df1af542f2fb2b4494e8c78fb61620d2515f6201c4f55eb06c759eb27f2ea6b56c1;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h137d6817cf1632e2490da4661aa27bdd48a1ccaa71beccb85f3370ce0989b5897635c96467b859893c5576a0a5f1a5fc8dcbec79a46d23f4a1d68bdfb3f1cb5819f8b6734e4ca55e7ffe4201d2be73f73815022ab7e67ca589e594ee0db5359f3342951552c5093b72a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf46d3b5b107138f5718519b81b8a24aa5d9caff4f1117cdcae39bd48a025a5f10ca979766728f5fd2b8f2b5ad744909fa61f978bdedf74c6f6e277094bf9046faf910d8172e43d04b4666cdc47b3b72aa79923cc839e18d59f5603a74b623b858fbdc675b0b76578a5;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1acaed179093385cc9e682a2a01f29bddb3b6dd9ac02b3a26523a665351edd9cd246dc4112bee0640f78bb383d19757c80db1a1aa3b608f4b36932474b04918f257db7e774a4ab1520e2f75d2ef10600d3f024f1aa94a776904575e4b7db5c97248e69a92f7376dac90;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h9651697259eb1f5271cc913a58ad96bdb382f52a4050cda8823371cd42f57719f5714bd7d3418891c23b25cc35300a072e23f50c6ca35d8f0b6123223f56d81d3bab1781f79c9c4f53ac0f0fd977559aa62383f89d056501d8da0448f4422b57be674392fbc3bc4172;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h3283b7aafb00cd8a5e7c8884c0abdefc693e78048f284869a2cc5528fd445e67e4fcb1c88607d28ef3f78f59eaac4827823d9cfff03b57ebc92f7fb4c10d2a023d819daa78a62ed0459509a59b8b4ae97b28facf2490200b32200dd6183e69a4f7f19f4aa9b4dd7c95;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h14a568a1dfb05fa1b0d1953308b034575d562b7b0371cec75412c7da76067f753b446f744830231ee4c86f5d79b905bb5f9dafc2e6986b3cc772976ee4dc8630fc4df9695b466b31f124f2dea118379185fcf751502ca70b9708e136d27237b99c7f1eea49232276914;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h38f49b872e359cd189aa53c686d9ffe38d156c978076b1008e4c538cf452ae8579db838d68893891dd2f7ca639de026d38d907d1f4facde39aaa69a416d24ee6cea3653a65a7f7e30a915b002a685f275f2eacbf0ed86bacedab6fa75c51e7f3b2e05b3eeb1316e5a1;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d3bf8a99e5f90a8a0b9f0b7933af196a9c59fa20bf237c7cab821a7ad915c98930e35a354a1c5ab2f108befc07ddd892857d025b5e54d61bc5e1dfe8612c9cd11461359c06940c276a287ec535866271b48c76123aa06e3a3c9ee8b2f35355cf2e65cc65b0654c27a4;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f4df036c9e275c0f5f290021d698d59aae06892cdcc4a8ec55095c3f9f18574e2fdd4e90b3ec35520f5c89a7fccc899ed3e64bca9894a211bb8f120f6dffd963c1db17a6442c3ba9c662b69927729d85f34f0e964ba7644146099e35d0933c6f985f6ded3f2010df29;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h13f75e0151922296d2cdeb1819c383c9d70889d8fa946f11227bf90c32a015e793f19226c26c46d2bc9adc7c9bffda6701e9443d8c5a77f388996187c30a227f4c7e6a662facf7558b51722c9b622fcd5264fc7229cb6943ba259a8988d156063bc63a0c5a4d909f37a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he749e78a2b779c1580b10d5bc86e906cc35cc88733debaeb9b2280586de403cd67b761cd35c378b8ec5e9d829d2122b0c6efe60593983727d1954824c20cce553ff462be8bd9736a4001681297ae823d1b294a5839f83a78104265addfc38b085644ae2bc221b9f23c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h11d1999c8a66e4ab4aa3a6bb73e353d07b2b01ad7948d66fb50be740965e63ffd8466ded34d2d6edc3f9917e1ad20d1cf744ec27cfadbf2b28a4d6c64fcbc334e14ef7db8133bc98b5629a3e0f8715555ca6757af05085a83ed04db58b33797af57105bcd51ebd088dd;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h17fd609d4656bcc17d2ce05ae6dbaffaa58c02640783c12f220c968d5d2be42ae495f6fb4b25350fcf9749099a98032ea089bc139f9b35827f53c681ffb070e7912a9cb60784e10f203188e86e3dc31ccda97a492e7019be496fb235b4a982d63114bbdcfc4381e413d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h16e364105ba39be644830aa6528a5ffbfe9c8cfec103d9894e69de3313f0fae9e046ce2882373952f2430ad485efe512aba5c0ac56e4639f6528a2f41ed52b588430624b0a930afee631de1902d754f3ec0d6432d1a16bdf765fee79a01ed21448f919fff8b335d3b3b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h54176e6f4698dc879ef4023fefe0a1e38c40bb2ef77469b1fa75d931540f3e3bdd6ff8cdafbc0da117330786c0c4a377bbae516885b5907eed112a788cc59a8eaf1e59c780cafda0414f8704c098aec78903f3f319994a994151948395d7c6bd2054259a5fd6e10724;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h5dc124cf3cdceb66fca3e5975b566058a1b68975ce2487b1db679fbe7cd40346ca87e19d23fa297e859408bc7936aa0aefb47df20add6a4243b9a7819c7d7b5dc28e0b5cbb4fa291385d32bccba65465659475c36e75b880636f20f3dfc274bad3397f186cdfbba0ed;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h448d826da84c2eefac68b40d3c7a9a8d34ed639900c6c2c0bd8f9ef3f95df3474945db153f4f384f3a8b2b3ca2e5ffeba30cb1dfaaab86cfaae1bdbfa2c7f6b41556d97c3ce35aa9f79545eb5b4b4b7f8aba4224391e1b566e3e1dbc3bc9e4442e357231462af3f753;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h19e1b685940067e4239d0b7021edc11b59fcf14a8fa12c7f21ea46962ddd2bdaf7a1ff9e6bed9f3530b574006119f12a5b723de6067447f3fdc47a47f8dd0a204b013fe56a23813aa87f8f5042d840d672ebbb377ccdf2cda27dcfc6a0fb594993842110a42104607bc;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h38dc8548930bb478404cc3a1d5a69a657bc77e02b243714e51321eaedb826668a82aa27d05a18936bed8a0a22fe06ec22f1850b057e5ea2b22d10d19f5216afcb404ae0fca40857342079d5dbc78e7261803d5f20cc945d3cae1ebb1aa31a318b7f79a8fc5f29b486c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'had1a1bf583830410f8423a387f95ad0219f0685e092c1d3c9b5039d7fa68bcaabf1a06182c2a7dc95da1e62aa28f53e0e4547e3b3a4b15ab57fe81bcdb6e215f52ec7aa48f3522e002db8ac380ec64d132f99956a445b0ede7f2f301a59088cbaf9a55f5ca5c55c5fd;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h289e4073c775518aec82fd4f86c82008e6e93bca19c1354ce3559f7efa42492fae5624e3537565d7c55527a299152a5292d76017be503d47e27e9ccc6e3802d7c5cca0ad07d337fd0a86a98558ccddc75e10bbc4d8b36e27f89dffd3f58ad261b53ff1c7237e0ab84d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h48ab7e3bee06c7ab949846e094ebeee952cd12d863d3163cbefed1b2354714daf09d75acf208c0823622fa89a8cff72c873fa97f6ba068141a19fcc550fde8dead1e610dc40cc780de676184b29666c5554ba67eb33e056ca12a8e6eb03ea67c94e3948dfdb725a994;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h2ae55a7a01522fe205b6c554bcb24f261c8f85e5a3947fcfdf1485f36325b7a4527b9cf20acb26c7337f0c9893a36fd45b8ef5641e17a16d7256a80e17c6b433816515319369756fc897dd48e1df0889f9da2e35834417bb96a0681c1397a083f6d8379a10ef2a3ead;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c9ff614958e03c139d5a144399649ce7b90825c96c3cec652b2c95e47d935aff4c1d391c4d96f3fc67c06599986272244e1af0cb630eaa850bab72822dcac9cf94e034932c456e4b273aee84be6e9cb88ad774be751d852c492b085a6687d86d9eb6576d2e217737ac;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b1876282732b586984b8d68eee810f3a35312f67edf71ab5dbe71c5839d813249d74f0b9aaff5631fec20bab2c7970a9b737d045233fd0282741fa7270f3c134ec47d2bf0ec461aabafafc6332b3e4a950b0a8f2c5bff959e3ef47d9a72ebe32cadc596d4b5b526aa5;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h536cd5a50596b01ad1e6cc91017c53474db3c662a8c5497afb958ca120b6413cf64e93cce74d10484b2ba23e2a6a9901d03f75bb5e145828cb45956e0ae4635817c408866640eb2b203e80edc92e2f1eb90b4587aed667d1402a583151c3d8ea39bbc1b377e9bb2ecc;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1aff09a5ba2f4c4c14be702fad945f7b7a0f7eadca9d8582baedcac7a070f5c76540cacfca0d1ab5a3398f48fa371a6b9feddf1afe82ca6c5ac0bee2a4396b76348f21dbe9cadf06a3c1d62ae5dbbda68bca933475057831518952c7abdf33f349b4e7252e2f8c491ef;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h15d4a6365909eaa564cfaf147d90c542b8cbd652aa4e29396d341143d363b3d528745aa64cc8041845223ebbfd11b17737deb5a70cbe8ec20558dec85e58d83554927d2dd54dc1e1bd234df4f64fd7cd6fe1fcc532c53661148288dc4fa96427dff53bb498d0912dc9b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd874f7e0e777c8f59bef1b0dbf7fb7d11474bfc18c4375add32c2430ed82521f9bc7deb633bbb32526c20ad8b3cf696eda6c7293994250cca58793aed8edbdb4344a9c91f95a55fa887c63e6d3565e1055722f1aced8b90ae5b79aa850543162523457412d187af50;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd01e7488fbfbb6074a5c93f74e967a1fae6a098f22890f09d652f0ce0d9423f40f294bf8698d35fb8282b39b813dd067137a881ca6f9637e4fe646e4fc265b485a812d76daeb2b6cf8e63d0f4e196fffcd01eb0f5196c844c5306fd75496e3874f908e8581a67b0f2;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a501e8351fd8f523d9dc62615cc86ddde3d9c222cb32e7a718d13e0199d1dadf226f924174d628f57dc86cd0f6f60371ad39ba890f51b37b40c95cd593501b4a119bac0689c696cf7e4638b06450c9a0b5e62a4a04e13155d31e2baea4541ba7109e1ac2d7eaf6873;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1926904d1d55cc9d33e3572e51934ea63ad2e95b76c8a3e4a2cdc413e5abbfca4c96f94b29d39023cd3835be8ecfcaf669af75950fa412980e272a51730bfb7d24e8a5ce2644be8aad0455ffbf6eb59a3cc96187b4f52e2297d9e2b63055d4d526565defaf88047235c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h13d5fd3396f1f3ff39acd4706c1782c0a0594b95b5b1304d42e3c5cf9c1e958b1002e6237868b17159c7e6f0c57924786caeddc2455137b887f80b82b3104c7c9bcd4cb9babfe7661f3840e38a7b6d835b58b3b778de731c71820d85996317b1005d5945e92e46e3447;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1918aca4fba4aa1c447d5a7859aec045bdfd986c49829e62b14817c507df9c47530eda66870de4e4cc1aa4b9baa84db839219596441371f6cce04478aaa8960221044854604c7a73ffb52ad4c994529fedaff0b12c104ad3432a5637f5e7cf1357e1f11aa847af77809;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b8bb08dae3ff611fd12ddb5dfb2433ef01849e7b2c53aad063d743129bd59c9381d6ef5309348c5698bc8f1d2eb0202b290acc81f27a2e2c43c46a30e59c206c6222e903d14b54b9922411b71fcfb6ee7709db631e8a9108b973b050b201a7fd44140f00809f8c77b0;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h16886ba3ee6de808a62dfcfc73b8692c6c9412a7e30d598d5517a2e1dcff0eaba137fb1e83068001a9525bb8d2de7089d6edb8cde301c9fb229b539da2e7ffe6b288ce14afab8cc7a59f4755b37aa9b81a0c986084ccf19c3d178cd52aeebb5cd39ad9a5cc3954ec4d8;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a7fdcde4ec8c39ffc9e6f0835bf7a65c28959809bee20b9613189dab51a0d49ab6efdb26f4a2df4d59aa8909451f4d8c9be0079d4873f7058044e687c7b0965e67950dd87481a5cd22181b234f2b14e96e33700d0e2343c5c2860bf1c8779032a78e4b53bf7e02386d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h177b9a6d9701a3483d5ce786d2380e56df0618150127941b6fae7785b8c036999a3bfc674396d427d06b56fe45907d6ffa35ea670dad77296730668b3d95a74cc87d18a9f4cd4cd0c732d3c379d4024790d08e8014faa86abf8af1ebcea88a00669644ba16dd2992b90;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc3879799d5df823862f288aebc8a33a4d23036e3766fa375702b3998a7f60803a0b9447dc996383fe60ad9f140e80c833cce56945d491dccdafdf62def6145bf94528c8f3ae5b7d22e520120a1a9bd6518c9b5f5d7e1de4617b12c5088fac3c79f419c5dda97da068c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha592d652fa124dfe7463eb1778d1f0e1355a5f557fd68cf5f0bc65ce6b4380b6f94dc4c7ae20262aa658a18db260a842c7f727fe5810c1d518fb03693fe83879ec66967ba8664247967135a189c66b4cd96015b743148c2f9df88ca9a7846b418adc32f9a144b2645a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha513a23dc96f295fc330accef707030d16e70df05eeea344a1efce75450a9aa7f3e946776b66701e2e34674b68c2f8b87ff20a425e7f1b3af061ac6e8853efbd36c4281cbc2f3e3e4a431c52e4f68cce1a181aa5a315d4df22f414715cb07196b91f8857ddb0a44edc;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h5d248b6d60d5438f50d90111aeb7a37f44e976b90eea4dd0bf28b681bde85b330b843258b2cb76c49304858deaba0c7127eb583db505356a0683cf96d539d8497630ea0b1ba1620391c52612312ffed3be2419628ed779dd91001ddba8259e705a709c30d066acf43d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h138ee4fa52d35f9fdf1b3316dcb4b42a10d636a0f43f31ee41348e79da6958248db2bbfd27f43a2379a1602026a8629bca093e06d17bace4cd6334b73066cb7923c1bb90fec7c14eb90fd7c0ec6debb4fda7980a0ee15ea13b468c16a671cb0a34687b5b5ed88017d3;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h155264522a13e2eb2a9f7f4a5874899964fc7baef979b57a546d5e204e9760c104917e42abe64839f4b271a2c17e9b76ecf88a26b87916305322265a1b95624092771910c3b8f41138ffa6f83259d779813b289f3cb944271d67456ac876b010bddd51091eade53e4ca;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h17f64ee61b65fa5b296e9eae1452039a7d596dcbed7ecc54f02de4213f6c058db66647e24de4f12e555da9b29dc9372e91b8aa251bce3090bb6b3872f555f894d36671645361f88ba63776ed02ff19cfadb8549a81f56570538dbe4c53dc12ac6b1eac188f4d80d0f57;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h7774d47d47732b23e4084cd5740c45da60446a9875c99d5e2ce28039e392d9bd22867d7df4af3a3574f4e2f442ef46a6f245dc106b186796842da9779f4dd4698a48e52c8cb0ce08a4c557dd309d866cba4e442029e4e2fdbb2e8ba5627b9bbdcae5fbf01be80882ee;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1105eb4611171e2a37302624c02ea00ba3c1f5beb987284694b5597ad97b084627d65320203b19d99a5b442e3e64eb16f60b84d56ef395cc37420e212388d64e8c66a387e84a6aa36db92a2703c1f93f6233248aa08c778899da324e4b6a95ed1b52981b2f9d3509023;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h134c54e5db9eae6b768e6d3a76961664f4589807f6ce8b54ef3ff05084b2b68760a0876e54361da788ea6f89034345d123800511c0333621e1f48e2e50f1b28df84fad934d4216ffa14c72b8101053838155e3977f80a001d2577721dea8d927c336ed3f612be6b6374;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h5c15c75d756843cd9aa6ec5a9de8b1c921bc73d654733336d31dffd5d4c7ce6569ba94779214cd17d11d914c4ea2e85a0d386350a215dfd246226b8459fc040d37dbabcbcb497e0f615dd24720afc349d22afb681e8317fb6f5bdc02ba7dd4bf129388484b696e921b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1bb81823c641daab59db461c942a47a8a2f964b80ffd78af9f4e1bb76e4921ba7ba8a31f62fe0325f94df48f93f7fcb6e29cc35b3902f874722b16befed8c41c48ad4b218135c4137b524b69c8564212c628977f387f1a3765662dbafa2b78d21717951c083e8947537;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hfbbe202bc5bfc073508368db36f4a7736f861d0e4361178fc0872af3f0156c13a5d92032419b8d721bcc8c3555c57320c135188092c48e23bfbf43bd2b1ca6c680ddbebffe8eb617d024b4dfbd5c9c5aa3dc3ebf02ad026f2fcc1310b7ae6bf652a9142d968b7148b6;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h186a0d17f60824ba80fd754bd9f103d2c5b0a0716fac1a3cd62b78d49ddfb61254692a4e7d725ebcc7398b75122a848e3def22bbcc9272c463ba1ec39d5fd05d2fd435131820b2c06339ef56ca4b22e6b39d04a184087f504fd6fb3f294f07153870d7926c54d692655;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h12e2f3a2cac32d7106bbee87da27fa0eae6052acc8ca4037c993e9e296c226e9d0da2b16d37df22bf97b0d2e5d749f9c49e0628366ae79e8f79f752c1cf5c5ddb9c317a1e0a886b4822c2131c544480e28434cf5fcca29b72b03b5345a00124b89407fdac8e4a09161b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h12183994a1e665a120ce9ac6d94ff039a72d7ecfd868cf04e50f58689d2396a674e68c98d6c92ccdf7beb7d70ff014a5c789296086f21483d38756be6efb43b5ac6e3e7ea4f2030a085a2aec0a4d01849d2044287356e1dbbc7ba253c1ff9114d1b80d8b251b8311585;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h51975140995394497d93b5cdefa3cb50e7c65d97756bd0d31e74423a9366e8b16c1d1fe579495842bab4ab4f5a38fffb3544d679f1741327d9e70eaed08928e673822afdece8c70eba022e2f39771be71997d87b1e9a700e6b4bd5e6cf96a8f9b8ce9b67b0f44954ec;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h100eae7f95ba3ae55cf68f8610865238fa7e68888121be346872eb714fe33208975119a85fdb4789e84c39d3c47990ffd3127cae00534e2fb34a5ed690f6774fe749d06578279f0b18264ba3b0d673d0bb553333bd11c94f2df5047e819df7d3bbda45064469df7b8ef;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h132b2764dfef1eed7c0cee513e8a42c2306b58b291b8c32a8575b69ae6f54d679c10aa95e5b4fa6f4dc4ccc0c73122563aca916f5d95fbea8a13d6a2879af6ef62fac0bf2da45583eaa7399c374d357e1b697d36dcebd9e6dcac4770b85dadfab9e977826c06369ac69;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h9c58f58d1881529da67bf72981d7404de49a61a70518ab5949893c816608b167095fc6021ea253528c9711cb23ee672c923791e9584713bd030a3fc5033591ab961ec4b33e2e828132dc0c284ea6379dac037da7c8523ab1abaf32b0ae309fa121c174438ef2b8b6f2;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h4611d5eba6ed5bd4d117fd9fbd31c00eb6cc257b69cab7b73236f1b3dd8f48a22f9301013eb775aa53b7e25bd438ffe0bfb8c6d32a153a6fb6609dccf9ad812a4baf5b7e293843c328c18f112d69c423a922097293322fa32e2b7b7730f85dcfadebf5f2136e7115a9;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1bbbaea38740e4ef1437bcdaa01143af773e30219eff8d889839d38d141f9a37be4fc02af930c1407a4c90bb14f470175701562b86161bb4d05ccf447cd2a0ecbfbb09f0585d25ff11b385029cbc65ee162e42d3f4c006efe80d4e0ecfa4ec5607f8c55f37507ed4374;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f1cfea86b50c97e736e3a33b7979930ec71ca6e8b657cba04b320c9004c642a3afaffc8b29c78b6624c7951f7d9d6d40381c1bdf10418a764ab16acf50015bdcaede4d11874cbac9f8fea8cb3b46b159ca8891aca9193ed1757556007c5f6ce179a4b3a83a78a412de;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf48c90cc6af730e277ae4590357d823660b8368b5a2c2690cd5cae7bb4796a70f845849971b9815a07d98125fc38b73ec93d4f2dd138009b560e1740bac20ba52d44c9d23981300e6c32e84d1dd82141c741bdecace3382ff29436e20960f6f2c58977a17104393ab9;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h87934ac2f53006f790e55822cf65b0adf3e2524d8dd0ca34d1481938079c4ba3262f43f0ef74ec555743c9c4f12355da20a88ac8910baafaf195674cbef190eb049bcbacd24abf088dc5d20e57edd3b50bb5d764f0814a977dbf82d61a17f31572c64a73dab7b2e393;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1966dc0e8b0fdcde5d24ea03df18029f2ea2f4e3d5c3cece614372d6ed54e151be23c3c526cb1938640fff5a78b842ceaedc45dbb522fa43fd6f3eeb1b1ef53ca76f572dfb98f9a80b788fabd8a72eb7719cada7623053cb27436a036e794260fe693a7d676a1442252;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d8a20b8386b5fd38615daa972d8e8bdb5e90e048b329b83218f7db47c8bc81998a03d92670885d26954dae9de1860d64409865972d5d4ef69a57d1add3d1e1518dd3cc99581421c422f957afa581383993ba5afe60cf6dbd1323e11eb4507bb1aa9122629858cee498;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d039f41d0717f8a295047fbb27810eb511af24b8085364b56835b97db80e7cef7318201f519d7083935bdffe9ebbcca60cdd69a576bd6178270427eea07eaa20bd38d75d0ddc04404d2e23a9adfe6aa9e184488fce1035d221af9b0cd1e7f6309ec008175b3e5fde8a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h4bbba4f2857be70887b3fa590a8ebbd7db641633ae656b59b6e60216c3900242802d4a8a15e8ffdd469b77437f367a393bf6c5b3d58960077b034a9be33db9921edf9c22ca88daa750108749ff1487d89aae8f07c1a4613780f03ae043abade10cf93ac74b866d29a5;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b855ec2d2d61076e57d38d4de83a88767a6f2a532a3ee1be4fd2098cf66537cbfc779a030fc29768d671b39f8c96dce2f404ed6c6c620dfc1ab083625e71e4308de1a1c7a3560e7a7f2dbea974fac2e0caa65fa0c89c57a3112632207c5f6e2953696bf594280fa434;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h19cf29bed273c62213ea4d4f9df10b5a99d022f2aa6c4b4171adbf9086cafe81e28e0c565d446e3359cf81bec9dfc5b2b2e19d9b492c23c487825c9ec1662fc44d4db9e22fcf26c804f7d3fad75525ee0123ca622e0caa83768cf85d26d024c1535255951cd8c23b7a4;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1fe30211f815a73f663b02b5b3d79f9750eec51f5c5cdfd1982e8fe977a58e5454ab91aaee5319831756f0e265a8d586d54e59c87b33e862045c9a5420c9e9f20c542d6a1633c39f22bdd6590c7e15be86e40e3848cf3b9ad54c31880f44ac5253ea3a3880a648fb054;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h12de8e3c741cb0f755722ed703dbb1a52a2b42ff7f93331c1c6b2fa7e958b7b5726d3cb229521dc4b549634c3fcf47923e212ce2f02bfeba695890ce5bd48bf89533bfadca3f8bb24e0ce7510ed1a05d80832e58d461306312de59f410f16cc964c8bdc0f9cb8500779;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h144843341218fb60fc3dc01e488dda1a83936d01429d996563b0adb44348dc805cc772a9b72fb3b1ed9e0c896309102bfb5b4b7fa8973971b810f65fbd77f783f1a8ae480ddf97b40da5d2e71f0b2d8ffde95b8bc5855950658d2b69ee54aa8bad8a4a1b7b3fc7be280;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hadcf668ce38a635671cbfc0568e33d00fd9738e4d94d102920cbea3383d5bde3b1456ca885924cc41c3538e41426b42e5b4fb0d2cec3de18a9f287a208ecf7e0a8db8b9e698db6d72e50cd02946c9975bde7b50e481538b42e68097838998b5a1c89e5d3da8019dd30;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h60e0ae90f56336b26be111d198712c63ec276ad2880e5701dbe89f311fdf6e1a510b6e78f9e91021093218abd49a43482d96ab09b2878ee24ae2fa9c314fe591e7fed5785e4ce9666f1ef12d9fad180edd24c8eab0a584aac0a4ea4665ad656db4541c797f50cc0d1e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10fe816576b5117aea89b57c6ff80279872fd54cc382b8f06c69c658c4d7490b3e1c4ce30b0eabeb268f5338ddde0086aa6ccd8129cacca1b81b2303880bed682d7e9ee1c6938eddd0c6b93384dc0c07d943b24488327dbf63f5effd5a2118fc1391ac35a6a61c60f6a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h4e1fef39c3a1607598c2f002a27a525c84c4c27b5f4977d41c8bba1f190ffb0a2923c55d76987f62adae2cf73a0399d8faf5afe9733701427ffa1186ee22d1d2e7cd4977f378ac441adb4f500f416b501364b7e476f5fa6dddbf1208353c7552979cf2ca06357039af;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h29138b4510c17af46e993746ac67de100db5a8a49ec53e275602bd5b4026c6bbfb87958a7ea21c0ebb5e6dc1f581522eade765e17746a78bff73852230583fef97b3915cb95ff72147bb2156d7136a1cfafc4a3b1e10813dbfa8ef146c5b4dcd8f091cf421927d85db;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h14a0f5d1c274e70824cd095a7b564b4018ccf3635f9a1d4aa8cafdf1ec98bfda085e243381595ed1eb515826927f217b396ca287c2b456ee8e0cc1c3938b54c7c648f0d792e5d98deab5469dac8ad7b263887db1c562af91f3c7d626ce98bca767f24c129cc2195ad56;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h128039b36dca23ede65916027526623dc50b042b64b1c81e66c2a0e4a2bbfedccfa7b7fc447422ff2ad85424dab9bb8648556afd584ea6002e7abece25e78ec18e23075ee43f59e58a659d91ac42e7546da5523b433db39ab44acd49f577991a8c144fced9f14b5fa24;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hde2ec9945458c8d01964779e7ed10d155ff00a813073779e7550f07f6e899ccb47b338b6d68fb418ed10bb8abf41f24ddcf2f995a5d5979fae023882e245e907890fbabdef861dec3ef64d8641ecb6fd531deaab71a8954f7add5b81c024e92e605f43930f568f8a4a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h361d4d1b59a92b6aceca6f8717c111aead752b72488fcd7f836a80cfad4d52fd967ee3573b2a16b1097a92cf0ff9f183ce8da1a3e68a19f3b3262f7f4c68a50920d4fa2f85c3320af64ced8d161e0769b8edfe6c6933fd2b4a9528799ca2bf58d71ce09221a609cf4f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a71c2fcbabac89aed34e83eb7a88b434aed703ef13ddf1baa88bd3076439216704b18fea909403ac32fcbc986e7c8078e9edad81d4bce5c030b284f53d77a56e4d4fbaba5101f6a0f87671695652a37d1d26de5b1a9440a8a752491c149f450cd0443ebae28c30b042;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hff2c3201eda22e1adf3cb1e6aa7899a5cf62591f9ac06414bb82aaf7986c775efeced4e4c3ddbff123b8f8ea2cb54df10fadc556e2f39385b3c6e592dea616e766af96c10078ea81c19d5dfeece8ed0201a20f37228734046e4249df6ad5f51639fca663e2a490104e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h70369ef9d98e499e7896033bb49cf94c0305a27fe5db9a8fc9e63f7865224c29716d7295ad661ca474f137fa1df70325ca96e04115e857debc682557b42cca8213d8803fd1dd1bea6ab6b564c3815ae9a9fc9ba9f1a79091d8e94136780662cfacdd870104ea6f8f08;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b359ece53a57935b2aa5440caebabf9696de50b581a86915438e784e1ecfeeac827c1511cb2f730ac6cabb1d982688cad62a0143b1618b381d0037b6358d772387daabcdd9fdb083a293198d5bbc30f88ff15a5d05653feca350a2403a55847d68303261d2469ca1b1;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h62ab968ad4decaf612d937ca8ba9a432c4de3af6d01df6573a4a3db2bab30f8b2804626486467012f9add16a7348632140f90628af6626d9f2b135bcc54d8f188b61cd9de539747e52873e82a8cd690013ce76692a07f330df76b4841b0b7f50acf26017b4433034b0;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hea921b4d1f71027c619efe782bc26b8a0d074b8d42b79293fb0d637ca65918a7b48471df36a22bb47537b6b5e17c70c44195e382ce6324a2b89d68dcba79e03afb21f9dd7ffd8a2ad3c4aee5bcb2f3256b0ff8e2b70396a47d4f8b5cebe7fd78496d6eb012d6a87460;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ec854c6b462e4851d02666e666e3d04e3a8bb8d1e09a6e1c4f3aee3b762372fcfcf4be88922e6c8c2d9b5cd3353657c4c3055c2150edbf9eb31b94576b2963fcd7d65c7365d3b05a0ec8284442faf370b5868bda5b8ab6a0043ed17e6f9339ca0a08182ce67b7d224a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1372ba00faa4c5a8a1293bb152388072a32fb31cf01e3f9b09dd294968317f0e1208fa589a983626c6c2f20b63c7a4bca266d17dfcd25ffe5ff4d8e9bda9e587cc7feea217cf5b6d0fce5726357712d41e17ec390a05d64bfc51188b9366482bddb9c2b792d1355c951;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h58edab502e8c87c724c04029959aa36a9519c527d525b76ef2bfabd7604c1aa485a7e8d987fd55453afd59da2401895992c6f707d5f7a3c8faf0ced4023e9326a1f07356263a547e7cbd8661bccbf90e430c3a5bd8b2bcaf333fa27a2609309ea544df9d1741752a8f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h19beba2713165e1decf0438cf6f134c1c2edc323eb244c09c52726b38ded224aec0526b2030158bfc9cd942fd2aadd582deea2640250d836d17f11a79451690503e3001b961b8e5bfc4f38c3a858fb37194a4c20bf442aad1bc5925d6b788c7d6589bdf058bf6c5359b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e38594b6d74144f1e5907ac948703580c7eb74153c2b1b4efa630bef8f78a45e00ac59d500e311079d243efeba80239678b448aebaeecc98c62c7cefc3c7e265e9b6c5b00b109ef9d51b8b21bdf86b7dab384b72584f124088021b63e6accbeb627fda15d3d7771009;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h190aea4965128be394754b8a69d3b09b8b4aa4e42da7468ac6669990765a79ece07d62ea42d3e2320ab1abdfb6ecc23451175fe75d96ebcdbd232b44c6a5a4e082a6ab1f9f84e605c488f66e4e7f487b3a6fc8163787c10940e4150e2e0d28b5971c2626aaa66539b2;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h112624c07ec61395e1d915654ab526726c6954eb5965d6203726aa20fecda378a78c350a6a154ca0dbbb3a24c17477d0ea8afbe207b342630bf8bdcbf1df20b1649bb4dde597e0fae28ba15473b4f6f3f2231ffbbe56df65477b64760874016cb3611535f7b006b465a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e9c4bfc60bf1b380451a4ecbe7af266ad6cecc74b8e9a00f6b0996031fb056101771aa4c937a1cf4492100e65fc3f0364358bc99ff1d3a260917b33302c1cab4c2fa0bd63ce83bd95d579829e1182b29fa69b2fb7ed184fdb7a97a3b5a16f7b21ed7a1e2f9ec692bbe;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'haaddda031fa222ef8e1abd02bef65b3488351c412bee638a6f23c3a35d0b2f5f9ca9f9120d03d2cc0678837cb596a429296c8b22044628a5df024c947f6f8a619bf9f86902053d594179009c95546f0a4f51c10b7a04f9c78b06b8f90f23142cef4c8fcee6a1a977b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h74503204222205dbaa7e67e4d3f0e70b9b965c1d7974422461466490e05f62c35eb932895e6b4ffa9579cf887793be7163fc63b95dba72424c55ceccfd2c6e1f71fa640936287c7b368948dddd4cc7d5ea0ec962e60a77534aec3527acb439fc5be8a2474da984db68;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a95adb4e8409bbed73e0163b4de415405e00c4c4e656fd4bfbbbd1513135299649186f95dbe81c6e0ea917ecaa74390578e692b1ae0166d86309949fbfd4b524ac6bae6f8f1d245dd4337fdb0c0395749a60f9bdb8200cb52b12db016a54aad0b154c9923adfacc8d7;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha2e47dcea154e14f580b2df1c74317897fbe3cf3ba527455dfb2ececc74159b3d63a9421397093684048f2c102cbd378cf579412e3cd561fd184b863cf8e9252990d2933a970dcfafea6dae6619927b852e07258e12ab5cd546abc567e0efa73d5b33cd5378faa3a27;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h84ba88e23485d6d9b60275d044f0e1b88074306e9dad538becf4266648d720e1fa8260aab00cbdd9a358a0c6c64fd708d5c4877ad1bee6507f0daadeb6c050acded5860ee99794b0c0d3f37d83cee6bdbedcb853e6aa21ac6945c733cb214cdfbf184d178eb0106f3;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he1f73aa6e5a9ae6da6928a8ac8f116d0e82644ba2556d837f4998facac0ab97671e7e71d4f9e361298beaa7c7f210b227c422453c66bb526c53fa1255ea88d045498462c0fa61f7c4aef8ad60d9007954fc7c957a2e5d3998e0aa55f4550cb270e77f36aff33caefdc;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b51690686faad333c2faa3b59a41a952523ee0ade57b70ff3f72e742a3ca4e5706aa4a66550db5f5ea83d3e959769c36ef5312d98f9a6ffc42aacea7aa8138451d7f74ad377692646e689e86cb41b8d3044cd2ba11ce05a0264e6c074ae71d5539ec1f41dd1c441e43;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h6d73a79f7493498b0dd7dfb0d5d6a15ef1acb9028095dc52fa49b3e4cc4c5b02d27da0a289c9d295d3e229e87ed85679cd412cfd75e9814f3903b3f28b01d1aae13c3b2d7571f1a0d366b3a98598c48880f975d74f4865d9ff250269c1ce04afdab8378b7b06f5a009;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h53e7fe1dcf4196fb84b835b4230cf464ef3b1ac3cfb7956d5ccfa01bc44849773b1ea1183880294ebe63c64ee25771fdfebe4243ff035e180c1fe682571b31e03b8b96323cbd32e63242dffa50d4cb5d0f3c934d3f3071ce2380292e669f0af8e2c9801223490b3407;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10aba3d5bc102ad52da75534823e6ab0d2d39ae76773a6679e340d2f72c81804cf054589d65ba61d4dd1963b2f499abf17da0198c32e740d5d7716588ce0ac23abfbb27a8b31418cfb672ff79d09aa60be9590319cf9e16ebfacab77eee6152b98292d622adbb12c287;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c50a20fcc8a4808c966922eab0982f77aed6dba3d9e78d935a2dc8b83b5f71408c11d37589885e64f1ac0bf28518b54c57af56be7a2ef981453e52a66ab82b9f469f1ae3a4188bcf2f77d47deef1a445d9729c5df0b1f5043628b1aec74870a7ac6f9e6e5f8f735487;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h141f00610434ffebf98d2bfef973040e7f18ec43fd2c95a172523b45190493db046eb156dac09865a1e5d49fa246334ff0ad169c05d95bf013fb433a2328648a4a7ba748256f6e868961f67e8039476acb11b5c9e3c05010c25cad2d1fab946f162ab2fe0f2103c113a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h73fe6f32b5154aaf735ec2ea7b09bab20767ed59d71690e4271fd56665c517c7fddcf379b38a89e45919160429b34e35587d9b4d5ba06dfe484115796282f8f1c2fbce9ba29cde507c3abd2a42819a9ad428444010873e5b4b8ac63c800ad018a2c715beb535e7a196;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h4184363ad3a81a77c48b590acf9d3f309316f85a50a4fc401cbd2c5fa62945b5472bfe89f87b501b717cc9a6b5ebfcfe89f1e4b3a472eca183cd3d27a6a9691264c93c0f8f25ac60e037e48db4b792b9546e484e3843224918cfa6be004fb48308cd398a8eebd14e94;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h28d327ebc5616337c7b65644f9a35f4c285364659eb5b61a6c6c7bc4459d21543d3e3827afe214ae80dfaacd09998c0b0ab2e68458fcc49455260900d6816942282a16e91f7984b062447a00e682040155553fb233f0bc0317c05b83c2d70eb1ee568bea6d3dc7fbad;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1fe8ddce15302e6dfb928732eee73981601022e948c3df3ee5ca00c3715fcf6d39bbe203ddc52c427372c9a444b6cde5352d73439ede16b4fe78746e4f5787e773bf1a08d54a52b429e8190b8f0d5b8761c12863985d700bc664ae30fc4fc8f1d120325521067d701bd;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f59db5f2e07028ee84a0ac15f63f4a65281fba4c840b1f45e47343f8c7b4ac626a2db90a3092d5c243d431059498303917cbc53742b425220b976d0a256c5b5cdd1c6f362180995fe375bca34b6946be99ba9577f1a87b406d8c48e7c81915d982aa97e83ee16b8fc8;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc9fd1c4d762bb863e312eb5289ea499c0953a77082248a135a4cc96ec870cdc29141823187b82d0fd255cac41cbb0086b1f8a1afbfd964199c5a919acc912c16c1bfd6904e6475ae9f7b339905fb15dd9b1c815e239bf6029c17c6c847a6503ea203f7c9f544c4c491;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1410f385a75662a52c30a4c73ea18b86f16ef329ab73c8464c9db4db6cf8aa32066619754deb24ced2634755e0504a204f9d1a53d0f8ee89fd87eb01bc8d6fe9f9426933a1bbf164c4dc54c08bb7a0ab6a2e1e40241f316f91df27c166cc5aa35341a12b9b2694208db;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h177a0fc863038dabed86f369f85d976924da42096a6df42176437504b3787d555513de18573168066779592fa202f00c59914fd59bc2ade35ebaf0ca3af2d733b4b81c019a5700afdd6a7739554538cf32d1cc9cf03462c637c931a3af897015461e32a0d0656c62bab;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h997273c5e48d811bf327554f758c0e6f7accd52b4d1d0d80778caeb736d76c2e1c8839c2972d91718779841a4908b6c8ad6daefb34ebf2796cd4ec837ac677ad2fcfb1e13adbcdaa054eab55afc13fd604ef902c7988797b2b3310bc7123f7657c76f600710328c8f6;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h12d5babb40e46bdd3bc4b1ccd9853202e70f8f6dcca15c338c015a4f64ec729fcbe007e483150e30e36586a54c5572083b5c7434ec93236ff53216c1a6fcc4f02eacc1f1ea12265135309d9933c11d22bea710a5b98461142a03b2ec70d5b49f2290ae9338fce2612e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h330ffd4e1ad209fcc373da21596d238e82be314e5bcff754ddd9364cee6267199e6163f6e98d926b5d56835e30ccb1219c2c5d670fb1566303048d6ac3ddbd988c18a605d333443efe2bd0790b6eb38970ec737b783ed0211b3b2e02e5d058bb2f8216cfa7e604307;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h76e05c81aa0a260ad12c7b928b122780467beff20fc1d2aca823fcdb6b7eb1bde51de7104062ca0a31b154f9e80cbd62b41325c6fd78a87067749254a77471b9cc90524e84feeab7ec667eb5e25a53f6914cc533491e32e471903392209d522d46ebc3f3edddb512ce;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d641d6260a7634db6d970b59537f9564395abdb1e52160fc04c70cb0b7cf391c6592efef2ba8a644f695a378f2bf12ce654b05810281f3d5daac5357b048ab9941eb62ef9a79011d5a5a64a7e88100310311c7121c741047ea844f65e3303af2839ba1bd7bac8fdf3f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h100f74fe78a7a1bbf06c2a0f3f84cf6d7caf1d4bbefc2e417ef1c454a6185ed4501e71745a59e57bbbcdf534b23b04a4310e1520139ba55c7e5fe222166a510ed941a06427777cc3863d1e330bc923faef00ae484e93a2ae3ff21ad167c8e358c818a76e7f3301a1e5b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h71725f64f556c91de49ca3ef2bb2b568966063f631c00c70d2b42858f555831eaf523a9b74e7041f4e9794027943e2eef82902323b585530992c4e3be5e57e057935b8a570fa43b51227110d31c031249dae1bf80363decef19b281e375c037bbebcaa3a4b558cd906;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h3c5988eca97e9b355523070475e82eeef34bf2e404960699c876a91a7efb24839046ebd5559cd62a9d5ce82f4327059d0dcbc251bd8ee180f534062f3de5906f0ab04c6d121816fb85bb84f4a1c4a0b2f8b5fbe5bcab0d17c334ce0787b86944327caec3042ee24677;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hacf00d302eaee8937872533bbaff4ed8d9963dcf7b92505fb728e4be3f2eda18c08ccb73cfe51977ca45c3bebd1c72bd8219c6088053bca5021ce5e29ef05d8fc2bb7e82fd25800d47ff071ea5b91db5ce6d5ba9a16d5eff3a689a32e26c409c6e92e760d5965241c4;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd9abdf65af95357f743b8a45cee28529dcc47d2536f54562896a1c05b71c77ce2f2fc64444d5bceb39a71fa870b7d04ad3eabf3af9cf0dd5c23f7aee5c2a8d3e083183dc971aa673c8b32c37854ef4ba212411364e8a96d668aa5a442e12d03ad9bcf67b23827549d1;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1304a2df2e5880539250d617882f4692b1810b9549924c5e0fd6add14f87d1fd350d1b46500c31754dc19c9c98788e8c543e57b4c2e20faed174ab53c58db8bad1f6743d4c1bec0050e58620f3b541a96354413ad40b9fbb2b6f55dcea51a62d89a9cd89fc5846b6b5c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c3ba6684ce40f5973c074e5716bb0541945b443f90a8acf4ac27d4ba33fab4d605989345cc9138402eb7d6b3626606847f9543933e9bdcaef67c99ee67361c72a3d708d2e9d73cc7177fd35738adba579f37d2c3656fca11622c8764338cc13b5b5a9a8de8cfa8a233;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h86b56a8e92408374da7e73ac4b826b33750ab48f8e6329f6a6c961906c0c2c9ba5316851ce27b366e0971f64ca94631ba9bad3acf33514f245b2a90188347ed26b986c38b63a9dfd2404bc6dfe4216c14283758a4a86a21dded863319f231679b254b9361d29db751;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb891c31937db393afb5638fbdf38b92ffcd8c892d3efc5854b37a040fcd735d00546966e52b1edf6f4a5434036200b6664b1bda06c7896b6c526777ed0d64c5ca6d9995f09716c92871e05c774324df21bca411a7a8dfc0c6412e8a7ea284eb59a0dc7c748de5aecf1;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h973dba9ab6cfbed0f0ab9d1d0e9a929c520c47d34fd8861210add18853557705d1fff6f270dbdec4723f73ab493bd9db3fa5868eb96b4209521ac0b87763de81b47b86bb4a078fc533868800308e97f5497c2548e9175a634c902267e32d4472953bcc1deaff2ad84;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d663d8e167c4180e364afc84096fd8ef4f0089278d72baed6b2bfd4fe4b7c4e5889a08b5092f281bc23a97c6fe640973021cebf517232cc450e6faa6ac66a52625d266bddf6065b074aff04394352cef9ca1cb7aae5300a321d1974ba90a140be180531677fd1774f9;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h174cc62da2e6add46b2425fe0fea387a7607aa6ad24c12016e7edff6dacf482ed67ebdba0b826f0e5fe52f05b2a1ad230aba3da3729dba6adf043f404033059912b257959cb995b21539102cee21bd75bd7ff0c7484137fb2407b6ddc3319579689897b7c5301020e1;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1af1ea7068eef587f3b37a0262d8d65ee73dee743367cf87c0df60ae7df773e2adc1c7233d9bb503eae133eb2f5ead00ab75953ebc685605814ff8c0bec59eae213f158aa92b447be76779dbcac4a459b584d28d1e08c2b2ea36e9745c648301488f6feb34f3b5211ba;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h11aae9a0d8ba1754805b3f1ad9d7de7103ac2adb907e3ea61e8aa6cfe4da4eeb7c4b77277f7feafcb02fd3fbe47e0166f6e8c48cf3f02e8cba17c6ea6cc7d1c9c4c56a65d640ccd8ebb5a46044be4a366ce31eddb492df4fad65edf0f7122c2fb613224cb4e43d3ec84;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1620b312f987f652cd2d837d49a55a9ae2f95ae52df5180a2e0cf31e47d4d0bd24127a89d749524b4558e581e4f53900687a7e4d29c3889aa15ee55030b23bde3dff078401d148ec4a7ac8f41dfc363753bc267779ce567ef0a586a566932590be419a0e147905deebd;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c0a0496c95c6c46c7b8b776dcf48dccb86d0752707e59832a5b1147f1cf07d74ed8fab84704ef8308b31b2862939e54d97f92a539cac08effea723cfa36a21dc12a89d6b0689ae06cae23118498a5c6a9a1945f541f8d1a83e3597211145e4df584ce8e045c35932c0;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h32bfb2812deb6a9363e320fe4ecbc099ca1dc45fc27adb969ef7aeaefb041b7be93e444ec10f882e3e8557b649b18ce1e919ce2aec2c272af99133eb36524cbe5bae2bde36031dda1d0b0464329f0f12647cb248ec3971d087c475bd3b601d9a22d3fdde0cb92493bc;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1dce499991d383100c42bc7003cc88e1d080afbb4ceeaf3a9593daebde5ee5ea2a0a148a0b508f4f4a6c1579bda35f771b5231361d7f3069f964b367ee81302add61eb7565522cbd723315c9b49acc3d440a2cef20f269c45768249225edc4e884daf9e8d0350dda08e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h13af919b79afc9be203714ec74b86971b0fb27d4e271b9538389713dc39fdab31c3aa072e53f889a6db70b1842eecae6341294d1c96b9d83213294ee086fb37980116b61ea2388d2527ec637cb70e194055d4a83a029e9d0d5f3bf7d4dfeb70d57f69ef07a07f081630;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb0c6e13a999b4db9fc22209dbf4478818362ea9d25f9440a65616c1c749a62a4ad0dc7cd12cb33a5eb7258c412af00a09c732e84025e70d522713066fcb3e52bc41710fbc845f23320c402efedc22b8110c8b77b4d2ba2524d26be1b89862d2be6df1feefc90a66996;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h150110526a0b643c3e50f08939b3ba17a5822ff8a141873aff4166bc3fdd3887821802b5f26706678a618aecf0ee1360562d4e6eab5cc777a35115f77be2325dd19fd9c3bcf6b30b07743083cd8c0181db6467724c705356b32ce25a9be28a55e77546ce584930477df;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1994df98bc55bbf0f86c2f175799478d9722135a5475fcc11a72d126fe0c9bdf4187e2ed07542c7afb0f7b6caf60e6fbbfde03dc0c5daf05fceff3e6ef7fbbad03ffae4d4e7d92b7447906e238e24ced78d6611468123752da1832a1c48d095cf8d5db8981c688712bc;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h37c85db53bd04922ab0ba3e715fe9e5dfb47769cb26f3350e613e8c0dafa1b61b759b66ca87ebbd70459bb32e659d93390aae47ac970a2729e4f022953d081ba0e6795cdee33f1bdd9aeb95c622cba12bd9cfc6dfd76d5889358ed5071143a9da4f5bb5902e84a3bf2;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hddfd1f45ce2c108192d03407ce9cd9213059878921cc52c415f48de78d4a71a0190ccadd80a60c77d378a6dd489b4a37a6dd0781c22e8f808229d007dab0d2192ff7b0d0d6aa50017509fea75d5c41df52b38fee9cf43d52f07cb272205422ba10f0fc0df40ac1fc49;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h172c294d9ffab47987a14974c3ef43a663dd19cbcbda705eda7e4282b5bd326f21aa35fadb37ed8e80b95123114d373b34c507a0384ffe6537d3b578241c4ee2dda4a3f8afdedb780dd1315e1a4fb54cb4aa49d3948baab76c77ed62fe98328c8817e42ff4209080bf8;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h173edde150f74973624de480ebbe825146f954621d65f8b2a00f014217a0efc5b415e2f6df1bd1a4b2b6d069bf8be93f60de943177b5f80c00901d26a86f51b2a71181916c33e613989c243b797af2f084e87cc9000823b2caaa03c83b56e4ec578dbb038ec04c0bf35;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1fb0e0b89f6cd5a31ce71714e05fbac3aac277fb0f8c2b3c0eef7afb94d80f4d26e4c81a60c8ce94ccab0647315f2585b894718f60d18ea22dbbfa9430c4703b08a2cb1c27a8fa15116d2dbe2e646415a42c447bb77083ad21fbdf5b35b5c13de68c1280f82fd1cde79;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha5b7610663b2e599d5f5af38c4d8e29e99d1fc089f819d5cf888f71e9439b4fe707d9fa4e944fc652b5cb992679a41c1f51df0c8cf7657fd4b6fec0eb151ae70342b1ef942b0226bec0a42a63454e1c64ffae899fa5519896bac8abe0e920e9a0d73659e4a5536cd5a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1271a8231eae2d55f3be35607276324a00750238432d2b128d94025047a7045b6cb97784a935e9fad182557dfefc1cf1293ceb8bf71fc170b0b7f06272dd86ccb68b1b3e7ec17082658281e56dd0740660a0bec435755625e8a32998bca3bce02753567e7ed60b3a7dc;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1988f2965fd68d8e4889933186c93f8d5d142c13d6f8241985edc0f8c5d93e914da39d9e07c870d6f093d9e4cef87484dafdea16791f90067f3c1a0f8446d345dabecf55305bc434390aea0bd0ee186dadde0723c138784aba4fb609b633b1db5cf97c5973c0da4c765;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h15e86f3b432445fbb34be01f30a40588db6f28ff45f7a43bb767f81c64938f2fff5f0d03d48170422961c2110d1446e42fb4eb3d7e6ab4fbf0c1ad1a94ac475b1d334832c5123d68a87f64e765c01e3d429fe1943864552bc0b3dc72744949b32c8617e8f7f588e1b0e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h9f0def8a0c3fa7c043bfd7279fa0612cc5947bd6ae7b2e1b2f644e6359737fd96f127d7f242a862b0773491ddb32a74af852d3ecdc5e5ff56ddff73705fd344a02d40b702d1a24088740c0f91368a35ff0363bbad20d9084f2e2cba9c3a7adde5ce323c8df591878a3;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hcba183a53e2562a1a91ac0d88084d221842f3749e779381616c7ffeb0e178995edceb2337b0379aa017193b6c7c727ac7eff3eff89a5d3d81ebb868e9d9c53c25998398c63f2d8e1aa70d1fda1a6881c892f07a83b67208337c56a54d38800e5b8c347747c6b23010c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf22bb0c5d5af33f46123eaf07a6bd76440d122d30c956fef45b76ea3c195ce9cf734625a71e801de9f942322e7371c34e4cbc9e0e2216d8f8e3d0d0638fa8cf9799c590b8895b09a56d025d01b3287caf876433c4d5971229957f540fcbc1e37946cc1a118976aaa64;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc086fd29b104b26796b7f9b736b164ebdf96e77aea3a33fba7a6f2d1326c31c89b990d93c7728260aebd5c22325e5813772e740cfca3f5f53d81bbbec3afec1ec4e3bef41ceee830cb9c2697f3390015a5b75c27b7ddc38b4e80c7eb0c2effc23fe107245028625ef9;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h12edeb4797789d11b1057ae4120fdb2a6e7fe1444921d7de493a745b5d7bfefcd7f2f0beb647cdda60663fe4e5a53880c545e4a430466ec97834b293d428366a8d90ef8abcf201cf322d925759e446a7e1d58fb9fb46dcf9f4f8e21fa9c67cbb6b35a969c0d23723e58;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h11e5aaea4bf681e3df51374592ecf77a7ede1978ee3b09c7d87ff311453fea58f0b8d9f9872f52d9d0515be752574b9f479e39f1f7c2bcfebd7690f89ef1e40efd1b01185eb8a90806a2cec26741c5fbaee9276d7dea99c655f6a9d86f6aeea1127ed7221cffbc12989;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e31cbdde1a8ec9a51ab1c99132a680d89845b4916dab150a1be42bf8c0f5d9a3fd0e2963f174ec9b5ae5e72ab9c2d11746ac58fc246c5782dfe3bfb9ed88eaf763bccd880c47bbbd3f26000b03e8f4a38c21a68dd0971545621751b0c1d77a98cea3f84d96ef3aecb8;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd9fe9cf611df3c752001cd1fde4bc65d8da0714bf72899d9e213051a689f0ac7b18885447bd69c808557350cc6f900264d8ca82c2f3c853939bf3f0ae074b418e36400ad6b6f2e501d96290be34768883964cefde1c1bb84b7f30fa219abbadaa184fab5bfeaff8aa7;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h11c35726c4dc8ccbfa68ad86ea79b0872a320bf06081786f5d8e95460256889a9bdc1c8f7a82813081c435e066c22c37d6a7c6f818650ec3cb66439aaafa53dad015d879a31b5a4be91dd8229969eb1615d5ab44f157425278d7231dba6e0f4c8a48ee039b8504c3935;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h4967dda158655299b11a16c4650a4624d295deb7d396050a4499710497369829c014e5ce35c4e56d7c579e7bdadebc403d16ba199731100aa24560748a67c8142e45f5437990ff4c3d2c566d58ef06e6522b3bd7cbaad9383a1832755703c02fb857013bb475fa49f8;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1626508dd15f800b873af669ed12b8b06380879d11fa479ec5c0823dda02c04341f7cd1c91ecb4c4bb1dc9e51b8075e2117fa459ff6042ce9987a602dde35ad2fcdf5248cfe699312f3f0ea153292cb9f787bf04f607f6e1d2395ab8d373bb03855471b22b0e51b6edf;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h65a39d53eda50e67336f941f6a91c2cd6aef1ce81add02f346c981e7660ca8ffb5c8cb5600655f2ed4e92531c3e1f2de0922dea2dfff6768a880c6e7659fb6c8a2231402bfc1d1a4190dbd8ce8121d66f31e60aeed1f47bc00d47127b2aef59e44d120e057b1eadb14;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10b94ddd3f7e18611d14da1be49a7b5276468ca6e07f4cfeb678b298bf55a02ef9612b401d60824f2cdf79e46bb7e9747d7d7b3f3bca69e59f23ede6b96450993ce7ac66e225e43d9f8be04fd4d1f5b96150ff9575690fb6c24a1b7fff29d0c9f72d7e4a0ae08b32158;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10a8c9fc38a8151888f0f20bc5a03fa591789100aed5d823afe88788dac8e64f3db3619e9a6fba713ec8619f32346359055a8b2469c416e28939d06ff82b3b0716ff3d51cff1d5aa1a14d4de9c254d7da87b48e6bb4ff25032c03b18b6dc8bd17a5c749f6302fb3c451;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb9b4d0a11330805348fb271882218f6e3d433c86a526426462670d883cfd8753cb0a7ffbf1f6f231968b3f10a361add68c4263ff31194c473b04b5d177066adcaa90753c045411e9286433e615f7317e8b1f297c4b7d4fa18f437bb5e5b66b99b3adec9ef1101582cb;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb381cf2ba3e80c3dbe7da94066b614f117572f62361c239605e67e3a4ed710e6da19e2bedc3fa8c3378913d9258c5fbc848235915447032aa1f19462b7934706a72d8115b61517d4d03e270f8e7acbb919931e6099b6edaa9e6dac5d0fcfff07d888812d92d24544a8;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a921bb2947154964b28747c85cdc475d53f1f5aa34fa40980a291324c10e3128f4828e048dbae70ad1796a6bd29f22efd2d035049e6ed166d81d553590dc073d1a76734a9977a2ce8216483aafae32890681b29976483cd7feb8ed16f892c7df9081b6a71701f7b3e8;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb5eb499a76417aaadf5d9f6f1e6087ba53fe5ad0ba31759596b628385e128d6c1aa85c9cc5afc1226c940a101634a6678af84868a4dcf88b6d72f5d44539aac99c3ffc56f028358d09f06a79da083fec0ff77d24570d8a203e15ee4ee2808a70770e92fc2ee4456a5f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h3bdceddb611abdb318bfe7244ccd33cae8af1c781f95f5905dcd4c98bc94b371e6eea2dd6c34caa105817a592e2aa409fbcd1e2fa23a35f36523e73da4d8ccf31b7da9cd3cc635266ec154cf1be7dbdc5d8370a3608f7ba7055802b4b29e01a8d1df5ecf124981a63e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1369db165b29290e8ec103a2534010bc3f3f125b5954f700076ff50677ef6dd8885c37169c5a184d9e0b284b021fb15744422bffaefc8a821074b61e95d322b1b07fe50d1cf380783cceab8722b4a37f1c6e38e6279b77b1cfd07d1adc327fd4e770039e662ca33c793;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1554c2f4d313c1d8937d6b627259af571253bd1cf9200348cd1aa12e371330a526802cf9a481adbb776d3c03dc38ad7b4d9d41cba092e421f50a86b942f2784d0009e4cf7e43fea62f90da5819b09be1621e2c422d7c31aff298bd83ddf6fcafce2b3c81e10ca57eb28;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1be22a59a8b87683cc6f6691285f3b19f2ecdfb13da2d442b121f8fa2d00b28aeb368564c0d5fdbd993e4722e0e92359595ec8d71f3a5d3969dc858c4a4581286f7d1be1dbae2a0c72809c28e99dcf3a3139ca752ac337e0c5b5d4cc24ad5e073a0c5f4385d947862d1;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha77bc8557ab792cb39d2ed82e1823f6458f5400745b19731b0474ad4821c3eb7b5f25925b217415f577767c16682d6a52c5f1822f460049009f12cef8142eb719d0653eced15c1cf3905af14d8861e93b66a4090ea778f942817cdb164e60151ff9dc1cbe6deddc3da;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h196f364a57eda2614a024a14bf2fb165913fbfce0be6f5d1bbe749ba23ce6886e9cc002a3b590484647dc6dff6c2eede029190ee660cd9bf6aa117fe858fd3c547f208bb72acb234c475a141623255f8739e733e554521c7b3f440a0dfba28e509b3ed87cb191b4fd01;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb79aac51c278d2b9acd655dbf30374146b31e36b23ced0dd545b0fa0e25c3c19e3c350b29d51ce4f8b7474d53fe447ad61923d5e848e1f4d7a790305acdbe5a469b8f0b206543c9b3bedd224ec33f93058b076ea1191774e75618afbb5d57613b8bcbf8bd0f7ca144c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h38ad8462c274050de6636a989fe0b24a671be0a44731928f1736c5eaae516cdd747ec42d950826b98682c9c202513e0f19a8ea74b2d14a025241b21ff6a621df8a8ff48915e6635ce36e0b3ecd19e1b56058ab8e099b7db5fb3ab35d62689c5d2b52e89ece114b5f7f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1aeeca045ce3572261c84cf025ed3f88bec6da8077f638de84adbc3b3149cb8234ae2f0c57d7fd08b4c5b2bcd1bb8bd85996bb49162db8c1852f206fbee289c6076822d2dfb220e22891626ebb2f5d8e346d4985497cbddedde2d70582f7699b4723a00fb2fcead00c9;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b05bdf193f50e20ca55933beffc315ed1433f92552bbd7eb627d314bf8304e1cd1ae3c024747a5019c8213d728631915fc430f4c4b8efe1f900e70ad9328663a6fe6e8776d3fcf7af6861e4f37d63731f5fd089161330b85c515a9000995c0c4de426f1ba03bf8d35d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h16f2b51c552cfa8930e9ad427a50d1a9356e62fe50c36f67a37c5337eaae9530864dbbfb5f26431cc5c2b1a64c426937fe8302deeaa8eef7d019990ba2e3745cfa77c3ba9244a156976fe8161f5efba68bbeb4adc20baf636954b2b5b8d9218743736fe244dc4bd342a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc6bc1891d660575993c039715b611ab8c353169bf234864db012f534e454eff74a870b73e149d1f9ab6e78880d0c5f4ead98cfe7a41df450a3c5e080d9f0646dddb02993173b86a67b0441d319fd777195bbbda64a4e9b737ec91ad72bc1eb21c2aaa2d93a5254b8d3;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1baa79bcb3a562fc92fe5e90432615b9c8a902e23a48dd1219bb2f007bf40690117f0ef80ab766cf06d0edcd60bffab71c0cf58e99e1e3481ea507140a7a93f401ef9d33c1f27682ed97c987535b8b976df65bd7973afd8d9cb8e3da6d04c4c6383f2ecbf88f609d1c0;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1744ce5834030f8cd78d4a6fd262131b3acc898d896dcd81649d9fbbc6f3b7a468200f35bfcb071c6a43acb5d372f63bd5bc23d82b218f9aa63811aa9cff63d3386f90e136837157e7a5b04bc6e40f763b228d86e3167b0f50ecf5b8350697768c2d4a6b0fc0263dc35;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he461622c4a074930e5df45c978d607fa0cc7a8e5bfd59f33bc359d94d1ac476ebc51f9f48eb216ea4ba8b7cfa723b4d350132604b73b8a7b0fe4098d9b6011f1d3428adace9a31e18f88c80bc9d2925b061d47b263ac1fcb29296400abd6dd85249d54e10e0d46af01;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1972f1a93c0e2f874686587599b3609aa9f33ed7e6eed6a4c2c91b8ae3f922ce56e7d47a6d218343ddd784c794c895104f68561bcf9175f42d42319fb501cd8024d74ef74feb3dd7828b2bdb2d8b13e0fb8fa3a9b633914e460573df6024b4f028bcf0c07beefca9015;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h13f6b2e4472a7af107322cefea977c3d8f37753f4eec8ec9cbaa86d75a58b4acbec29b4c59d8a440647c4ec5f8717ee27f73578d47608d08fa393b9b18942bc146fccb38afbb19f677f96d8b8cb6533e6997223b57ba7505e6c00de88cb6e6bebbbc192273d0b4b2ee7;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h311ce3469a0fe113462472c97f7b7a8c083a3d7f17556211b53db7efb6fcde76a72243731dd4bd8004eb30dfa1b8ea4916249625e32b7b9e74c51ede227d53e404aed697820c0816350025c343d64356e0de9dd48cd0789e96f72edf466f39627d41b8ad142ef5b95f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b1b231f9b158550f850e82f4173d44f810445400eda969d6de5e9fd184026eb5e38913dba889d98739cac4266b220e71cd745ee257ceccc08b62ba7e1ae1cc0d905c355b09efc1f74f606b62033f9dc09baffb0f729b44b27c69bdfa14b4133b913a622725ecbd9222;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd4f2f0065e62145222a933d3bf342d37071ea44003eb08c000a5f927489773c5a84bb0581d5bd9a3eff55c1ea0d987c60c1a29313a17ad22687d14b74857b4ea7ce2bbbbf04567c3b3d2710bb7cc7f31416ff6465018c3681179cea836bc8ac8d6cb0665eb6b0f27e0;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1763d83d57fd2ef9439c25c9bccc4907771dda4a47407c1b22db208212217cd3b2aed717bb2eeb95d451b0bad5dafe61d86ee520cf618143c898609d3a8bb6dc51416e3f4e8ae1457f4ce3ff4145b11d32362ea5afed493067e6222bcac157bce25ab89af654593968d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e8a8a01c0648e2cdb80daa588123ee20d7b7e6be3a9cefd3af176c0b1f4101d153a1a94a293c75adf9b43ab1720a58e8fb84e9cb71f81b36afa65f0f3b643bce53bf54768a1ff2bddd04608ed3fd5450342e544701e1ffa941b8bd6bd226081dc4a60c9395e29b0d57;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h175a75dbc3b0712b4db6c4bba2a7d30641e24bffe74a7aea847bb6003060fd9eec2f1c75adffcdfb7e5c035891ff458009bf25774f083d6356d7a85577f8514650944eccf94a35ea2c07140bfea847e7df81a1c5e571bdbfe2273cb05e471bb1f0e88efde4680722657;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he36088baaab1937581ee7beeae20d0d71d3862b488549cfc0efbce7a438d8ebb9261c32acc1bf4b9dfd2fe62dea9569f230642b310d31b6783cb7f358ad75d052677a2acae7a91a1c5703ed951b8c2cf7be00ddae1b4aabe50892a086cf08535c695fa6539902e3413;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b985ebb56d7fd57110603b53a3bb8f097b7feee1b9cf2285ed466ae5307978e5fcb2dc5e8ecf41df1637484e9f2b1502b21577462018c734a7147ddab5ce357443c4e48a60a6b424c9ce5c74f6e1a90c536f48326333d3967ce4594e4677b4bb54566a4ccd64741f7b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h38e9aea6523e9050acfe1f596b6345dcbe7ce438c0a145d6628abc05650a8eb27f04045ae65d0358a2d5acbbad17f57a9624af443326e0e73b59082e2ad0c36608f01e0f79db47848097692d244934ed1b174fb5499d25945036501ce1b0e66a8056f5571fea363e85;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h11a1480fa0c9a6bbaba94f3e2191b98a19993d7dfa9f7767d9131f99ef4bd5f2cbda2b1715b9070757a5f86368e85c50a75d67b2f492ed07033b3d2141dbafc45a4a60a60d3da7e4f3e07dbd4e6d4a1547f816c34c255dde2e5baa00e77569b34742cb49d842909141d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc099e0fa4b1b7aadfdf09a346b551ed2152a227c720e58c6df280d2efa98d89530c618208d676c8c39e12e66c090d7a70c8bf3ed1e8c0d10266c3841445cdc2b8e2ad52fdd33ee9ff748614c4dc4aabff3a64a0284f668bd54c5e8239b6af896749938c9daf6a4d67d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h6ce08ef8256bc8e13d44bedc763fb14558d2e68ed3423999bb2ce8582a26ee72299f9e5fde62f8ee637f1dae2cfd9cc64047346d6c2ca1a5ae4c9e971068cab4775f1d41e23a9c64a339ca153fef0e8b762da8542c62bc2401e26c4d989639198da9d0690a693bde2c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h162d782d79be08daca7d7f32fdcf109c2b970dbf010d25b2e497720ca3984ed98ecaea55fddcbed1d1d580c6a5720320cc91ba481164e0753be21b9044b6b7fe6c306283290fc0cead52140a696700af6b74056b545d5eecf6aa1ef5fd22431691a6059bd5139bba422;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha320c5f5bcbb2d095909534efef20edd6b0b08ff9532c7c0cee7afc9c65f7497d36fe28fa8feb069167a08f5aa20421ade0c3e183dfbe4323140e6424394d0c6b737d9027c99481ea0f5ba3fb4aaad36d764387041d194cebe915dafb57eb858526c1faf3032f65e81;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10a6fc2164cbdda330c6addaf5fd7e15abc932c816a4d1a82b57f93a0a68145eb3177c39d38bf1edb75c91f3115e689acc2cc9409b228fbb7216b9f01b55391639b6de9929ca4e4d129b372e9d53635778df862ed6b59f4e98998a2f2c5a3810ae9ef518886e716139b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h361f66f844d428da54ba4455f7ca6aa234208e1cfbf3364e95bf935c5f922b813f933cc33eaeafd71b918453616f214c6cd0fdc997283678561b2bad698ed78bd018810352dbae511f319c215a9fe9873c01ee0cd365c8a49b906f143dcae7eca250df3a2c4446c5cd;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h8ac1bef52757114be143e079ca9e74e2d40539def24116f82f13a1798bec6da8d2205fd8e0577700f03dc2d1e744a4cf566d4a98383163920c21b8c65e65bf52d7971c1f3ccab5660f087cb4c0e2703b782e07f6a857dc070a5c0f2f34c4bbc4fa298da77f756dd0d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h16b23b8c2b17357fdb5483a35e44bc40f339a20e7db04a430e8f402646af21126fc42b81c4d6c4dda5c80aae81bd28897ce7390ef90fe33fc8bbfdc4196999d90bcbd97f9df93fc523f36d921877a7c276585599b7a690500169d233d4d03d3ea59342ebca7e6d3ff58;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h2cc3f9ed8880d326aac062eaed129e4b6b977b647eaaded6b05f1e54412f6a829da86436e1bb07f6eb811a0504f8747238d3aceec41a78ac816ec59f85152d4b67300c7a7e9f582b8e52d07a19024bf09f9d11874aac348bdef9c1c2269b9e57680b95f12cce7fa571;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hac8ec843f108dac83a87ee2cb482b5c3b45fd094b2e8101bdf2ec56d9c66ee241bb867c2313fcd4bb7eaa4dad7b85189df9ce59dd692f946cf9a44fe3e0958dc9e1d214f90c1117c2ccf752afdd5c50b309ce422806756f56602ff1c2d3051a072c9f729bad92c4a64;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f2b167db33e9b4d3a7132fc10214a802c7e5d441feba19898fc3f26fe2737dfa239d0da6ff7dbf8bafc6c327e57e76554bd161d72483f4afbeeec7a474253ab09ae405ed49d4e8616b904d502e4d4e32354a4489792a5ad991a2d2cb4a7ffdfcbf6ac84b3218eb2978;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ccd1b4603cdb482b9002961241f692ec8f04a4e051fad186aec6b2904dfbc4f3496eb38b3fc8ab03df4502de2aac21aa1335dab56c951e2dc6a2c652a7adcb38ce03777723fc7c9baefd26ee3bb321c49dd4839e06ec54e818f767b56c1a2fe2d8df69bdc1c92d3d55;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h17d50a0039130b40bbfe89b9b5284d6abb702cc4a80f140dee3ce9ab49fd07388253de217a882c9b85bf07a089d3396139ecbaea390833a374f4d7eb7bdad9f67483a0e24781591a273886d409698cf8715004ba9792e42b1e6b16757a19760cef71aeed58ea898630c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f198863ccb5970d5683937a7d621ff9aa38e9dd1cd7c96dd4811d8c09ac3ff6ac61c88e393359d4051e689d618de647d7843f5fadb9b62b565eb0fa4a16b8e79b65c9bde0ab2e66cbab35b199b96e34b0acd6578148b7de8f1e6e52fd265dbdb28da23c896d07e53b3;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d626074ba651e5e9022fb9f297a028891cfc1c53e8a6328919e25da9c2bb45f737c4a63e822eaaaaef649cc8b8655fd3ab227314cb5cac98018a796b8da98d8714e541e432654575ed76685e11d253c27dfca07ca0f38843a42072e269a588eebe6875c7573e635f3d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h3feeeed79138afe0bbd69307f08f895ac2ef4bd73063ce229539d11b69d20db416c3dbbee2ccfff489149809d24486ee1cd8e7092f55173f12e485a53b932c3c09129e58fb1ec35d3cc1742d0800be8221c4ff570a47e8b35ad5c18d98af792e7a43382844f5165542;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h19837f47f3c6598c633afdc4c8023b78bd60ae3d114659c4223fdf2348aaeb462e59c8f4bb4abbcc41a104b04d2342f3ec9851c9d46bec0c729bac12450a063790537d93a31d2e287304e6bdc122d0d3b909773c228253b7d6b8d16328888745003f54ab5fafd6383e1;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hab74b1d7cdee020d83371645a4d08e8e2e552cc53c233ba09218d98778629ef0c3a7b92aa425423472614c5a2d9cb2d500ccc2904f44a69230eda521cb1302b96b570d847ed4be163ccedd273e41e720c534656e769cd30e973cfa559ca391b6daecb58aadc04b4bbb;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1cbf570c3afb396076a1803a71388f600c8f7f6a0b29efc035ce0d6756d1f2669e7a6223e4cdef0aedece625f6e37ade6dbbb1c6dfbb73b7f1ac1d4c2326daebb10d76f6f3922ba509c1fae0ceb0cafc6c601c13ba9c56e411bea928d439a63d73f6a90846847169da;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h16e0ae9df531025de0058d4e001665f6aac2113d0dc63d952634a91828fecf21a228896fd5045af46867230e06855dc69a1c2a10372f665e8c577c26cc46bea548485cedc588c18f57507abbddd8fb674bcbcfa06e1e817f8d2b1e4f41f30ff7aa365915ee5ed46ecc2;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h5b4f90d296234419ea4af65a70517e5c402be6ea361486a36e402bef70397ddc18f0399ab409c7f24cd1d134b4153dec793cbced6d27dc0b6a7c31b15bfa39dd22b7bd259d514d55859dcc5975916e3af26123d6c51a56da5c76912d0c5f945c9c76e194ae8b5229f2;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h12148004a8f0ab641b6f69865ab9d6708dd1a9645de00e7b1e250825e5b1dbd46b8633180ca2c710817d3a3d356cfc66185d8dddf146c23e14962e942e872082de6ca5c9767ccddb000ef99a7912c5b09f05c266b3cf8416a5a86c844630a7e308db7e89afe9e093eac;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h19e5d523ed535deaa5a17fe540a4d329028b51fcf77f4b4f288f77e264b4fa2cbcd403985b0696365e19a6ec4d2a6484b715db29fe9b4c6f6a397f679a81083cbdb4c0c0efa37bd8a112269cb0c39d124f2f2e09ec7c8d1817d69dfe706bc148f10bbcc0a808454486c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h48092932246c539d14451b1f62f76284b6f7e0348abaae4737212bac627d4e08ecb5d8948686a0fe9e442d1ebad600fb2ae32d91eeda0bb110b1a88874cd5cdc32911287327cd5339c41c491a162c54172dd5e463885aee9fe9aa6501230df34c2cc55c792597183e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h4e48cf3f078723eb07604601f396919321bfebaf606ac8b30e20784ad403c3556cbc11c052f59c046228150554f0cd64d91d7f4d93f07b9141fa123b7057a0329b357962becc4824c0e6ae7eb0adc8127d43611f3aa8fd25738f368a8fe731dce0594ebe911a88f49b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10606caaf9df22c1e6cd558774b3d4fbc9a9e8a992a45652ecb169d5fbc7c5cc02b8a2c4c02dc31936b7a6ac4c88be63f52e226b00ead3f70d96b0f18a4df96a22dcad170903425d3553fe34239cc55c0e87c2410f01c4176c98704cd82b747c46c29ce9a06603df34d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h4dadbc7c1d98be83e664cded9986a8dae49f2449dbc618829b40b7800c5c20c551a080d9935f4d909d33fe55a3f1851c61359a4e8419af09a569992634a6419602b1223ec8e40ceb7f26824ea36dd81d45f76c4cde8d6d0f212c6c40e3226f31915b0d90260c91d6d6;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f3f07888fc14b3de8586d832a3b425faf5a27181b39a20d01d57398d6aadc40d1798a307cc07b38ec23f91d789261aeb3e2000dbc74f1312c25252cb34b4b38f856eb319dea65a269e4d1a28b88a3c6723123dfce3def4f10dc64bf890e8dddb9970790ebeafec1e09;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h64133fdcd9a506768671914bc533865c1f19b39cf5ee07145b23668557e9dd89c77dd30b7490de26e25e84764ffe9d4cb9fddccf5b6fff1846855a655ed01aa8b4f2493bd844e30f25a5b61d021d769fa18077a5b92af40783ed5a233152c38990f1a503b8b9db0e70;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ba20229989e0679147b1c76c5f882b24def26b469cb6daaa9800671c4fae59e80c992eeecca1c8355588fd89edeb58767ebaf4d8c4b82a829e8c72263974f0e431eef5b82ac59dbb2f89bca5d77d75d0882b8ebb44dd4d753d9d96596a2183483ffed62bd0cfc9576d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf841267e32be22147ead57a44d5dd382cd0bd81056e5f58a10dc2383b64bd4ea85eb458c82e61c74aa43d142cee91201b00aa2539b2ab941854d8bd9fa0348b58429e2f6dab7c683bfaa6ce67c0fccf621e6a8de847795cbb15235f78b0c630e3832e053e522b4d25f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1fe6c9f9d4a873607d0d976bb3fb139ceae46c084264f05a6c8cdbaadbf2d0ed2231fc236db2f58cb46fdb01004a820722bbbf7e678e16ec6da99b575b06a69c89734650526b2f83c29d8b60af063233f97ac249583eb289e01f362c17082bf076299698fdd6d106063;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h8cc5129ada58464710e9c06024d5638525c880aa1daaa2529e9ec76cdfb8d291f37ac56e007c3534c5e4209f9d5de8ceac7c22acca9fd681c559e33c299ee56e899d741bf1e5e9421009fc340e82eb3e3ab5acfea873f0929cf871ec6ac06f8f6974e67cc1e6f2ba3;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h103e84a96582fe53334094cffd0b7971f860c33d12cb7653aea81e6ff257322bdd46347951b085882400947023b91dcc337f67cb53bdd7e4f3b9b3ec0662bac7322d9c0aa2e2d432bbf3d66a61d2f952ad643017654b244a6ef6745151ae29301f38aff6d3900669249;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h181412a05e8c4982e9fa8cf49db54f900b988e717919fb39a6a7b4b036934bedea8e5b211218d0aaa2ef1187ca7d5c01136ecd7636d59c8751b8191bc37b35bfc9ff8d272e2f9ba0dec9806e8e197bf187db2461e50d697361de5c1de9789f882cee3c3cd6caed6c959;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h5c9bae8b51800b729ad786eb1dbf25c95606cc2a0b932aa4401d229689e9f236d27c4dad04b09857c1d90e5d553d041a25b488ec45bef5fdd1842931e1482a7b61dfc5d2a8135b9c3e404b4db24bc6832025cf352d877a65272ff485b6d4d6a4d5ff7457b937952;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h9a64e0648493e042010f6d0660c6d5541913ff5229f2a0ec8530d8be39dcf972dd200650d6ee539f720b4d9a7175e2f8e4edef94770f880e40a0ce018811d906382c83d768f164f199273a76c35c8951d152c562aa044b9c80317caeb725b21aa00129a3954769ffc5;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h111b5b8e1d914992935e89850c4ea4510874eb28044f0c1add2f75b965b7a4853023140597f678601d533dd87cf64ba57fcc7c7e4216171ea72cc9cb85970cab0b61543b054fc499f5875d952fea1287c2d062484dc312f7236c70bc07337aa85d23b43754d8f5bf700;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h37b31d68ea731aa6dcde720d1878f4877f11409097c6592f82fd69772155395cc125387007ef992a29fd5b1d69202f95f9a04ed911f84c60316e9a66a9a805ca517c2e98add4b0829b1c924ef47f8cdcc25509f182531212d46fa9b7f91a415502652b5115e3a2a987;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h8cde4bd640a95fd9b6d85744f3909d239cc9d1b9f7379af33045d73ef8b5c46cc62e4234cab2d41cbb5f041a99010c6ae0637366aa6eed57c99e8fb4e7fd9f4447e78274dadfb06bea140ef9f33458ead9c2803fdb0685a2bb495ba405d46dc077eb9135f60eabe5a7;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h196197d15e04d388ccc6c28cf9c23b6d940b0565ceeba124ea2ca6b6152b8a88df985facc88fbbee1e20ed6791456c2e6e11892a0ab02a90711b837d57c7e72f593d7452b417b54fa051cceb95cbb8d85ab28df0423d51f468f30fe509bd5840af1d5862e88f421ff3d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1095ea23481d8a501e2cc6f1ac6e6bb5d5cc7da29a9c30a542cd0d9e8aec8eb1e16b16491bd7e34366abec5c48040f8bfd7227224aaa94baa3891f1a8db49ef444a23d7fe8857a8f23464419e12c9b8cdf750f4f83e45213beba9b68f55e0af5c6ff749c894b37a0c09;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h163e1a92e1701441d049a0bd6730a9c4ebd656bf9d105e2c90f6b6bf6168d2e6da1aae7b9561d99d30059dbf2108cd1e62d24c5978f815de7caa4039e4fdeb399cdfb48806a73bf145f347c26882494fd998048aa1237c25342db9b4def113f2f06333c60f48e6e0e96;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d1b0494200bf635120b229dc72bf1dc342c1abc7646e3c4bc032e26b3c048bd20114bced8af1b1009913793cd228c48da712e5679fbf45ce8896c83014309de2c0b282b6fd2ce3731760c4ab3a6fa3fd174ad6a60e72b50de86302fc520da367e536b7abda337c8707;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h52e0a580eaf875399827109537e5828b10e2740c00ec29062d95c88ce7cc820911f6a974df6db70cf74471224a6940df0526ea2c38fc1acd2fc82233586a2dbd164474756a6c0698d3a9378b00646141efb64d3718379502c22395e2c19c13776754ce674ae9359660;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hacb21beb89ed72d47a51fb9c901f6a27bd57d64a4a0c48aec7069704cafba0993df4c358d2b7f4f0d43d4aeaa22db8efd1ec48bb326107ea63db61e67cb30af07d88f3cfd915a89145f605cbbdaf07bad3475f54dccf487aa03178a02350bb0b2e74327d04cec65cea;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hfbeb51dcb4bcffcbe103e510cf80a6090f875321d191801bfc9885eadd31220daa5909536404ef1fb8b72654b4c0f5c55e6c16ac930b57e46c9ea33516ad5d5c32bed67ae331d2a152febb3ab8b703d9d3935455fb729b4870639a604dc8f9294564f48b11c5726b79;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc99b9d1b4225ed1ae22ff84ff972a64bca1886d79f9b37c7d0872a475917929e7c365927ec2cd7fd74e0426a0f4e795c01b9aa01bd0948f3f8e67c98a9bd7b09c4f74af7c9e8ef3728d6c6a793e4625cb24df01db0b8a09a2f8665e1c7a735ec4f4fae1a2b9ab1efcb;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h18eaec2eb471f1c98ac6ef104a2a283ad893100662a92d80c199782af84a6a0ee4b4441d1d14aa19c899543df919a8ad1599d01c643c2bd60e4f1d51a5a6acf6fbcd01a190834a374564ae899f09a972484761453cfb4a45479153b6104942b25504b0b774f95e16b55;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d1690ed0be821e6deee6d387baba0cad34012762ce08645821f36a5aea9ad0e5173b202780376ec6695f966d5bece7978237f630946cb05b88567a387669a7e5c4d92cbbec8ebe7d9b1ce5b253ff006139771a29bc928c6ce0d18550981d6421981b20e48203b3d9db;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1dbbef96ce5d0e6a21e0310cbdfed42a243ade89312aabec17714658bcc27a8280de91befbd4247645d578593bfdbe350707eb7b681e9c20ac2126c25127dcf6c88ca5db1f272b48299695a998f700ff583efb2e3eb56076b27945059685bf7cef6c0f73206c94dc7a0;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he75cbeaf463c24c40a649a0bd1c904f21e5435775ddcb5e631343fbca5e85ee539160b04b5769a9842e978dfd0cb2c6d35a23afe7980f0c8bc7c314cc767bb2d44c5d059d32b10e6059927129cd193b96c3c2f880de0f0efadb27dc59fa7e958859eadce3b03c6e004;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hcec4bfe43208e80c7b3d000f1e61a480cce1eec705db52f9e6e742eaf1deb2ab48ffb36f56023503a92928eccaf05533560988461802e388f64bbaa588505316ea885277cabc849b128305b2fdb01e198cb310feda07744589f173705d6588019314bff06aaac5049d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h13d991a1013922f9e3885109da92b2ef25a6e3271866ceca923b69da662fd0e2c73d74c7b63f66a7c64b8524cdf22e9610cdb90f92d6e70f94982a7a8fa427cf094e342533d51b0e9303577cad2b1cb33c924f9c61c78f95c01a26030617055576f2f2f15533a9be9b1;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h9ee1f56e00e5759d545b9f361743db84a294610562e4e8ba147b45ceebd195ddee44804b0de8d63ea5189c5743a8fddb430600e1881783cf659232ec3352d7ff0c959dee25024574afea864e492d057abe7dd0a3313fe5e8345ae717bc5f8482ab6e22a2baf0f71e81;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h17b42ad5d805e0b707d806a021be1dca923afed595aa2900465400186c83c3746ccf42feb7dab42aa8c9d3c44b617f1256f2c60be8361013e7c269a782f0b137485d4b0309011c71ee26518a2b8e2c3a6ff6bd0ce138c91606212d6beb8494ce46095244654cbabb1d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h16a976d8d48249f00875424330d14aae8dcf6cf0104b252c09593d77ecf98b1bf8ec25260ab5542f389cf0eab11fb2c94d4f0ffe5442b294946ca649a499bf5115877a2bc67669ee1ae90efc204d4bf392c9939b86fb9303af935444388d2adc0bae598b4546aefbef8;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h152bfce0d446da205c26e0467fda542bde267b43cb7969e3756499da9bfe61e69a5a6053e9dab34641ce052bd79cc56a124fd251178ea97ca42bf582857d4a3b7fa04caa151d71a1dc69ef8c50bcb29dea7207d965213a09d0f98c4c60fafa754467ae44b2383655810;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1235d59b9b280b14f5f3f992813ec7ca68545dc427c830d6bd5bfcff15fe1cb6f8c96109c3ed27eee1746a35c54e24cbc5a4491e763145278bb7f012dbaaeeaea5b614742dd51feb450c5f41c3fbd439fe5329fc389db23a6b33ebd1da91d0b5b774b477b3b0b4f9320;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h17c093443e8fb9c6cfb615ac316b210c1cfd6dc5049e235f643fb2673088891d078ed86069086db0a723d26144cb13b3ca6a60d663f7b7867dd0b5d950a79a5d267f12321ce248a10100206f2c3f9ac44203504b1c65552abe26171d035d5fde444e83e23886a02eba3;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1942b2d8dbef1bf7006ead98db40195cea612bedd7429f3a29c87428dd1646943591034e43686a422760070f564abeab0b754a5e6f0393283ce734abcd1295e74b0d678e9efc81f3bfd0f41f08d2909d3c50f2c54a358083cf3b1ea7fb0a331d866c789b9bdcc3bd58c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ca0ccaa8608d3707366fff1c47beb58691dfc8d27d501ffcbb7bcf50c7e76d54827110c6e82d60063dd75769bf8b5158d48f245215d114890332f0100df5b7107ba3e138df727d8fe9a87fe3cfd1f9528e5938ab8253a44831248039d301be01653d64b94a645f3bc7;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e3ea5bf38ae4f8c69164d041969c5053c9387d2521b0c0ff1ed582dac67ecbda3e464da3635ce0b583d9e8eb37a06e8235274b5b54504934bb608d8cc7b2b297c49efbe05f71823fec294ea9f2fb2535db70a033effc330bd1e4467c3bed5e24561f003f1ba7721a68;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha38ce4b34b00e976db295cd2d0a566b6adb4ba89d3b693513f46b1899178b7ddd4b6be8e5dba6eb3ca82e3c678dd50a45b0c6ba60a19f5080bf6dc91d739dfdd7547bc4a5848ed47817549aa0975f6d70f9ba4b81981ee8f66a0b7d20e013209433c6be70ca6ef1b95;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc39540b0d26f2868275981c2427e4bc6dbb000d3b410b8f3cad20efc15130bd412b9a909be89ae45514cd53d3c1ad40b559ca2d381174893726fbec622fd1583c2ea208120470fe290f741c7854eb1d06d289b4d8024238356f59621773e45feb3b0ed26ae3b9bb01a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1963e2f80694aeb7138a83285b1fb15b5df7a5761a2e0ba932d0abd5ac16d52209b0d0a5ccc71c36930839834aa6c709d71a005da98e65d0d3731f7b59070a209c94a9b971ddb7b3ec769a7ada6c4283e22157833a97340176ffa4f2df906f06df62d188264d88a1b38;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h12bbe1052c993699b47e0915b2cb57260d0b0e5ef38178fa5cee2dfcded65419265f21db4cbb8d4d78e341911aead640572a0c16b79a87c82cd04e855af58ac42d263d9b6d92a9d140012117e1a7f8fa32c026c104bc42df48e25b6bc0e59991f02dcffd9dcf0b379a0;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a7a1e10f36ab56219ea81ef0e8815eb9e68f5614c6bec0b81eb415905232bf02b516f93a0e21db450ffafeda597c5e0f77d22a47ab419bc7561550c340c743d0761049f4a31ef6b38dc4248b45b34075eabbe4b405da164661ba92e6d1efa846c7bb4eccd3a77dbdcf;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h293b9609534ca2b9b719ea524b2bc4442d275c01c0b51cc1153b993996a21e3a280cdcc143baec1079d143b2a7f258fb34bb5f78132ab11dfa2f67f58c6b9ec43506001ac262fa0cf735f098194dbb26b600499c5772f57154078dac9685f3f166361039c2eba65cd9;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h7aaf452cf8cc7a4cdd978c45f9f4cfc254397ffd1a02f0885254231325ccfbce426541a832006bd7e37fcc8620d2ed46f432c025d1c48da18b4bf48aae3bda54a73c1e186d0da78f3c4e86df862fdad2f7efc2fd0987134320d5b3947f19ac38e4c8fe9b677f4193c4;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha137e922df53408a1edd54719d3c818147e1d0fa5f1b0077bfb160ff7c3d079c38a4981a60332dceba695ebef6a907625897a62e16786e317101907cf683ea75776888c3a7b7ebb6ad2969679891d42e5b4d57a36e8faee7999cad62c75927732e7cac1994282ef043;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f7cfbfd3683c23d8d827b57d4e7d91e6400ea5fae53906f099075247d252b826f931502450d2433cf52c9f43c76fbda97b6ac58f024b05dca74b63ad6e134f29591f08c8b24d788f87d717e880d8e3b7fc474ee9270b8b89c26c1469b1990cd0dd7e1d97f72e170f96;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h2fd1b7eab7bddda352073d9fba9e1ed4d171b0eed59941009eeba0be85420e32c2bcb6ade93e55120450a87b644848ad70136cfc4b2a3405747aead3a57acb8c5368a8214639dab1b872ba04f86d88775aeaf2713e888501560e01efe6b3b5e6a8be38af37b00cbab6;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1746fefea62fee86f1b02e204e03b1c80940ae1439b49b33fae317c6d19ad182306c7d83d33f655a402218b04503483caf23948a6e9602de079f8eb084ed5939e8719138d1c43eac22f64643e9cea71a831c24161e29353cd1a502ad295305c18301972f61919475101;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h197318986e790cd68fcb24f33a6033b66f35a0e90649366c133e298468b6c6089e2637052114051f0a7f8aa50fe773874c6168147c2384ddef46f90981a8abe2dd068e6c70394a7c5800b816c5e2dceb4a33c78b62487e3456717df713482e47f8fc14f5981810cd273;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h9e42dc3061126aaa0c8057ee108c6b1dc98a120a0c4aa7d1a0212204345f55b54635361a5011eec7f6fe7d2a811602e5f18bbdca0ccbc38ffc9b18550993aaaf5e7459feea7203960e2af8df1cd33535840bb47f9aa7a2e21e90192ac6c003d7a301fc6e7984a6e271;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e188bdf0ce11df1b54e7e4793e53c2b62b5bac6554f867b8c9efc67c0f2bacfd1cbc718044772b7e0f088b62941ab4707098f9a24bf9b8c29f093221abedc98a3546675e73ca2e9ce274711ac73e461132861c0d1a594c8dcc1098b3ab21917fedd5dfed2e35911e93;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e8628210a51933fab38956dd3567441ae47109d75f0d51c42ba184b4f3808a384e66b49026af4000d4cf4527132c3c7fc0092493d8198ba497cbceebbe7d24c0b5e9554a70aabce0d307f48a268af94213b9505713d057e5dc15715fbc91ad07e147963fdcd50be67b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1988911c6b18411c8cbe23257c4b70e24f5a1c67bb7b8b17f68cc3198967d008fa885c6e71431451771229cbeeb2ddd61ddde7662d5add89effa7fcf8d8ed523dd8d8a2e4fbd69cabb87a348e4428beb62efa458721b792712152b4c1c8ca2b6bfcd3cddb9aeb2e5d84;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1775b5a07239b385ca2b699116ae6f9666ebaa6de7909519c3bbeb9a54f49ccf7cc5f0bb0df3ccb98d99ec23da23aeeb5db2add1757a19e705dd3aedc2da834a6c2792b2140cbdf6f319c4ed25f631f1e89352605e6bff7e92675cd2dc3d932e7bafd6f9bcacf1a6675;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1cacc0a6806fefa8313d9490157660a5f36a6f4261435ee5f2b4f5eb3418d460504a5cb4d9076209c7c89cecb8e5b172174825613bde895413bdea275a33d15f2e3024bb02a8c34e70c3c66330f221b4f50b6875256602394e3bf9e8feda78861c60cef4b228afae26e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hffdb574f1bcf45986a9e58dbca63a659f8af44d886920a96e42499df1a4619897eef0e089b794827aefb39ef7d1f419d804785525e591647e384e6bebdcbf31bda145df64a0fcb11c1b82bdef3d3dcd5dff659b27b32ed201d76d81bfae913558f9e8c6fdce971fdbc;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1455992c791bb8d8e5e3ba92633c571023079a3fef68f23b774827e0c2bda18cf1f67c4a329aa97905b2b6f341521b29b583b8fe1686b8f9583bfcf3a60a41928a0802a3555eff705225656a499090a459335b21475321a5be7164791fa45fec28cb02984fb6d352bf6;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h4b204401e013b179d76f683b0fcaab910055db6e73acbded874a7c5a5b946bb86db9f2b442e37a1972174e905834a316622dcbbd96e5adbef64537aa0f6a32a553c341c85d5bbd09d9cb892d98e3938c527345cb8075e40e5f5ed4fe6f5a599ca6cc59a88e770a174a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10273dae26afc2f5aa11a85c9f63799c89af48f5097fa7cbae03b8fb57a5aec3e62a5e9613e1f91d73bc666ca20791b93683a4183f62b31b1a3fd32a37e8b7d6eccb341db9e620d4e8e713d354c7ea8db8379c10e008ef64f13b7fa63860c4ad48053649dfdd429ef47;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1285050a3d61f0bb2d21013bae02e90ae7957fae651415f7cf6d5cc28841614ca682ebf04e4dd74c3ba9210c65d8566ba2ba6b97a216506526123cfca031d2145dd3c2f382abb527060c9a6503895b8b33f5d3e725af1243ae45fd493999fca44b8c7a0f26607789161;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hfea545b741284d6741dc2c59899410cab23fdb641c89b18b1882e9a5160889a5ad8ac1af20bf8503671b386049bc811eb2473ab8e35aac3592176fb1b5c90e7803bc4ca21c118aaad3b33d768772135b6bb85972822afdefa508878018469022ddc0810440ca84adb4;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hbbcb15f0ef92efdb8bf4fae25ea782c31c54613fd9a3d4d3d921631ecdd1b1780a49463c21192de24f5ee9a2cd31f47df172b7f73b323028b6f28b50f6b66d125c0f8f0876887058b64fd6f5674142bbf5209669a6534529fd55a2508934ce447f22bf17e6632d5fd6;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1903451146a0c55142ac13f870251290c0d6b830dcb2615b589e91760d962b906eb1682f21c5fa489e996be638205273e38761a8877ce7f2b7733f25b77f7730001d5059d1b15d10c08ecace9032b0f6db7aa0819eee6b939e1d014eb81596a14d9cfb75e79d6f4b24e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1704a229c49ca301b18eb8a409f15a8b82b1e2aebc74102738df01576ecd485e021e4e952fe2b69ae43e98681cfed8f26e47f39bcca121825346388ad530b13739f2316bbcfd3ec2501c7f63a2240ede255fa5ba8f14764a0bf24c75ea61634e509d8bf36e795e5ad36;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he5b45503d2112708ad31ee0e0af0e7066d40654dbc9182144e10bea70837ef1b78e473f1bea9a3d54325a6faa10586c714b4d7aa4f738e1582ac0e43f28c068b9508456420b3fb060994d9638c787c7d8bd08973dd080429b449e99d172d4123bed59e1cc40edf1fc7;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'haad8b4f325f7f0b9577d59ada13afdf4f96c0dbe6c0d042c5e2a536dbc3ff0101000d858436e2454122de8459b5eb38f94af83da7cf0e6c22d4ab6d13bf034fea55adebe5571f777de4a2d88ab23213b32b46c9576f12752a8382c1a0ae34771b4ed13b51928385ee7;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h63250450ceda3f19fcc77202d6fd4a9fd1df79892c74fb7e70e79eff581b90a259f5bbb707b53fc9aab7d1eb514a41deeba0abd2934475496f4255e83a7bf2f7d39a6a8cca872a019698039a17418f4384394239989ff1ad870813f13bd63b0e390877a9764af1ab95;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h175aaa99469fc83b48c6f0cbd4c0c3fa7e93cd196d8f4e90f54e03b758c16bc62a5848d5e0dca2fb11a527071c112cf7ab91dc532323d05fbcd1abc34bcdfc2c2e431a78bbef83a4a8e13efbbb4a4f6ea7b4acbb942be2d9149630791519605e4a4effec12a1290baa;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hcf04541127c6778bcdb0f93de15b5b51bc4cb34df08556be6a21582516a91f904039e6c9e5b469253db879f57d3f8d885d86d63d333ba4892bca2d04ba448106160d0aac4e75a257ffd49be9081ac70d2a59ea8d391b2b04991135260d03498be27987d727d8a3760b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1990fa7c55c50967cd41dc0e026150864a36750a1de196ce753c1a332b63f02dde52a9f374ac16604e76ffc7b17ee744f1921acf2a119d00b663397386fabeac23480c2d977eed25e63a738b2e5e3846b59b62332936742746ad7c0e15a76d9df6093b8e7e4333447d2;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f09ea456a68cc1d6bad6174f0fd077f3c413db23a93dec5b18390cab1a38246be56358482807191864d7934398e2a3f7228c985d3b065ff93e21bfa731b9a279b032f67939c23807055ac65b8512d42903de92dc538507234d4512f5e5932dfabb795253b4a48c675f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e48cf37797db2bb45a27ecf0ead6d10b13414c35509606bd336f679380ba6b0604e62958e6cb5fa01d1ab2593d514fd7d01bc9a8fa923cce7ab0573e099ece4a40e8805504b8e206aff3edd2342cb0e58914c0cc9da0a210621fd91fe06e4057ad0f279b6131599940;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h93f439dac6d43b04b0edf2414d8bafa45ab8995a7d8f7d5572378d94c55fccd7a4abd5a5e077a364fa65aa8a78bee3c3419660e4d25c6c6a1804810207cef27c26d94c7de38c7f70495946e7f8e5d9da26b1543fec1b79d754d4343c17849b921d4f6e91d27351c77;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h131f3ce8872c854ddc13dd5425068b34287399dbfa2efd44b5bf62cc549bb831fd19eceff5e731e161e64a80183f53362a0b33126b394c3b46ba6deed564b27d6b00105961b5c68d44700dd8fe965fc0d955dae5ad37000a116d3653a55529af3e38661d73c5b434089;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h17cd35ecbffcf84b0ba8edc88adaf569e1710df236e454b6cdfd76a8e94efbb0cfc0c87646d03fc671fb08d3bf557e32235d95350c0af30758e902b0ec3bddaf2884b9ec576b9d77def5c4ba1a3adcb717bb459c8d8236f3d90dd82e06b953f7cf6f211cb989b2794d4;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hbda5f6e35f0181ee66c70bdf8270bea2b541795891767974f27455a3678fab07aa61ce7662aa3b33e66426a0f3dba95d4bab1cb0cd022b591bda57fe693683ae9246be11efb3d0c74f1cd3290f56efda97409d24ec4d994f8a847ebfd021641e8153b225852515ad3f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h14d68a461d275fce1cc7dc0fea6c299c5ce32ed0767b70ac3082eafefe7af632a9e5e510bcbba1ca30514d313cfcd24cd3590a3c582f6894f23d03728c91aff35612d7e9647f2930d2e2df7b4f33aa920fbf4f5e77b9fe897c13783332f64580d31e9f014d984390b8a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h6bbfd9c60bcd7cf684c2a2ca4c0058cc1b6ceeaa8b862d43f9cc1806646923a133ab8d91cfda134b61fcc6c768715f2dfbab1445efc75338267999349de90bd782a860090c528892c11711c8935a457d9e6d43444ae61361ab25c41d6673c1b4ba019e3e4f12b40dca;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h15cb5685edf5e6adb0ddd27e4576337aea450c8f5919224974995d239681570389b88a8549b23ed567a27e0cad49ab69032e03bee86587ab6b643dcb39017df7db5f9ace0c697868aa8f2f8e4c734b484c37044dccaab6c3c82ed29f606f9c5400166ea03b2dead498f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf6da5a1ca712f4fa9974c4d8cc9c9ec05e79dd5ef16e0afc3db51a129c69277169335901c20c2d5a2bb8bff55f2e9fa2595b194c6d56535cb5a2bd691cabd7c7a31f64207033efb9e1dd8ec17ec7036c1f47a9efa43ac001ffcb52573ccb8d11710106bcbdac125ba6;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h5d43fdb3ea13449f655d585f483606759307d000ab3bc1f7eefa15684696b856efea0a85f61c1650dc237a38572121b35f6b0de6dc652c65bd01348a659137692fd4ea98aee0e62248c62f77718f499bbf5a908c337c28f20fc4115932fb36925dd183f331cd685e1;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h800f0059e7db4644ea584a646f6a4e0a8d0ea83ecf5157038616c11084ffc626707fbfe5a77c16505df35360c8bc52276bf8694a93dcc342b3a74cbc010fbc27d9bf7ff295dee33618fe2aff9d08eee5c3fe9d616205ffcaa8932377ee853b4ade906e0c513d78e5ad;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb1183d7e923f2276aac3ba8527109d6de2b4c56b6305bdf4b45965ecb183a1eae614ca0e0a28c856a846a863fdbf8de242d5f6c8f97909276724b70a092043c41e5ce047f2c91025ccd8e1e21c8d5f145e2c3ce586367bf5071ec854f8d2b211083d682a8f278cc87c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h2611df682e2afbe1792e8ea23da648617a19edc4f3c1b55891621f4c54c56532c2c454609033d59f290b4092326d607fbf989d34a38968769cdbdb6de125c0b5bc97a664424d7e436900c538bede9c50d855cc2fe5c53df0810c8eb740dae1b2eff31409b1ae7093f4;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h63155c66554bb607c59a493e789ce3e08cf897611921bd6d9e8038a11e51514cf4a8c33e4944164f1200c5dd74dd784859d821cee20896a6ea91a0349c785bdb3f3901fbf400bc2e8302f9133e515ac67e0fec15e61355d62cfa340fbc25bf5195954659d1a6d905d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he9c75496830d97cb8ea38c82e99238e193efa01a00361d02940d5cdea56fafde6257c7cc13ad407b4a91337cb378c7bf0e3c53b27ad4f9257896c28e4bcd284c6a173c5fba84b267849719751a728a1ce63cf77a6971e490b1c1683b26b61a81a67feb58548cdf2996;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h16f3e241d6db25d29c27104e060cccfb736b0e844ed76bde1740e177713249c0d55d20f02266caf93181030772464bef664b15be8bfd7ce168cf196093b739eb67297b944d04846583e2d3859d49064b8fc497fda6cb349a25bfba44637b8ab93794e06e5c00357ae6a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'haff35a81d5bcc7bb8b8f3ad1a9b20f60a3eba7aada44b3559414c77ebeae2acc47ab2911d49b979f6227fa28c91418b8768c2399627638b5db637b9be50ecd4fe0888717a32e4e4daa08428badd072e382f51165d294293762c9a87948a9e218740915dc4372eedcaa;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf13658d73e2b682b789ebf7d87e543d1e76ec14e14fbeebca53d0dad8e39bb889a69dc3b090af5e43c219868ecf20a61c5988553bf4ed1354c3203b6824b38a53bc8a0d15b8f188b8c880053eded47d53c8d6f0b7e8e2310c9349ffe499e2822c2cd8d0248530c3358;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc64585cdcd2185df8405f2dfb5baa1d20afb1dfeee85f9aebd3fcafadcec37a4d954f309179efbd6d884774fcee89d8385f69a486f25ddea94e1d7d6625d07d2f7a51ae5297f401e98aad9fef1452b8337edca730795ee03eabe9fad0fc7ba8a3b4580ff1be530cb15;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h182f5756a2a7922b53d0e2d6810ba66976d0987cb55282366e6a10fb74c0c82afd434a51ec325f8d5589e543c5496a7d2fb04730c07968ec9da7a3b292ac9c3b10fb0153a0c35eeda8f739c238b7c7ae1ad3f39173b9d3bedf9abb365b9114f00e0ca4dd631ead551bb;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h852004d3146b9bb79eda3b73c821c5713659c351aad1c1bb20a1def0703a4770ec05bf905267ca022f1c24b420151e6d37bdf9d5842b92dd18dfad2a2891c7002a92a90121bc668f1bfb3123123e05bab21aa18e3f0e91f42b95f8b6849d0ee11cdd83d051ce6ab9ad;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hcef46a994e2e2f14515e2722684b85feffc8c6ae3702d35eabc9521a5af845488ccd9871d6b7c5efd228eacbee361cbffb44b2026e90698fdbedce3b5efd87b16436eaac8408f1d406a9ad53465f4e7f7538341010b26efd17d3d09af73c3296c463a5dbdabf7d4d50;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c1846c8a220dc355960c2514ae65dc8190f7d2d55001dec034c83439fd9b1d46a6d13e358f5b612f3d63063c140f6456372896eb825d0167e113fd2b83a1f42dcd77bb29d3b361e53df5fb7c7975f25db6ec1735269b9fed51bc8e308c08a6bad39f46996800fbe450;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h7dac6cda539331676fa47ae2be769e5b0cd15688aee173940c43788f8c89c4fc9c23191b7498f9509445213c04d53abe74cabf1f9482b0bd26965eb153c586a8b6f89706131dc6aebc17d35677b9a55d255997e4b9be4fc81337307b47a1f0aceac4ee5865e5b05cc0;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h114507d474a70eeb3478a5240b4fd07ef497574b386d58cd1d5d7ebf7382042ed8e1f5df15b4d5af25c848f776e0ca3981975984aaa369c40f77e35630961cae6953ca55e869a81296493874527faef7522f8c821629dcb852cae19ea355dcd541fbe53945c56ef5ef1;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h83c66b44a376e6518ad92497b679575e1eea93240013bba3ff7d73a96557411eb97dbe23d8970ce2cc95d1f35b3f976371fce56fb74d70a4cf40d610674fe087357aad1a2bed946b1a8bd19bfbeb13f6587ac542043a4ac3584094b650497ccac1f8b96221bdf8b9ef;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h18b4de32d5af16b6b9012e3010fc09cb6929b02b1bed198e09e0ef2cf6ba92aa7546b78306822391dbaaba0b2e3f4e44a6d299a5a875f8d3ae5bbf7deb8d7dc3a3c7c99e6de24d34718bbae41b3126e592f7a235a5437f491721d268bf39e672b7aeae87a9e137bc45b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h13e1bbcb0ed59cfddf7342ec13852161ec8ba7db2492fa3e6569803c85716afda636670da34c055c2beedfd85be7dd69e3e04c0a691eb36e6650d38dfe4f0ea64de2c2806534f14bdc7fc1bbbde2bc7d20156dbcbc67bece69f4cd4d005d1fad2fa729b94ff1a73702f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h153bd3bbd8d566276af9ba9caad659dc81490b82a68c194b73a941a6f9290cf12168148c02998361b362e6d3a93bdc3cb7524ff145acd6bcbbc6549009f5c6f336b35b26dce77098a996acc793086eb6f4c433cf747192cfeae9ca023efb14a23602b7d2c1ea10eeeb3;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb52af26e9ca6f3b816dbb2e4f0b6529681e0a6f260d57dbcdd3f3513a27258e8df36a123562720b5120140aa4d7b015ec8c3f705538f6ed4cfa3cdc72a1e166cee0269be7ebc98e945e2af2ffeaf52ec3f9b4628cfe896cafc019ef187769bec5a25de58391a27e138;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h158229700b83de1bc1edcbe05da338b5e55ec2d5761d78e9bc31a102c65c07fcb8a6f3e73f1d3e809ec298db92856d3b6195fa23b6c88191dc86d08c3a62ed1e5b2a61bee0a9b73ec3d0ee32fa790ab170e295e826c0bcd327ca771563e298fa64c6149ce51a14f32be;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hac5e55c77ee2382905e4426d20275ff50fb417bd007e568551fd5563661b19bfa4ee475b94e876053ebfff520f99b09f50382b19f6045d84b73bf47b9f9ccbcf21df7cf90d577a2194d054bbb78f47b7f7ca5c2bf462890bff096c8723e350997ebfd6e1ba38d5fa63;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h137dd76e046f11678a62635f48ecbafd1a544930342f52a2eaa3db2337c48b27e2d1acfafd7576eccce844ef60ad5e69a3649fcbbd42d4c06492afa8112bb95dba5a68ccf05b1522cac0a251aaedf32767de7bfa77eaa3b541f00c652cfa54e7ed20bf1bdce0861c44e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hdb9220553713f562c141dbd900fc237dd02df7d30a45365349b645b78c235b231f2fc3385d128934db6148f04ba28b4d0fb30b8eaddaca57d3242ae0f2de2eecde3b1ab15ac033f5c78bc9670a57028eb9156c21d5da4416607465c8842a74911d2fc7404678e909aa;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc2022487601e91df9342f253a1bbfa79eddfa577a835c5a18703c6ee2c1b6c4d5735a363ecd3f113ee85b526e63b983b7894bcae9b7c55756981ca4492368f876d253d1b2efdbe5126113dbf568509267928ff513fe6776bb5d94b0cd2777f65dfda00bcdebb156096;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h59246bb4508a2f2fffd991ca7a46b41f874fda5a99d7c9ce7ce54e7d6cce326eef6ed217af99b253b9860a45c6639293f601703a0110fdae3b5c54823c25353bbd910307b29cb1e65b486c6af29b7c10457d5921c3c218614366644ca8786d8770ee0a35eb0c5b34ff;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d7cf3f312fb1e20f607f79b2a0fbdbb18fe3c63c5fa6d57fec5b5d93d744d743f81ed8f13a6b0318e4f31249ad5c59eed8f3f293d354b1ab549597c324f0cb36e0365e42db12907b041dc56495cd17237783cf3fb715d6cb546b35a688be0edebb1a97958026df78d7;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h79a29d45fbf551c14c77b998efa1f5f330e7b1b554c09d8bb89cea826b02bedd3af91478de5c6cdafd91a963e8627efa715bbf8bd0be3ffe6580b6846cfe8533e4c8e304e3cc2da188512b2b206faf80bcc0986b837e5b24174d484f5a6dd6b317880642b96eb2704c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf8b9b0f90d7b0efa133ebadf449ce24dd1d9e0e45336ffb07c3f79ad712435c6c4efb42ab432d192ab37ed45109011fb291273b9e396e13bcf8298af275bf4a8b35de59a2bacb0f0c09b79c815311fc54a61b80ed13ceae8feb89075a31ea2ef66045fa41cd0f901be;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b5882c2ba72e371e3b08571b859f9e8b25605346281c13af88e4eb53e12b8df1802fcf3d88b0017b8c56c2ce7e105cf4641a4af5bc1ce3882deebaf67e0cff27918be60686e44014a98f454cbf5ddf68ae67c91ea606deb99f0780275804f7c504774c7e741711a954;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h4f10a8b73d136a9f9379478e8baa8157be6f25d3f0948bf58ad6a843de9b2861f23be3d1ea41dc3f56072901329b2cdcda7ed0a859c7de62e998dd25bb8325bef3fd65a1367fdd17b23b4201f639716544f2138d3a61b5b1a1d0bd807ce7680669a1cfd2cea681cbe4;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h49bcc10a3dae8af7ad47bf03ef749e5a40b12720461b15824ccbe5ec8736e6408e3e06991b56d09d532c20123282a16c1ab35959120f2a3803401cb67f9bb8ac1fffb6994517ef69518a78496d8fc11cf2f5f72a70cdbe2e2ff754eebca543f1ac97a9cc6b2bbd534a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h52875b93e0a7a52627f1054d774e3e3b18d352af421e9cf4c239f79f4d8b7b20b511f784dc92084f331e818e96e05abc57e5a54f47896f65bec493da926fdc2ed02c0464fe7b72b896dd59cfb1522b229fa69679ba0cac31a18430f2fa2314a81996c3c75da3122cb;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10b6fa6efa0c37267690138f4a7f3487b5b284af6c59146b8a4f297fdca5dfe231ad3fe370a19b64ce634bc824573f7d422f978af15e95faf73d90acd5dcfeddd0599dbc6f5038402d2a2ec8066208bb945ad2d584edccf4da7b256af4cf70abe7d3a5a32b9cc84e44b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h3aa112f62fb8e2cf076dff463540a312107168180fdd73f99f2c6f60bf077304acda3b57ea50f33eb15e34cacca88fdf533c32867b92400523471358b629b98ca0bccbdc86c2e233d42dbcb3c77b589bb3205e9ddec6eba163087ceb6acc05f280acbeaeaa66d5ef77;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hee6c1c282b227d7e82cb15b9b041c6b17ec38bf9c66c5a830ad09274cb22d5ec54102c5cfb5df15be76d2bfcdf6878da7a05c49beff8bb7ff4dfdb6e4efaf85c7d26becde4fbddbfcc5181af55acb93020b669faa697d8d226c486da972b4bf319c735996e8471c632;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h8230dcca9882e5b836711e68ff0b69c5717648530b53dd06435e0497acf0e845988daeebfa5cef7957ef0f4bf8090f83b2af9e6856d771da60270ee002e095aa94ac6de865937536c9685ff36a70cb0b8d101f2f4a963c54753c99b91fd1d5f78729f83d9a40f233ac;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c1f65459c5a9fe3db5a956e9f8e26f9fae2eed5ac080b6a802c611b4730cc5d09459f272a8d78c77732801bfd9375dfb89e811fc288f3d73d286194c58164a86cfb5d819e53d16179a2d57a92f6337609023155d6106664ae4667ba6624da78ff857044aa5aa46302b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h5dcdbbc6e7b87b1bffa9a1151373169abf2f3abc38c8b9512253307db9f8b724eb4dd4a972890bced9ef551b2bbab1b53515d0d5740219f1ed48a771421a28904d2a6867711255ae203d80ac7df8109a6b9f9d95199d340f6c31b492024568b9aa4455571b0b8b228e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc20778cf30b6aaa95e13e548618edb3a2610a4c53183fbeec6fcd695a2c187375855711fdb07b887e8070e5b71fbcde136decadf76adb5dc001802c3f413b5a330e8e94819330552a35b0a6fba8d02521a0880d9eb259f757a52cb6430e2793270e561442170bde1d7;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h144186a16e64dc140bfa22357fd09560bcc2a9dfdab61ed69a7c3f398f1e41b52cd552836b8bdfd8a21fad1b57f60cf13157bf9a30c092688a6e89ac441ec785be7491ad2fb67b5f5f208c9f242cda40ad9758f0eda56c77db1bcad16223b0fd80f956c3177d5142e94;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha2f503b1510249de90a11af84b7d28dae79999aab619d9777ad4f6a14c0fcfa96ed23146eeb103f54320865a6f096329bfe74fb01cbec6e7796b95a9b6ddd730166ad090c9049c244d59a24d14b4ba336ebb1b859dbf4c6caeaf0ccc48f0048f32c8bd16ee9ab533cd;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f9268511bef37c2304ccc3fbc6d23be84e40c721d10af5db8f0870e0a4cfba28866c2ec5daaa780df01c9ba7579d7d87b2b92d4823bd712bc36f861d530739fac140f70fe6c7393e2330b5318f5d9172e7cb30376a1e094cfdc15616e9e95a82c582be778b22ac5994;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1823ecd3914e2e4e3aabb900615ba0025a14afbd3eaaebe6e63a48e62c1c977dda2a699d9383cc558710e848effbffc6175e1dcfc535be2b90380321422ee81bef5e389183bebfb55a6629b57dd96166801f0cf173e812c202f009607e8d519c037116376b82e70efd8;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b392765f0820d92dfe880d0928b0ff96aa99c8aa6635f4067aace78827cf790b5b06190665b9cd27842149591e5ac47c60de8ed80240248b6e5af4bcf8b5ce923e26aa8131cc625f8cc5464065a7f5686899be8bfb0ac5ca1b28dde4bb26ea9a02cb64f348272d3a09;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b207edcc92f55968472392d152f4e1f5fc6c6f07ed844dad7c281319507c45476a0a0a41eb432d053bfda8cd98c5bfcd50a7c351fe2da13887c0828dd6ce77215500c4a8dbad8a915fecd9baabe4f1b356303915643555814d8d60c4b05b7aa5515e47993c0571aa83;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h27cb6c411bcfc29772791551846cc6996bbd4d2d2b053f4b8e2a8d90c368d582e5d32fbbb490c0ce745e518273a194f9b006397ae034067982c7839da8da6f8df9329e6f50eaf0c8b9280924afc8a2cf6c9706f14dd8919c021f412e4b522d453f49dd38846c518175;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h5c21f779900c688c1e2b317725a5d0a5a3f803287685def41d13b1b248a53c50bc52262f753863634281860b540681df061dfff0ad4c377d5606ae51b79158bced3b3ddb525145c82e69aed546a0ca6d4181524b154c8f800d0115b0ea940f89ecc419ea05f58d974d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd266f0fbe644a60e9f0ad9930f17e7eaf49643fb506ac019bf0dc93345bcf1e4df2ea4db8fe41122fb2506189aed7ecdd111a43722c2795da7ade4c31e284092b6690593a4f5bec88ab98cfe8334f0702b6dd9c00ded917c2de9381dd19b08388ca1de3c8d3e0aa52f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h14833e31fce21af5690f49e3d9a8d3cdf0459f37f06c4c9f33ca16f66db674261b25a002df52655080d652a5732e21a2220f1fde2f1c080e3ea2abc19efc63704ff9850fcfb936fa433f16646133755b2be7fa2e8dda1847343a1f0ac45caa11d0972d1e51d6bd4221f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc6fb954c6f0d62a661e77b4cd71983b7810dad2b6ab20fc2d66f1338927c2211b4c9d9eda52ea931c4f31a14957ed673b206d9fea92c885329a4792d59affd69f668afe2622ec85816f21ddd98aa0beac07a138a8d9a253de74b44619d1a054cae4f071ca46dd19003;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h2da1b8745f6dcda5974b8c9e366a2728de5992f9bf78b43ccf247374d2b81396beb37a0f27633a05210eb8bb81199d243064f3526fc4fbd4e64d6f838e3f4b9287dee33d057de417566b246a31c944a862089c6308248131b8a01edcfa615c665fab4936cd6bb1629d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1794caaf380a8ca18e1b69b91bdd7661f8e2d4ad15aaa4390b066c2a392ac1f20dc7e2780a5fce53ec33b5ffa6a15d926076af99c9e3d29b5da15a7c3fdf34c4b3bb160dd9573ddba836aed87bdb1c82b6fbd9f7173bbd2c251b0b08f066f390f36d04f3dce4d093d59;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h12a9b0f0d3cefbe6574b12621932e8d656b92ede16cfc691cc05720e8abf661c3912642b2e1dfd23e0366d9e0a4200724a356d8186fc23c46d69ee2093977efe49d422d17b776ba145cd238be05e51c54e8a883f7ea5c6a5dae4e2b6f4326715ebc2e682db307bb5392;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1512adc6f3c498830e16381d6d4d2a93f0529cb70b468c619164f0c14ff679853b7284b0a2f7750c3443aa978ab7cd2ddb23f96a0033d8ce0a9d740e2bf1ca6be8a8b9cad8d81830d3e8c13e3ad3ce8f69873c4ed4bce1cbbc4b8d543f8a44e3ab37cdb559127f3dac1;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h133f36f5b1e887feef2fb0a115e2a6dbe75d2b1a2d2867b29e44c6a5fab45b185ead6ddb16a399b20ce0454973087d701b82d7383f005cb8a42040a09454ed1fdf40d2d3a9e601747d710eeef3d0437b936e863c21444a3efee099ba889ada705ec165e86693f8746d6;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd63f6f056a4661c2308c660f0dea31a7d0acb6d8ea677af79deb443d301c961426ed8d1da1d918b7712cede0a5deb695d09162c2e837fe9058e90d65a1b98187a008d734ff02e091a4466174314285925752040651f773db7ec5d89278136d81e667b11bf322c8ce;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h5a2106a39ea4df4e7eb0f042544bb933ac3428900a3aef722bf10c148575bc738aa155726ca20866ea8dae6adc722683a0c2dd85b9d75c7ece1f7de64335bafdccfce622483a9395541077def448665f77995bdfb14c19721a5f240c2cbdda0c09d6f9c580170ee2a2;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h5f60f234a834a492c6c6fd4c447a2310d78da2e0d4867ebc80703d742b4b2ce708fcf2ed3c62fd312ef012478f07bb4841f67de979a7b448b215b0b7cf8ef20b4d2a4cc9b328b882ac3addb6a8b8650389b3ada5b54c12c7240ed4b6b15e1addf8f4b81e828b09de43;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h3eb7efdc806639e5c38f485aa301c0306337f0934407e33be21b274b69b6f40f3950b49555b1cf1b1af7273ae3c908dc62358c33cd3439073498785aad4c402fe059764cf29109b1d4d4e8e0c16fbd8a53741d666c62f5f850863c765828aa3e03a55eb0fe9b83abcd;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h192a9ac50f74464531bd9b7e0114439e68a695d981045c20118354a235457acdfc04d89d92e70d606e35b952ee731cb8ab53c99ce8920a2ea3f0f56ddf1c0a5bfec29b2c6795904363f0629ff3a85d997e995ee2d15bae6dfebf9f5388fdffe8259a68b2d12ed85d10e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h169590e2dfaa42e416d76701437bf27e87d85d8deb7c7f5811d818a13490c4f768e084ac8945367189652e816fc3fa043ccf88cf47e2188c18d08a95b9eff9ce5ad8aa4b7944ac41059f644959bdc777e076734d01832579ec05136a313fc0d65f9682b0bb913deefa;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd312478e31a80874c4cbf88ae4f1a7c60d26eaa81e10e768bb1f7a4fa1bfb0e1f04621d447fc39bce3809f3d7cd91fca73cf572d29097999800dcdfa6410e2b07b4d29b6d3f3b078f6f5cd4280def4493f09a914992beb0b3e8cfe07266350953a1682b30398388de3;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h2f79e1d6cc2f275b4eae807ffcff69d168b274dbf47e3adc0deeffc9b6de47141a8a292b8e47c4e22fb8d6f54cfffd0425c21bd54fbdabb81c3053579cdb464a515cdd9db09ccb32ed5e53d5c693f0c32921c0e3c151c1a0e5ae6801930968d8635d1b8a257e87c901;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a85ac484861121ffa31b73a5f844f7c56f8d3081e7ca9d0b677484e62ba169167f9efa84a57badc3dfdf3b4d5ceebbec6741846abe522e228c837db30945326457295e7d78fe0936ed8b6f8b64d3e5b67c1168e8f50e8a49151899d1f53e1b6429b9a57446d3a506e4;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h43728b573b845842a724d48191223d98c65dc1849f1b0ae2276dd603cd61be1d9edea9864d7f3deb3f1a029e3a776a060fcfed8c280dbf878e36c52497e55279b100ce43651558b64103338facfae09920921b5d13cc1330038c3267d88854e98aaebd765b7a372d2;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1345249da9dc8733b1b7007c59b9801528bc1729069c9d44b42e08b3bd3cd62a1a5466a6b5c0e8bbec758e651450099921b4801d8acd90ce0acc00b065874dc43816cb9eeb16d953fa9eb7893e1464b99045e6d8cc9d1fd472230c2f398bd7e56b9b59932f4f50c25cd;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h16aa87b5f0bbbf908797a21cbc2718448d9528a01127f5a68f478ee6e3085c51f39059dec469864b66537e8e0c7d9ef2c5a8184d2dac4f8c4d31ead2b4f20053acc1583046bdb8a1b4de71ff6a57b5eaeaefbf901bd24827155b922b0160df34a32f2aa9e01f8c6a0aa;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd231132699b89f09cf29b06f15b8511d4f9fa48265ad345d0a89d3742c863d73c8207ce3178d02a6d2e96ffeff1afd7e8210f8db05b52a8f957599bfe484ab9e4e73dc8b29542ec00334bb3ecd4ef74506ec0a7c629a6cd23d21b5b6b523dbceda46c514ad514d3317;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b54d19a6a22608461cc32a4487672eb2ff49d17ca948aacfa5ab18d5a08663aa85edf4c2d3c516baed0a975a551b508ca5234314e77465b5742221615681fb13f85c432a8136aa549fdef387da6ac8c01c6029bc713b3735ef5650bcf488b8ff167120c8b89ee26624;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h11c478d24f64610231e81590e7263eb7b1fcaf82590d1f9ce0e72b16516149e2038a5e9255123501043431226ff8d1d299c7e48c3129828013942bc2985acf6795a2fd3709910dbe29938b352a3899ccb93e33e0b06af9ce80cf12eac36777be5af6d9762992dad2e8c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h13bffd50a9898d6e0627659562fc2163aeb5a6d5283bc44f3b7d52336295c4363428cc077cdca0c0b9494459fc03e01e77b6eb89dce64eb49831f7910235daedc7510fd5dacb3622ddeb00fbd2f033d3667505ecf6c7037c6d9411ccdd333c419f0033af18b45bf5475;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h576d885abaf22082a901567d55691bd55294162ef0f90240ae48f7cb52b5d928c08f60fdf7e45504de73c114ba7c94023e7256b19c11077cb473e17cb28778de2953d9689ff6fcfb1bc3633809d0f675985c17c326e73b97343af6f4125b835fbcb8151b390199c26f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h158989c2225e4518f5b3429c46cb56a6fdef68727aee4f259d363926f7b9b9c85c4620c7a734fa45f28419ad52fbf8ea22ff70d5fdb61ba95ab23a90407f4febbc818a4cf8001cb570d64f4b93165ad164f77cfc654086e93417cfe4df3e947c7c0e6c0405d97f7567c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h279a93f7592f0060f08a795e5689441ecd9279e2ee891ea28a2c0562456fbe4482e432555e1d2eaacd28ae51be722410a4c38cade515e4ae372e35b3bb1f7c6a9e682616ad12b545b11a245b1bac6e487d099c5873b8101bedc73b7108c6795e89b22e7478077e033c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h4fa4c2fbccb1bc0123cb89a35dc827185ffa1ec1b72f3b8118fcebd52859e63ea9415130976a869889adbc777a0224c4cfdaa6a7936fa1a5f9417ac74ee4eb5e80ab1305c06acaf82879b7feb9db2b9d85a32826e968318b2d14d8df103efa4de18e5ce0a0dc2c7105;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ae174767efee85c70a1ed7cf5ae8c875681bb233f7da8a659746e5d1f9858ae160888d5e8ee662eb7d064220b34d8a33516083c9a1235364166c03d609270451899c63b1f620511bf23cc5be99e285c95c7c9d7826e612aca15113c6d1470e0288b5b346265d4f6b1f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h17bb8c309ccd097dad02a3f8a7376e5d604502526846f31cdf0ff2261a71d79fdc1795ab0823434305bc9d0ebd6d90f45ba2453cbc1b01fb41145b93d9c1e9bb38b972183d1575d3afee3eec8de600e86b5e06d44df9ab36b6d46d77c74750aa9e7804edcc6ab17b1c7;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d2e680529908be2f56d66df7931deee2512675c362be04344868bc7d718aa6cbdabbf1971355ec0649f644fc9aa1428098f0eaa1429d7e3fb852087a81bb92ef17fb1939b36c71dcbc60c0195c26135946a1f0372901e5d9a1f6b17f82cb92c51d3be1c088460691ad;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d3d9ad280cba670c7fe1d55cead6d00f2e82d666b103b31acc9d9e05cac65cfc35f21853667e9ae16ff831020b4195af8d5d52252246e1c1ac25be8fd2b849e25f91209ccc98af6f1b79b8b5f989e1095494f755eb05197eb79876959a604b7b4f6b108e0835962968;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h100e55007ae699453d07a37a97ef5ef7a8f77da78d554fbcf139d2ab310eb7941c653c03567972dce68857d49022b903d29377e54fae8c5fc7f89643f0d6ea905f7e9d438a931a97d730c0ac9e8188d007f2e3c4751468e3fdfda5b76ac1cb44f922b5dc00956db9234;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha2abb19ebfa33d1440ae10162c69025604824139dcbd1ce435897539d5249da85d31127a9fb2b652dd2696e0334ffd2449f4b3fb6212a39a3a02d8d2f57bb92ec384bdd67ed5d23285383c8785a55a9879ffc936b3dd3d5b4b68405a988e82a9d73a880787deee5db8;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1061378692d93b038057bb15063632e3a61da9659dcbba7fca9fbf66887f4903cf0d8609090f7cbc9852d9801f13f12973e9daf8a66fe9fa60139d76b2e5bfba0b6ea136594f1e7f8969253be32ea2bde7db773385984e0509dbf3118b9a8d34c348dc61d3ad8782ba6;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h16a9c7f7f26fd5c940c7f8e3dfea4e514d8b6355c04c2a38f48bf5244a9593577b808bf41c69026694c976cbdcdc93ff8340c94b2d88eb2e7d0d894901c679ce32b4d08e0561bd1efce7bc90f1fbba8460a38abd7c9c149b7362503bcc7b477477a3bd1424d1c2bee28;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h86fd1a29746cda618cc94b225ed5272b5d2dc75733b35da6350f51eadbac719bb4d6f1db846214ad69ff46d7d05e5108b3caec64c7349ea6ce7713c663b60929cd3a1aa1d27a0083897b19594ee9c92cee366e21e02c91e827a62121e79a1d5525fd71c6dbd1dce504;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c06377ac347df7473561440d8a94ca5d55b0fb5f048bed196c0a5f9f47eaf3aef3decf268c31620e35fa3f6b13ad99b6148b903a05cfc4b29a3b6b4da932e5017ec236af790fcc03e1bed2a4da3adb8959780742c535ba8de3866842280c4415f85ec407c4bf8f04bd;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h7a25add3664660e9fc19eba2d9ced997bfd47dff69b2825691fa8a74c85f279ddaf26dde32648e6c00285ab5ca44b841fa758fbdcd67b01525f6f23d87314d13e00cb49b812264db9fdc69f4892cba5a74ef66244e905c3f5bc59bb17da7359bc45ab986515df69de0;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h8bbb46a39e650afc969cecc4721888b73277c1c8083336f3bdaebc0d0b8fb4263d9fbdbd4e92d980e8ff98e786a8e1879692f489d68ca9f3c28b360470408b34d26e488abc75deb744519a55a5a55bb848436be0c03cedb995b40a2fc2c2433daa5a454dca47514666;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h933999f1d2d611c1e131a97a4ac5af224160830df12fc54f1d13ea4b18bb9a1fe50d983b4aa9dfd147f3496dad1bba5d1fcc166bf2b6543fcf6c044d1d65d44eb4c61ee2f7922982a6d6d5a852c80a1ae7f4a2ac20e2f576b11b5741f580b4768a0a38029ae1220cc5;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h86057a857abf440b95ffa4c9b7051fd2f77012a10e9ebc968912cc06705ece1f97a826e83ce655f6f239c7b05d2053eff91f6659131654c6b0345a26e954325d50ebf6a7086e9ebb1e3fd99d7d74dff33a170a2db7a7ce3fc36ec43a31aaff1dd145a9b01a004b330;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h16401db9dc67d9ec0a364cf46995cfe0d1bc31d15ca5a02bb45774cbc46cc001068696e03a4dddd09a7fa0f592fed710daf09d1c27fd5432b83277ffbb00f3915556d1c3c66523bad9314f67133a527ba130b793cc50a019a7b0881c5094f9e8d089bbea10b8cad612f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1354a40e2ca0cf44b931bd202cd7be781845c1f59f4b97c38e23083fa6162b89d194792de2673905a2dab67e4f82fc9bc94966be8ad8078607129a97d9bbe539ec03e0f1713b10cfc2b9139a67ee04179f2147830ef90080e516c3ee50d5d4cbfa18d4a8ca56c2702;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1cfb387d789c4013086252bd933eef7b8808cf384cf55f9d4f9474035aff093f26c9c5517b83d56aed92fe7fa56fe0d2e03ef701d803f50964cdb2439133463cf8a722b98b4c3532d5fba4a30a18c9a35d88cad332fd2dd026a8b1931592246efc92e27163014936c37;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f16817e736bfbe90c3803a7251da50120032e20d500c41f8dcc2ab88eca8d2a381bfe5a2c195ab71138fb4d3a7a81e84323c658695b8785e202b7c8b2d7d0cbdf2d92e8f83fd68cdf25bbcf678110f162f6785350eec7ad333227c7445e16e5f094859e4f5f5b1bc5;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hcfadf23dcd5873ab9dd3cabcf0ab54f553f05389dceeca873d5d9c4376019ad2d32442c41c819db0a7dae8b7f056236058fb99038371825db211012686f11a5ac59841463d62a4e5c12a73ffe06bf651ce27ce86692b5ff614250c4df397fe351d8e3a8a39858978a8;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h17629b2cf11a9c1c16ae9a6adf572432e2dccdbc3de1716475cf9d2e53945d69b29df7087b4115d67fd013a9912f7976a552534ea60627cf01f16d777c287d419e091a8c88aa0ca03bba1f289ddedcc9b3c538a0a2545ef2c54cd3bbdc061b51bf03b62681c336efac9;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb5c6f0826a5320b66ff702f939643e0a90ad4a2c898de81ee62c57024bba4328a06eebcd13aebdb19c013a68de1d0262623f397a580162dc25860dece9d35844a417b33661d68eb29a734c9ea3de698e1e17fb7836d4696692c41a59b50f6bd698e1093fc7c4546cbd;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb4b231050e55b6e24d026db662e7f33df807de82ee0f43091802096b66b925c229d2f690f197126b674492f1cb0fd4af4cf2a6397caea4e61ea2cc9217ee503a71b4a4d7437ac884d337014fe2ad1f6b846fe479a850b8be3bf77131c690b8c136ee172fed23cfe39a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h19f05418e49cd53f8d76362c9fe07ec621e597b05334aed666428788c7fff0c5d0e0f08a8626e60c34d7a8cce736c21266d68c430a0a5aec0755cdac057a21a9234bff9a53fc23c5e876fad632fd6c67897be7b29c20bd417c8e12d43aa8ccf292f9a836b78491ce1a7;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf55c3f8aa6c6a5da8b0b82906ea756bf6b71e114866488a6b2d53e17f4db8e891194b1b44b224a6ff4bf6837ed1c3153bdf1071bd62b11bca7f544bb2733ac8319ebdd6618ab4abcfd6d006f84cd587119ca28b334383a693e95b755cb56075294abfae6bdb05f581d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1781d072903d3976a2116a205413487dc071988836796a9b97fc27c89604dc5fa3433b2d8edfd929cbd8c5e4770e7ada657fc25c16258ed6fdac94c432aa7e6f2cc05def05749109b2c1320fb7b62f72e8753f5259424be8bf1c2b7b3b48a22e01a6b20f5dee883f66;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1fb6c855dc85266696efc5a626f982012e8497f6154aa0931b4c542e5f64d3a4aab931d0f20f4fb9343e7155d91472f5e9b190631ef99eb3967bfb825ec3e76fde99069f6ac3f02dfbe6195d119b64a13fa5530a1942e1f550a8765513db9ca344ee89e77f60fcc454d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1983455ec282c92aca14e12a82ef5fb82810efb2fd332f69b2cb5a061f8a508350ff6ea63dcc8c3bed9e00f8d9b62951fac8f5a16bfc1653755d34842cf8859dd0736b8b975b2c4ba0f61189f3286e54d6f8b9153ef4995d7ced967d67d73068c7b4bac75a610b9dd5;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1afbb390700ebb63b44976f6186e62d2a7f75828b2d199b26a111cd4395ec304956932473a386a33e9e20d1956bcff86c22eddd1bcd6ca1d90855d033c7a6060d7e05dce66c2af6053b185a618bc5185636e9228d4f7762e6d4c870d298687f4c1d641d4751f0655132;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b2227000a3c3114eb30156349c26a261eb8f333e287dd4eb8760932ebcd2fdf5e26dd9201ac92680af5839037b6c203dcadc55691eeec4c987bf6131147cb3875c1096007280dac57a960af09bef4d08c645269021c063f9e4c23b4e50582c561f66e8bfd7ba274a70;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h649a97820a3d5915b5217709bb8460b3da2145e706c4584cba9c58b923119070742be5860f0beb19015d9d187fc711a124b6d60b1eb2393e34d1660b69f92769b3451f1c90071cdfebba286bde3ae74332ee14f1695e5c8ec67aaea5fb634725512f91145a7aab9428;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h32df0371be1c2358bb9c4cfc120e220095fc70c9ff7407522d939935bb818b9e1aca19ca342b82cd98a36c62430e39975dbb6380e1548aea7d80a989de681ce929f474e8eebf73444a92f96562a6ec4a8ea4bb137fdf22e13e69e5fbe359ab60a458ac4bf43113c028;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f5113afdc04ca8707c30264cd819b89079956c42c8a7cace74a2fa34ec6b750dff395ceb41478e768541e76ef88bc71cf064427a523d003a73f106624c841f57216c639028f2f120ac32eb9a29bb9b3818bd31ba8068f6c5858c52f5d025eefa5e8124bc33108d0664;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h12d9385105601ba082ed997e19f4aed6c5a589c42a564a92604439763c6e4e616f88ed579170fc2d884c69daff1cba1b264bdcece7c81760acb0f90d7e1c333a43eb389f7ea785b21bbed3d3d1f21d07f15decc218d73e5399c934f2fcf5d6d5911e2f7db787164fe02;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a327a167ffac8c3a2d608ea505a7516343cbf1d916492dd0cd35131d1f63f4488a910d2fcba1321f03b15ba9efd1abd07296c3071f29464957606e1c05b1afa4a25b636cec584b525af6e197cad381fad6168aaa816cc2836678aed59e3a401026b7a1919d40bd3731;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h181671361484e12c4012fea0209c90fa4736f12c16d54c1d48291c6dcee93d84b4552b1e99349fb2b9f678bec7c27ca83c0ebb457a7a95e8bf1b79435c29cb54324db990e9d0dd96e4127f2c5845cdba191d3ffa362626161ecb1248c72fbaed3920563e4f3abde6979;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c00ffd75c7a164d3193edfa0f9bcc188da1232a771087c1f88a6132c0b33e73087194803b678961a3fa35f645cdc5498275e3b17d4258f2bf2218339dd5bb5edbcddbca7d8d78a63a033cff77eaa996486ad29098fd8496005f084d38ab9759b7ea8cba87509cd700c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f1f659c15b6bd10647c41b34999904f3ebb0eba0672f5de758e56e7c4beeff7ad5506a45ec193fa182f67f813d630c61ff6cc3ca249e6a2164bf5e182d93b650d9bcca8c43c0f49b3c7b7ff4e2d98bb2f0cfec3ea7fdc783a58df6151b9608812f699784bd8cbd4bc4;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf7009b6c975e64794dfdfcb75c95be417b40ae884b1699a517350058c79595fb6b98f4a9d625eaa92d77f0b8bd86664cc7901df6741b1e5bd94f3ca13f31b27835259fbcf5e43fd4cbecbd9ebd4178167ee8035b05f026db85d7564ff8fa5bc0ddc783e584bbb171e6;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc958806561e3d42c5e2504ffc5110c9efb3939dd540b4d04a02ee3483d0ae91fff2d84ab0392f096184975a5f587d3f15ba99b9487ad8bccfdcb297726dc632c22c056b8353ab49ce516d936a2877e77880daa16de5bb3bfa3ee07d4c67743189bba3fa3b81532245f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h16bcda58421d2407ec3b607e63f18aba349f079bdf162ac07818a4e91658e3f64acd642c40888657e0bcd7e5e246f16642f148e6680d9a41d3c2f367402ec793a095243ee1e2566174660c2bb6ebc337f318e6f45c09a7daae5ff0f87e6984520ef4d29a2ec5e71f5ea;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc048cf65880020b1d57178883712840ec383f3f30a63489e107bc0986bdbbaf2df949ebf02b071d070a7d151f6282eefcf4a360e5466b4abfd763c8c809a360c7845e39bb7ddfd7c8002437c79da4b17d4b8844d7262a0f313242c7eb565160c3ea40246d3bb7fcbcd;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h4602a401c1c429ae339b0e95e575dac03a8764252e5d7c5404d8fa4c396d6f41cd6df81fcd479fb97e594cc74a8fed66cbb76276e3b3a99feb3bceb24b5c5b61c02ed3674c1fcb9f04a5c1e89141ab61158e9ada393522000d9378a6a50a6f5b4f778ae8e84ecaa917;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h16fff3f6da03c3d439a67999896b62ae98ab232cd077afbb3ff515fba4b70ca57e3b770b16d964ac00fb7a45a0479d22005e7b6a59d40e155b14c7975d926efce53da16495bb71c459932edc88abacc3ce7795d66329c3109d146d49cd2b2f7a560c88afa56974951d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h153d9777093bd2d677e633aa5ec22a636dff994a39126f37995a7771d474445c7c593dded3bd786cdf69a9a37bb15a747e5e33c51fd95d7b480a76a5c2e72ea97c7c8ad94701dd46368206fb1a72b233729ef59a6fb9fafea676d2bbfd0cba4913d640f1c98ab0698fd;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1183ef620d7e3514d970caf81bde9bc8bc1d72e458a7746efe3cda88e3644eb841256c61c7362554d9f8020d6c3278d964c91254409c659c642acd00cf3aefbab5e09c369959b39798dc1afe62253e72aa10cc34fe38ab97984df13073f9029208d3b1b68790c08cb76;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hec2899d2dd3784053e0893f9a0082719e8bfc0006f09297fdd510215ab1ec9f1a948efc46589c9a2f1f31aeb1ffab5dc7ec609774d12dc1c01748bcc3ac45ab25854ad2c1adf9948f274d72756fe8e904c28c3f34d42c02ccd2f62af4d4cdd32e3456341c8f3450b1d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h18081127109778c9bf54db86c2fc2ae2bd7e722b0c5b6f17f6d5ade3e91141e341f463b79ffe467aa93c2c4dc5982cb866b66e53ecb22bd5ef129ea41f8f1235d2a6639b7aeb56b0508377ac834d828a9f2614a3cb9bed74e4965cf09dd1f1830aca661ae699f60c036;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h13563aee9561aacdbe7f92b462e498f9585bbac9f31031e7ec184cd2e72daf171d12a12b87442f42d3717d452c6df88ce7e754abf097542b0ba8f521c8e26c128a35e40e2948a3064151e88dab7949cd03e38c6465a44d4e5154ceb2c078c66c870ae64eb499171827c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h132a9ee10f82819c601626cfb6790b5a3b0b0bd7f20233cbc47e208fda922ad8e730085a33bde5ce799b7c6552fa66650974fe3b33a76f991e19b74ef6837c7b6298e778130e0b77fe20f9160344bcd40d72f6d561ef4b794a706f268f5059edfcdad35a6a3f96d0438;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1950c603d8b231f7d800f1f880a03a7c8348b75b00fff70e7a4dae82558a09e77949be6f0788ec0cf0ce89fb6c44c2b12c8373581d9fc2ac8c03da084b04cc9b299d33e696c4f0055b4b885d825ed093ac43500d6ebbd3cde49fa37c9002b0f8ff76d2aa3baed9c65b5;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1892a657c33b7cbb11a3caacbba647e1854943d044bf445426a6364d189b48e4e602da9e625a6acde931d6afdd98cb59b345b5392f17e9c2d928277430f9de992e1523b8633508717344b346e22638a588be7134901444675bbffb5c39e0fe47ed8e7eee8f9adcbf9de;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h178cad63672fc4de4d16f05cc6d64c1b4bbe4a500cdd0c206a81d869f78624558430edd909ef6ea6679bac7525d139f3e990dba17bfa551aadfd220037cd7b8dfb39f67baaeb373b17465f3e4fc21e35151bbfa631150614ce83f4aba6988898b8417faa0e4d5201a05;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h8068c3d8aa9e3e7c69fafffa8f63510358d3862b87ac11a8cdc37a36054fa1bc27fd46865085edafdf88637e4e65c6ae0f481fd0c9547f4058f32950bccef2c033b4a69b3b95fc8c5d97ee2f91bdf76495d4092cc9cfbc1c0dea4a887cf1c9d559500470ec40688976;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h12a61a891f16f437bebfa14d19908bfc16d638d739fbd71ea3ced81995de2d17b17e0c213fcb9090dd919c4c2fb6a9c683e8772cb97fc031672da9908b8558c1fa88e88131cdb62c8b316803cc40a36fa0cb7183ba9e50562bac8989f5b873ad20e90acb68f7a9a60fd;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h517e3eec4f09dd096a387eeacfd7774e48bcfeaad1e4790bf5fda35c863342130cb74aa1a0fe8735703305877f81bb28002ec4c584bc2d5aa7b422007223c280e451bdda6af6284fcdfb7b3f76f26d401d1adeb1a213d22aef3459f9de61e638b501fe715e523809de;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc992953caad6d7fbfdf04f2c4a8266e5df4ce52c487a9024ec83095cf00a28caa5579d0139b91ae51c8a7e0335bcb3023285f6ed0efb77b1ef398cf02a8fe13e1b1d181d9125a084018d499c070920db2311b1f67b679b47f8d3d2a1bc4b017c8d0b452f0e1ed19873;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h14d155d09962c32ebee55942b16da683397cb7f1fc855995b599bbac14d8fb5d8d66aea71b441934f26363404f10d78168a281f5ff6416c132233f5f3d8a6c8b4313aa190b972f25bed5e873ef4dd81b2d5dfe8d3109ea159a3c28ad0c2878ec08bbffb0b3860fd5c35;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ee021b839b7891e7894d64eb2396f54d5c4acb306732eaa02ef8ee5fdf897aeeeda4597de459b01a0f174f69b8e77485005d5acd03610624e4545a38cd83a4335e57a7870fe749284c74083b741550d3a821dfcbdbe30085e3da23844583d7ccc05b32636a6f43e280;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h18d81d164202bc405bc98985f6a8e08a8e278a7a2a5bc43dfdb38180a8b5533ab44de0d7fe8f9831192c4dc2f668a87f385e5d22bf968a11a6908f05e9ea2e5867eaaa6d748c871f71c7a928dedec34dde248a1d12dc1e7a9701a1c702e42e9c2b84e8214f155999515;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h126b37756385aecad396c3dba8725d2a14ed485195f8e48577d13c391add0a7272d2f5770a3aa2077be1262c1b182b80f499338c1f12a411a0696fb1eaa4a2f33f57d04196e01c4bb62b344b1df022a427e048ee088c272f1c022fe43c77191586ac4d63ec6e15b8bf1;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e39bc0690248c1e24c40789dd6d18457af71fae496f4b88654106da65ea2c2962666a13758dfec871359784a418da4a07cdb60ee563560d1cb8efcf93ae6b4724e70eaa38416e4394d4bfb3c48963c898bf9e739d23df47ca6281c697f93c5b83a9445b8e10092a123;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h178aa53543312f551365200ed26da3f858e9ae7a93d2e9cd738421f72261f25362f61ee03f1f48bdeab49ed532ce9d11a2cb98b5dcfbb634e1eb971bcf42a1b968eda770bfb9a4dacc677e51aa25971eafd51eafd75d904b3cfff1e58872169f72a5b2ea5eda3e819d0;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h18ca11f9cccb9d798304e01c96e418900fc6cdf552ac90b6c5c1d2eba160d9dbc745d75e66c64a36668207bef5104696a077f8b74695cba4bcf10b91807a77ec1997892c5535361e292c1717252d243bbf5597cb5089eea94b58c969203a5e6fcc2bc76a23c383d95d3;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1873f35587d0a1de6d1151ebec735b9d6c2ba1c5ca93f22aa652cde36566da3ee5cf069bbbfe26c7c7cf3eaf8f1bb4f726b274997f208c3665069f1f2b5c5426d903d8d2638536c7349223e7b34c31e2abae61c664241eba1e4c151402f3f7414c1a2f616b74d1e5988;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d4f57e68ed18ea28a1ce387dbd3cdea4d257a35560a2b867b9a834afa36f3fd33e20f619d3942e3cb912b825c5a5df9b66bcd45492e8a707709e51fc8e202a0cb2f30058c753ce5b384d50416c42bcea35e3918be2d8a94eb3770cf11207aa1e4277361896e09732f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e3493ab116c67e2048d1de4d5b6b55172d215c9ae3e3f2bd7b9d1f677b8ce855a35d0abfdaef6400284106260747431ecefdf226c4ddd59f13600acb0c5a2a2b4d028eeb043d82f6192d7766652898ac2b9a07b6c6f32475bfbcc2ff836dda04258a01126687a0ddf6;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h128a8fd62dba5a62124fb4544326c328dfa067bd2c9c42e7b21c8c7b07c20f5605b1ec1042275f5c1c0e7517c639234e857eaa8ac8a8a58a1b6645b6982796cc4b22270910e53d7e855d29c8b36623c8112f0a71d2be435837fa9969341bd7ab8bdbc0f78947c00069a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h170a14b948bd4371229146bba26e3e3eb91c3bb779612f764920fe9cba21d76bd4fd4935a9f695be837886e037671a79b201807b776b0a87b6185058e7d33d31689d95e8c67ec7adb252e6759a1197b2091d247b2aa3ad85ebba2c913f55f8a005944d3ce34e027d169;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h12073e625cac133bb968dc74a7c4526dbd9d577d6a6ef9f5c632adbc1388a95ef2e005897a4f221d4228fd406a564ba66cbd1fe446b30d8590deb56ea655b419e0a93539fc97a5e90763bf0e0f75c67b538bd226e7220b191495f9c8827b384f06501df74d413e4d174;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h187a20c6d13169003982953d8012c1c667f9c7115042b37fa9781fd1cd266b57e2a3e65fabfe142d8badcf518124f299f64f6362e008fca644a687408ea4550a663c9e2afa65c5a6b6ba71b946c029069d23dbf234c511656b5a8ad28899064dc4019474bfa2867b55a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h164a316c181397a661ac30a79efdf01a16343950e86f83aa4d3868705436961191d4ce8f0d1590ef6c2ad3cf552e9510bf05d1a33ef9080d67135d8a377d37083243219316ea0ac19b09bf79265487ed42324f60a4ab746fb7fb4c8867bd269f0fc585f5c08846fb977;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h5bcb4eeba603cdaea6a23e0a5fbd2f1856bb9070e4bd847190b843d12a3c0a7e3c190e59121b63d84256b02243fc35a0b7175263596d99113e88aa07af8578d299a596d339e0a967f0f27c8469a3de16ae5f9b525223b22f9a90061362d20881577c599934ce619ee6;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hff27a86d9b3b68e37c7f62cfe1d4ffcc2378cd4d75aeacc8a581c3f5e615aa30a5c523939a10fdbd298ce66235b53f5ab4389c50a5b788bdf32c7678c142e50eacd352de76fa0c7ac75e7bb19819532372c0924c11dba548ea80bc34aad6bfbc9b523da22afc07b949;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h8888850f42a093606ba993f17345ba19b598e500fc71a5004105bdefd6869a8c97076cca5a1c3d29126f686663da30c4f0ba5a40d033230edea1dfd8efe1b623cd4dea06467cb50c1353f2879f1d3222e3f48cc84450c4be657e0ef5489cfdee589f479443735e5caf;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h654f6a8a27080e7d075cbd231c42fabc8f69e7145e0d9eaa8337c0c98132ce009d8f239fd5a0c455776662abfe61fd9b3ec9cc2b7e327f5a7971976415a7a910c73648c3cc749960ec314ea550a36a14441d6887011e1dc3bba8a5f1b4dabe7e7896b24d3d38386894;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h2ed7ee9381e484da01b235abff2af493eac27faba5f681d9406a9707fdfa7cf047256374f9b3fd3f90e6f9a52452bce48c360b5f29059d28bd1253cefa2f15476c5e4306fcd770e8041ec07c62dbdf72a45f29c071c0119b840f7ac9cd8249f4b363b0c30158dff29b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha74daaf2e4cc4f784e1f9a14e7a7dcb372ffdfde41929a93b9f2d72bb37555fdef3914bc7a2c151ec5765e2bdb5966d23e987b1c8e9b642d3cd3e6476c515b11df3b4f97c5a7a4c2edeff1518131c51010be4b0ba2eeaf88649d8c4516f5a0dcf6e0cd08055ce42da3;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hbe50fb985638466e59261539e882fc089155f33ce63daa840a44637b1efd1560b98c8f434964e482fab1b131ed83636b2be7bd7edda89e337fec92aa81378fab83b94e1a07d715cce6b26731ee746a525693c4c7b6603ac67a82c7d3747645d46018e518a6a7d30844;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1401bd3884dcff23d67384846f0ee0e9dcbc6a17f610c77e18d48de53bb17319ec26312f2d1e6f3f37ee00aea2ae6c05fce386a8455ad413f24d83592fe2d8f5f3aed315d5515da829192bdfe78d72bebc33878c3c93906e7ea32917d1e17b6e3cd161056f9e84176fa;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd66d48d060c829611290d8787f867ff2a9f153463c253d56af691e28dd3e744437b590be1c4a4426061238e66e5e9d9e468a2063e7d8d9100c69473bd11b6df9784c25650b1270901a6afcf47cba0ba00f4f47388ed13de3686a084480acc4bb9ba57d4b61638bebc9;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb0a2d3ec409ef55d4836a3363dad081c063ec9d6f6a176e06571e069f53e1fe20022350062a2d5d5ad9d4e81af8bfe5ba4ae58ee32f2015f55c3bb0b4315808c8223b688c165d1440363b0eb17c482324e6c1cc39a7181cc110b26962445649ddc97b485bafe8bf48c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1cee810d2c24af9b9327bf837b789bcc5833c2e3669de5dc81bf0133326e083ad7da238ad428aa4827a745d85f61551a5a4198d7e5f28b019cfa2c44edb2881e35884bf4bbfa3449f7bd3d7e9c78a53ef2d7746269c7759f1045f36bae7f8956120c6d7e475b0dab854;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1efdb67a140fc32c7cb413d4152adfd56773c523e626765df8e9fc1b889110651c39fd443a7640b1592e980ac923286b0b8778515e2003828cad562face7dc1d6c8e4f56ee646cfe69c0d9faeb7bc647dad006e9d352511237ec986cb72ad0bb1d0245be1e791a794b9;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e5a4a150e8c4b55bc56894c656032cc73a69b256d22bf509e02079c770491ce2006032d4b68203a88279b22e04aa5530f21630c6a4ad07b415de6879d68e1f19b8d8250c02b314dc7b8fb7719c9f12cfb711e5fc88977ec8e5180d5957846e312a942c18d9fd5c057e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hbdc0a778f6db06d52a8bd970b91f4a7ade0346e919db556d2182990e51653dd4f9b6eeb3e71be48a9109b211d3961013a1c411a0ff08571b0f9524a2585bbc061eb04f10e2649bc4167bf2a57cba3dbf3903b55fb025871a1c499a1335c5d39e72427519153dd3ff50;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h3819d39a52b64bc0862574a89264eeffd35637db2dcaf30b52701d81c1af6400921b48fb8bc6d92c7de454d327b4f56801bc3e897da9e20cf97802c15356643f315e076579e9a981da839572752fbdca7b038a982f86a12a442596ef105ce41f930efe2a5539c55bf3;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf3707f34a45d21aa909b7c6257e58b0c551fdec0da284c5a5b56e88790d4d65a49c1d98f53496b4d292da7c118806a09bb32f68ff406b6b1bd9d3d21fab43ccd0bf7dac8732b8d2b01c51bdce9174572bfb88b478afdfcbf7d1397cc21f7b3391ed2ae2793a4c60c7a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hcf42c95719becb3916dcbeefa810a289f30f3fd2307e1b418f62666033bb4644eb538a353bfe3691b3f3616eb9827520b0561f6d54f062166013ddc4d14e4b2ba4f76a029e01b342bc183b740a0c8b7a178ef8908fa9a0c981948744dbe156e203199cf79468bc548d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h706fae00ecfc088b1953adeaa0d8c1297915f5ee90e55d833d5c9cf685fc9dfda55c0e1acdd05b30fc1134c4d1a4c500ad7b506f2a77f9ab046ea976f702be28399bcccdc0c3e58382b82fc1ba5b4e3e73e6077fc0c20c1f8cb54ce85820dfb7e14706e0c2ea12ad7d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h13eede48acf3de013973c542b1469dd8fd0974e049df1c0f2768abe0944e9eb2530f0a6ee395dcb60e6ed24f7ca00579dd7a9e88064e693d9e315127ab4b1dbe2c207a022fcb13940c2774382ea34260023c167233f29fe998a6fdfec11847048254fa842a9febe3ce0;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h850700f8394f45f845aa55d101f487162311b45a41a3bf9ad233e148b7888bc16027caeaa5042e55ba47a26799733bb2e09642fa23a814033cd078d055c32bf13299b1a46bc4bc3fbfcdaabe4a6c1c3b40eaacd381d45b21d14452b10ebb09113ee17c500724a4549c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h191799fbc882b6a39fb86769cef951a9a32214f0a3dc0b128aa6fd278b589181b4a031d77f75e7274474b44daa0cabe8a5b675e57101759aca08c7e5c3d15b99fecc8a735479df1522c6a3fa43fac32cf35469fa9148006ca25acf286df608174ce7c5a2bd4ef3a9c74;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h19a282aabe83869cad27a35933885d19872cafdf53e2495fd42a1b282fc9c099a12e7312510f4b7cfbae4a8c5bcf42ccca70c292230963d00fd82e674f2e8befbe77b608a53746859c273d284b2b5a6b9ff8a5450ed9779acda3c8e946a9cca4126fd43389c03ce947f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b9fdddcbef1c7a225e1180aed1a5de6b5d607ee7fd78f08fbd3bae3675d044d2b2e2b50859c746f15b10e04809ccd20ef38c6267be4639bd39ca718385d51668c463f92f3ee80cf1123140260ce5439837d824d10e146fc58ac25e58dbf566c67ea8d3fcac280a3764;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf6e2ed0c40f3cc643c0ee2ebd5359c4f0658a5fee4074f2551f21fc2078c1854b6ff0f8a89072a0d78464b009f6f2e319f6a3baa47709dcf9fe5876376463400239641c7f95201f0be9685bad37b0233eaa87f0d7e90947cd38bf58d80e353df1d0873c30da7dc53dc;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h237f96292cb5748d6822a2f03c796affa2af97b5efc9603b04806474a7db72e5c81b28629297222bf98917a2bff5b7557aac38e673118678017c25c08476c665d6ef840e2b4e1eea6cc9ee849f5319a765f218c9babee60b3000378c90d49a36ba64aa77f8abf247ce;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he786da4d2c05a904d9fec85994b36b63c611ec219ad0d8837448e4b8cc213168d9d66ea83b8667a3fd9dfd82e24e3c7825216e7fdc66c5c56e7c0ae88d688549107d71bea487099ad5c98c419889e4f58d6845df0e302047a9ebfbc78d670930c1ff046c67911d1410;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e0a4e70675d2a818593957ad2a6ea335bab6b3faead0f3d6d7978b33234fa8833274eb923223bf067e994b9b9b67f25993fd13da910d91fa3b8862ed983cbd8c011ce3cc846d0de8f58ed272d556d839780bb5100e7927819ea869c516fabae1db77398bb4f1546637;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1365792f05546d68bd18d7c5c518043bfb2ffade35d11d0f29583fdb3a6f75018534b02afedabbd2909de592a1ff15d74d724082d25d5dbc5acfecb89893c165401f77e7daaccb7116b07d52d9a5fd8e8af93efa01104f981b73a27b4cbe0a8ae315d7f35c096da03c3;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d5127c88004d6b5d583125d3dfb027f583bce5edb66a4be09c5bb66d6c7e58a597774f87a0ae7dc57fdb3538250b733616bb1ab94c7a10e7f42aa1f620dd986f15bd7f6fef265a7d47c75d7e4b548ea600f9626c0cab38bdbe9e44d408f27849f131e4911aaa432695;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h7c2aa5ea93a10969c15c5d90ec0ee743f8ba25668a004914f135f3ea480ef9f9faee614f2293d25f768f741380d7cc732b9f43577caf845b1d52991b8e02c4464a01eba5111867978a444ad39a5c0f770d292964ba6869029c26ecc37d50d8a50a8e20e94c1661e400;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ec561a7c11c1a8095fd4004eb159dfcfb434b4dee9d1644069830de7dfb9df7c7a725e1522080a6d8a48629eb03960090e676fe2f8347bd8cb9fe49ce37dae7e7439f935e3a115d6a763ccac6925dd9d4448d0db97ce3d23415907a704744097c2c16551b8c95188c6;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f562ef1db84c1e3768328d0f269936b161e8aff2c801c3e1243bb728c040761a6a5412386c580e9937f80e9d934333d2524ff4c703a9f14156a0ec3bc41367b4b8d41bb8d019169806907959f1e8b1e1016674696e07f23855e2f7977f7668b638c3da19a2f7d5971f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h75a8d5b03bec00ac97e3ae04d4350c99383850ac6479b221454c18270d0b5d5fa4a16a26f9ed4b3096fabaa11aabd7d066cbec977419b7987e5eb4ad6b1dd7861dba1b386fb3f43d8c0c6a79c4606c2ee2ce1ee10023f371eab92097f08186eff235a28c38f4bccb3c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h74e02a8091d3b25fba82720bd48e4602d05fb87652b09ac24efeaa3b48f0363354636774eb3ce0124f3fe0935b9c80da6b6a74d33e874a0778ff8fd806d7001ea4ab410cf46c83b8d66a955f9e5a557db17845b06a2e8661840f779e2e5d3f79b92247b604d5f5ac13;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b3462d8ee29e36109763adfd5153b31d378c2b9d556d4ea25f7e7a6b59b3a7b2aaf361412d015f1c97aaa8f240fbdadf26524c168a6899cfd9015173b2af54fc49b51e8b0dccd5f9ea3dfa6375ccc2628af4770aa93ae76cb7976646252cca31ea8f831426dbc6a668;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1eedbedad2f80c5f833c34f41353a534cc54138a7f0e7804df50196b80a1e7e51288a71d0050268e1a22fc929a544314db7d1f6e41082e5d95748f007fac57ee11cb57426b81264acbd50315823749b03a81db7c2ee340bc8b5f4bef9da41f8386a17efd6ecc78f0d9f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h128e2752dd4f6c67ab04ef6125738276aa7f9a2f73a64b6bace84cec3db2a677d3cbc005b3e40629fca742acb56171d47d01252f1008873b3ddeb10602b5598f527665d79a977e92f6f20c28cfa5c8b38d7c62bae59d91d2352dfc384c7313a7e9b7b79cd14b56da94b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1069ef5c28d63f273449faa6c83f278a2032bd4c40636608f49c2bb237dc9e78849f6d84635cdc1598f5c6bfbfd9ea24512c928a005bd8279570d7a4df7ca58b5f48d78edc5198bb988badeaa07553c1e968bf1078852c6998d8bd1aa8a603907f0ecf780c0542e9f56;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hcf6622875872f247e654a8b730edb3a2be18cc2ed888b2f298511174813bae15e6048e680e8ea48a8dc46e1a6ce9997725643c3ee251adffd760994da7b61a642e8339a083089b0466f9b114cdf790690cfe5fa7a55b019f961d72bfe34d33a5bf179b07e56fc41e72;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h45d43faad8c928424b930832e66336dd5210966e559848061285efdc72afca6ac3c7c4aecf206c6ea6de25bb1d6e47b4808a5bef935984986c2bf4871ed81f1696915dbc925b20ec87ee7e7b0196c708c136846dde4a03847c84e5686920c82d33cd5f8122d5e800ca;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'haec82ebde96508ca36345a3e86eaba19116ee8b847e0577c812c4432d814faa26b0fbca195bcfaaa980173ae6e3da2ca87f3fe454a37b676356891515b765ebae11fc7f42075e7e24c526f4838612aaedd0449997f2ffecd195dbdf381dd7b56a3e2faa6e595512f26;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1bc687484f1b181610304b7c304b644c68f0558deefab5f479d7268320a002682085673eeff035e5a625886e0f628de98a08e9ef7dbd99240e1a584d7ef7eae4e06b6e3df0f5cd298941519a74ccfc8bad7627d3ea9ec1dfaa19ca4d7c273c2d4cba57f6e8a1d61ab6b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1365638fc1cb409b6ce1e61218f7da8a9ba43a1ffcedf573fde97136a1e931659a06ba4f51c223513ddbcc3e67e434dc28fbbaf8115eb1eb8c29917fb481ea4baf8ad17cc4cce8de24fc2fb8d59269f4ed9cb461405543b5d973f1e119b8d87988523c8dd8e194863b2;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1bd70a1f300d20a7ef092a0ee62e21bbd9c89ab5eac126c25a0fa8a10d4d535abacc8344fdf28cee78672fa16469c07d9a2798f49f3e201dd45cee0d8d03250d81df574b10e4db204d359c8d5c3ce2f68534fac47d4da53853c8ce426cd87599780262c564cac875a12;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he0bdc81c8957db5355a186b125131d087e5d039de986e0334a47f600c5190f94db3196abd46c8c991eac4b27c2e04abc6d9d97442e101e42fecabe32974e854b0b29e2b5bfa7374f2331a7093e71376d50aad32ff95122ea0898c2c01b6e68eb62b3aadc909ca0a4f5;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f01d65d06ab8259a9563fce6ed53ec50086794a7f0e56eb800e1bf0d568aa92692957aeaeada5f1ec46f75f66a12f9cf80299c68ee136bdaf42c57e87dd3a6253e37b7991b2231276a679914c223723731c79500210c2fcd6475e8feb9876b13b8354f1bc12864c826;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h7e524997c65e6b931c950c53148706b84c0e1c0277056a299df25bfdb254ac55b82ffe7eb75f79ac370da1c9cb4dec676dbc2d60a3ee16686ac0d8de24df17ed7c9a87561f03e3de0dc2d3b45da2a68e7cb6043dfb46bb04b754acbea06547ff4fbc4678b2131ad3b7;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h7ca648b0da5607bf1b6ff473179213e40f8bff61447a3e0667440a23543471dbd2fd892ce9862703b5e90157956607b0e2794665c68467faab012f260e0961df3f61aa4b98c85ed3debc68d410cc31991092265a8f5262b154008c2acbeb5c44c017b00338fa97c7b5;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ab663be6d5096c925d47424cf5c13488106169a90ee86f5fb186f0b45784aeb9ac3eb84d1496442ebf3166c5d321bcac273703278ffdd499e7612ff4610d2a382359990b10451cc1277ddaf6e3423bd70de4d6c2e04d0e4a1e6dc8e3a5af4ca7df9a49348693393894;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h137613f435570eb7c49a6b78e585ac9a65139ef588d8ee40ab9fff319ccf420d8a60e90c7a892eea265a8e0282222124c9c98059975d861a1da0aa39314c4a1d5af97d6df8824aec49263973e076e5b8e21d8d675896f8c33c45c93176c3a0cc9c07ef30608f017ba61;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1fbb0405255a20a7eaa784285883183601d660ad0c7fffa6cf359014438ee8ad231b4a7f1291a94dae46d156799e701facbbd6ad1ad5feb10748c83be73d94ba2d78d11a6db2e7a0b25702ad4ceb775f43f05db3ab9234aace2db1bbd6af736d853845346d85b66f452;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1606adc3b2c7322eb09a312779e7c93612533ae777026c315c83c2f8c28153d497d0cd118d37d82d97b408c4f8cd77d068ab13320d283e93b8de328cb9436d2dd218000bf6a34527eb548352c86ab9c2a7663eaf770953b63ac123d453e66b48addb6f92213e91eaff6;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hacad8a80136e004718a22d0f48ed9cd86bd8a3a0c254c30a1a5cdbf4e008fc12627134551ba52431ce8e73d4db6d7d57f190e4441fe61bab5a7e323bbe60457d71b593abffe186765f609cb6c60305ba7b6678e8c6af1671c28149050cd26402d241ecee08f5fefdfe;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h11ef25d835a855764fb5abaad749d3d24e9f19ea66d18c63c0f5e14351e0289f5c74c1cdefda1ed5e46b44260c67e14de52eec112b91110bcf86c307fc39c8502676af1472f32059de81e05a70431610527f9d5c5e20297427ff6dd5caab7f8d03030ce16f19e2b2771;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h11e0ae6a9171beec3a66b11528cddeba28ee93d6aca8027a5e1699e537e171bda412d857d9fdfa15ad45a44a56ca5a41055fcf5814566d00d1c53561b82bb910d1c557392f6cb210b4b7885b8eb68c5ebba326c4a2100f7b64affef8660a7e87867f02f69e54706142e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h3d487e4a1aac50a46f6edbafe8b8de59ae0e34010bacea654e90e2b9b9b2872a5983c5dbed71ebc60434765204feeb05f023859165a31d50e5cf24947f36567161eabc487d6afcffbaff51ea7ac893053723e361edc8b1f2f39e316ed18206641f98bfea3fef4b9808;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1977d56d437da2dc83fa8ffb51fc49fa963a8d681b3020613d2cc8156384c08b00d9a958a7734b8e09eb5031b153cdc427232366fab29ba3ec3a342cf544c3021bc08b3888ff2623dc52d4e9e617f2695235de3de9d580cbf2a6e9bedd80f2eb5176d9b70213b06d2f2;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e0bb0ebaf17e28b08ed0260356db5a2e445898ec9226f65657b279f79eb4fdb620f83ddb45459bc829e76b618123ccca4c36b2ddd6c4619497c07097472242293a06ae22c53877ed45bf69eb79bc1789fa5e058184485c48ae314e7ae603d0cfdb905f6a219061daad;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h16f6153e9835ccaf61f604414e4de520d3a5079a63331ffb3d0ea6e1c807269034789c1b4daddbc0e2a046ba341f954b8f2c03b6d8f1607d4baf03c37c3ec69f943ffcca21c3bd643dc724a54ae1881bfeff61ffc58fef641ff123d42a9b3d4cd3ec6c382ecdd182ba6;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h5840eacb4991a71f5362505580d30a9eb1fb56954fc39135ccd8108942856b4ed82a3096e543952df2213c1a1aca567397a5f6ed8286cae9cc29c9b2c7b1ab0814304d7f8d6a97b24bb27e05e7a3fbc71066979c7e1e9ead956d4bb69746d1c144f584249242bbfd8f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hcd45a6d4a13402ddf74b348edbbfa256d628fb334bdadee1de93e725548dfb74016557e460b0589de9b811689ce9e31c9b5e9f7c571e5beff00e61b965de5dd83b509bc5678b2c2645327ccd336ee70e471712222af2b23d3c6d81ed15d6a915b793fc82d8b7a0694c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h43f3576f9a4444a20cc427b5d0cfa6fa47966f546882b274999c829f8296150f0675b2dd012371f83de4af8a803cc90ba5ecf3120dcbd327ed2f73719bb188389316cda10605a5a17c064ac140afcc9a0c89673ca29a365b2459eef286f995857426558582e0623d19;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h497a54e8889d6a0fb5438e490649274a1f59c473cd89fac25bd7455c6ff3c27e37cbca5df6caf497a0ee151e61dc6a91e4dd0d4621be1f7c8558b01af161e75656358c376937aaa29abee20b002ec02dd6ed3f955e67b92b0ec52cf6c7e1a57aaaf210a378681799ae;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hfa4e4af43323cb336b0436b4587629ae679ca3775b98caa68dff827a38b8e2a50625edb2bfd0eed30e9dd61375e16bb611670fb3fc7c9983604ce736bda9150a938f4f654c8600db770bd59a6010af88ba1de4efe267af1c0471992a8a9b82d4f21aa0c3c3a46771f8;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h8c9a71b921e1e3a5f7c261b7e8f042eb0748914403a59b23dc06bf95c1f03953151618fea2833110a16827d0a46146dafa545c971f37707b0230d8372c1869a51e42bcb4d00d8aa5aa452d1e036aa2f5398f965ed850debc3ae4b82a5308a7c49cd27554fb1e746da9;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h112e2030f796a80790aff412e80006c27d49c7b6a148bc465ab200100a9d9bfbcb75dca8a73f3f3c155e342630c5b9de001d87096140fe5b851b36339fbfa00c6a488438065d7b336fa9651fa27b58c9791f097a11addf1e35d40fa9400e52ca1cc875c8a38f1dae050;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h16063d4d7ee220f6e22329a626209f57b9b19be28720d457c2c24fc6d3c9b085d522f305d57ffddeccf9df6968beab635c146831ab5dc84d3c3f727db47a529d873e1a9c29d035653ea06f84841f684f7315e3ebf19a0b84f2fdb80cdc466353f90ef886228158d8a31;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h418c580b75cd6f12f70835ee8212b7ea3f2727dec46de4d6f0c2b08000c7728a347e5d1fb58d59a9e4fda16d418de3630ee2e65e2260b3fbf7ba5274fefb392b4f03335477824db498b36e7278a1998029cadd3f17dac6f4a4099472d51a79be7d12fd4128b21ce264;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h19bf535530f1f1cf93b66b49073a0becbb095cd4ba441f016d1ce32b62afdcf1b8b3be038ce984f112cd8bdc8f29dd7b8d84a1b795044326d81cda3e4a9583e0a694740a2d8a9c3113fb15d641f8fa2613ef21ba0096eee6ed441c74c104c70f42aeb6d9b57d62407ae;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h6a8f4605a515f24a9c44f2307ee4c4467f2f08473090bf5513b4b1352d9b0bd0b259024661a782f8d49e2bf6ecc5616750012bdb480f8aa2d13cc6bb33a22b18a4ccb24c69f12104dc36ce8aceff5a94c90d5dc9ff72a08f8ada32bb55414004588de8d6e2a002b2a7;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c464e1db13efce09031c6b566e512aca8e107445beecd33d1b607a9cb754f02b247195f4deb6bff2ee587db3b1061a9b55c53d774f6663ce3c67cafff92723530fb8d000cd68baa7c203396f99fc835846376d6a71b7e6d7153c6ee6875a335b8b8fa1ae22a5294ad6;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f996a9b47e504826aac94be0a7475d6b964b71fb079a44562f76dd88c3a9cd15584ea32e3c76e02772d6337af3e293d07933bf41d3a86c22b1d44fe41b2f52f0ad383595ffaf339d1b7dc7e20813cbdec9594b823859b1d0d91b36544cdfa12eb84738adcd528be6d4;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e991afa38ccf3e83b21a4cd62893bb0597457bc54b4b91484e1afb31084ead680b6b487c51b4f92354ff7ad5ffaa5a56e6633aba875b62eb307321bad216b8e6e3288ee46eb74359fae302f6ca66685ac218ee316f20ed3ca1b7f464832a6197583ce457225d70558c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1652515f12fabc0bfc62cc6c4eb2386a5e27e6d20873004636e27513f8a75c6943136b81c9619c1d4fc45dfbd53258cd3ca9d4c7e3ec0c2fbca2e5a5830eee1bb07ed15a68ba790ad12e5cd3453b04361666dcf962a2c9cf8257b9dd03d46a5434f8af5f0d5eada5081;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h13253bef58ef40a0a82815c0b94dfa975abd2d753d763207a529db76378550a68072fbaa8c84eb5e0a61e2541f7544bb2abf897920d81017e52481861ef780875f059735034bb09498746a51a7829c9178e2bc0e6b3690b693421183db57763a7d457577f2fe2a80d5e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b37866b86e2d1c3ad1889e3debc1423acc2890027313063a0652fe13a9d4b6b75ddfce90ad7b5c442ef26186c691e6261510baec9cf77d0e78f8730c50486dd23f3984e24fe63862a854f28698cc034fe1baf00a9488b59e2fdda148893b0f8bf9f3db0c7cefc62794;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b50dd135f5bff683ff95fc8f0df71a32011b06363becd406357de38a895914ac70af7751da000a8b8aa674894a7d2158d94843d6dd746e00cb44c4e957d5a59e94a5a2ba513010d87df10fbd68ce16e9cb2ea743c51f8a9946e221d106aae82d8b05b800c17d9a9344;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h18518b7d565058ccf60ec2d16f4bf7bde1c1654dc771c546bb746506eeb64a6a29dc3daf0273dd79596a71b5f896beab4bdabc49a4610517627be4ea9def77589cbadd10f8ac5aee0ef81f8539a7d6bfc73487c5cdc13dbc6963c1e3486f1b3205fe23d65501bce8a07;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10d2901d73a96a911ebe4aab95bb4141f4b16687fc858ce2a6139912fe87b806eb8352c2005e8fae5c3fe0921af4fdaa287bc7ce6c64f4312e285b07452fc1aa4b2cb8ca0d4a3b674933a3b3b23196df29097fbc0f92e6265fbf3ab3cf22d83074682e05e659b6433e9;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h6bc3d90d2af1427448ff47900f48916ecdcf4a429bddb5b50a92970f089c9632276486373e7fa5e87cd78bdfe729508ef3d47729892440a918450ace9cbfa6328e642f61b658ba5692bc3f2d1db21a4f149bceb52d6651caf9c86f364b5325def6b7e515510e659979;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h15838b27487c95109695a30bb34c2eeccdeccd54f3737e0293c9dea32cc2af894bd3a2793330ce865cc07483493480297719c1508e92fcc6f0c5fbca7a021e66477b65fb6e055806f7d878dc4f20cd68271f6de1e08a4228840b9bfb58f703f7621bcd61b0dd6fecf7e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b667ef86d3d74eb16b0ac8d22a270050d21c224d049182aee2f8842c77750a98f9ecbde761a314e090d73937c52e23da46b9fa89edbe76b0b87dd15f4db1ed70731e6d853ec85d5fb702a5b015a2ac641b8df850bd1806d05366443da6c1c86fdd3ffbab6eadeb594a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d763fc3ce6ed459caf53a90f21f1729cfce1580fa216bd70a0e520b02f9f4f37e4e8897fda88ccb97921921e4f600df10bd297b74b5c3cf8450eb6587fc4c7a8437d65f2ef3c492417011635a72643f9433b5410d2556ba6b5fba85f59dbfb1c90163e21696d88f369;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1bd2d355a0c5b4a1fc3e5160707415ee67f03339aa116cafb94b9b82bb3d9f5640e1859373c554047c5726da34187f6fda1ef289b1a7bc0ab1040d902c4021717f6d30215fe69e6c1de0bc4cda1178a1b2465b91c8212f517861521be22288cabddecf59c6d998b4706;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h998aad86a9852e568ef82afad84cf3b6ac193a28b3e77c80b44b6e930c80103db95f004cfbfb9f293f70f583a2166c67e7043f16ec774efd5eb4b26694f4f0536d3ef2aa44dff81ef3a16fc8e3385ce5a69ddd2fb9b33ff83da7461b1ff6a86641b9c55c1df13fc5c4;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ed49a6ed73d681e1544656fca36402d33892d162a35e112789101259df9a8b551f94874830830f7694a34e6112660de66aaf50003bc199c272cc44aae77ed6fbfa235ec0b0ede6a0a15b5d208c58e45491ba782ba3b35d63ba7c49d7201e648cf25539a755c33e3e9a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h14ea296a2220622054dc83523ac90b640e501f95d987562881e41f38091e8b4d63ed5c8a4b632aa75b1c24a4a5b7652e4f49ab94e75f1a68dcb8a2f8fcae1538adcb686446403f4f9b6ff312f8de2adeb2195c7b6bbf45e3dd3577f709eadcf3a253d3246997e361fd9;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hff310938e599c7426b07d35fa0085ad1def39b42010487ddc745517b82b773ad11545d4688dc584665a4c14ec358d34b8a451e7e14961b2cb99e6b263c1061b7b2d501db75ca72600dec370cdae499d1d0dc40ed5babe7cd43e3861bbf85dd3ffa9982d154277b18bc;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1fbc79df51698ce9353b619f2130ecd068c937cf852c1138b25bbde237b96361b9de7b10015c1dccd30578c3f3df9f239490d633c116cbde846c88e53b9ed7d8703b759dbd6b1ed5dce12085ee6b29edc9249c91dcc0e2aad1b1384bfaa08cc97ac36396a70f189aeb8;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h28b2702cd4925af53cd0d7e100c5d1f1a3d7e83f46e96a6c68762e6438bd0220ff9177af125bcb17567d8f719147ef318ff203cd7bc9a9bf8088889d8657128bf8145207c235a1aab7ec6e9ac40cfd9bd976c482186536debe698c4fdbfbf35c7d44fffdf4784ae5b1;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h8eef98277c98bec4cbec59ea701545950352dde9a4d90dce833a6df4f001f7d1f9150b265c3538c8ff74ac91004d0624d563871e65a65567a248194153d582a2b663dd696486665bf11df9f66171f9e19e7246b405e9a14a53c9ad8f730c12b34cafdc36c5f3a8b3c6;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1913a9db8f755a1bded60791bbe0024c77f903483b385e39945ce01e1d2e9ca29edf20ceec926dceb02f07a551cd25f5304f87dd0c7707bf3f288ccdcf35fe394d0a84df30d8349fef9ca759e3010adc7e94469aaa0c41ce7b4fcd3f7f445a8970f7f7da3c656596cb5;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h5bcdb4d47bf5ccddc9b8595e8ce4f85fe7deab1214fa4a678dc012682e2d18ceb65e7e9bbb09562235146e850d111bf4dea859492621724b4b2da3a4c38682f276ff73803441945d45fc12e593dfc8d1b3cae3fc6665168b9174ec6e866364c55734e5ce72f1582448;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h445eade3249d5d40a35e71370ae0c2333f4b0785e47dd5dd6c0d38c3b164dd1c5e1d8e49c38b19dc75cccfe4250e743993b45854849218f368f95f9ea7e71b7102c42a681b6053233dad29a9a8feda81c679a8c7801effc823d4b48fee689d65e546e34929c049f0ad;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h19c7bdceb9111072209f73bfa2a0b26fbead042ce58743ce6b7e43dadea151a80aad768cf0fc313dbfed4b716bf929440cadc662cae3bca0faff694c06e0f0e7e90acc19100b0d07a490ae05f9e7ad41e7cf89a2d350a3bdfaae010f1e42eb783391b9da397b4bb82cb;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h724a77e1e1d1a18d412eafce7f11fd7f346891159c61b2d36f2f0cf348479d5dcc3ee93f0100564077ddbb8cd64fb2d77b95b83b94673026d569860f787a7f2a33672fa23b0117f04a0bda66b3be86df4836f66a4dd31aad0b1a5b200e6d561f0b2d69a8d9ffb0dcb7;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10dc857ab7d8533aca4118596bde56622e84df1694e90727202739405ddc270c5f19b35e4859484fb6695b8012a5bda651c8ed7ebe670c321d40bd5aa73bfe311d25b0486dc4998d86a5d51fde8bae63c7eb18628f0e07b97281167176fc70d976d2679a874e2fbf041;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb8d7f2e4c5672dc36673059e48d675a7c8fb6255b99cc986cd5bccde6c620eb6940ca89a931fd12afb0b299440d2e4718f47d01f9a2cd0d27af5bca4492f087bcc50b1c45579231f7a3caa6558dcd9498c4c97c5e33c317bb7ae55536e33a365ed7f9ac6c1a00f2218;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd15045461b052b89d544212a545b42ae227c0b9d2cfe66918eb3ada600cceb6a5ff3c65603bc9264b8b1463951d23a555a9f2599bc83ff0f8da676d5f9a1611710204bf4c346cb0173306b8ce38db31ba1a7b306f81a5ca4f54d5615601d36f15c2d027d90f2b5a169;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h40e1c89658d5f50ba2b26dae648e7f9c8f8e16439cfabdebb18ec977aec22e464d6f5551a9861967bd4fc6ff2cd3ff2a5638182545c183d4bac20082f76be38e09e8bf64a52f1f09b13fa983c95f8276f4d0df852ba5d2553fddd5bbc8d7afd9c80c0904a8b95d0218;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h14cef8501ede12d707d69a804df8b78f0680994431eb3e2bed0641d829ce602c231095080fb5e5a99e5c135ad0eb4bae06b22f89223ba40d40630c9f3b297952b6dcd810e3720aa78f8b0726164b8c2ca26bb9f6570627f5d9add70f94dd07f7d4ce6d487de7f49ce7a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1435d561b7c3bec29f7a86e78f9caee3fcd3b20826d660647dd32f9d347e3430846c05f023f3de265336ac78f2aaf866c6ab5310ae643e87a3e4ff8f548c56c68e1cddde06e780c9fd23a8d80a1d0db1c89d4486dc082e40635434a3b780d2ab4296899c48f5da3e9df;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd71d2ac5a641fa3ef2ff841bb87f4274268676f4c300484f3df6fc5da3f5febedfa4f0dc7f02728e2922ecd83d36d3cb3a0cf45ceae82b747aa4db17c66ec0827a24324002f78190b24fe586b1ba290a026384f1460fac31bc0231ff11418fd01f5c42cf8efc561f6a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb9ee41aec1a785e32f62139c07835bdedc78852db315c5b8471291f8198ea6688cb52a557de9cf1f32f4f0effbaf3ff2aedc3e22d2340dc346e8ee052437b20af356cfd365d70018432d1f3710455009eb6a9e477843f9a71daee822ab6a7c6487478df9006576f13f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1da4ae5ce83213a5ad3eac7373031b10f24212d24b6f90bf79f29d728f5036296fd0229534f3ea9c20253472d64a8ec04ad49a5939dc962e577c8ad663aed4b52cf0ff172c0487468ea0290e64f6d2dc3c2d76a54ea2ec7719450d66f2cfcd748eb87b0b51ea3a3441e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1384f562837555efe3ff16882406c4839a631f6ea90df59a18e3f407e4846110d78e37f6d741d6cae89505f445c2579fca09c76fe421f54899a9a5af3ab4334d51096b1827db54e5c33e908dbb4c0d1c4de7e6ade8db79dd2b500382f737cd89b0d9b2b9c88fd5d4aa3;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h4e0686e5600bfe457a493c194b5e963fc7f252293f6075ea64232993273cb4f3167d9d0694531b019016839016a8d9aff7bcd46570423fc2d1ce5aa2d70908fbe43bd80e05309a4188befd498446f6e69b06c330ce08a7b8b3697bc6cf2f3dc26d563e0b83c58bc0d5;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1dc19ac9affca40c3418e19a22a9e4033435fd0d585fc5f1eed48e9a136eaeac9b1a179f1386cf008693313aaec7475a001090c7b955878caeccdfe9805791d264c4a6ae0d8a85025b7421d2c044f629f09278f2681d401697c3c7b7d1b9bef3625a1c247b6da8331da;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h15e68a9761fda8eaf7b4d142fb6099653358908e2133d75f0b424fb321d33fc07ecff6e568eb2662a22bc6566c14b501201521fd8dcf03e1babe4aaf4241c727a74f2514525ca9a703192c3c092811596bdcbb901efcd3426e3ce3ca1bef1024edfccd745f4917ec8ba;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h6a137468f5a9b958089f3ba960ae8559d8f343318622caa7f3b6c61115f613158554f9f5da553d7a7588ec3fbb94c4f786183f6ae68ab14200feac6b8e8a46a2ae84d107a30f1098f694c2088a5d7d73826c4ef42ac763652b77aa9f02e625c9c148feaade47b0adb3;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h15ba8cbbe970c679984416c99004b271005b45f4d17401573d086096352bf54f350e607cca4a3432d7c41c32dbd310bf4ba17a21a6939a183a08924a3dc833b7d5e3e2d0407444091d8858261ebe81cf7654fcf5d58eb2999a7f341535c3633d5c7402daf2dbf5a2058;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb10b39de174c6b8bdd72fa2368a92904b1276759d112a0a08f24ec897fb929915f8804d5c9246f89794487ebd36375051b8ffe874e5c183ad16a75d76ef0dedec1ddcf42eab4d8cb4f0f8288e5c7dd91209bb5448802b7e890dcabe0dde99da8705cddcc9738930dcc;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hfc9e253462abd558cffad2190b84e570a14e364d5c4d7da43a61b61fe8fcb81fa7930b689198fc18ef728bc6ceb43cee31d9d07bad8850b93265d766bd9256f9da7c42d8025dc3ba8ca67d982fb924ba60f1a27a387b0b5d58b366581297c098c16afe99a6c0ed0d5d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h15babdb31a19f0fb2be172e9de2cf81164d0a1af59750d2997d45bc9cb8b6e30d0580ee80a34b8bdff558d700d3c7adb565470e67723e4408b4d0bd1fd8525a97fb3e48149cb55ba5ddf63283c5623ade8f2a2d6d9f6503de233551e3f02b945fb21c2102666c256f06;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h177a8a2261f9046db9b6c14ac89ba7e0c0bd1bc6525209bc074f0e09e1c6b264160ecedc0a82c860a415dc8d15350e312e45424d9c5b59a63d27c59913253e03834097884332eed08b9ceb97755826c10110797c9f99ae7b354cec8433fa4c5d26682968a07f49acd39;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h9977752dc6e901eaab59016700bf27cb1f5fa22ae0a725c70badd38ce9e2c3c31abd1bf2acbb0aaa55450628f0267213263e84c4a1095b686358b89b068e659a46a87cb92bf4d0c2fed7fce2731335d39434ff32f06cd2422da09534e797d7b71fe1fe2e60a7c9528d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h3f526c569576d6baa0c76a68887e30509c8f0911ef6f40628c9c7e5736896c12c6e13e2fd488b3a2ba0253af44b009c0f1665917c0123bf06efe5f6b4f15d67949a0c5d8eeeb601d5af0aa50e07a18e9544cd45c816371084d4d087ab9860f8f5a6728e3de3433921c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1aaafb822c3d764335bd53cb67761bcdc4f138fc89a18d79bc0952dcdc5ea745e74c13137b3f499058deba4fc2c991848c8bb00fda90489b4e61202aa81e463ae9e8947806edcf43df3e1b1685551e093dcb9616aa03864529f723b357564f09067f5dd49ecd267cb5d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h76d2e064f8986b090f92aff6ca3479a5f1db8370fae974f438bc2c5979e25640016b7d7e2bfeddede06051a71e6efa224c7233f89eacf4edb3f139da0ba31fc0972d76bc540115562e28bb25558ba7490b06fc898a2c5a7f4f8f4e8030e8fc6697e3f5e32f3dd9e9c1;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c7988ba90861fc3e4d57008ed1d77f7393a45ac1ba42b2aba0b7acc21e0a5e5a81332b3ec47052ae39b0da5d816b35c3ee9e9ff897da261d90e1a29bb528c1c926f870a0fd5ddd144a06b7e27d783df0fc46d1e8c20b0aaeeb7c5f68eb9ea610c7af152a54a4d05b39;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h142fa72059fdb06443fb40458c055ffe61302ee5c9ff7fa7921cec7809097e293e6e19bca119dcea8a49398e69a7231daecb83e729849838ec0f225530161ec3ba0e57294a51628d1e347f3ead7b476553c9bf4e9dab58cc661a788e76d0015247bb086577d1113e4a5;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h25905fe821d42ecf53d3752dcfbd5da25367b028c07ea4924de97b8fd4f8ff0639f6d820ee84bc483f6e2e0451dd9c981f9bc0a9d4415382034e3f9b6e894e87eb4c4ee465a13c7e2b0de5d7c3c046dd9adb270b62d5a367e5235c42bd17805280f5264b8f4e06fd01;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf7be1ba81a5b8297bab946c9fed3813ba7e0da68f6545d720be0730c76a238c9a53fc0701132cc901cfd2d18816172903adc69c9d302dcf36cacf7b0ad6f5c995f82fe7998545c1352f4252bccb663ddaaee15d3775d97e5ba2d3efa667d25808488a4f0cbd4781842;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1fea38fc2152597f31a5a180899c696d056ccf00e896a22779081f15dc9419d32e44308bee4f94db6c0470ccb5817badf8b7c8da76295fcba08ca540063b3cc4f07882f8d1228d1c5e25ddadd4c93af87a2101b27d7a92ca9a86e547e2b303281af2e226732ab4b9767;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha56710a4b34676153bdf18d65e0be64289cccf3647d03be2b8d536423c5295743e99a77a690dc9cc8aa139b37fd46c2835fa08149e3f8136878bb71ce781db68206f4b24f68149994e7aac3a40868fc77460b7552cbb6c6a9cdd7d9a1a34923b3ea5d4374b14d94254;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd193f6431448ebd8b912528f6adfd38984779212372c48e2e85874a95149ee5c0e1ca7bc4b49d94cea3e86aa18f054c766122255579bf00631c9fd655513dc182dbc7f5d945968d4c7fd9e12322238c375a77af4bd3636dd4bb6eae5e123c0b870a2e9b3d12bd11fba;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h3568ae2209c39fa6514ded4b86706cc8abbc4aee66bd83ef3d49ed3a8ce2259880ed02b937aae115707434c3b25a81662d1afd11e377b05efef8fb0ba023b9de6df37749a9980542541964fc549d8200ae1850716e2a5512b215bb33d37b87e587d2e1235bb6ecf991;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h29b77c872bb31a89d1764864b4adb1ab4ad2e713194a0864a11afad328b4ce1b99f816304ad5c2ed1ba72bcb4dbc786b57a17942069310fa85f527602f70d76a3d1f12288ae896ec244c9217dddc8b153047b753c441eb21f1742928f3804758807c24703e007c8bc8;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h151bceed9d4f7cc063c0d91f9d52f19cf569609ec9f21ea858c009d1c85672f75429efb9e67e595f2c16c090f793a20b878e773fe1c76012ca83787e470b9dbe196388e55325f087fb95829edb233b0234df1d5b14517e721bdb921ab30773548221bf310ad7afd4f92;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h27ae79c15dfa39f9669d674770934058744866fd3623465d5142db2c655a18dfd4471216d6c3f417aa8da9e0066a4cd0907e3d665cb95403df384d5d5b575b95318ca23ef5cd23b56e9560f6ce17b4395c19b21883701dae24b087a9e6c4cf678701644e7a3a163dcf;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ecf2e1480c8082facb8dadc7f43cf5b198ecfbca04e464806e7e9ef4886d6f3dbd13c8bc39f04cfe598db8cdc05380609aebadd6a6294f28d1daefd955f537a56eef6b15ef1ad64a90fd98b60d7254d89c2dec392a207e21b1c2ee3abc085920f39d8c71ba053d5c58;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h103514dc48f27c0d479674413e3b6eeb0d97894fd1935bb6abb1ef7365014ea969d9b6ce25715b57e9c224b8d2d269e3f01948d8ea5aeb0970f9470ce632386b369a6bd65ceee4d08142a05bcf79f8d0a9249fba3b780fc217606b8b685d6ec1aa45f77c56d0236cd9a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h16c0d8fc7d62ab2f5df76f87f161fef29c7032567377fb564f8f61eed428f853d62634cb5d0530946f466d451bfbbb7d435cb245c48f3e5acd0f87ddddb3b7f373f924714471c4883d5c104819ec7af5d628447c32cf10e018fed7f6a71aefd5ebb42496b5d5f122434;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e815cd35c940107042e191731ca36f017b4011a6d9f508fe51a0fc74840ba698b4455253c9b97a5b4a53dfe22e7c69fe03376243a1a383f505a893343489ba0daa7a68b05d6c3559394c353872ed27e5fa2570a8ea2820bb74681febf3268e212c4c1288dc810bb843;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h19bf79d3d81170d14a911791fa985e1c83608896c15d8d9782396dbea0b87b5928cf928022fb54b70598d514ed7d83cfa4bc2e073cc378731fb303aff818a40d09fd759f4c6100dc4897c0000ae0a86c44ee9902bf7e19b027b33f77c75c415efd2a255f5634c1262;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a568c90bf410e38a1e6e8c075b5e623c4a567a444841ee3f298373162aba061034060292c1837c322e5d34c9374a63e2862f41d1f6df8c9636960320175a5e28c954c5df28fc8aef21c4dcb74a7d4f4a0b26dce58bfd6288387271d8a90fe22f679334a69491a9964;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h61fd15e0fcc81a51bbb86ea6d23ead9af71a47b412960740e09340732e3b70b9e208b5d27a52b460f782b6ebd43ba471f4c6bac80a2371a0928de76b3966b94e04aee7965bc4614cee0ad6a2f205a7aaf9fcf970276732cd4efc254a0c7ef2e7e184a456fedba37203;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'had07e5b6f662e58075ad14e35d31bd36cec14af38066ed3731a721dd1209e7a6dc6834335bed1c22a40ff6b43773df800bf3238a26a124a7d67f4114ad121bc257343ec266c069ac8225a570fdcc7ea26c22c669078fcc14db97ae98f33447ffb0dbc0b7f124ec4fac;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b864d14f26b24de0a2ef3b1203a8b3c4ed0e15f32b85db6a027e18a46140d15def3a9023722359f871ab7c8c85d58d5640e8291eb9f15f063fdcc72f7d6e86e60c57d292eddc40eabbf92d8822b3a1eb91db8a586da93e3d07b06969eaf5f873792e65dfe6ac0a9fc4;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h12da8788b0e3bdb5eaf816d35fe22ffb9b171175531fd6eb3bce1dab1741bc0c6cd5be49b733125f7916f6f42b66e65279c57b1df7b8af3b7dd7ee04eaea5b962d7bd0f61265477fc7970aa1e7bde48f4a5abf306c345e4872f462df91d24077fe9930f5f294c542ce1;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h19a6fc5b9a934b5ce8103328fcaf857c5e243817672f022bc507a5f5f0ca017a6dfbfae3f1c48f161586f7ed7add602723bbebbce332dc6f8a212bc668331036b585e230c2d9c084deae7f8ec49af6131b081e4841c716265e774091325769bba5b2cf1f35c12ad8558;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h14feb1059b6a777280f7c800e2d5f68491a8f3d3f520595a5b2ac4158ab8d9aaf54e180df28529f8e37bac190b1acd83359e876d5bd91bf4f4ca122963b758842ecb97283f7e15cc10559860832b42df1365dd71deca113fe2ff73bff58d433c8ad4e215e8c0b98dac7;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb17667444924719300100ffdf2edb6cb35f2e2556a0e3ac983219b3bb5e47af400cb28cec6ddd5329ff8c00d7971152e6dda50218c3604be8bdc52c6a8bde27ee817ce260f2518809b13b02b46834ece62d5ce68312de767b95734a9d36f24438d583fcb8097f8c8c8;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1db81321cf2eee0bea05fb1ed699666ca53b02871ec50a1ee15ab86d3652477fa401750ddc93e15f2ca0c359ca15383ef7318a08d7ae36bfcf8dbaaf3098955e35b3bfb49636906c9f94567509565cca84edb22b28d069f51f6cc02d01c3a1a8bac01dcc457bd4d17d9;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1324fcfde5a04a3a536825e07782b072ccdb8bb8df79a27eb915a86a597637902420f116f1b7bd3bdadb8ceeb69ec901e11d241ab644269c166ff158617adad660bed4ea0a524ca161d2a57ce6634293966db537667289546c26626dbf883a281495c148e5b9cc19f63;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h618943118799bb28405160b16c65f9be021a5f674323b93de83ce3710aaf36a36b8e66cea4314ec2aa44c193b0799977ad3df44af9c3ff69ed4e51cd0bc151fb2eacaa065c76a6cbf3aab1240b71eba95114fed1baa7451c130431dcef840d5cad92498a5de66e011e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1dc226b32179568e86081b2489e16f1d488314b30285662e7db95f51fb90d337fde7733a4bcb6d9a087d62e01101565235973447c8e42c6e9874f9ee814b697ff8875deb041618abf741136d95382c15b3771a8875827cd13a5211633b7c13b7b6bc40e929978e14157;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ca384a49ecbaf5c1613f78f6887e685ac67c284cbb2a411d90300d328403c6920b7a475a6204373c131645ce6398bb9ba8be674214964fbbd44faadec52e773eb47fc7fa85752bac2bb7378a13111f6d50aec6b9926d85c5053656d4d19deb27e5d7a019d0b093da17;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h466ded5d55bb099fd541314f34c23062e765715a2a9bd6b5920fb0bb007cc4c2b64922b50c40f8ad86c238c25393b384283a39de397286f42fa28ff3656807e09a4cf7dbf7f4095e51bc6eb756acba614e56d54d5a2a72bb38941de1ef8ffb1ee6010be97d789c383d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h5808681e0b3787c0c58563e48a1d2d95840fa20216d3458b5858fb8ad250cbdd5f311c2d92eed867ef930b1daa813820470fcc46960fbb870137aed32102806bbd32f933458b1913ecd59579f86d494c41c3e43df392ef671d49c445779163a2fdd88e38d7e95458cd;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e21e57d2d1f5f5b2d0add92c235fd60ec1169aee881316b663b75ed8299168c3b5cd2eac69265e3dac1363fb83f42c3db9d76a2b8dc8eed2b3d0151295fed43cde03627c446116ded265c6e77759d5b5b423100fc2ff5b5c064537207b9484e55228279bef24ef581a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb7db55bb4f7c6ac1e5db8cb03549a094cf00eb3322f6ce0a216830149ba03a78b53e29e9c205c30064152802c245f5aaebfa94bd5686546da34a67ec474ca85ffb0197c5dd13224effbee0e575f069375e47c5baf64d9f079303451068380000fe284ae46c4f99ad99;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h155afe1a972eca15b2afe64d7c3af3cf32691bbe2323b585bbbb00e490348d719f24af28b4bab9b79ab2211bb0e5971a915d06b8a6362c27de174ceafa05ebbaec608cdadceebfd6cacc5e13ce2442c678a929d3769d5d779548494f6daf13c203463051f9e678e579a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb2bcb6bc42280fd5f7ca8e80528c42c7e3b536acc0363108ce2dd39d5d724cf126080b15bda8423ef5aba003a47300d6ff89c647ed2870023587d13b0678c257919067dc3e54a4d824ae432a900b50afa0a972b2ca089d3775f928273c102b44a3d343a3e2d457b029;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf289e9270ac47744d2666929318b7b40b918a5cd90debf156043ca0714e3c0158afb8d241f466816f51e5f4b38451d89aed995e9a355791660d1548fe5cde3502b2f96928f1878b63fd46666054e94e6b3c860c1db15eb90f4fe1f1528ed332887d6dee3194885d289;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h47199da8d007c136a86afa52982bbadbc5ae0a7197e3c64d680ef8479fca7e54e852b8d5b6daf97965e50940c5c43a4ff42dd853dd58026ec9664d8994101ea27b444515b37b2ea4b8766ebce5f98a6e774f2ecc6bebfb824d8c1769a27823906b27361bb2de57fc56;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h165c9e074eff3689382894b88af8b8c31e33cd42faf748020886bb377d737dc3c54120ff3c323b2833f8ec4f48ecea6f8cf46c1f8a6f9678424cf15f5d7f2d4a56a4ca31de0d3db0caa73c954d3ece886255281ae309d191d7efc8f86533fdb1ebaa3c6286e4da9e8be;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h55776a7e1d1d63e013b854097b8db9c92a80e20555030a90c08fe3697fc78bde5d2c7edb4305fc8aa2bac49a69cbb9b85e8c71418628e8900ab2d55d1081517b5ea821ae7cc8e51e16c36406df3c9faea2f187b4c8e41cec1d24d1638257a93bd46ac3e676b1734ff3;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ba9d8600a44148bb9fb02053c8c2dbf7cef206a3e565f195dd972beea12ae2ba4071f72748548338cbebc62aa806d9b13fd9c5d117817cb67ca8867f0e2e77688b777fff12a681bea026784515e0e2c78de22e9277ef4fdbf4044e20e1d3737145cd0fd06ce38e5593;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h198ec596e57d0c4c3ab81a9adefc7e35ccffe6462235973937c6bcca118e0169ce9c1547e454db02169303d5eeee111b4cc9fffcf3f87109d0f70b07c220b6cc72499898f18b1bccf5b79ae8fe10b92b0f705934f0944015cfdcdfc9a19e95e0c30210d59ec881ed9fa;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1aa3cd37d20886b1da9956d8baa3c146be96eb04207996f5199333e67bad1aa3a33972679f5f578a4a46c27f054205aeaaac0523e82f37b44ca7ae2a7d39f35e94bf14d62f98772e64647189f26bba1a6ee4978ba9fb7dad86eccade26a5c54276d775e97431c5ede82;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b1072f40b5e57f20aac3aeb1cf875af9d822cdcd67fab65230587e5add4a9901f52f99c69320d9cf4bd0303d8218d88d7f283c2cc69f90ba33fd241285cee65589d839b31533df3f55e2b6006a41c0168e524e934904e707b822a689f1fe45e888313fc39049edd034;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h3745056742fa0a16fa1061fe6c0b9cdb016648c6c54b328ca7dd86d8e3e4a3e7c70c794d86660b806bd014895947836a5cc5a54b7a564b12f25e5fc74f4b9f78e0c9539d76010623ac2efe43ff5d433fe20a2ccd471aaece406b28c0d96b1305791092fe310b3a3194;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1deefa897afcebe95894c9aa06406c74067d69a0bdaa01883714cdd3dbaf599ecf55e9eda0cd2588814bd551fd4d0510b65ee2d89d66d81cb62f4555f16adaa84f870f3f284823867afff52209e322c2e59044d2eb489f3c55851d1e01087d607db535ef70d847af4b2;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h197c91c74c11f632468efc7dbcadf6e41c8b2efe2dc6a30a5f06a15f718ac71d6834ed374758d4b007636f8c13b7317f2efb920a37f95e086d6a71422d86678cdb0e9c617f3c9b5b16534a50514ae4a4a16c2a4163bc9408ab440d68125a81ca0d89295a14aba6388e5;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c70ea317fe193e4943be52bede102718f8b057e5ec3237ad593d981aa4cce38b05e861ec3ada8d67f27d270573365a8c9355fd4706b26cdf7affdf286542b6e82d1b01cae686dbd02ed66adee5afe6f5e5efcd510515ee7f70d2fdf208e7dbdb98bc81b139d5fdaad0;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h5ee8c3e027a67cd0eecd6ed790a673dca6cbb115fb2136362f5b7ef63012282dc120f1472f98b31f085289bd9946736a2e2db6218e39f462c058bd005256102cf889f135a90749294f56a2bb1def908d72778ff910d361d6d774f671cb81e4da89ebd545fd2f75fccc;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1db498fca7db7341d4d13250b6ccacc9d22927799585cba9c914d2ad383a00d70801a7098a33e1ead499aa0f37aec55ca9de1783845056f1c2f95ea4db5b40ac301044434492648c4c566a0f98682b79a901bdc9276bec979d0ceac15d6a92adbe68cb69dee6339239a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10837a932997b53d4e1d670d49885bb28ebbb6b06c550109737709bdc94ee175a9c3cb44b1d9cf7b6b5ec0e06b83277037952b33bb5e2321aeb778be97b2cd3d0287296a5297e39b212e36b371aa1c5a78ebdd6957b29b5090e6907669c9188af265b9bad3404f85c79;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h17275d4b68378541bd1463bcef55eaa9c10696cbc06a8604da7ad4c1825eec849f8f09ef23405b726828bc1047727b081aa103f6a4152a0542e7edd78b6c0d70ca93fc128292326ae7b9809138bf6e32462d309fb73ade030f82c44ef9fffafc90dc57e63f5f0c68543;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f0fb3f63e0a21a098d54f1a04fd70d9e83fa77e0b46a931d179c85a9b5b535cf86b2e3127759444a1b8a5730dfc25ad7a73481b7e35ae7471d94cd250030b6b0b75e8db5733b94b54564aba170b25033965ca0c709df0d2fabfa7989937686fab3aef17df6df3a2066;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a06a51ce25f06877e7effd288626b10ef97d0673dbd63dfbc08b3a8ac55f4c3b8d126de1cc1e3cad993bb668994b023bb70c637457cdb416917903ff2949d79bc3aa299c10fe99f7bed7573f24ab95f97402908df3428819efbde9bec0f5b2bd0df77bc30642db5bde;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h12515f9282baf73eae875941910abccf278a9a15b4ec5027bc3009418475cc10e26886e8afb83b08c78afe09d1b975fa34791ae620d68c0c384dc0d8da19851e711e377262eb88ea8de2a270949eb385e62f74ec47b21964506fddc4369e7be265e4a566f9e810c6653;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h4bebd54f548c36254d07abfffe274423e40ebe10dc79f3f1a2a56ce851885ff5709fa63566875e412a7b48d93e737be653eeb1eadcffbe1741bc8790d3ddc8f3895af46990fbfc7d5a455e2e4ab99a6b1d653e45842c1a8b3fe196a42e6fc588c77dc1d119a3b72a82;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hfc0e2a00aa9115ac778622810b792607e5da0d05f85173af81e2f062e2d81a8b76e1a3f4bd8246e6778802df4ef1a70e8b0ab8e6b24908d9242c6c54025cb95fc92b146c56774ba4e97b3ce96507477011ef5b39f3ade054a6c794527f439c377fc4a83c4d61fca5e2;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd9b969c6060be4dadd741ff372bd953f88abb52c2f4ce777d18ebabc25ebcb957910b9099b6ca1c6654bbab226b5dd74223ba8b6644cff1a45b387b78a90cfdb25f4bde5c092165b75c359c8dd02060f7583e1fa590b58e0fcc07a132b401f08d8f428c51b803cabcf;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h15725dfdc1e3d9fa0ed006930d5e82750470cda8ecf4173be0da2cc2b8761f9734661197df291cce480df2a7881fa6481833c3ba61782687a1ab06b34b4d98be9979d04ab62197390fc7edaac7446faf68f275b68c44819f3cee9ab92cb4cd29c6b29c427a48a1a33e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb608457facf776493284fb9518fcb7f9b90c266463c7f9c75fe24ac60f72db54500110fd4c2cc7a41bf3d9f89660e9de3a7b58070e3cfc71a0ade28c01715073f44e3f8a9b2db681cdfcd2fb4e788c43649e92753846994216ee710eed0ab2aee4c23e69176a2897d8;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc9f685a2ab8d204ebdcb075970ab9ed91b39dbf59557cdaa7ed90a9b0859a7d842caac00fa9825fb2292cc573fda514f2179c0ad5690d3e967749413bba23b83d2419cc597e3ac6b2f4a97d6c5f6db080edf3d60db7b3f36f9c7babdc0ca3a536c10359db8206c0fd4;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c1793489205e518ac864e50f3ec993a6a7ed81ed6d87857684cfbe917dc96e4b5adda482eeb52e7e7f3b72a292cfd5cec0c98e7c8e4730b43bdc198617f64a28bb4ac2b8844a3216c9f9d844335c9332319e47ea3ef3df0bb896f1658b66de691ea6aad9346d6865b2;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e40c40388554998559ca3c339f45278fad4392e6f89958f220071629b33e74d125fd78db84371caf718c661f2361291bcbc9ac9358d4923764c4b193fdae77c430989c700dee8809dd04146be27962f3c1c6a05086c5d48d7711ca25961904e5747675e5790c4fe30e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1390dfd880ecfedf2df2266483a2d550da2e05b45fe7470dd30b72ab16060dada971d477e295a2f444fff965d3b24313be954888ea18033835d9fa60bc08c41aa1e066961c3dd1c0ca90414203ae6acbe42c823efa4034ec17b44fd814e5069ea61ad7224061b6c5b0e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h12896edca9895e3d2d24050915ff7775a37acfa960cf631cb4c09686a57abd53d70775f7bdd2adab3370a630d4fe7275b2fad0a579264d3e76a7b987549f784e888fc67cd68258c570931ba1cdcb2d69389f4a5e2e4c794fb90fb0bd68a946a7cacbf92c426f0143bb8;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1911f1001087ad39302f364026e682da6b5301bab3945bda8b73db1108811efa536d6b1f6ab425f846cb3eefe1590655d6e2bdce68c41f7d8046e7896f14172b46bacb23e1a85f9bc09c2996cdd4aeb01b6b7f550a276a80eb20aaa59ef7e3e97522bc8143f23e0eab0;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb01d72299726459189411564de65ec233006d010206d34e96587ceb4ae86af69e224b1ff3475125d0d759252d2b90fe63a97c013afdab69e55c1dc90db44bbb58ca1c774bc953bd3bf3a849d6494f7fe7a907772c1005bf992179705603a1055fed73013e339e44c28;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he83ef85cbe808ce4c6a35f1aa3cc87195e9350f3d62ba08b33ef512fc85efe27ab710f0bb4951c30d119b5cd6136aac53456ab681a6bcd8aed56b1c238cd8c47c7d07d656e2a525f2887d99fa355931e819eb871a760e0edd8c0b9edcf9697472a8ca30d87d1281ccb;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a8d728200059e04ab964167f625b91b72115fa7978c02cf09b2bc1ef7aa7f55fa7e3f1aa36fc599f4f9189f45d617baa7c889d4652c38463c4ce07a90cbb6fad496693c09b5e3784606fae4e5ad05be509509e73ab053ee7d0ee60b7bf5254b839df6e897e5081ff06;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h4ad9982c0c1537042c310af77dc93c474983094a61a86550c022025a2751ac556aed09c9f2ddadf9ea874583dea4fab94c6d38422c01fcdcb5500e3a0676e454f1962ee7824625a9c5d24276af9dd4bb7f8f22ec33c79d17056a5118e32e77be29bcbf8dc24a47271c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h2e0b87aa7d6fe1f61ed6eead4d4f4bf209fe8c308627406ca4a46069a17dc990267a041490fadbedd8c21b873466ba29dba05bc4d51d0a568bbb8e09a0a1f5baa05aac9456f651864af68498125b16bceebaf32f8eb10fa0899218e0645ad6e1f4aabb95d659217533;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h17454c77ec070ab3d4a8143f2cfcbd225a9cf9f14403be4071ffc8751bb7ee9d54f888f5e55ee0fe82d1d5a1e0fc32b4f5b5c67b38181d4e0cec568c9f315e141ff3e707f305a7748872edc8615e3255a12aa6a04315fdd926ee3fad4de9bc079d1f37f54c0a00a4186;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a62bf5d5af0f9ab6344cd0441d0e847e39e7469cd23bfa11935808219f475e941cfd046bf6d18abe7f9bddafe02aef421bea00d4eb03a7436ab3ea811932b57a513cb1758aabf0bf3890fbe4f293e98be6dff5dbf6c1aa74138f4bc769a84adccb10244b3ce49bddbf;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb7be95582bfe1b8a1e482098e5f5bc100dc506a5ecc3353b73691449d9ebc637b5d2412292c26c8193e94b102249359ab562f07c2eb7bbb41a1e74bc3f55c3c995fa45c7dababfc0c9c68cb5102fc6445c83c863ab28bdc4d9ce092e50c5c18f603390f0fcee01dd88;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h134e769031c8a6fdccb003fce25ddbeadccbc1c8947d125a235552fd7f7cfe2f590334c0b4e22dd8aaa613221a31b0179bd5ed04e8f79bdd0f04d4a25a853de1c17ca570af52be12b68058be6b11043fe44826851bdd0f44812c7475134a09a96294767af4c2df53b89;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h17c911038e0eb860795f63dc9773d6bb69f550554f0219d454fae8c685c4bfc31192a59f87ba8e4da918f116a540b08810037e3d876e59ed3f82e74ab57f4f01505676bf98083e6d744e9892fd7c4fb08ea5aa0e6d55707f22022880ed6d164f236d45ea6c61a6f6fc9;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h18a052d3022490db38642a6d3b51bd7e1ae747156f3e54b60a7cf85d1216f7f12d8904ca6243f46ba0162179eca2a32157da7c82e02f032946ac672842b4f3b9771719c010ab7c11972ed964133f485ab8e3f2a6a27f2910b12801234202f7c0375fb0b963578953909;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hdc498e35e7f801bd4f2d3a65f0c58d21af4ec2dcb50a17199a9a1a247bd8bedfa6e4887e258780d5cce36c171df00b888f6406e20899f1acf1ae40ce459a9ae2ae6cefdbb4a703037c3da545288c3e6d0fc071033055299da6f6f80738ae782025b511f2637e85cd36;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h44b569587a83a00f884fab99a31dea0087dc8c8d13e4277c1b578a1b3898a5efb12c77951605f9c215c92424f7963348ff0588812685d3586b28316868159d5ce2046967485ebc62a89b945a18a4edd022d97ccc8d98a929550208edde19d15c9e1145723f8ad1a467;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h4846515e8c978bb7ac1626d90fcec51b6267fed110c603162b60095f5e3d64f40a7e9537dacc8d1fbec1d7463271d9963c4bb205bdbe1256acd46ac0965eef2409cc2bb514d8df9131e7f6d8ffca51478c10a6a1e906789e32131f523aa7e96a2091483382403bcdb7;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h84ea62f02c1c9130754809dbcc835d454276a78903880fa425fa84bb57f139443342de5a4a5a5c7b7a207d779091d75ef2376039f87193b0738042cb6741100ff2b51f90812ea8ab33f6ec82ccd8d7016d2c61891e388927bd441553a9e49443bb503e19dafb56f6d0;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1847b595a20279a0c6c33d0adcbec28e7e03c0d551afea3ab58df7df80c204b334041b935658abf964a72e5822c36a3283958f0c9bd19be2ee18de9ea0093edd186fe7e2a64ca5d4d2c4722494f126ea9b98c65b5423fe1de81ec1860ac4f713e00a773c342957fd333;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f7133fa027bb82b5eee9c3359b9011f7258dba870d204c525bf3e6f92e5e2e06013424351a3851018ef2272e24f03d5a6841a1545003e7de4c4101f0a9e8d9ff1fc844d860c99345a6ba692f23454cecb1e4acbed58f686a782dc905b5c8ff1a4ef5b9e42c97634a45;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h52eb5e51e079c764da5ad7a3bb75cd69a7f6326bc1c1de8a1c5dabc43352b5ba80af08755494bb12dafcf5ede258a4b934e46f2bef89725832bf237c0015e13c6f7c9675951fc892a407a2bbea87e6586711ba14fad6b4730121348d76071b01c29bf9a643dcbaa66c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'haab94322710cdebd868f771a531dd94db2a204db710732744fa86ee46070a62c58ec5c925e3f27ade3dea63e9442a89662776ed80bfb07667952753101a5b73ae1f190d115d7d6c74796069cad4ece862c8c0896d87f489feae2a426507183f8cc9a07bcff1bfb89ab;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b6e79138a691310f4060bc8d09d2824a7062553773916d5f59d8ca94e96d038ecbbc6a1d068d28342443de414073260e42116eebd9c5dd3297133c5143ec6f64396690d67b215b1a36151e872c6e3d7e6a03cc8b997827beb782b4f8a2b1a9a407ef14d82d044a73b3;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h124d5469717dc6175a57f4cbb5c196fd27dbdea28df8e63fee34c8d8d4a28399dcac9a380599c2814210298ff6663c19ef386e80744ea5f6f76482eeaa8ef2ceafc8168168b1cc6288403a2289ecc9fcb903b25c7114a6d6ee121493af97568c10ce3a68a01bc445836;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ac668152230e4ced6cb314389a08faaab324d2ac9dae3c7153ba31d6679f36c4257419af44e00460c8fc821b0e9a2d4598cc0d2d5e963861339f33df8c649d4f05d77007092434b21344b157d52a7f3facf731b226a1c48fcbc11e7960c055e1a2515f5315352910aa;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h197ea19fb2301236ba3f47ccec1b9aa000d3dc0d13c086968a72484c6356ab7d9df4678ebd22b179eb65367c4bb98364099f2177639199fb18f8f527dc5adac8c559436a0482181fd3203656d19895a64e5986723e63fee30dfddaa00189eec518bfe99c429d6e83ff8;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h158132e6c45ee88a8286811bd8690d0dcd46dc129921e2b3c4219c2f9aaeb45d4978c6bbde54934c9e27adc70c252a15a943f777c724f0a79e48b768f36662108abffc794ef1fb7e17822cd5c9311fac4d865bf9b0548998fcf0cb2dbc27e26eb06a69e2e70dd0e65cf;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h7513bb2b3aad30923bccd5b999086674a4ff8fd3e8817326aa1448307e03c041a993408b3fa639746ca74da6edd590d8acdd23071802cf64a52d0efa96b40c31e02b5acf70298a6c2326d00476dcff1999ddae258c8cf816d32a9268e8e26acca8f1f7597c3c3d43bc;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h888c0ccc221ef54e87f3e4248c70d97e59cb326df5f64a010deabef33bfa0bff811a97d155f48638bf6adc0d2fac87bc631b298a8f1e8efa6454a7f7207a5a13f4aee10a35f3acec541720b6c81741e6842ef85f5fd81a2f090b4f5bfcf8c1381af8bf7646ae9922f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb30dcd9b0ab2213f9257c8db06421b3c4de0091027d9b2e4d21a8fa9ff0e471e683b7b1fe45b7d4c11359a91ceb6d59002c865147bb6643b4cf36fef697eec2fda7f9b1ad04e1fa79b7e499262942f1ae449ccc6f9dc705d90b264f3db806f5629fc1fc458ab15c7db;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h12b2567cd2fa8f3538d3a18b77482deb978c30617aec3eb4dac49093256f951424c1de21219e7e0653f24e22d8c4ba2bfd22cc0e2bc4b0e385dc790b39057f8b85657296ac026fe7ce4bf4d4e7e45493846b38e73a775d5e7369468f6a21118a537d7ff0a9f3bb274e3;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h16673383193a1ceb9444837999fd6b17d500b731c5b3519c1c5f4df8ce240ce657932c71064b45490319e463451817c4dcf0af3dfa6586f7d5b87cc254b9aec76e1141abe1764f9e4ae4c1bc5e387ff971c9c15cb33310465296aa7af9645291f92fe0118f776b34505;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1375b55dc4039610c2cbb9e9124792b5d9bdff505b2c871ff2b7f0dbe34eb2376673b7f2dc1bb3be18c72e1c593989f67c4724b619a5fcd19c302e0d4c7f36653944807433130233385869e894ddd9ba0c94057ce196cbc9573ef472925e066202afeb47d331767047f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h4094fac3045131dcf88be2e2149288636a06fe79153a26274f036fee1d61fac4fd40cd0a371441ad760ffa9538fd44b6c62b61a8586c42903ebc2b3c3460a35edbaaba29e12b84f9854079246b27c0e75ae4bb3769efea66ebce1bdb8cc1b8dcb2cc3f1d61b1f6d4a5;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb3cfa071189aa450c97203298a260420ffe058c7bf094ed966cb0cc409eb43c00df7161a382b24dd40a45e6543a099c322b74eab6fae518e1b70effafb80a31406ef28c8857a956ab05efe31980763f0610b48b6eb2d133f6f4bd9a78692312d7470c056c827ab2ed7;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h2d1bcf622d50b4210b6bc9dda7a29329db8b4c7f6a9d83e09a4147798cf80dc6b9a28946f79cb2307a97f53ed511b9d9bb35c2254d2f320d5a04b35cf2af0ca13d25d41f12ad660dff09022d6f5943f73c7aa6683af9b288f0e0d92dfcdc4029ec6d3b353720b3174f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h2c7010a1feedeb2adca5d7e7959fe1c36a6316bb8ce39094da4426b3c7ab69543de44bc20721af27f207bdc87e84e50a3b90d0b289a7185dd636d0cec6678ad0fda346f72bad51cd2cbda2eb591032b4ae735cc1e2b4a88bf20c7590a9f2fde6e35c7f44a1dca01608;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h12203e9cc4bfa996d4d287a1bf8e2640b528b4def1efc0a00bc510e0d8c3ae9a6baa2d23d58b3f037d524b4b9cdf8a1d45878f8dcbabf1fc03776228208e82f3820225983db287eeb0af71b0019d136f64aeb822d4eae21fe3330d3b067d8aa2763e2d35f6bf580a7ad;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1dd8b8bcd7d8894119c5eda3d698384de3be21ba0511f63e234a17609863b2fcbe0263e3816a76b58caf63745c2ceda326623c9ea1be1e0230e31f264abf9e65e72ac4c02a8877ef8a36dbfd01e567ee3175d63f9302a800c4af962867a6a38da68e5e83346ce7494b0;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h46fb7fecc4d75f503c4a7c61d5f8ab66110319a21741c4b7d2d57e4f7d6688e9f4e7aa424c818a92bf870699c2bdf4f8cfe72b1d984a339b8c46c73ddfecf92b39147f400d0d22a066bedcffe80942d367862679057978944816143983430db390abe25f3f9235992c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h2b763bc003b75bcaee064c0d841b2be8be61afbb8bda4202b954a20121c46c8d41074ed4677e9c770e7d9b88318cd167c098ac833cd32e7260c421bbe7beb51b70a910bb617640ddbc3a146b8e1dfefb45182ea09e73b749629d5b42282c7b693e5648ead8c0e03a94;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hfed65e86ee068ac671fb7f85197f6c44fc097665d0ad45cbc5fba731d267574e6b0a312341124acbee062cff519378435e25ef45a9755423e467d197a9c12fd36beb1bb99c7a2f26bce62bb8eb8947c6eb622ecd9090d874a2064e86ae2b61d7ad8d4e4e29bd79dda9;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he0f3b5b6c1a82c513a62146faf4409a92483e441f2575242be3fe10ea737017d0f7faecc4abafdf8f703d92d63975f7068cdc6672cbaee03821de8b65afc400a4746b01692843b5cc14ac9dcf0d0fede43e99b1bfca4674c0eea80c62af6abcdd9b67de8edf5df516f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h146cd7562445000eb2f0eaa2af62b4aa00c3f3dd92db0a761659ac244b2940566528a0aeb09ab09af37512eb2a154160ec799adfbc568d7e01cc56539ff665e5ef102e15f20404849d58c897cd784120f10fe78b3a2210f70d3ac6ffa51aa29903f9398c43173064474;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1cca90ea1c61435578ae1bee64e855afd798da1c350371ae6a0f8da61d0a27031499d0bd7b3f8c2477c05142d146bd1269e08f3fdb1159ce7949953de007ac5584df94611aca65ab47aa6b29771c6009b122716530b86692e94697a6066b7cb1a153f14e87a24c9519e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h13697208c0d7922f6033352239df63a8a90572a6cc0798c0ea4dfc15ccf0e7af9b657340994e235b70306375c29eb7c077d1fdcf78cbe44ea2e69741d812b5130bad7ce6d3718c321042722e992c491afc029f15330742ac8020c29e7d5401ba6138ba97a3b59e0c3c9;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha74ad17c499fa92003f5cdd375f3300c65d39ec07a64d0d0424e31211e981aabe90e6c764be955509cb25dd5cb808fa5c0ced80a41ae0bf1399432a659e51c4ed9690dcae97a90fa1cc84374219c117fa5f4982ab46067d2f6081dfede8e509598941541f0367079b1;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1764ace5d27b085d9f39d17c2a47621b6f22980fec8c8300b0c8a983434cf1e2000d42d5ee1c6ebca9bc732943ac088de12c22d9d662388671cfdc73b47319e7490d2dfb70f59c556f64966c38a33467147aa94d9336e73fd7abf70cc25a05941fb9336ca61861f7df9;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h8b53eb60517b4feb7c29ab8748ed11c6ab3ee97c92a6cc63cb50323f2a66c49800b2f7b6d1e89b35f5c8dc47bc481be037371003f0867187f807c1cd37467f31a3064f97b0118cece0dadc1d47f7addd1f10be881523ccc5ad66b18e01babb36da6ed574f7bce31623;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b27c24fab2021c33ab6b63af9dc573f925b9f48b2338e25cfcb2a6ae37be86bf41d7bb1d2f7b9cb94e9ca75a40e66e69903f852b07f8d6331fef51f7405930373130d8f8199846bf830f84b44d2a9c25c369358bf971280affefb6567a8460e189170c20ac7cf7b2e4;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h16ab413efe5205dd5bcea0083fcf76aec81fe768cc4ca3ea417ba59354c9cf4d5f49c085005426fd679352e23d09cad0396c870302640330879cefa6c3eb49734bedf357ec3e8b8fa8418dea32f6919b2a7d7c6ac009654e9b007a056d1ddb14ed0465f22016d3368da;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hbfc1d64a2b00125ba2ece5b4f8aa4ef27fde4ddbdd6bf6717065b44fe04ba1e0ab3b1ca90dee22b1569c6e67d142fb46b988812e72051c0949a7ee36c2d78c7e09aa4d9080f35253b77c2ca1a269984b32b53c6c0d263b3e5090906b4c21062730ef90198050d3a0d5;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1dd9e656e3074df3487032aa429851007bc86becc2681ffbe823b3e279f334b02dd0ac9add1c81924039e6441cbb1fa80587b10fb588c109a2c67b2f1c2b11f9efb1274466636565b7a00fa34da96cf9b07975e34a5c4fee497a64f70c20cec68d77aa1fa17cf5b54d1;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h31c132aab47ddd14c4bae25d06510ea16680215ad2e964fbd1add68156e28f118d3eb6c8692270f43b4fecaa5a5cee66279cfdd7bc804e44a5911d9ce3fb194cba123d53f55d65d3afaa3f5aeaa9caee489342c0d4a6b3c4e1b6c8608d6af7e2dc9df821f76795231;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hefed43eaeb19509fba2e30df2cd53ec53dc15f5a03aed51bed03571f5cbb95416243376b4816763a2d0c1aa3818ffc1a372856057e7447aacf345acd1173d2cbf3566c0d0bbba51cef4d02719fa492166ac75d303164fa366a6a00bd3f239041f7a5df6c14d318ed1c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d07ddd9b90a97cbf91b15aa125f46da7b8d09b2574ea2dc809efff1e58fa193ac15f3e6777980e32e99cca5e6027152e1fd6789b33211a7176871989abc29b0f5e3c61ba199209c282df77f8f3a1f5c1326e3042bba249ae91488072ef5a63966647c7a4f9fb3f3b20;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h23fd8eac864038447b2fbae80d206af2498793dfecf3990f3a7774e377f2f4fac6a1003ce050753bbc5f99521fbc130d1ce864acb6e42dc3546067f31f6e4bcbf1970791f66c1720ad4a146560b5a658a8db299b6d2e61571e6bb0aa24b89d7fe024c78fddac7c3215;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e683b3a8ad471e405197e00faf09f0348c42a808b7993c8292dbc79a86a4598fb62e00adabe896b2d0b489bd7052f6f9d7dbb9944268983430af752eccb05b7dcc6324ce07cc816b599b429ed4306fece43a95d230466c981c8ce13477099b5c7661a6078f613f5dce;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b0bd4d926aa18c16724b5876559e9235e396e76b9de73959cd45034ab25fcf50b7b0129923b8aaa2261bb4e0bff15f7bad0e378ca3ad51bc3cfc0ee65ccc44e08a3704619b9dafff4a9b36c99f937a45b1e42c5300ddac417f4740d001b7f11e0c3ed43ded0ab4f8ac;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h15759655aadc1b1b20fff9c6ff3b5109209998371d1df38747d00fea4d44f74131b9355d04159a3ae7b863e183e59115d23a9b9ff4ccbdd94039819ade835945a03ed2e8e5d2203671c90db0d30da93ec528616ac7efefa24e573226e20dbeeaaadb1468e1bdd657c55;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h16a50c62662875ee5d937588056348428b8a247d3a44d3bc83960b1f594021394a7c500ce5a69b923ce8d29096dcef3b38f9310a9732b6fffde9be064fdca2f4c6c56859d5845e6fd9a4ac0317ed41e4f8092ac36bf52ddf4e7599b1126b134fcbec7f168ad6002645b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h14ccef1f29c995e4896fe61b26dc30e1cf168f8aa669279960317ab5ddadd9d4b80487880f3f53afe26139b31791c295595f991ee7bedd081accbe9835a7470a5adfb061344b927418fc27ca08895e878ef2965dfef59ab226a254ba6c34c94648652a7819f651b6548;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c11cf9570537c97653e802d4af44ea7a968d690c547e26c96266866509dad95801bd6a4ac3ab143eac32b2b8f9677bb9f49c2b74f14099a98e127454211da5b03e07f2d795d258b3a27f77bb1bac052f1af09abddd2e46c8b6e83b1d312e3c2da4c74efc7c2000474f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e07344c7a772cfcd7a858c4532651d28af2d390ecf6ce051b99c0d0013c490324c6d365d38a00389c2f8072fdf91bdca2a32a45d3cba2b5024289e2f2c0fc2b914da764c18dfe3ed8fe92210a9059231c493a02215578ecb89756cbda716b3a521b7930629fc0c9271;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h135d95e806577fdcd2d66631353770d21ee4d16cbc54fdd1ce80c518f5b6c76a57912ee4b087ca3c3ac227c5e4be36f30ef93288d7922835f11f5e89b2a7bf08e611a3bb6e539ce586453e0cbab87b78153c30f1f81bbe1f407a95f28fb841d2f5454808d098a79c7f9;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd2b657c18d5ab794b63d514a5afed6fe88b9554c48cb40fbb31b4f8f9bdef8c378ecab9cb193d3463aef88334c4ce99cfeadc90e810dce899c19b9afb86ff7a9e4c2f75f634cc4d95ceaf8607a214938b8e513871b7387097d8a8f30eabda40b65b4dd39cde404d628;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h444064078290eb5711f798d86d119550c3039b2507454ba135b68356bd034a5bdb1e984aa096f8cf808928cdff63a357998d2b501590a97a30760b576be215fe0bbe9b807de55abe5f9eed3588570f02bcc7cb82ed6abd2147f6dc1b9bcf0d234bfc4f034f06195f34;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b967434d14c341a10a64e8c1d392fcdcbfc7ea6339f078088acd3c50a6f637c5b269f0a63fc6dfbcbdd93e0ecb7615abbf997c6c25d6c371a584546d0055528a0cb01c4f3a9d5d14ddc0f6bf8bf64e5117bf317dd4e7afdf052cb2ba432e5bf68daac4006ba8670eab;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d98259e5a9cda2634805855c1e03a1c5ce049b9391f6210ca5686683f36fbafb16013f4d3f48d94d43683a69ee5a1169db506ad52c9403ed4350dc44b97e5267a20b45b2df0987bbc51696f804aaf33403ae827a687d2eafc45170f1d6d46db6414c698fa2f928feda;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h63b62ec710f100958e16cb5fd7df0cb5419a2b043cb61b88615cd1ea38e5fde2b25efce144758cc30b025c01377c8ef9c17981909539c3e2c80bd9a54dae4ebd9e0c3de15d603151de3295002093f90a18ebc68708dfb31ccee7a69e46d4f19b986f77613d940ecec4;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f04ae88d972843c71a42b3e737cc19cc33ddf16865511d876608717dc008f27bfe9b73d7e19b5cb0386e8f6b6073a1b02b9cd168a44f88818899e63e1f2aab9ec55638ea573cda45918f5bbef4e2e74bfbe17c23c1ca663851e322c5a9475a0ad3bc6822e2aa7e8103;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1caeeab78921c78967c17700b20ba090035ff5ed628b1c65f67bf3e81b4ecb2211406362aaf5cceb7490704c36b22933241bdb534df5be873daf0b641975b9eae68a5cc4c414251dd2c94da97f1fa53b8565556790d5a4cec23b40155e786bd3a205baefa424341bd00;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h3edc7c975261919005e4c91da52239b6db3be6813ae50b73b86006572f3fe7e12c22844159b088f9cd0d5eefe0dc3c785f891a91dd9b1cc3f96747719d8afbb3f9b00b933d29bc3929412d711f389f05714d6353e0f2c453a891a9eae16c86eeae051dfc937c1b50ae;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h3697a9fe1818bd069fea739c4c07e168df2a656c97f0f8e61f318f7ef64c56b3a08ed7e393798d9eb839c031c7a9c2846735306b2493a7bdef125873c560b21194642cae924575806571097864da71b11de70ae1131fd7dc5394f9ae41f6d204f9ef9820f7f59304a8;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h7aed01b4443c3ad0b3e2f868fdf4c1aa05e2fe341b9e0eecf58e4f85e930ea915e24e961522fcba33bb29d79b9593e9eba89d812983fbd03c38eaa2df8f3f4a7c9aa3fe7091852e5ffc73e9203426c34ce04c51d7a2e3932652ab8c29b6f2e9fd091221d370937fa4b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h15cb04caaa82cecb5fd0953981af40aacb51b056973156389b523b45052adad5ee54f4b0b7b4b77f0efa6a611234b903fafce5482f1344608aec5bee1ebc047e82191bb9e878fc9df9d97cba1f3365f4559d4848f355c07fc0a568dc82b40dd2e5a568cf5375f8f0a06;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h154ef9477e5fcd91df9ae5dcb1a0edb8b4c776942275002c0f2ea31061c78a69724317a180a25f129d18af1a12a4945d82a5016b19b4e4aa2ed769d7bf900e338993c869c268d06f5c3622c57ad0454bd8d59fbb56d9b57f12cfd4cc1e763746af8ca16194533aa3a05;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hbc0c8abc6c0ad94f2433871449c26cf5439a0bef475a3b098e63e2fcda949d31a5f0154c67b7420a650a65a84a4bda9bd54f8a51ee7e8256bfc7d089d99626e85f9062962e7cc30952a9851496bf32da9bbc46c73d862e08573b569709779fd4309306c99f303a6d3c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e185d9000ba033a1c11df465bb06c97c258e9a3457aabb040ed86a4b6ba9968f4c81f90b33e895adf588829fd1025151255127a24cae79b4d15238da24e1ed1fcb96398a823b2f0b186722d8dfce3a669eef2b664489e69af71567ceb198e73cb69e1f72dd9403f233;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10364bb42a47a7185612d3dc3f866343340908a5e2a20f15c8fd8ccfa2974cab94d6a46aa7ddd8ae1469a66e720b95b3282d329b91665dc1193ac63dfd08acfcd18075b5ed63aea69325c793a1e1a63a7288355390b23a8c0295160fe4fc8cc36b6d610489853e623fa;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha935e9610acc1536e91d316b61aa7a7129c01c57b11a5600da4e745d06cca815569241048e119c20cb875fc5afa875f880d0e24001511a9e944ce5eb7541fb5fcf9ef7faf24e2ab78d30955eda0a459dfcebec2c4805fae11313c9f2b1e6a155a628f0abb2898205f6;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h246a5e4b7c14b67331b1c88ed9f195de4f197b77db1545d8cdb97d5c66788b42655d7c80191bc7c744a28bf5b3509a693bb9c5313d1e82fb3db44d01f2e41970ca6b3d3b976070295d878ed55a04e06492bc95213d32a33d5c134b061839a7cf9057b5e5efe7297f3c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h8def81e80afdb6069b59938bb7b0c854dbc33fdb58f38679c1b01f123263ce977e210c99a0f36077a4926852829c97518e0e5544eb798b26e3f14c8617edc28ffb34f38a4c879ef2c69e703d3ad17aee2cc54088df9c7faaee3c2801066de195a1a948cb4e899bba46;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h743d440ffdcfc44f8c0dde332530bf9657c20ce0e40b29c446d82f1e165a11c34fcb55fde9e758628ece8f1bdd1ce66c88d6cbd88e155ee2f0b17c850432c3b07b6622bfd0305c2ec85a93e1ce35c9c936a19273884e1efb62e026697570f2c0f945ad3e3c69e2b82c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h120e9a6ae01a0dfc79ef9189f8fdfd23490a47b28920dd5bdc7583b5a8c7b7e3419004dd36483bb871cda9c0798e4e0ebef7551368e357fcd0e28f38354b7c0c2d00b4864501b67a798b8726f4c0473be97a177bf83a32d7853fd61a51d18ebddbc129e1375344392ba;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc68f44e830dda99f0c8bb37cd27bb33f3caf615d50d906665dc0a77eb7da983b66234a861ed4d97bfb7d672b888cad85e885a74d982a825e9d84c0f25da09a359e3a17a72f32ce2b1e59407a81e22036f743787def8890cdd1cab085d662095e5b08de765091780f7f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb6c614ab19f2d774fb8ce3d204905ed589bf32931c13b015af9849e6f6e81691f716fb9dbe4ad9be7b71ecbab0b0d05fbfc30fbd8816cf236c88ffd3cf10ca9632c5685535ec203ad369d86bb4b1fba081b63e936569342e75665a26c1f128ad47ee36ce7f2b641f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hde337a2b86be90dac3976950e318cb09bb36bd91cbe0c86885e7d1a04a70409d5776f2a6ac9149bdffb2b240a46ec4b3b52c79a21935abc086b3b43b4c4747d251134d3ae3fba5ccb9bb5e7a1abcd205e8e8829222d33b5ac9aae01f8c4dafaace2c62c5bf251992c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h187eda54ffea460b91131a386aba2567248930c9e1f2bf1f37aaa4dbe4e423ff098e78cfb93a5452810b0e6b87de1fa74e5227ee1331d1d04f67b5fa2e6917500aba77a2d6f94602cc2ed43013c50fd6906db718286341afdb184298963db0cfd8a01000714b95d7e9b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h2688a3718cb3131420dcce6aa43943192310408d22db87343edabaf1380d3ed1b95c8bf77671f5dcd6f0f7fb240f6eb96a482b03625fe303bd50929ae76a0d78c8cc92657989b7031ae29b29e74484ad0d98cca175af80f162977cc585dd84c9988edd57513048d762;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h18a7f27601c67d6a4df0e2143f1e7352733200ebbba7bef1c933bf0e69a4c1ac4ee208dfb70f1b45ef19421b4127160e5b57bc3b94e1ac77cb4492b6e5d8e91f11ef8a672d7aa606ff69a6c16347b5d9bdcdbfdc0ce614617609757e6af36bebcfef4d8c9328063aa65;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h9cfba095bbce635c746f7d006d26690e1d50875e307323525ca1ae6bbe1970c9733a06e69a399fe5b9fcd54c5dade5e357f78af8c542493b017c99deb630f9a6e1a0d5167b2d82846cec140e97245239b8a912159690f2c7a4eee9145b7a6f3b91218b17d272464d39;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ae60c27993c479aae4efa6f33ce23151e3efbff7ce22f653ecd94971423654b4fc4266f986e5e2c902afc5dcce4825f4387d244eebbfadcd19e73d273a2ce85e89f3872a013fe88e5ca76937ea305220a58acc9f610cbcb2506465aa6ca12fce69e3cec828fa62a9fb;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h19b1996d3ce16f123f9b9c8f97586e491e131691d06f81b365eed1d5b3989df2c806087fefa440d965432efac1b8969ffc5ca4facc75df37c2c6c5a03bf70ff595dba723f36a95ea99853b2226eb1721df7da99395432925716aa023da62f788a0fe4bcfff83b6a5619;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1896d469d05cb0a103420259775970f222699107f5dcda15f02bf8ba5ff6eec6f5ca39f778cf26d629edbb2f91e3fb04db64b82f519e671c30b1dcd5a87d5bb14423091087226f8eb788d5603d4cbeb44675ee3722df6085b3f5a592766aff7851294792b47a8ba19cc;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h118eafbc3b0c7d06d41a52604f481cce3343db54a667c42bc73e6104d45adad7165f20d6e799276e37d78f33e06c28798f51fe8f97e2b120118dbcbff405c6a32a9d212249c45e2d8fd8d191488c94addb89797ccde202da5a5a1d8334ed83dab7db21fdbafb8bf54fa;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1bd61ac5a14bcf2cbfd508f581c0e195ac9978f635d84dfdde6e0fd2b5c4c7db244fbc0cc2894a79cdc0d2828e923e0a29e6a32dc11d97753454fe1a505b06ff4be6d9f048b88e52e6ae178f13c613d56be590b97b226bf25f55c8f65b119db6a5b8ca6657cab200c53;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a2a6d52dcae529a36b9d03c8aa54581ab0517fe073bc2a848529c32321ce007caeaf6d468668546c7f7748fdfee3e3c084f82f4afe3f1707b78bd73d1a49587c6ff873fc8a2a3bb71fd7c4a9d2fb3aefdae53180d3811c04349bc0838bee9f13ad6919e2a9c1f5843b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h42a743ecd2283743923fcbcf60485bc6bf09bd4331d7a034a1a7445f0f3268c79a007a8af2b678595c2c477e545217b87e2e69c90b459350448e062791505f764b9859250024164abf7a0a01c0c07f38e2efcb208611943f2ebe722587cf1054299b4e5be6576d86e5;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h79899105db7bff4c351e5fd768e4da308a85c4d981dc04cdd90cc346c8d253541bf5a99b19cd923574351f926def47e019c73671d817c46301adc20a9ee3fe514edcb2cd0883fa8f6e9a0884bf42dcca1a68c9f8346940ed2b081ba35e6b016e8039b3beeca63a2072;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1714411ebd0c536a3633ee118c1b604b8190c8bea2f4ab581ff9eaec0eda73fbb2bd96a918cfff13269d14ad3b662aa339bb7d6fdf22955fa8fb6e9a27d61c3c56f57df655ac38aa155e735851e3990a320922d8ad6f348289e5ab3bb87d5a3e24f9f8a22e1db2176a9;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha584ecf426b244b26c3405d33953c7d7270c4d5859471ee677f41b280ed294e3f8a844072936e8dac5d6658864bef37e744207f3c2f6876366c751124d3592b5e9fdd9112221db80eed446275a9b3fa79356248f7a6a8d8566f1abb69bea3d25c701962f8b6334e7d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h831929578a545fb8895009ec5084eecb3e67346acb7f94726f0ae5e989d248c3933137d8ba59f22cd078d01354cc69fff51f07f1e4ff51cce7006aa34aa46f535cc3d54a3edd2a0f5df03f5c37789890d331ebade27f832a3e1333a4e79a9967da6daf912861b849c6;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h381a2727fb9a1f6fe57473e521b8fde49d811050e4d9dfdc61f1154a5f56d9ca476d7f4e4ba0c62d6388c0ec56d3dc78746124cb7a34b22757a7e009cc6aa4e6bb53fabb9d9cfa3400f4e527bdc1feed37ea7b9bac38018c231f9c0c9e95ba49b8a3f4418f1cbace1e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h82ed579fb8622e1d592237680f8b70f5f9615c53e243427f279c07653b3cfff69c2da85ac562459007cfaff91afaf4b46b56b5186f4c826fd9c17037368e360f4628368f9c8d47a56bb500a05790bd65147f5ce3043caf9060a01ee83d0870cec1cb79d52393e20b78;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h142ce45517a3206b80757ee20db6660685d4823edce8145604ec81855faeae6389629acc107f5e64d7b22fdd6ff4175487972f5e7fa3345abb9e43ecd55be472a2c0ee755875e8dff68e90a18ea88c8976c774f44105d8e9af03c7631835bcb03354981454ac32b7ffb;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h261a6229a31a3978a1ab74d88d4e81f8e89bf225b28efa5b2f5d43200ca4e3e4a060ceef9c756887c83db043a15b74630fae991e3b03eb5b9098128fe151e95eced524d33685dcaaa4b565d8e7bc79c87450269c21aa9ea6acdcfe29fb49561a43ab87083c84f70b29;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h124432be27e10f08bb6984b893c32a4c72dc87da091514179fbaf47426352da5d0a1473c22f9cfd55cb2013971c9a01166461b74d72a644af0d04db1eb3cdc05e5f6b7b2c4710a38769df232213872903cd790fd55657978ae382c8301aae5d6dc996d9e29dd0f6602b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h13b7dc6098fde516c12f0ce01286c7bb3641e29a0df88a5944913039268a387649439614fdfd8a14f75868ba0a2768f6ebd01c459c65d520a62c9bc28320495bfdac476d0dfe7709895c77e9a012d97df5401a4087bb95aa89e6922b6a84d1e6b8d347cc93501cf111b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ba8535e703fcea0a0d50654fab4efd3226510110f060d706b0919de3c2c3620bd0a3b2fb2ffab22595e4dc9c7651ee5dbcdf6a29d7896cb8b44b6817ffe813a66b53fd8c7033471114cb81be6ffbbc8864d56c601d616381b210641d2c1228ac3b524cff0c6bf1a051;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h18494971e2c23dce9fc4cc622d389c0b5a8fb21cdd7278946a1197065d65fda6b54835838e2de5ae6bd2caf2938d9e34e9257700ea34bd1a4d928d32de7ef562523a76def3a9cae4d9b219be150123ddf31253f37d0584c697f1aba011ccfcbb40e0b5a48464b914bdb;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h83c5687949b1be467169a2d06d493389e1bf61889ecacc91d17d66175b5f6128378ca444c51d303b29ee4ead4fa836e994618c9f3d4b6cfc65f0d210c7224e53f7ae4a3cb6d3edf433c44dc36f465c891c9a5b0b41529e35b5f4d320e51170640ded0a0e311a46d14f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1bc6c3ee573fee010f9ab83ea9365047c280faa68d5a55e9ba891aaf15cb6dc1888e73644ed416f650005c1af29c3b11f6b14be84beaa844711193da6545d8cde4180db2225d00fcf1e7cc67d2581c02a8ad0380369b4812812cfa08a249f7e424cd36e3d3a7ba6afde;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h14463191cdf22a3d35813a17c92bf330ee3c6e61f496f0ebe6d3830b9d1040c4b93e41d84cd64be439630217eda8b6018e121d974a3da3c2d9f41eccf027bf9b46d79b27e5f6cfd98bca7797c1d1e54346f263e97e8b46153d2b93f0d778ba9935667b7e57c86acf733;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1231ca8a793485bb23463c3d60d90e4f59c5251309288d77b36e94dac9fe66eeea02fd53256d2368ed1d337ed388f7ce0d3117fc46f0464a3e4f4dc074a95b95d014f7dd6e68677692a3a14bec328ff9c1c8731b085b9d98c5144cc5220435490e400fe23f8392e38d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1475806530be533a3380312ceea3a7b7f08061aa6e8a661f4b94be08ff3ff4e37fad55fb0591f58c6fef0f94449cb7ea034c5cd666ea3393bf4b901dada8ba274a83c9a8cd03262b5d14dcaa78fd0899394d603e55318bf2265d52daa319e4df62b40adcf2c81d7a008;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1de65d5737af12fbf0828150f2f0d63c978875b4569607eae1d61aa8260b52c7bdd5616330e598284a5a7a9dab951c85acbfa19d569ff00e5cd1c39b0b14829c9496f1cbc6e50c0af164844f048762f259afac8cef3ecc88ce5472eed1e457ddb8228dcc2fe33b8b11d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h172618c14307405754e669746d49b6e0ec2c9d65af08a84ac127d758688304853a0a823e4e539a93b5ce166f6b43da2d6f3e14e573e661ad02027448e7079942a563b941c847376e9faecde0765c19a824f62f19c055ac5aa24003a362d64c7e7d6aac5654c0fda68d2;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d8bf5f7ac23d00e814c1ade7b09f702cb1b728a73c1099bb3e0925710afb18388d7efd45e52a809fa07890a403d31d32017b104a03b3c026347fc2ecd3a42ce8f57a14d9b7e235c89daf692441a19a291b32f6d7d5eda68520bb5d84188f640b4e8daf4ed86fceef5e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc316042f273f5e2432bfa4a9968260efe57740496a3844ec4d0ae01ef5902e72827b00f97cfdbbcb70c9a79d071a6f0982914deb4cba9e46459382f8039740412164f1a9101acb8fd7fb1925282d4609a32511c05a0104d1856f31391bbfbe223bc5e555ab4cd7d30e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1dd4d47be4dc71b512d6c119a50f3bdeb48d317faff74139369314805a3026b22c93e068b316cb133db503224fc2157c21dc8d4aa369203e1853fb05b0c97a8c573fb45caebd9bff5a03431c9ccc6ed99e7e317465e55be35bebc0145f4dba5ace1b2233e2fca33fcb7;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h84b50377e9cfd4d9dffd239e54aaf9130321fe79ae7427e7242fc189f7138b8767b779372fa8ccaf5129714684ccdb9b54d4d89439942e1a355f0d67b79d1a1e97a8d95ce26a1cb77355aae4350ceae7ba3c7d1aa2e497ea98e8406dbdb8a9341c41f5333e7ad75ddd;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h12907f5fb0a182a59675e3eda0930d6c88223634ad5fbdb64aa8e0dd155c1a61d8ae7e3b037de7c9d453d48092989e86be24f2f846c6fa027605c65ec51a9fc62629a4c3276c5848c503dd58238f0842ed62298a8bfc2278b4606374c1dcce1b525168861f7436970b8;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d8d4a8c65bce8e63efe4e17dc29661a7cb11a2058820851577e0582e4ee503403e522629d25ca7141b46880d78d8de980404eb5e746b36f172729299cd4eae6cff075a8dd671303523f8562259eadd538f75df2db786cf85691dd75d6c9db43c21493d89bd34b6446;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h8110ab734b7b21cf6d3c149c89acfadca8c2a05f48a4aded64f5579ed8804ef398631bc838bbfaf6a66115f3fc316cea9a3deb80bce6100f8ec2d8d327b78cf1685e1f6ddbf03b35e4875fd887b98235f769cb57b66b9753cf4dacf2342b093581ddd92011ecc84a5a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h11eecf9075201f8bbc776fadf07ada43e3fc0e1768b9c6432b406d012e074ab643212674ece07a145e485fc319a77b8ccbffbae7e43e6328c501debae88cea8e3ea60586dd7268286f7a0cfffdcdc34541cd7e599b4b671b7262e1ba6c0a84633911413e84ea0b8167e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h130af105122ed25ec42d6d98618813d038708075a4324d3c2b02ee88a457a0432d23c03108475274642c0169be6837182d831496792d5fe79d0e0b2253cb50723d3f781595af9500122e39b260a05a17a6647717b4eea398d5919e519624451df747cbef4f147bdcc1;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1bcb09a3b05ea53de11089a8eeb30b4c98335ea58d20b2f0a61bdd5ba180d32f2641a00c836b56033ebe47dbf8a91d066f2e102a6ed0f915ba720f42c8884784174141100d78fcbe8d9417b451dd26a2e6e7bc8de052b6f958ec45c2e00c748e20d48fc0ae67d63fce3;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h235e1166d686ee54ea5e056dd50e7ef6789d67f5ca1f0c128fc878071105b8e993e9c009be7e0f5824160f9f42e2f4a94dc374a40f17c361a8879f0c03b23c71d8b023a59498d95609e84dfbbdff20acc57d0053ffd217460b2348f5cf18b031c07a84b24c1052324c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h12a2b595a04c280c09299c9e5656f67aa9021d5c46f33bc0295bbd84b51959b53855615e3b6c177206595a8e883bd29a2e33440966410726ca180df0c5afb140679b2bd9abc03723034233e781dcc54d03de04b59595b1214ad466091da74af6950a751b8892ae60c2;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h17db8e8c70af2826dba275d5749047494cfa58ca3265cb639faa1d128c8a05382d8abcd6b7939fef80db831e65f99f1359ab9c45e56a9f7c9d528adedcfa704c32757cdf1aec6af261660ad8f12229751de3e1d6f349d3094fc8216972904c6a82cc322a515a615a6e1;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c17ad11aee5dfb21bf11215ec4372dde59c5be3480a1ca0407e8d1f11ab1e5b125bb1a4cfae011819f1e90cca2e077938bf1d7cca0bc44f7f0991333c86d32b695dc15270fd80a13a90a70e0958bc7e377eec5e6635f400737742d08f5b8c514c436b18086a0190a66;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ff336295edb695dcbf6314abbb322ccda6f2e46fd7cde181f7dc32cfd992c1302472457740eeb8269cce1136a2a364782628d0abf53bd1d95b7e9a2a50cbf2608ef9be971b9e1b00979e814f231aa057d166e97cf67c805fbed9dae218e8d4fe35fa477181a303fce9;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h12159ec552bd42cb4a8aa511adde8b1f9bb4e419b385ee245917c112980b1051eeab7d00c155597a1faee90dc61299eae8b953cfed4930a9440b89dd4030b617071ae69b30c03fc42d8d62815a6e58d853788749cfc4b44e4f85f6a112d66450d0eb0efb77bfcfd1d22;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h17823d9e55f495945939d735ef627735f7b1a3e5f9b1dbcd4e8b90e808defce894120f7eaa3c0dcbfc0cfeef719ec04867e6e21394baf760c2209bc2f571477ed9717213f3fef8a9a336fe74b6e1865d3f5494b2d0855df6b55378a2ccf2d29915db2bef2687d985690;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1abbf99abc9f5b5125bd4f208e31c5f1505557d1dd4487207909c919ba9473e2f7a665fd870bdac70054630df1fa0fa8b1374bd80eec1750e438a4fe088fab65407af1b49c86a87cbe9af0e3ce18eab79221570930538ccc9cb5fca9ee1de802ba3f9d3208ab09ef077;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f498512a6c9dd622e60715ee486e0a76e0ef426740b38e9e278be7b280949d268af9590638160e55e5dac417399fc330b6afaad6531db6e63947450381a750be85f1bc3d65f378c1f07ff17f77b6f7bbda35a1d28810c95e5fcf0a97be2729bedeb978df60044d823b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1aa7969f0e40e130646d1fb3794434e963c72dae3821113b264bb73b79e8bfd719026cba369a8154235bcb419e5fa290370d3f41b101afbc9219ea300988023c2d3e83c33712c587663c300b558bc2397cb7ff95830fd348346516359217880bd4ef290da7271c60506;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hbf0c9489f9a2134df0dbdff3a2c6a39a96f10fb4e2f13c8d945cc8660936165b9e224552bbddd709465fa47e99563011e2f46629342d3f30c2940b429610b5dc1251fc61868d4e5dfd4be01779e4981b1f8a5b53d986cdc25b7c836d489fb8957237c19aa0336b28bd;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h5fe10f0cd7deeb60d09da41a6ec451c301bd51f702564e4ab405399cf4ee75a7be25ac654f826bcb5feacff077f2256b510de20689b06741e19ff3cc7f211cff8fa632e9871954c9ae392a4643d9f58a196caf8a421e1ffd15148dc91ad5e300f9231b235662d57d15;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c84c8ba0bd268a28287e963eb0986b1d5401e3bfdf4b8fec4f40df1902871e15350d7788f7d584459ffbef283cd1b748cd637ebb34e63b8245f198a3e2f583748572677078786ec446abe4757e09a6cc76fd9879c30fbd060cb4c798626841e0ecf59b12d7a25192b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hbede78880b1770f42f73a691a2caceb956e2f86993531d2d2de0170fab5ade90b6318fa7e3a3786fd3a3a907bec9e1e3e0db405fed4b6309f2c1aaff34a0963692d424e310c7c3d1509e3b60f1bf9d2d2605a4e2fb55e84ed8a4bfa17aed6f50a257ced9f3f9d76e86;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d93fd4debfe95885f002d91667479db84215bb315b9c18713876e2a08a27b38e83768b9569a106078085a5c4c228741e6f1051cd6543f2a888b556083deba9cfefbd0648a8ec25c3445193e9585a33dded37c63c4292ed2524eba539d46ccf9239ea2ee32f6c17c52d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1cc953fd701721cd2bc80e8fb89e0db205bfe348c3f24f8ffec5f6cdbd9d4b0a8153877c008c39f5ea0c1bc50abfebd6fe97b2d7db1560d3ddd67357317dfb46e775dea3bfeffdcb1565f4160c2a9b3b0deb15854aba47b4638ea71a9a197e54c4e1dd618765803e6b0;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h55a6cfb187121c95f6ddccd430ccbbe87539b2577e98dbda716a3ddedce74289a8de970d8ed3b5605c450c28bfa9955d686968addf10ae0a6a005d56ba7a76540b1268ea4be75a4966c215f2ee17984af95a0c6598cd588a8623ba641c0ad20d85e1cf8a69943a5a9b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h4d1aa8e19086873f3896bbbada4542915a8f5d4e8a22108818a3ea590de843a919cb49efb24060fc53ab0caccf673bcd3c6aa02a081462d9cb3097ea256f7ca72c0779b15ca59b1775682b3a340027792a0c3891c5d3ddd580a95774ef590d8631e4ac60933db56348;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h120dcfe14f47ee6f8b2124e22db7005fc935376c79ea0e43f99a54ce97a2de75b5b73425467460107f038082dcc373c10dbce7364c0aea7612f422064db9e5358612f2f52818b9aa45dcbc6858df2fc958385793d406f428cb7b1cd919020d0b26a0cc95dade084241d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h18eb6717cc6c6fa251e531a805b88ba60f754e02a4567d140a9f162663611686973178cc5a0a025738b070bef4567b011a7c6aad7c830b012a3be638ada8baca056dfb4140952b4b83314282562656760a0efe44d6dba8d983680b45ad40d6afa460ca5e2a273ed1ed5;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h18d25cbb0400627b238d889a6cefc11ea91df7bcfed29a64b804cb52a96f296bc81b72892a9090bbff837b6b227efaa3f021f010853034484495a2f5f02245e8c74fb02da9c1deed9bdb6c8e291bcc0fdaf12efedd780480dc1a31be79ad99801a77b592f1c93258aaa;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h85d81d0ff3c49e198f0787330b55d11a07d2b989d9c2a435bf5324d2ec60d344e8c6361562b7fbdbc88fcd498386bc35fcd7e3691537df0da6895424c511af047331bddfbdaee656f54bf44c0b377249d506f0657dcf161e2aec4a65baa6cbcb7c10b84a0cdd3dab6a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc7ba2467d57ac9382bab9f1b6e71b1794d3adfca71e58df929db029daaa0b396a841343f271f63bd05ab256b8afa07646ce2e590c1d768346e6dc216c44dd3466cdbbaea82a3299ad142f290b5890a93f4a70f3c4d1c13612f0da8fb7aa0a4fcd6d7d7322e19db121a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h158ac51f5dec46764897587dfa16ea3ade6ca082a03b8a7acee81b9894ae5c2390d17c2034af11170539c2874e880ef943a1efd80e60c93da71520751ded24a408038665b07be2bfc183162fd788d7bb84e8d88d643d91f60d3dd599cf05b22a131321d4ec4acf03ba2;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h16016d1d81cb9c72bb5d4ea45f6bb83a0ef24b21a3045af9cb91873a72705ad5299d3fbac61225f5dd5332075066cde4a3e202bf052cb95f8887e07bdc65a223020af8c99e7c2c912230f80530c1f104249c19b393feca7937ce5e066c3ab16cb11b1d6bc0ac1ce795c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hcc02e106662f25e70c39e05bda6788fc9dc818135a8591c76a7603c3cf8a21480b3fec0d157acfea825afb7737b0978d3492113e6c4498568c054475432cab2cb5116762f6c9700be5f9591810c57e63b99e49fba8a2874a47fbeb53db2a3a754b0c1d1abfa5656e61;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd79ad6d2946ed1fd38e161f399577b22ffe633768890c038e15f16828b634fa54c112390cd687d1f008f8ae1526ff19ba5beb254c33b507b7043fc6c57785e51b83fda8ee8502f1c81e74eb07b50dcad907a6e4f355eee5dc1fe4c954114d45e775cd1fc640766ca85;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h18c34543c0367ab3cae524ed549ad5e380f8a20d4201a10a53abe2f0e00d6d7fa24a8ad533705dd9a901c1953f55d49921a98ea114a0fc36bbdf940be8fd9ab864c8b0bf29973bff9d4a18962956fd6721272d0851dcd99eb56ab563123fea7cdd28c602df311e4766c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'heb66aca3b7e18c8e56fc5d1140acff91be8ea53b0c2137e0a22551c99e0e40b70ee7effa5d397ab529a9229ff412e97ab0c1f2779f30d8e5cf165b5eb5372f5314572cc4df424c5718b93fd68740a66387b28135454fcf20b008e7abc61e90fb9584fe3905e2f87a3a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h185a34538e81341e69d9a60a3a8aae2a441daff9f657bd587b90480c147a5005b9c7ba446c19c6fc1459081df962c03724ac87bb48b222153297bfc6c2ad4379b5d7a90a92f643ea9b92f174afa2614053a7edadd3faf5d8b469d0c24aa1767c24d61379d313ed42171;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1bcc4d05f6fe407a99d657dff2adc7f6153bf389dac327d3954afe6e8310b81cca8930ed6042d047ab1c74752284dc8dbb43327dcdfd2c330444c5c20e9d495c8f7e6f29e1052feefe598a91cfb346cd9e2c7113acee1ab1101ec8ffbd94f0fe2362c0ad5772c04ff07;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1896b1876acc8758cabab94a89670e7aa16de558def049e1d05caa96425569f9b19423bf95201b3bd6304d8dd74e6d9fe4d29c651b7e65878b5cd8dc7f6d027c6568357916e733ab5b55e7f51197cc8f3b6dac4b6bb6cd390b3c9b93176864945e54c939194c776a4db;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb66b1397ba50406f06cb24568a444550cd6f0749bcdea4980b9f4687ab30c19d3a76a48e4583f207f01482380fe84e1832bbc4df37a52d9c68dabda2b7e7942a75ab0a9ba3dfb565aaea348902ba37c3cf4d0c2793fb7cb5c9aeee5cd7e21ac834ce1039db3f3bf465;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1705a336d8324e586b335d7de4aa5203a57578ac2b8162aed9fafc4cdaee308e043fd0bfaad29ad9e187344a9f8e9bbcc749b0e2ff6d5e14c6390a4851a358f74e82da8782d7680de4b5e9fcc63c8a57208895f8462bb555e764512618096c1c3a78e88e37f3d14ec6e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e32e862965d39a2ba8214ab537cff5c6c534d0765b863fd127d36fa2de180185c6f38602bc7fccaba549cf05cf518017f070c895fc2599950dc13ef26dad17710da5663e61dd0fcc399f2a470f5f504e8a9950e4de26dc6d7f5abe04e9fdaec86acdd8cd114176b35e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10fdf81e54979a8cbf79353ae3aa5dc70931884a7baa2953fe71e50e239ede308401480bcb4c3638a243b877e77d0939a0ab3c22bf4500dafc14b25d1268855ddb97a52c77db507d96f62f647578a381b7e3345f3a9e78dfed2ced2f8fae6b571c57e9790a211d1af79;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h694523a503e130eb4f14e8398fcf1d60731065a3755f55045a610fe35fae54260924ff6cd3c43ff6bb2e6fce4c7ca9f1f2e7a0343f25381f9c11c188856309f5dbbb61f44c691671a0c47eb7c16870067a05e7589d5495016ce8767abb7cf8b4e11b331ff9318b2739;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he29ac3ca00777b1ddd8d792520af337fa46335b968126a3f0cf0d528b07eec8eb589ff93e414b28a4bb5b48c632bef0406ab55edf21aef8a0559d61a41c7332fe08624fad051b71e30aa9cd695ef54f7503137c382a20fa50a9e391023b0059f694fb07b5045881ff2;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hdc5710603b6a3546b5a23be6684dec4d32eeeb48ac53601416a3502da756a379a46d37b2e66d01dd54f9aaea18806fdb8c32e9bdb1acbdb24913d9b4fe70b2c43b463734914764c996bf292e952f78cf949f99d2415db9f186c263f2285374bbd4aeee3027e9aef8d0;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he060b3e1c1fe7aa58319c8c5d333d08fa8c6b176fcd0b68c8bf8f150d31ebbd7a3ea53055aa49be21bca867c49a0f26decdb70fc4086740c55f6b7758d615ca5692716607a3cd1e9840bb9bc8f9e5afbe230a8d9aaa853023cc0eb7171eeb2b35e916649d33a712f96;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a723b6c0c6577807e6427c352191cc0394ead5cfc3d457068865f513e1b25d1201c6b2f62852da88548d67924df3a45d36db00ae21e99e0276333544a7b693d193ff59647cd80b069b4dd12ea6ef8cfe8be90428146799f7d4573be72c0049bff99d6463bf352fc5c2;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h396738222973135ced8e6f169813e2b8837135c95c6116d6efc489c09e390b7cb04e52a8c5619e412e89839b6e6e8df997f74ec40271058f499121ac5b66cd236c972ec849a1e1a8e2ef3a4d9607fd5b44fbc1fc83b58c11e36d93eb61fb100c44c5c615b986c9f4db;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf17c8914445b1d34036b2e2c0cc9e5ce30fd9b3f7ed18f6bd63f0dd263c997b8fc6321c002e9e1c4152cbfe19f48c815435430b2ac898661b10b19e20a4456875eaf8c07c2846418829e364ce18d598a187a50d12d8eadd7cc006eee49ea26b44514e84575a0a954c1;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h156d5080dd017a8b839fa570ced257b799f38cc8af1c229d2030376cddc601f0f397e0785373086bac723d25c127147efb365e8531ba90018ce3db96f823892ee90c2d01d6e3b5ad96db4bf0fea822a9ad67f9b2926bf78511e3cde2374004ad6daae185a42bad334e7;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d4b97b99356829b34382c89c4441bf5d525d5240286dd017e10085ccff1dad23e85a002c2a90c34131c0fbf8381c55b0ab1fd5e696a6e02c5fa4d99ae9da67d28e4812625b7d3bc59e9c27427214337fe630c0f91b465555fee2d3164673b9c304e38dafaf838fbb10;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1826d025901bb46b2deb454afc0af241a4af2acfe56bf046c6680f0a8859cd5e78b43b31b0761a2e2b59ff131aebe335fbd3b69061158027a6ecaa2ae2d9f2ed6bc10efa3ff7f14719d32aa470736f855573ededaf905f1b7479af8b145d76d176f15be7f959cf6192b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha46d21006dd5ffb3af1b510791860c215c7a5fbeae9d010c07ee5b659c39209fff81f32ec01798c4587b0a043b374ff01d789051f2ef5934a87f09e928522aed6a870589fca8927a0bf36519d6d02284e109f21efd96de8024671224e4bbb6f8d5cf771bc88518175a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hcd352d238402622783fb80693d311337a94af06a28d8661aed33330c9d878f7fb8e3e8d9362265ccfe5d5274f85832553fa1e51e82d7563605e112701b5503a6e4e0998022a29e7bfbfe3f7781c0053a3c45254638c4b3f4ea52f6e5c6c63f0520447714bf41c1b3c0;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h3b7911c2ea34f15ab667c074df06f04363d00da7ab68c841fb348f51871020e2fcdaa4e1e8e3d3115d89759cdb027939907d47cc030ece8ff72175f7abd0d872c2926b5913766e28ecafe11d849728b6aeda493f594fbc4c75d503093a318c6797db589c3003311fb5;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h26478fa9eb44cdbc6fd5d6bcf2d2f517939a271429a169fbbe1df4dba4e1a5d8fdb0e90d79ca5da59d1e2d5dc2cac9dace1f4691f7100910ce58352c4fa6173a0b4b56c15d91979a4eae2807d6f91b3041a2efca6b8cd0cf3b131f8cfa29d8891635f6b9c623b0ed2f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf9a8f6e93f5382176bb69cc02da4234da5e7c6fb140e07f83ac1d3a0195840c91801eca7ed506e60bada377ce3b3b30a791a06808cf6e04fffc22ee61030a5e76419a840ff4eaa65a30b047180d60b8dfb3519b3eb8664e4962dfdd7975bb7435e6c5ef3950fdaf63a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h83d2ca5e56f43e2562bccc7622a2f7da77dc02a4538aa16b225a2a46fa846bb4d99611ee84b798d2d5ccf6916d1f390fe4bdb38a27623691b7c613f30152366c97b9ceb68ac057956320b4247c8e25aca41f010c7ad003af9856398edbdcac15d23a175d6f6aad6bae;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h2b8c67a5c8760d865fc1f87fb7a6f12bbbdc97ff757bc81cee099b32c2468a47f9ebf56f8d7f82ee954f2c8f0fa162bbbe1fae87e92a6dc8a932b79c0edb9e614f768d7875cbd987470cbc1d14ea58163ec3e2832f2b55b2c1d5b3cb00bf440393116054a5ea9899fe;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h684182874388562b497c89799ce02c0b8ea94d4cda6690a5ae28d06394b600a264389248e0bd48a8ad86cd4cc5a9469a241187eefd71507b3450e1e1e744223c5d4d77acd0fd4cbe489a317dd87dfb94860297d5ac799bcebdfcc94acd873e125af0cf47850986ce9e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h19e942876260a919cbeff124de015836d4f63852d9e28224a0367902b0e00528368891874f8c11449b55ccbb2bb31d05070e1b1df6eb397ef261d390df75e30707fa786bec5964d295224525d6a5009096c4cd82d9db84e11fe3ba7f054c9e9401ad560f271cc64e8c6;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h90b6aabcd9d5aa9177f6b450bca26bb082ce92f96b21f8a75eddde665147530e1fc6b0311b0b2cf9f3327376911d036058c2b6e4ae38afa7dae68234499d40946844343703c718e3bb416eef70f9579ff5a05bef24f46917985a0268fe145975ae90a3e388e1f4dca4;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc8c2f601abf9758cc0421b0bd82c1a96ca005c655e935056865ce09e5f54e8f30990d8e52eb99dba7fae4d6fedfc8cb0224b73bb02b422868ce26856875b0bc3e5f847f7cdff30a5a1ced9e5f0dd3e9d316ccba58cfea3e03f50faa2e576e39fe89fd88c4fc8a8dbab;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1fe4061bdfefad2cc19940c1a9cf6ead360a9cfe2050d53916bac9458f3b244a0f98bb5fbf6d823528deb69575cb24c08110fb26730dff7f424c6d11335e11d66c58069447e35cf441b7bd2764abc18dfc3c9d9d726a9f7f16b2f6b0679bf81be0ac36e20b4e9d679a3;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h11028ce055b8c33411967ebb1a159da2d8806978a27497acfe3f4252a4e91a3674fea8fdc737d5765cf2f328caacb69d13c2b3e2427afdcc04cc411480b3e899273faeb074a8ee1c2b03ca7700d3714c3e5bbb55f1d17807f46f9aaf9ef68e627b599043930569f8885;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1081e15af125fca76c43596bca98fc4f756e20a249d0cdc4bc142048c2d2ba1a39699579af3ba81464aca205f90df0803bd869cd677b56a0f182c36b8208fdc5892a4f1c88174b7116ed1bd5bcfd26ceaa9c50dfff15c0e2bb4dc1d8c704bafb0f8618c8081b9f05066;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h140d2df210c34e011bfcca506f57537105ce8465a381c4f1c829e3334b0be2429aa5e624d6e74d0f43ae49ec008f58953f8fe135d58b36946fbd05b635dd7c5b526820a9400c367ab6da8e0cdd3ecec1791dc1662624b6b04f24949a1a7d127fe43ecd912133004c1a5;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc2ce5eee21337aa94ae5f4886795a64378a7daaa5f883571f75f61858b58976e92febe46ac1080c221b3540e15d7df8bf7e07ad5334159791bf13d041afd18c8b1928a5fed9c88e53509b5380699b6472e649e4c6a8d158c76c1d288ee0e7984cd497e2508eb3dc610;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h16a0d967d022c85ec2cd3b63776652ba4004f08ba2b2e897d3aca4ca3525a057afc785c40568efc0b93d23e390553c00e21cb7eef511756f760c3f6fde354f11dafd225bb075efb4bc56bf2cc3e6a755d8bedec4be77121834b27e07e12448491c2accd61dcd33fa402;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h5f51b3fc4d5b7f93612d486552695b023f75a19b84caf293e6221b6293773958c6f6b1429c0b1ddbedbe2e3fc2dd8ff4aa6401707124a17634323aca072595d2ad719696293f18154f183f6744be88455194ac74ac02a956e4b7a3b13a1480282c47b189657b06bd60;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h4a56d94549e244cad4548e84cf8b29194b907e527a7c8c7dd52a8619a08d2de7d6765ee8ed9217d2f7b4dda0b8bc60df527bc2de35d4d78d1c8e5d147562cbc849de2e3893e41b9a1243dcdee35910ebabd6a81991c91d328e9208d1605acafb5fb83cfc1db1a3f718;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h13370c79223f0784ce42851516f8e73ce45e1373b065599a7de63f6097c0f11795722cc2e3d7f65659601bd1c5df1c935c9e854e113021a58e8d957c818fc8081ef91849246100db1fdf16f6ae5993c81b380e5c3da9514ccda5f42e24c404c2bec6eba8b7f4f6aba1c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h16ab17e3d79ef4d2d80854ecda791917f29e06b0b4446a72a45f6ad9bac79ee25ddc30c78993cf0e890d33ef0a3e0adab635b48e95d358eb8b0a08d0f9e8dbe5d863c9ed80c6562d3108faf540357c232d81bf70679ac8fb1caac54e95ad21a23b442fef10fa98d8cf4;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf2e23a46699dcdf178dcb198f04511cc2400566f3a3fb564dae86de0a2c6620f76199c1bdcb6fc3b642a3921ad9ff3d409ae47639e44b92ff1530c3a2fc2a41c9c9241b7b8d385e89d2c17cc63e60c623f877e6d3dd1011c07e4158a21fb09568c52bf19cb47cad8ee;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h3ddee4a87095363722f227ffb5c026c7884ee713ad6ec765e798ed67e2ec0a55a22b3d64802bdaa05f9919f536078571aa62d8950869121262419123c51c29311c17d30d4e1e64e7999b9c27ea77053ccfd22e97f23cb74d006f50aa65c69c7188ac341ba2dbab1433;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h196676e8b1e9914d5cde78639409b84ad8afe373c268150ead7652e2d44a99f275355c5dcc3ffe5e1e8263997eeb848873e19483dbeeb023f05b301d9f2dac5ecda45e0e71a8abe102b5b68f00566688b4c0150e8edb0c7d3dceb5fdc0b644127efd4bb3d7694d1cc99;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h17e3f1ada035fedb3fa2749e6b9fc15403b3494dbc3baafe2708efb0d382c67d02a88c8575bfaf4d0605dd8ac9daf13d694b4d13b8d00c63b3ae7fb906a51f1a7a0bb8ba95b812d12ad9d4b5e2b08b6b6d5257ab8135e519d2e5af7972254bbfee10f4b4d81d618a0d2;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf59dd74254031dcee7441a76f632ffc420f47b401afa236ee212c92662af8c1b5d5073444c885432417a28cbe136ce97f91bebe5b055d45fbde045a8efcfa92ac9bfce95660d7d32240a3b98f1b324dcd2a132be7a0d86a00bfd23b8e43cdec29f2534ac9aa4c1268c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h6f7e379970fd7872fc180aa7d7c80b2890f5301aa1d784ddf2e0b9059d15c7e0cded7c9ea9d2bbe58c2ff73045b4bab85751936bd2da5e2987b5d0fac9405abfbfabf969d342f16bdf7e979e32aaeac905ef9ac81fe5ca77484d73be2839d0e4d2c10cfae42b1f8a80;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc47939b8a2e9c570c80617111734af0908226a5959bc19e5376f3ec3a6967d1ef32ab237b70a0a8a756caaaeb744e4ea6b4a59d8e3982b885b0bd991d05c3a4ec76c98b6ef475fdb746c3051c6c8d8cb3c7b7b3f1770ce0404c56a53233c2b26c1912c33f5c69931d3;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha4077a9bb575772a93c193f7f439ae43405ef0f439e17d3f7b81e80d22c047de8f1abf4a2910f62cd1d18c4b5ca25691039e67e1874453f2ec54400812f6591cdaaa58a9dd8aef76b8e379938e3fb99309b451021ebab41efded7cc6e625b9140065037854511dac5f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h5609360d178263de4d376b18ca7592ff3a36b546ce5d69d804e96ac4bcb335675e4795ed9cd7388b9a0fd4f113d6f752713b34831cc9c5aeae5230b547b940373cd660a251a1a55e72a29bb024225f1ccb692906f8cdda435d075224c5bd6326c278214c25c314a849;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h18b132345f2957c883f58b2bcd19f2f7dda5f2da9a4b14893ad2d3fcbf2098e695d11c7725658e213bd572065c6413474f3f205fd089fd4ea69aa221776bf4955612c0fa5aa3995e8fc762ec1212038ce169b0577aada50a1a46fa8f5d479ffb30992b7cda058c6afcc;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h13cc2cf63bdf4231c43d926a05c34ac9de1786dfad127e5d7be4ee07e822ccc07456bb6cb9612774dab2f876214c51ba645c65f55553fe58c155947558a7f1231d33e9a7f96186137315310750052e9d0dd663c62edc5e74acb1999468b6039fddbbff6826aa6a0ac14;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he73cb68c5e391d8b5f46738f31158c7d1a7104b9a4d4eb45fdc4e9b455386471221b729587caf693e3d63de1cf4e141789d93ddca4ae0f585af312328d3385e33ca2abd0cbc73bf47ea499d46b0700dccf8b231675f88316b2ca8a727399b7ac024ef561bce38dcc5f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b05ea924d73f8da905939b18ed40856ccd7d6862b0af31e4c837e2331d17e0c352cee988c78bead5057b6425c78d0be2735a6f39369622c215d8c3545066e73860ab1b176b4e9e011a672f4fc88460df9cc0ef03573fdfbd8cd516f981cac015eab9e0a01a64ad894;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hece32a268db0e9bb70ed9ce274fb086d2ccbb59cc45cb576fa1ea18f4df012d25e1f0f329583a175bda33dd8620badca727890a652740540e51170643913f8d72e5207a8d0ed57d4a7a8bfb34453799c4d19cf82d675f0fea3aa81e08dbcc5ddfb9dab0fff134de499;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1cc21eb78ea9e193a154dbc6481b97fcf73252cb575e42c7975cc5f120a06b5b2d810e447eca396f23c08b21a5ceadfa47528cb06b8e5046208da9dec7ef03ce86ab62129e4f090ede394f8992a04f57dfdf5a039da05dd572ef2a736d8b5175b1799d22fbd41f128d1;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1bbc3b2987e92b6f5c6a0660b8384ae85c9fd58f16e9d0cc07245e6522eb9f68e2477b87559e036511cd12fe2cf475789de85577aaa4aacfe21560d9caba6735cb5eaa800b39d0c51672a313efe4e0782f85de067af6f44a680fa4d5dd697637af806b36ac3f8775349;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h150b604b3615c0077aaeffdff0b3a71b1d170f50a00d9c8f39e15f540437d5c95448eee0f7fc5896078b4c6b922e875885fa06f26a463ae2f243a178b21fae50647ac02e254474e8ee1ac5e000fc7ce1d0502e7780e0a4ca5198a5e6238c17e1a8212b8e348a8e9c59;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h119723c3e96d5d17ed8f5dacae6a55952569aea20d260d2adbca61f23acacdced3150c04c03c78712c19f751475227d8e26f67ab4292ebb63b94aa56c9e8617d6b3ee49f566a812c07d9285ab254fc641eee302643dc1990e3f1832a4df55f081f382d295f3ac34b468;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h143a1ac1ae950f0964490933172159df0bb622818985aed3187687a6accb3b8e5f33511318f448b50e59f6c4f2ec0858a58d7eef55618c7d7ad04d96bc6ac973d19a4cc6e8fafc4d010c9d08b9a9f1b22481590c3509d60fc1c767f510241aae589224813f15f8a6a23;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h8b4458b4afc25567a664d365fbec2049e735cb783fb8d70231e50adb12fdd742040e9408d8417830ddf4db084a56f002f8cfc6c653e33107bed2bf0d7fa08d3e6067eb4a411a4db0ec70faf75dc3d42dc5636148ebb1120f208fa0f0e750385e38894c728a0256cf9b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h97dc412961b580694c7928032ffa39e78c9d3ee4bea51aa843235add0d7139a7eb8e26acb0e42aa40e7ab88ac35db885e4ac5da4b02ff7ec69422349da35aa8df37b9098363feef590fdb38d41062f96d772efa219189b0bba0502b1b802b050f56f2378c01b206b89;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hedb37fb6c75185e242d9fb8e51ae50542ae70aa8be177cbe08a6e3418959e8772e02f8da721eac6f0c86a1f1b1792c599a61afa4a02f1137bef919ef6918d2ee9c44dd69dc9bb600f0ca0267fe6a1fe901562452df0ed369b10ea812619256facc9dee0009782a0d6b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h60f971bb5f01ff685a001c863fd8565ee3a9dd6da8b35a1cfa847432a686d402c2565629a6ee72fdc8d8dea78f9f02f61e694f6c243d795321bf56d995492e70b7e3b5ca6b01dcdd5a487669d7562556b27280c4411a6d52484927cfb3c683b2bcbfdad2cb2079fdf7;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a0c2cb3c00eff53556c065d09e177aff67ed8a655bc6a791355fd31af53bddda96f709e5beffc10ebad29614d11bc99998c8ba0aafa684a66255f5bca497f84d9823f5c057da7f83d24a2c9a427fa00ff97492508b79075ee87211c8d314254e79090ca927325c502a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c7a8c6e462a31f6d64aed73e3e7f4a75b74fa4a978fb47a31285564a7568826a5accb5d465824e898e7dbe4d939adf303aabf18b2ea7f91e197f94ab42f836f8ff3f67e19e539ea280ab3b0c68253d7f7cae6c4a75571c79cdb516fbd4b21a8d61e0f4f77a343c2d21;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d96469e3868619faa6bfd61f56cec3e16fa58185d8dd49fe3432eb515108b4d746bd11bcb48e92c966ae1501e8c6944a6492f5626e1dce6e8aa7cf2f44ccad2ed07aea385da4e0aefd0be031d30af6f12cec177bfb54fb5d5e3aa243427fd4244bd88173fb3baa7263;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc9741b0813282081fefe161a017108db8b732cbc97f8976619bd876b6db8d0cd60618e972afa65fc67ff3f863125754ab7e92fe0c2dfc63fd51a8f9525a91de19eb67e52ab577e198cbabc91653a2cd9fc23387c01fa5e7d17a6b53acffcc0216c99a32a3bb11934d8;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f824626c23b07def67320a7cb226996ce739ba3e661b78c77acb1109f507d2325dba488940b4871ec8de88af5befd83d0cd0675e72b321b8e2648ea3a2374e57253d74bced5e422dfe1078846eada7bedd112dbb61ef90969f6b3e5bdd640431ef8762062143a3b24a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h91bcb038e4728f6aa832f25b717f45957b562bcc01ee5e4f057591fd24257fa2f36003a11bd183ef878d3e4f603c9c3f717798a99eff98b53c628e293a44f95065d51020baa46ed07fc3c71fc04de7dc0ecafb97ea545452354a91e3d55ab475eeb8a4519c5a94c980;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h6161260c3e5a9468a351ab62d182398005b485a38830699a672c082a7c3a2be69424076047214629a4e2f3de4ba97e19123181efbca0612d2e76effc10545898068ab3f40a611579edbfdfa4196f948ce2b780e9c32bc4c4be6c7bbd6acd680267662321b2f2024563;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h18e678f9b215e90570ddd28328d6c0b35eade08820a7a7fac98f9e97f77683cacd14fb40b653d03c4d76dce4aacf006025d178121e2a6649078c0f490fb8db3f5966d2aea8603bd3fb29cda3146af40d83832e15d9aa2dec39f3b2cfcf851be2e6cb5f73bd2470abc0f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h134ebd83ccaa9092f8f0bfff42a9df77c7e00488ac086f47e9da82b0d2046acf466392a901c323fa3c9858019da902e10a72f9dacf43081c37950cd86a3a798133deed754a475dee0a41784b087c3399df2b5cf546ac3dd9cce409e64c73c82174a3e0dc07a9b72babb;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h6151f885ba5afe100b524f066fc8cdb50d2df4a445a38ceae013929f69b2ba00bbdce767fc120791030398de1122be145978c31abb1ac2a77293ba1d7aa052fcdf2140464f02efd064ea2de49fbdea77df42e1099cf3c0cb6559cc06db140373428500f37c8223dc95;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h8825b658dda883d620702e00629bbf16609c717415f5f66456e5a0e2049526dad1e6ed7e7403d8cd72908bd5d2085af952a07301f421dbde6e5dedf1e2bad53b1733eff4d075da31a36188554db9aac06239df80df1531a603e83f8e69d7ef75c1b5814bb7ad6b114;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ae509485dea0e02c8d5d086545041436c12f8ab830cbd8d48b6de85cd94c91c09c9e37c6921907d8883cfdf646d765d19a4a5fc07c967e5d98bb94b37c1eaf550457a16ed48bb3eb7319ea1f497817e7417eb29bf0cbf2c4e1d2f9730e14088d7bb9c3f781e5429eb7;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h7667799aa0392c45c9605eb62aa68fefcd0f49690121f0398eda71b026442784b7375c9a0d541372dbb233c3f1eb140feb9082748f11f73ba342f9a68345fb3d21557305f51fa5f85c746ab5b836f62297320ea9196f17f5370da8411c7ea310a382951dcddac70172;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h13bee0d4f630469c963d0dcc749bbf956f8d8297c97b5cc3457c7889aeaf21afec9d1ce1ad2bd58491759602eb5e5eb10ff136d9f19bf4679054a4baa16d2bb2a0771a036e9efc572a16055b0a4e3f0203856d06f8cb29b5407c8d4e4a9db0d50ad0d1115ee5c31f444;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h3600f5d889adc446eadebb01c8a5576a34b0970678c425e07a798be2dd634c516c8b498e207134a656489f58216a58e704bc588c4d2405f8648a1541e524b48baa5dac35538448c4c67cf48b105f20987fd60d049fff0591ec7119662074f24efa715445f5eec45b79;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d97bf13f670a7cf9925ca8957178433ebaf9289ad0110cb84351b0bd421b615a0a28065f33455d2de263638c256ba035e4be9dfc0cd86ce89e6249608f2f6d4889d7e44b7f1ec96a5de2d2ff0f2aba7310f8f46b49ae721c284570d9059ac1eaadcba6d45fe87415e7;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h63d4cd7192094604ff8ce7ede2d7327f5c0f65c638eaba6c906c57f2f6b16dd7fb1eb96bf79958fb9e132e47a44a88af3952af999f0856906c3d1c7d9f265e78b17c90a1bafe04f80689e57bd94a9b64a291904687e9b7c63e2aeffff1c2624aef2f6753b24fabc024;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h766df7e28c74e8ed8da8f5587aaeecc4e51316c1e8cd208958fc63c0f6006e3768e0213a9295877915dc1a3c645573615eebaea4f38041bab0fc1415b58457d54d5fefdd641122db421f3c512946f055b8431733aecb3758ef05f13429acf4ebcd260283d10cbd4a34;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h4380c2be288d31680bcc917fad4f4a5d2823f25b6a0add0cf0338a75d8ebcc0ab138c32d0676fe0f61f3c915f4563ed941623513bfd21320a6e736cd1fbdad1a7c2fdae1b65708a14ad761047dc09175e4554664f1be516bb85939d520e2431c566228d5393046002a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h123835534baec33f0af2b8170c545210ec512b89ce952a34988772cffc667b18d3d720c55e0d0cd87582a5f5f23a7167270b5bb0c3bb09b1674cb061bba05a1c77dae5ef0109ce00474954d1eb06510753029e7f71dac393b81f70caf89c999d9631060b24ee7b4a75e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h19767a783cab24a93b09ffe3cd720996a16c3f87c6450df885d32d6b50b53be8d0a420384f49449d4f0df51dcd9a4b1cd32b7eec63ea3d0eaf31f7feb25218f44570a588871c133c394dc3cbca32a8d7fc1811de0090e309b460b940789a45b54b181f9456a1923e1aa;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h390ca4a301bd56d9804db19a1dac5fddeed387a7e249f0bb5f283f7572a4348587c79e9ee5d4d77dcd43c3c21d44cd8a969ab3ad28721dbbb2e475b40e3d4c69a6f79c374aa103fe00051f9f66a0de7de953d48dd7ee8586bea09577fda2ba7674b4fae8960201d468;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10729dd53dc6b5d0592a27cbd9fe63e24eb0fdf60fc4c49cded12ff979e9a9330f3c6b342c633c07e06e63ad5d1b8fad7494f27ed2eb40b962fa8e3ae0602dc2d24653637d1174059c9d232348f54b1ddf6db6977f4c28c52bab77615cd83afc1d634732c190d894f82;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1598e7b90c21a758b135958b562a186da7842beecf4b182accedba12ce1b71e855c486afd6f454b15c09d0f1703e7f0aae72afbd4b75e91b3d3b99e57bce421b4de1dca28777dba7886a2229024975cf47d092a28adba1bcabdb68433f35b751c284d171a744270769b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h14c6d4321d5344c3b8b856aeb5efb8c65340bf50e2fe2a0c8f05440065422a5c18912847140c87063a4e40fa6c007ad8b1b0dc266d6930a3827891a6f128c990ff72de616eef5e09e4403ea110ca64c1268b52ae346b1d2c075aa093d5c7523ec86f4b3a5778718db80;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h163a3ba2c27e210791771214495fc0e4ae8c7ce3c6a6b272250888e83e3c37113947adcded34e32d8b69ec216fad6625d2042198d639f56f24af858a6c892c9eed7fbd22f93ea70af1153c972f559330753cd7271b8d7f06ddcad5924ce4445387e81a62468d23236e9;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he455ca21c095055472e4c73fad92f1cdd615208c60d9c54eca90f9cd1388e35a368d68fc7a8a17e8b0a335b445f7065d3f5af3be38fc478c1f17878454dc10f7349f9d45ce32c9c1cc0874dd28c744920feaefc8d4e06f263b5337c793fcb9eef30cfc1add1a2804fb;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hffd05de6eda9056b1d318b3900ae2ecb3afc123834452d1b39d5ff48938385598809995205bd5fbd47d899613fc246736eb67dfbb989ba42e0ea0360f09390aace30807410390a10bca8c7925c443f86afa7e8f4b7f02f3f9f015809b7bf1c22e9d520a68f66991828;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hdba2fb0e2912d194fbb1e7b121ede3f3e7400077426597312bd777cc465a2deac9709d89c9a077cd604f5edb52934abaca677ba2cd2d67633d381fa35116f804f71b026d786ca064bbe29e052b5f4b96136db2e3980bc1b7f0482ab483c675f4ee0e196bcd894cf15;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h2e3a4f3d2cd922509441c61782c3adc2799c056289f3835c451e6d066ac8ab199c53f7c7202a66a3b1030545ef8ea953fa9ac16042496a3b0b0d7eaed2260982d2df78dbe6d3d8bb77e5e2d2a7f728ef10646c38f05878b1e16af554021017b1b8f585d596ddf88bde;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1995a086fdf25fd6d91153f7653a99241af4c6893faf1c5617faeba0afe49d3c82fed8d8da610bf056704bdb3fd30966e8797160c2eb6d211b5e507b9c8881ce6fb0434a3c823a93f6653e09e7dc5b3099c49a6915eade37e643f4754648395c5502bc51c1d6d481e84;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h7bd33dbca1c0f3bdf21ea5bb18415675d0e36a147526a9901f93e450a0b979c38c82aaeb30144e2c175cabeb273a0b62d6914d0b27d387a7506a38111d635c25a318ad3cf939ff0754d9329e5afad9dcf68af461dbf72fd4002fd89d6d243b7a253cf616fdc9b11c8d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1aaa256a72e20dca26550a308c9bf372f7f32340a6bf2893fb15a9660eda0295e33af072fc0b070c4912d4720486b267069c87f8033ee3d554f6a0fb35fa6dcd8b296fbc7d0a9e6bfe893915096c330543c24e77dc07331b9fed7900b71d8e4e36601ffa76ace575817;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h8d9ea3171af5a125fa6cae37eecfa10a32481c39796ab9bf76e3392f621d4583d3069043078734ab679fec383fac91a054f7d4ab7b1a34bf4832ce681df13c04eeecc40b58a3fa5e6437c45bbdb057bb20c4cd002ca81df15f3c2419747f8998786b5997165dfead31;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb1c662d59a70ed41064d4d47e16b22849cfd293115b4a41f391294d755fbfc7455d7a220e86fc78fc9d8a7a1750be910a51442d8d05be7ed0d3e0c9f2090c98de5e4c5467d80608272619a4fc3d8abed43262801da3af9696b66f590fc4f88ba2cb1fdede0564ec33e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1bff43091b9c70ededce0be23c94dcd47d375254d5ae8ef0a233e748732d3b9b7d8596c284d5eb6939233a8173ecd1d51c905796e50854cedb1d3f4b8d8619350cb94cf582c868f14ca14101c04298db86dd5b3c7bd2ba3ffe90d913e8d2898be4783ac73041bfe73c7;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h103ff5bd91c1fad1c82d372854ad4b0cff8a1b5e51ba0ee0a8224d3faf2150565f89f7c39abd6d8066ff5ca7b6dbf0db49dff0b90ae562ba39eddd2f6f982a02702d7f590d53ceb4224a2948b109449418f7bb571bf2ff63baa79bc66fd7cdc93225f340afe4a85795;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h220ee775e4fd644ffbaef4b7e99a68da15ba770aa1f93a38dbe812fade768e0eda28f19b3dbbe8dfd286f91d388e4468ab0c050c2cdc00a1fee452a4b2fff786ecf48da300d2d8b590f1b74f8af3330e4a3c574570373537205c40e842167abf07b09b43b4f2ebfd47;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h18d31f9801c5afd4b99df2576b9478dec2e7d028bc5d022daecf4f7f9cc51768ceaca4be3279b04faa1f83928715b6b668c9df1bef6f4ac4d9dfa7b05ee4edc9f047fdb8db58bb54bffc5fe8f1a1ca5fbf22a16dccd48804b952247035f7e21e29a1079a2ac395e4114;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h13ab19780d60a28f7d450b4cb4d3ae325dd922a180bb946869e99cceabc799d674fb2d9d1a1ab6263370770fe07d716b18139c57502fde62a2028f371d96e9421fe092f0a23eaa1158c83ad1268a9024119acc06aee3f7c9499768913e07e43f755ae6c808df498983b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h19be25113982b3632b04f47479418e0e5f412f77cdb29a75feef47540571c82e3366760880247b2160e40d8168c2544fe716b7c8be5c4408c471da30b03331a8bd73ea89ff6ec1d8263cb79e42e1e9c5cc2e48be7bd6da5bbd46bd68c6d299d363a41ce5fc2ab1a0e2e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h16fa8a9dca51b58103f8667e3c0ad2d0d335605598369d050ab42e4332b9a2e8bbbdc5b556330bf6688c7b4a3f103a45e94b26f9118fd5a18cf6827bbec40bacbb66d8cc98fbe0d24766822fcfb4df2fd851a0ec2c164fd614cfcef4ac333cf30e9f7bc336943d969f0;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b06058b8cfaca177ab2e739385c345d8d8897841832c08d49b381dc38ce371a2e2c61e9846deb66ea44a24170518d657423cb154193bbae942d9199e55a2df6480ea5058dcd7ee476f950d66acabfa716897c36c6cc07105bf9e498d3bcb40e781a92838c4ce5a483e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h116ac06d7f3c5bcb36571f71f7c729861dbdbbe3a09864d6e4a2b726470dea1ec81e42bbafce4e6691932700edf2d5531ef3e3294ce6ec467fc9dd42d3ed71c85e2352896c8ce4e32c674cd08094f5fc2db668db18161cc7fcd23009c26630277ef6ee081d272cc7b8c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1be425631223abe26be8b35e7846697381eeb87aed8b013e768fff1a7ed8b945fb9ff6607dd7a228d6e0b206dab93f98152233af4d6497b93fae28741d47a2630b6959de71ab59057cd75498bb1d21be99a95bbddbf27657a68cc7350d0b702785e6178ab05e481eda8;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h19a4d187188a584b2563531dd992960948edc7e63404f67566a097c0ec845be5cb1d54b096d3f8ef2fe45156bb6e1b0ac8ee0c599d9a4f2683b8b18df3a7e39980b756c06011cc300d56c2a489a9c017e1acf33589fa945b32723235ab3240e2cae6ab47d997741f919;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h185ec1359a13988bba9b577a7c4349562725b47302c6593d352cb428a427f99c0666f142f201c58335cb382d0ed3c450ec3c2abb98539ea4bfa9b93159d39b5f36554d1723430cff2ba1aff0e5ab689ee6f3fea026a316f269c79e0845cf2e858cf5b0c8964801f910c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf02b38c7f78366795e5d6e2665e71a009bc0b124008b5869acb3314fc3bc9a8d68d7ab06647d24373480a8e84298b618c1b61a5eeb022eb990ac3ca52ab13b90383600a975f5289b9edde9c9834cfd18f82a8cce8852e93c1266e28784511e640df1e4a7f071789594;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1068174a0d4e77c9386ff7cbb0dfbaa68beb29cedb29936cd2fee760c8fb3781725b29d70398334dffb44215c0d14a422e575b100c809e2db8ed5c01a451e5cf0f469bdbf8d39fd720cdaed6ea2faf98dce9a01f160bb9de661b6674604eb3deb44fdd46cb1bfbc62b8;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hbf5663ba5b582ce92dc63ab8dcff3e28fca0a006dad351ab8c27db96e9a8319335b725215e8c348e1704f2c387265c269ea7822aba819ba87faea0a0b64bf4a21a95ab90b74ccdf20afb728b839e4a95dbae38623f72427dc89d13f44e413b30f32c63b2808f3bd610;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h16e55b95a99262a94773186b32ed78b4c04913e5a72ff4dacfcf2a5548c7aabd16da5e450353302843a6a1efe47b3364e361144c7a16c59e716e851bfae5e2e0d45afc413a4b3d1e203643cf28f6cbf0eca61c9253bcf8a6512a18415605316eda80688dd3c30f83c2a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h135cc4845206b2301d28597ab6f290b17842c3e0abc3c86a5150ec8b618db1f5b78af8ec13e75ead1f883799681ca070d26dca3e5b200e1492d883cb545a396fbe75ffdb57ff1010efb8b9961792fbd6702ca6ae04a4d79c2a95e945269f0256344af56af19b9ca1f17;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1bee9b420a467a6054006fc69aedf45e6215f9793ca0a6a67e7d6ef9821823c3452954520aefda7bdf256ca1dee3cacab298ac703f354eb186cb113957e745f892da78888c147fd0a0ae2aae68b7fda2fa96478c144b26db195a5cdde873d7eba58389208fa9d415de4;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha29ef1a4118a42c64e06477d3dc7b5622b569c06f14782001ed63d7ad1c3134f9c74c7ec0245db65268a0f529971b3e83d7048a29cfec1f37b41fa488984b021fbdcae7fafe6666c6e4d35b372f030d48c676067587f9d1faf17cdecc3f7f7ef09f0963e11bd894e32;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hff341328525ee3085525b1c679307ce05a0e772452e18ebed152e1c74d1f6309625e654d0d852ca7d4ba3ed73ae1a8acb9d0d20ca37644fbd05a842f827f89f1b1748917bd828b21834c9e4750a6f7da1b8ce1b7fa453a2326b1c20903bc4ae7bfbcbf1d46abbb9c15;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h6a253756b706a7eb71072a809ad3442ecdc895d6a7bd8e34f5e60624bc64ee1f61abeb0eac84a61772a88fffdf09be7ff78970ec1e2d31b162a2ba33a17c84800210c4bda2c2fba17ea724ac14286288b78500e3e739518933a2a2c406b5ce0f95d2913f64a2dd7f82;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h13eb04c5b1be0796e21eec0d5774174d372a03e6b3a823fe9a3930f18b4337c65788240ebcb5f8340e8e66c109143fac8822c218b3241d680bbd271a3973fc74df564fd31fba2a569752631afd5781b416bdbc15b53f8a8ef5a8773aac609aa7e0e06970c60d8bb274a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha275466e45ba22c804fdecc895d3eca72e23dacffdde4254a69eb138673851fee4ff2115959090c798b0e7533e3160db5cfeb750f03654ea59a48bf7fb51dadcb3e6b1a06affbfc1b1c83dfc6dfb87cda53c2f41db46c27692fab8a62d5e6640ef43f5d902b38a2f50;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h4cc08c534546d8aa7a50f358d5753844db794e5f7745bda6e394765d8987fad72a73f26dd44821557c7527f7d53a74280262b2a11e69f7e20c3a4a710219f8854660fc606c29244555be2ea6272bf92378aefbfcff304822a59322afdfbcf272edeed66c50a30c47d6;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ed85f868dc72dfa5ff644b6be46bd39927dc9705b236bdb12cc3f17d796cd614b1e1b2ae83e17b5053da4c6c17288c9acae2496aaa3c5e35d84de75d1d8d5e79fd81fd3ccbafd4f74075b2d6e13a8b4ba8b0f5532ba3153e9062eb10b46eafa290f481ab7491a89950;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h187ce50caf77299b688e344cd43ad5c55d9328b59350aa8f8064a5e816f896294c7b79f498a21486b3f376c770101a666eacb12cbefb511d85c0ae0fd29cb041840e85858de2d8f8eeed0a9e1401482043e5eee2a4e5e1fdb5d520c633b4b92b3003af5c36183be9d5d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1456581f5f755ec4c41b3ab812e77214dd29831ff5aca954f89ff2e61fa5b39a8881d871a1fff75707595bf338e63a82e3b0eb43044ca534b6177c384660b41633651ff8364d650a967825d8a11b792de435e2e562f9d539a84818b4ccf5625848bae4e9d2a2bacc625;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb70b9be178b61c00cdfe5af9795cfa275021ceec4ffbc7598cf57c7835563159ad981b1eae7fcd9a33fa7405424498491ab40235857e8a5b93e227ba84e88d98de9eb2edb5e9ae00199bf73e7f857c2f08e6681dc7700c5392e68ff9b810dc798abdc0d7e1549b3252;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h108d0c94eec1f54e0ac3f388441c1f950a19386f4ff0ebb546a95b43e74b919abb551cbea2c0885040e8a39dcddd3e7ea1efd28490cd19fe7f4873c8287623357980b16449ec5731d4a40f0ebbd4e40ffab6024bca8b3345891f77ec1fec66894de4e0a05d7cb2bad8b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf8311937e6c9ece328a511e988dc41570d0c122e4186882681a543fcc752d6b5cff1cbcb536d1b204e9328c290aaf5d09bcc87bb2519e2a5d5dfc143940e5ed4b491a9112d6fd1c502ca2d2b365ad2f824e6cf452ec9337aed469fa88b2fe5e6511b88e5cf73395e89;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hbbff543f79b8ac7ec6db99fc13e953dc8889df424cf920908e6c0dba7eb73e6c98f515b531cf8a09ecc8672ddf4152343ee77c85cae071b35f6cc038a40f0a1a5676336ff77df069b946abe5009449411cf056e1112cfa4d4284d51126c2348e23d2df8266e1e3c8a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d22451ed5d2b9861e62c54e963976c60da66fe52cd99803a3ca805f28f8672b2795f9df22ab0764f413f99dab76c0e2fdb8e82f615145f0b22d70addb60a165065f2995763d1093050dec42bc5a7e3727032a3f413ae1238cfdcc8ee2dfa54ee7b69b34921edb61c77;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h62cbbcedb94d4b84aade0e28f11238cd4820ae8f775b6332f87e55a97ecb1081a9b2fc6172de44506aff9789f716b4a5f447f3088608295e55f962a948242c882ae20cccb35f73a7487a8bb0de7a2b94977e54a47ea4d966b8210eb8c9a25aa26dad6c73796258ac8b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h3085e3f26e02c80796a9fd942914a04ec3bd70592bd9c7da4f3bd3d31b192429f0b26a8045a684855a9861ba4e0571441fdf644367d58106cb490d1759bfe4eabd9faa2e6f4f6a147fb78b133f9c2173ad3d4da31bab51df8c2434de71540265c838d3db422879e41b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h9afcaa231b561b2fa4180235f1cfafa4808b5d99226d47f00e4a50a9968fb87133456b8c104b13b0df5a13740d836e793c8e6f5e144e5391db221d92e92830747c14586531645f8a6439d1781b46c0c93df8237283f8387a01e821563d6b63a2a39e86aa08a140d32b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b032219f468412c955af1397ca20f95f1b7d27c692b0f7fb19969475169e3d8b07ed7877575d19e2f52ecc1f23dad7bf7ab212e9445d1484c9aa2845b56149c8bfbdb8bc3561ea8d058612619652194c5c6d09c9824429f599d88f31e8cbe9f6d3aebbfe120c70b4c5;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h6b0d31269554bddc51168ecdc46428e36aa34468282f1a16f358529807c9ec69f2576d639b6a99fed7d11e58a07e69a7377f71613101ea5003e76f84ca6bf3dc541820870eddbc409bea8b89baa25c5599d787d83ec6aad3628f15f67c962b4ab7c95c22871c263ebb;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h18b162c8b914f04a40f642bb364410ab5f3817856ddfdaeafec00b90f97b851aadf65a70646fe92366f11a98f1dbc4339c7842b00f6c031924cef529afa06ef95f10d403eebe50333716c23b4621a07ee4bf9b4efc7e5355a132b64338e112d0171689b72dd77c66ed2;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c67b8e5f1dd54871e6997afaf50c45b409c1dd84a0f2cf7b7c793fe111c377fbab987a31abc05caf79097abce14b1eb6a324c6fd118d31025c960e643ee17977714e94126b144ca3acc87ec3d76cec4b67c4dd2ecd4bc6ea34c9528adb653fc053490456ebce562701;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h182726269497338a124746475298ad872387008d7bd4b0dad90b209feb4a8d130df9f96fa42b208663d2c9e088646b8a6988fe4f65644f543093e567a2e9fe0dff98a17520d9d69d810999d36a54029e84a03983c32c5b5edb0868be4eaf66af9d32faf3eacd6bccfa7;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h8eb80cd12e0ce4000d6dd06121d7f7071cbc6d9f9589a7ec4ce0be3ae579ea74bb3002b7f6d3fb17fd70b74bee6081683e848d0f80dbf7d7ac54d96905d55a779d2d4ba51c51cb73b74401f71ee97e425432ad56699b7527120593baf4121a17ee04a2dc4b318afaeb;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h21eee2d423ad07cf01003cad6591ec4bfb2c08abf899b367299ce55c10a1c5c527f7c5044e5fd1d0ffc16a28baa340eea6cba1901422a0ff5d8db70aba92926a97d70989d7e2a3523d0927362051369ec24ebac9faa96e5e1fa95b4d07a3d755cf71ec822d6600a4ee;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h8e7bee2fbdedbbfba2bc076b9b37f0371e1a15e8787431983b3f248725385ca4a1b2060b48306181e99c822bc0d8d8689104e81fb2a216e05bfe8eb3b396a1a22bfef361356ce2bfc20712d85a92dd80a1f31d259ce92c24392dd3d0bb2966be61a431d52e2b2b667d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b4bae37699b6b38aef0ae98ad60848de6f6af3164b8915b4ca6ea080310f0c69e60036a7270c3830d4b8138e36e824f9a6227eabfd93c659f9cd2a62d3c5c1f99c62c6fd6e0093d66b18e8d3a4d2671d0efa8575bc999cb652746d8d59748dc9cf60d52c10d3369110;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he8daf483ab95d206b91b4d54bc36d42c3c43cd8988ae4042451987413d9b96fbe7b74527c1e77d1fb47d1999e1e7e9eb32d4e1906c811ce6f6c45904a5887a8ea58641f613c1518c97cb45af821f2532cb214642aea1b6dd947ea663d6d3dc6ccad4e26aed4759025d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1411e9ae85bf0b30e68e18e6fe8d678d8c604c80865f30f38112fffd2cdcdc0017bdc079596d2bb19ed70b8fa2030a22563ce1fce7f4ac98281d5c1ad34256acc25fc1d161e59dbfefeb0bcc0b2f6a4d8c8ecd64cc262c614f669b99a94e54b99250f367d2528625c56;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h19305f027f424a78bfd41da7c9a4964175f7d584b234fee04921fc78c4fdd64566cd75c4af123d1675b299a0555c06e1af4fbd22f8a4a88010ea1bd5074fc20c1c34035ce7181677ff062358a313afadf9acd497e2b2a1b74a0c9c3cb3890e49900c8d4d3202283d195;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h161f6691b295b7a65e32b70a4e6b52061de18c6bf8148cc8640dfc6f85799465b76f4028a1d1572280827287062adbe1f09aaa192e1cecf3db9723d00eeac176bda64feab3f7e4a15ecdc5e5a127096a627cea51fdef1f411f299d1f8ee5553102e972a6f428820d525;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1142b1ab1022885aa7e1443d0b7141727a9fc451122efd2d887a12ab8f365b19df78e9e9d336a7ef97c983975153b5caa75b1f9032a8e0cb6c946960555864c316b5477f2cba8654b6a7d766bd3ad2572fe35d5d8a344fc4f6fd8a5b92e7443b11df00a564542628496;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h53a0e083f29264088b54a8880533d82f817c13ea196cd4e5df242a8f8706ef7b691843f84493ba12ac17ebdecaf2dc36cd0171018f8cc5faac228037b9cdeca331a3ebd6e646935ad372ff8d8b7b0e5cd3e15037303496e1e4f85a51859161a487f2453e980c0513dc;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h15a3445822a0b5017f9b6150241f24b6afb0d3a1975d3858ee61568c7f052ba92cc4dc6dc8950798bf74a354142f3d754f6e4420eac72938825ef202940984bf611e40afcaf4acecaf7fc62c11296026dd04b6db8b0f88772700532a6bdffe125841f9ce964f2c0b7e9;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hcc162308dcb99b80f1437e4e1dbecd1e4603f4468ff5ff37879345a04444a5a45c45acdf71ed4a006d59c49bf227223322c28700f89cbd301d9e968422845dfd4d15b3a75b9fe73eb0ed4730bd05697ae748ae2eb2d78f3c4010c5a45ebd0f37baa3ba7a8e12c9e475;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h11b48072110a1d3279228d3f7508eab1232f4cddd2d2fc2d260526fad659b09351299514f0be1123edfe52c7fdaadfb1316e63348eba9dcc48eca4db9bbe75128d5b4fe98bebc7ad9bf438b927512b70ddadfb282991dddcdb867d3bd32dfe354a2871d433bca8580fc;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h16eb3d97e05aa38d80217f311148f3c18c099e819c3a9b220576c4d82bec71b4af4bcecc7a6ae834ce550b89ef8b5452743b8e146dc7d424ec66d8448629e2b0bc4d54f1b3f26536327305546cdfa1456a1533a1d3cb45946b803b254cefff271830e5860c99736dca6;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h64d2fd4e501eb395699352e6e985caffbe882448eee735676a9feaa90d25c355e5dc43e789f59e58a3f05b41590f5a5b3ba726bd2ea2e17c6c6e4a552ff2b46b3e1d404c4bd0cb7e66b983ab3064727bede43b321af859f801575fe45b91bdf105316dc32b38c7ab53;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c563c89d3a28157c176bf4fe8180de615c5fab7055f16735ee2aa9e0fc9f57fd869063f6ec3e02d77b0b9abd79bbe1dc065fae1be4a03665c6301e18f7a6ad50786d399cf2e6eb619e48748de1fcfcd0db461fdb230e8c4627d20b00c02c25886026cb7fc993f09762;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h67f6f4ffd8d9f08aa99c9efb94a2dfaf8abb514d4f913378e925bdadd011adc30a28f695c8c477cd0ce2c816d2bb1e09559b3719f95c8dd43db23f5294cdfe04667bb08587c3eb4347873781ae2f36b4da2968807122e6173214bfdea2d839fc7e37740d5416c2986;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hcea9222121833b4491906b4fb9ceb00703f235166835aeebe2396007a848bd0dc7318950e39f240a4ec4880d38c99b920594c3671b4e755fec91042e272804120e50974f99c4acc165852bcdcf897bdfa1f1dabfe85d3a9e205db8ad1b27ee1c1b4118369e111c7657;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h195cfa5e530df6a5a70c35625c5d0e7ac17be8d0478dd24fed7aa51d4f52566fb77c38fb0ccf93d4a78a7677e81c5e9e204e87a77abeacf2110e2ca08257805f4c4e9c44fd1dd6f7495991f24b4b2a6427611ed63746de543e1f29901033ed5548e37b2e752c737c863;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a91bbfebea9aa3d192396303c9564999a8b75d51654532087c4d199a41cff0ffa33f4127c19b750b43ab18966a28cb3243524863ace0d38804bc9c1a5fd893781da52749211b5036fcdcb48d265ebc2f607d3522be68e050287bc19f86196436d6955ab60ea3bdbf7f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d5efdea20c14ac2b88e19ad18f6af26dec95a4fca31081ba59d325b86686fb58239bd1bb97be9481648c0de47b2713d95f99ee78309f934ee080e86368df5f931b80c000d5796a63213765d53c8df5462f62f3f0117e88e85ca3f58df8bf66e8bb3f315cb134e89f8d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf56568291cb2d7dd0ce369d7910244b084187c8878e00c746ff9cbe35ad3e8acebd5e00dd0874a8dc76e95fe2b89a1624f621b14ece5a2fb8c80d63e9f444a331bfe588b492946889859c9fdbb349f2f96ddf8fc65bcb4c10fe1e6c7e539b155e597694a0ba9470d5d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h5ed948efb34cb767de47f89d4a932c1b257b43688e6baf212534ece196a3e092c4c91278468bb6c1261c5e2b7b4dab59d1b0050ede7de55ada16bf0b21e048e8c30154d2f885a1826d3ac46c815fb4a899cd8413dc54e11786df64ccd686b43a44fe70c9af07876d64;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc8d0c00fa056bf61b410ef7168ea05a9c8e874978f70535049bb70261e96692ee46db00160b60f27d36a378ebb41b45325b8b215a7461fcbeefd477e873e121c23cf68a5e6349cd20da9bd910d341cf6052c1063c72f279f33752dd412450c7d49ce465f4d773f4998;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hac3873e989a0650df6ed26d96b1c2ec420723d4ab0f77fa1a1393698a23eace3ef833525741d8f484cc1fbca6622169c25a9b5fc7052d993a7202fe0cecb70a3385ede4ac7f528ea9216691ec0bf4fac24a29c128ee23bb6936c19ce9e591b56fc25f051dce664e86c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1aaf95f52f7b2d165546dcf60f2c8cdf40e68f5bd26f6674aa343c3642d313ce3375c07e122d61293ea2287173273aa2ef20a88888010eafbd3a4f9a10b9faf19653cfe011a840c1df8b8a0ff8fa2f0c5841251f6c6478487bfbf2472b9f553ba73e6c9dc64ee976b23;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h17921f989d7ccca6940a6395f8469dcf1aaed7349a68c593f0c5cbaeb819d30ef65eb12196a10cb50f393a25f1d889c86c0a1956cf96e43cdcbfbdb92bfc42513e0b5ccf3d5b0788025d4fee755f3a10f5a510e302f7f831c3f18962db99ff5e1e7899c2c2912e2e1b7;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ebdb83caf847416929182291e2035277cddfd73c9f8f65eb35e2eef1f81dd495293aeb2b544e72a79a40cbcb681ca34218a729fddc922a8b86c16e483027238933cd8ba3be55a7c03bf191559efffddecac002f71db66f0c3636bce5cbb7a4d22035918bfd4f9e1b5c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h94b78b4b8d9cd7a934d31ca50cc45b088e41da97dce2cc60b38a51ebae88a4d6457c3e5beb6e624ac54165b0d048c438fc21bf88c9f153b94692e1698300bb799f98773778767b8c901fa46b18bfabc8dfd3efdb928e2b987e0c5dbf2fe969afa35647d429a74770cf;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a1726ba057cc5b5de1b3ba9f870f1098d3276593fc70417542dfa28182444eea8047cf4f7a96570e0509c5e9703a71c633251b56ef5caf72d43740d910fcb6fc8e26587d0d97fb4cec4dd398680d423bbb05b0c054c28dc2c1c2b0cdb4fd96669e66e04ecc67bfdaec;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1230d4dadc392668c58831770054ac5838a3c74a629a7d3476cfad23278028daaf8d3965ea3c7a97c66065615ebd81a953fcc522039a052b3a676b4f55fb021243b6426d27ebe4ac38f8e4dededb13e44eb744ae2457f7f804371c82d63b1b3731748a55b78b7c47f56;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h14d6b240bdd366412210bacbd57c66ed0a6f666b15fd6e8af49aea4f83361f2276b4589ffe46cdabf6a0e88e88746c0c48595982b0807354167bcaed23c6c439a752b0d0bf2579bc79331ca9e078267a7a45532f0e8ef98642b5e843c5e7f4a15597f33341db0926141;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hcf813b6dd97b46a21ed304a0bd02e464ee5c36e2054e49f75733696a0961762517d790938b017c502a196a620c5cfe6068b1c1aded99eee2cc6f55b7c35cdd744475d56814011a10e01523d5c2796f287e364da843332b69cd9f692161fead9dfeffa62834b4bb99e3;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h113da749ab00f61a85013ff30ea87f4a036eb930d7274392c7438acb306b043cc98224c30f65bcdfc634179a34e1b28cfe38e12e6e324f1db6d682e8e7ff60cded32b959d3bd40fd904b4df6541ffdb32fe9f978c73f7b72946d4808083c59a78bd098817f8f8fe824e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h5d43e2deba14ae7d180bc22c2b400c73b89c187d60f687d676f71c16ba5723987193ae0026d2304778b570c67a8534ac6ee3729d245cd180ffd7a2e36b036fdbfc83194526c2ae172e69e69c443eba76f74cfad29e25bf39a922e76fcab6fe36dfbf5f24f6808b256b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h113f1919f1d5b4f9df877ce328602f76e1d848cb6ae642294db05d681b782e648346da8e02a8a3ada009ca19ebecc4e83e14af4192f791948d89f58a29526bb651e31bd5e04c72416d4a8e14859cb39be8be66d7658e5cf34252ef4c21270a862a20cf66e2f1960c33b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h5bf7d5782adeef823893c496e8e0e9dca5386e664c9b782a849ce7859feabbf1d89e991b3721846db7078415c86b5b2c4b95c4f50a98484d340d23be8333c54b19376efa2a22bf21a615b09ad243690ca862798d01ab58614035dafa6b09dc33d6a8fae3721ea5dd67;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h19421682ca55d0a8dcbe7e89f91151929bc2431d6bb00c5f18eb2ef94e7de549fe0596fb41fa84c0b711c52efcc0228774c5bbf7e0a3e4e77d0dbb1a4d461f36184abdc32f667b14c996241b6a511b56c5f081771ffb9d0f2468a5d1b3a17e3497bf682c51119a75cb2;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h158e2d159d84a926014e8b83cae6b774e80f396ae39a0eb9a8fa76bd8be6ca94d1260249ddb190dcc92986d10927f5fb182aea078dbcd9f5e5e8c45ff790d773abedc3b3d8733a3df2a54321d0a345a0ec3a2d5b1c5905d0c7f6e504651cc99b125c24a43b552d281ba;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha748bc2bb27c2f5d13ad1c8223b4ebf99522dfefe93e18c0e8657a944906dd9b49ecf5eb0e97e21f4a3f38e18b6520900c5fa7e2dbb994734c906e8202d62bf84cc826011215e78122ee453a7e40fa518d3802a1c44066859c3664120d4f9eb70464a49e9a21f72530;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ecb062ed6bdd618ba5caa98716b7fd26a807733c298b81a5a5a950d6672f7fb8b44f2a6a1f28f09a1c09071bd0853eb589107cbf082f22769a1d6e94a2b33fdda154834e48d2b6e02ebc0473203039bab50f33be7a6c5773ff50def993a19951cf30eb4ed39288985e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc373a4455e7cbc1e0b2b36e91d9e79f0664a194567c129f4266a9d302970a6f4028cedab534b17ee162d4aacb753d962bda173e8945709fd5b30a94266273e09f1b44bc6db9a5ed8ca9ef12a0a07b826f0e6c6e239f4121e90a14cbbbfb039df8261ebcb909ce139d9;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h9c7fae4139321d650cda5b60ee137ae5b7a59d658390722567639692925d0268493fa2ec3cff7bd202d8c4cf9326a0261cc646550a29c2c2936bb1dd241bbf09eda5ca24a5d0abed08fa830d54678e4f86ce10ff3982861dd9f147721d0116656916eda3fe81254f69;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h6b8796bd6e633a566304e0ceab2a77874c44f6f0daab8a8f695a2c138a0d6599384a3d0d882398964c6845f98711350414282193408ed2e9611adfaa28b5c0c43514fba031d490ab09d830df66f1afe288185a5f1113894117eb087c89e73c7c9f5ef5c24b3462cba8;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1380affd01f1105bfa0df7ace0fb0bc3918ae7da7a6f623ccf0bdd031216e3410d241b4a19980b1f93c15238873130860cb1e97b56b29726cc44f7f317caeb766834f75bbf98f9d45875ef1b3ebeb92d0bbadb7b617b2277136fa690ce1ce8cf225a630794d4992953f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1058287fedb9d98d5bfa93f4de2dfcca781657ca679cb574feb47c12a1527f61d687205afd0b1b8cdc14514d40717d9a0b0a6535efc2d8641abba1dc13a3fe283a4ca9497e446d7580b6ecce69f1d6eeb5b6b07387f357b97249a7c098b0595f7b85c91d76c3392029f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h17600565c20967c9cee92e1c9c9d66edcda8d2100db456cf3435ea949fa8fcea09d8740abfbf4784544c786bad3e73a4cf0b6785862c923cb225c421ff59d17c3c40f23bf586a5dad05a406ea0a5b5dfaf425bcb4fd3f48bc2a3aa7f933ce9ce7ac7abf76eec81f3ef7;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h4e2465f8b3bb4551437cf3418227882bb3a79fbbd78755bdcd0bd9574b402079dfe906b5aa5c8b359e81b27217485bd135bc7b93cffead47a184d9fbcd8bf9f034e4da41fe100e7e7a3fbd0a181cce8ef1d17b1bbabf2d0deae47f7e28f9293a104759f59d932e29d0;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h668970e28947e17fdf786182666ff8a29be0f55840272a88d57cd1c9d8f877e0aeccf0eb57e88c4f83f802a07adb641df6f20449cccfda9867546ad3b4c859f5ac9c7eb64909a0d39fcc8d2d11065bae53b22c96ee36dc76930cbb32bfeea474bd0c9879aba314a3b7;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f89147b456a70007425b85d48498f92696d48c4ac0390a36936dda3abd375563e69489ca0c29e3a23cff15b6bd703909c434ca5a7f8e161f983d2424d5aa98371c5896e91c0a24a1785ff611f6750eb3e7950f0fdba885b5d370ce5ae03e5a2a98ddbc89e648cde591;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h41c0eb4d2fbb97956b6cbd05584b2dacf9b46a3c8c24cec14e7e65cef551006f0848ea3bc49cc53571530705c90a7738c52df015407937104f60d62c7419ecb28947296d474eefe889f6b53193c926462250d5461f052385ea1d58b8871d1ba4a84ffb1ef55c18826f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hcd49e17c06775d4da1d5de5f0ac1486494e7e8526a7a5605a4b5d9dab835e7a218284969b8871e76be0360ca68f14f525a037af2ba28dc2d50a4124ac8c518b02771683d1d9dd794a18904cadc40d2521b6a67209085fe098e5a1f8a74b54bd7130a8f978c172bb68c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf79e4c6cb12cda7f4aaa61cd124abdc5b5cb9b3a9f3c6be80ff71da5afa1f70f9a50296856937783c894da508077afcf5d8637283f12a5866a7016f62f3adefd5a2609bfcb936c690821b71b677b87d8a3097d1c10fb85a908d91ef8f0dd8285e66bef90f6f1cdc439;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h16d3f97eb72aa61711a1d8af28bb602025f3d7e1c79826c41555e5cbb362f243caa955a8d18cc4ddc4bcb96daaa96e19e1139584bf43fb632c5f7f0e345bf77b52619e7be38e737894047f3ea7b6a37301985db982dbaa09405873ae028cfaf0cf72e95356a035b56bb;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha928c2e9f30dfccb5c91dfb14ddf4b1d1da50b4003bbd676d03bfd4e2ea5f10b160f87e30800801d9bff062003298f966cb142ff6a3be574414ae5b5569402e39f183516128ff6cc39972d290d76d428e42cee14e4b9899bf5f33dba701c6807e73e8beb3b02ef35a8;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha5843c92fc8e471d6117c52f46f9afabc6401e25e1626ba62a0b70511cbf3106a1df5f22c09b378156f2318f779e53c8df327959b1a4ecd4923a549d3cfd9b86c27ffe77d3ce9652db42e860bc246223f7c87e3e412d59010c436d78ebb1ddfae65d79947b850db5f8;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h13358fdd9c18521c1958b16468aefe51cd0bad28755eccebee40a9d9fe92300afcbb70e8239a2170855a063c6a36dd996c268b6c042f3423283613197ed0a266ebbbad26aa3ee9930dc71cf16e5b555f34cfaf780fdc5bb59442b4cde77bccc854b563c85c2c6b6d16c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hde898d6c5d21ed5ec130ad0e6595e02a5c00e98b9bb56702aa673b115b9553e7f1014b5471cb884f02525e806acde4ed3d0ca48fccd101d27a1601b6c5877908f51d7957329dcc210a2fa0b9183f6bfa9f595f4d3175d44bcb3ee46902f2bd04feab769f6340c30ff5;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c29ca1982e4eff522d94d8a3f4e0e08dd2209b7930fc220f2e4eb3122bd4bb5e3dbdb38e76d4ff4bc53d24f3332bcbfc6718c8d5403bd73ac7b36baa8e3516f1d09b623b3326fb70c48afb4f5d11f3d419e925efc388e6355f8e6318426599615d929f2172397cfaee;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc08678e67df1e5db445e7bd52272f12ba904f357bb63b300afa7c6b83c89192f810a058233206dc3484a54256148706d60251d930e876e98a0f894778c78b1fc7591cf205baed2a3781675d7d31b301a55496bdee6054e8d7ce2d540445053d45a28c27a9e6a169cf2;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h186082edd0697b7c66675505da724bceef802a99e2bcffe98d7f128463530aa0da8edf269a4f2e2c4c79eef938a6652d204067927ae4753e6e77e0ab74d417c4cfe1869827fce427b60042442287bfc5aeff1275b2564b449b33c08ace62e261919a35e01de89c844b9;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb17449ea6e112509f2ee7859c43dd2b67611832f36c3f85a99caf50d4b8827be55da69c8225d3b17a19d771ca5c67bff143443b4a434d6675e34e678ef95bda7e08a9c298ff5c459c04d25afd227c0ace4cbf47ed90effad27685dfb19c4b4a97f8679d2b7b5b41841;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'haea819f01df41052574168d099d7b1b875fa20466b5d4fb985590d83fce898ffb650bd2a7e1f6ac5676679cbff5b1d74c0bfce423ae9edfc3210dc038d8558324ea8636167fe818251a4f43643c61609d84048f77e353f68efb0434808c2033eaa18260050f64f506d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10f305c77e727feb53377ea933ba8dae107e5a9c99023af71e4f18d50b71e5aefb63c600e0cffb16edbe4fc5c464980bef6e38ded538a69c2612f6dd7a0a77ee5ec80a772382386063f808578d7851e78099b0c1aad622425d7fb4ee0688a4da77e21d0876b5f377e85;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h19e5854892fd57f954b17a6ff53b85cb6b72a6d728be9d85aca0fac6e59fb7c2c7e0b89dc3437f73905226ac9846f92eb0d3efc431ff01b981caf2a2c55373c7d95e91cf299de9f10ec271e1b38c11c98807f053802ff758b7598afef5b40891632ab2a32eb88c05833;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h131cda5d2a42f2d64fde496043ae8a5d6b329a8a981cf5ca7102df161b5bbf49d433f1d020809751c38c2672092e4ee6cef7db1cfd3c5b42ab3f5dbca978568ccbae846e2f0ea097d4fb8c8a52431516167a4b28bf2e8ae53d18bfb3d93acfe3a62602246382b700d76;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h200c372d3734e44313ce3ed38d7a8d59be5ec863d49ea479552c2bd87103e3af12877b3fd413f5c4838fd1b074fb8353c3afd06ff9bedb4ef15f104c3917b90fbabc08e914e7469da202330f0a200051dc6f98fc9a1a2772548f30f6b125f64be0807a558322228af;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h166a2140288087b5088af88f0671dfc3a9bcda453a18035a7614985b2f94d7de6d424538b15dd216212954c7368d293a8e3b0647f9a7e894d5576059e1183531095c96230ff44083316d25848690942ec663785c1933cd32f86def596ed7ad532a69fe7526da15b89f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h9a9e988f4e0b2d6241da88ef20bc8184956779d6a696bf7b635eb7f36f368bc4d245183e36dae5fb7b2c85f80560f89dc1c596d2da6b190e44f9860427e8f3c5ee188e39dd4e2a3598dc4281b80f5dd6ffed702c82ba4d97e7c003144d85366c2383151c22e68b22cf;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h9beb67e1dfe1b720579be07f9d200770d099c90716c35f8df2b8cacac0d9425c9ce68e35fe2f3f401701481236220b7890bef368eb17a543ca9ac7845c3303a2b8c0a55d390e41211cfc5e00b722d068dd23e6d4b849f680805751c1f86daaac0d8570083c3b4e5b2f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1dd381f71a37f342723f79a347544812cd6fe3a9ab3593fa797b09d6b5a9059c669d9dc7e94563728cda855186d877d3db9d42174d8bedf9a1e6c3751c8d0cfe30682b889a4841af452f58d39b60c9d9d2b86f3365354e10a5d24639900561896073bd442e42c8fc71f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h84276509d4dff7675c618aa91a750ac3670aae45c39e37e134553a3410106a8f52d286a8d3346538567054cc2efb992f2aaf1f62bc77bdc549d61bd758d86afe8920ab5b241b3c8234d2bae627da296fd8ffce5bade2600de19a6f52744cea46ae3aca665d1e0985f1;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h147b320e5f01b427219d9dc0aa4a9a1201bc76ce030287e9b393012a61552868cbd3d90d33bc7eb507d3b3c2d293e6cb5185447d46604da56e2f4c8e564b51ef9f80ef53b9df980fd2c2d82a0fd9ce2d39df98975fcb82bdbeb29524e2e98871d7ed95890e209bb5a16;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d8bcfbe6cc8e58f8731e7d74734fee4bafd7a30ec227c5dd29acfe2906ea0cb1ea968d7af284f93a76e1208758ff6caa2d6c282d0c562231db6cbdcaf995d63b1700b8279ec0968628fd3e039b4e8c52b202df9fa3cc3a82bb058531ebc77ddadd3a40d9c5ce035635;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he1d163b59eee72623b4d9bf8491de166d58b4b6f441cec4b1cfd908377552130a3c286d125a171fd3d2aec431daec01df490204a05cd7d88ee11cb3f7dae4c60b111e48faadfdf7fec16b941512ab0e398317dbaa5dfc77531723ba43775864841f64468260e8f69df;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h164df1b183d855b08725c2d37501d560e8f6107987e5fe4b3c8bd0385426e74a45a806eca85980df114dc2db1d02a824bb6749fa8b6b1eaea3feed7df3efd6b405614a6ee9dc3d59bfe38f4c7c4084522ade8dcbbfa7aec5dc636dabe7fa6c5a9433a67d5e7c6452f07;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h6e8246b06b9e8f334d265ab15725c0fc5fdd797a931d6efcf14b005c6ca6d07f67e6fca2a45df2797b6a8f7a72225cb58eb665c1f5cabae4292db875acff2695cff2aadef2b354a061bcd69fb5b3fea8e9c6c6f48807622ec7d5e70ef56fcd5b5283c9fbf10331edb4;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hdc6835464b5231599b2c0e92195860628b34dd5a56b6d103864d7705f5151e2a2d7c3ea4e0cee481122bb9d30ac0ef460bf7ae9c60cb3f3432bf04476a28fde50e0bcbef0eab2257e68fd46e31f7a8982aedc58d391f8aab8c98734d7a75d64fbfaf801b39abea253b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc71e6f159e0bfa321430a1b77009f1b1a1376d9af7b2375d2a85d35e7c7bd317ee11a68687c44b7a2cd200b6351c37c9dd10ec3b2900dcbe0384e849fb9e827d4e7032ca5f2970778325607b6a24b5b47cf66674991ae1ce757c86f38f013454d8c143db990e5d2567;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c25835a6b05c8bc7aa67fc6c0d6defe19acfcb6a7038f27c1afe5335ca3790870a97bcadb38fd8b5e1d56da6da95f15ac0d04156d898755baa78d7fdf74fcfb16c2e66b009f65ab8f9119a362d3b58ee637b543e94d4aa7b81fe056fc7a9648310797b76e5e9dc50ea;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10a278461a22dacc62d7d7054fa234e0d93ab1d20faab16dce78de3b26ac2fe65af9a21ef9a1ed93b1d8b0418769d0ab9df068ef4f1b42bc551215d44e63043b355a4811fbcc9e8ef9fa8fe4ae136fd975e1be038dfc16c0d61632ba9522a20217175ddeb08b7999550;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10493f2ea42246eb4f40ecd2d5ec4599ba3206b4c4b3d71c1ae7339f762c3117138b10990418bbdd66f126f19ff34df97ac798537f9d9240dca1f608080e29e3900c453a8563b978b0fa509c5f39c54d1a1599a453e7a71414a1e80f041a66815e01e59e4b52cb531b7;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1acc5a6ffb4c80480e0a3ba4a12238f31f611d5d38941747cae73ca794987871ca2db02e7da0d7ec77a62df57f404056369262a255a8cdf2713e9ac82649e923a55d884ce15072277ce4e4fb7f18e0e8a13dc27cb463af44410377ef292b2a65e5407760396f1bdf1b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h141f6c03eb4d4a7db52a4673d477581b31ec777a9c15e46bb716010449ab5c92bc596c86664fe930de058db123d7626b3d2ba065c13a0ac17eac445865bdf51eedae6c1781addb3a691c3dd71df21973ce5c8ef19d1002c4070ec07a947523c7f61801f0c08fadb8410;
        #1
        $finish();
    end
endmodule
