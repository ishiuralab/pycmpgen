module testbench();
    reg [27:0] src0;
    reg [27:0] src1;
    reg [27:0] src2;
    reg [27:0] src3;
    reg [27:0] src4;
    reg [27:0] src5;
    reg [27:0] src6;
    reg [27:0] src7;
    reg [27:0] src8;
    reg [27:0] src9;
    reg [27:0] src10;
    reg [27:0] src11;
    reg [27:0] src12;
    reg [27:0] src13;
    reg [27:0] src14;
    reg [27:0] src15;
    reg [27:0] src16;
    reg [27:0] src17;
    reg [27:0] src18;
    reg [27:0] src19;
    reg [27:0] src20;
    reg [27:0] src21;
    reg [27:0] src22;
    reg [27:0] src23;
    reg [27:0] src24;
    reg [27:0] src25;
    reg [27:0] src26;
    reg [27:0] src27;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [0:0] dst26;
    wire [0:0] dst27;
    wire [0:0] dst28;
    wire [0:0] dst29;
    wire [0:0] dst30;
    wire [0:0] dst31;
    wire [0:0] dst32;
    wire [32:0] srcsum;
    wire [32:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25),
        .dst26(dst26),
        .dst27(dst27),
        .dst28(dst28),
        .dst29(dst29),
        .dst30(dst30),
        .dst31(dst31),
        .dst32(dst32));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13] + src0[14] + src0[15] + src0[16] + src0[17] + src0[18] + src0[19] + src0[20] + src0[21] + src0[22] + src0[23] + src0[24] + src0[25] + src0[26] + src0[27])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13] + src1[14] + src1[15] + src1[16] + src1[17] + src1[18] + src1[19] + src1[20] + src1[21] + src1[22] + src1[23] + src1[24] + src1[25] + src1[26] + src1[27])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13] + src2[14] + src2[15] + src2[16] + src2[17] + src2[18] + src2[19] + src2[20] + src2[21] + src2[22] + src2[23] + src2[24] + src2[25] + src2[26] + src2[27])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13] + src3[14] + src3[15] + src3[16] + src3[17] + src3[18] + src3[19] + src3[20] + src3[21] + src3[22] + src3[23] + src3[24] + src3[25] + src3[26] + src3[27])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13] + src4[14] + src4[15] + src4[16] + src4[17] + src4[18] + src4[19] + src4[20] + src4[21] + src4[22] + src4[23] + src4[24] + src4[25] + src4[26] + src4[27])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13] + src5[14] + src5[15] + src5[16] + src5[17] + src5[18] + src5[19] + src5[20] + src5[21] + src5[22] + src5[23] + src5[24] + src5[25] + src5[26] + src5[27])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13] + src6[14] + src6[15] + src6[16] + src6[17] + src6[18] + src6[19] + src6[20] + src6[21] + src6[22] + src6[23] + src6[24] + src6[25] + src6[26] + src6[27])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13] + src7[14] + src7[15] + src7[16] + src7[17] + src7[18] + src7[19] + src7[20] + src7[21] + src7[22] + src7[23] + src7[24] + src7[25] + src7[26] + src7[27])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13] + src8[14] + src8[15] + src8[16] + src8[17] + src8[18] + src8[19] + src8[20] + src8[21] + src8[22] + src8[23] + src8[24] + src8[25] + src8[26] + src8[27])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13] + src9[14] + src9[15] + src9[16] + src9[17] + src9[18] + src9[19] + src9[20] + src9[21] + src9[22] + src9[23] + src9[24] + src9[25] + src9[26] + src9[27])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13] + src10[14] + src10[15] + src10[16] + src10[17] + src10[18] + src10[19] + src10[20] + src10[21] + src10[22] + src10[23] + src10[24] + src10[25] + src10[26] + src10[27])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13] + src11[14] + src11[15] + src11[16] + src11[17] + src11[18] + src11[19] + src11[20] + src11[21] + src11[22] + src11[23] + src11[24] + src11[25] + src11[26] + src11[27])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12] + src12[13] + src12[14] + src12[15] + src12[16] + src12[17] + src12[18] + src12[19] + src12[20] + src12[21] + src12[22] + src12[23] + src12[24] + src12[25] + src12[26] + src12[27])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13] + src13[14] + src13[15] + src13[16] + src13[17] + src13[18] + src13[19] + src13[20] + src13[21] + src13[22] + src13[23] + src13[24] + src13[25] + src13[26] + src13[27])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14] + src14[15] + src14[16] + src14[17] + src14[18] + src14[19] + src14[20] + src14[21] + src14[22] + src14[23] + src14[24] + src14[25] + src14[26] + src14[27])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15] + src15[16] + src15[17] + src15[18] + src15[19] + src15[20] + src15[21] + src15[22] + src15[23] + src15[24] + src15[25] + src15[26] + src15[27])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16] + src16[17] + src16[18] + src16[19] + src16[20] + src16[21] + src16[22] + src16[23] + src16[24] + src16[25] + src16[26] + src16[27])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17] + src17[18] + src17[19] + src17[20] + src17[21] + src17[22] + src17[23] + src17[24] + src17[25] + src17[26] + src17[27])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15] + src18[16] + src18[17] + src18[18] + src18[19] + src18[20] + src18[21] + src18[22] + src18[23] + src18[24] + src18[25] + src18[26] + src18[27])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13] + src19[14] + src19[15] + src19[16] + src19[17] + src19[18] + src19[19] + src19[20] + src19[21] + src19[22] + src19[23] + src19[24] + src19[25] + src19[26] + src19[27])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6] + src20[7] + src20[8] + src20[9] + src20[10] + src20[11] + src20[12] + src20[13] + src20[14] + src20[15] + src20[16] + src20[17] + src20[18] + src20[19] + src20[20] + src20[21] + src20[22] + src20[23] + src20[24] + src20[25] + src20[26] + src20[27])<<20) + ((src21[0] + src21[1] + src21[2] + src21[3] + src21[4] + src21[5] + src21[6] + src21[7] + src21[8] + src21[9] + src21[10] + src21[11] + src21[12] + src21[13] + src21[14] + src21[15] + src21[16] + src21[17] + src21[18] + src21[19] + src21[20] + src21[21] + src21[22] + src21[23] + src21[24] + src21[25] + src21[26] + src21[27])<<21) + ((src22[0] + src22[1] + src22[2] + src22[3] + src22[4] + src22[5] + src22[6] + src22[7] + src22[8] + src22[9] + src22[10] + src22[11] + src22[12] + src22[13] + src22[14] + src22[15] + src22[16] + src22[17] + src22[18] + src22[19] + src22[20] + src22[21] + src22[22] + src22[23] + src22[24] + src22[25] + src22[26] + src22[27])<<22) + ((src23[0] + src23[1] + src23[2] + src23[3] + src23[4] + src23[5] + src23[6] + src23[7] + src23[8] + src23[9] + src23[10] + src23[11] + src23[12] + src23[13] + src23[14] + src23[15] + src23[16] + src23[17] + src23[18] + src23[19] + src23[20] + src23[21] + src23[22] + src23[23] + src23[24] + src23[25] + src23[26] + src23[27])<<23) + ((src24[0] + src24[1] + src24[2] + src24[3] + src24[4] + src24[5] + src24[6] + src24[7] + src24[8] + src24[9] + src24[10] + src24[11] + src24[12] + src24[13] + src24[14] + src24[15] + src24[16] + src24[17] + src24[18] + src24[19] + src24[20] + src24[21] + src24[22] + src24[23] + src24[24] + src24[25] + src24[26] + src24[27])<<24) + ((src25[0] + src25[1] + src25[2] + src25[3] + src25[4] + src25[5] + src25[6] + src25[7] + src25[8] + src25[9] + src25[10] + src25[11] + src25[12] + src25[13] + src25[14] + src25[15] + src25[16] + src25[17] + src25[18] + src25[19] + src25[20] + src25[21] + src25[22] + src25[23] + src25[24] + src25[25] + src25[26] + src25[27])<<25) + ((src26[0] + src26[1] + src26[2] + src26[3] + src26[4] + src26[5] + src26[6] + src26[7] + src26[8] + src26[9] + src26[10] + src26[11] + src26[12] + src26[13] + src26[14] + src26[15] + src26[16] + src26[17] + src26[18] + src26[19] + src26[20] + src26[21] + src26[22] + src26[23] + src26[24] + src26[25] + src26[26] + src26[27])<<26) + ((src27[0] + src27[1] + src27[2] + src27[3] + src27[4] + src27[5] + src27[6] + src27[7] + src27[8] + src27[9] + src27[10] + src27[11] + src27[12] + src27[13] + src27[14] + src27[15] + src27[16] + src27[17] + src27[18] + src27[19] + src27[20] + src27[21] + src27[22] + src27[23] + src27[24] + src27[25] + src27[26] + src27[27])<<27);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25) + ((dst26[0])<<26) + ((dst27[0])<<27) + ((dst28[0])<<28) + ((dst29[0])<<29) + ((dst30[0])<<30) + ((dst31[0])<<31) + ((dst32[0])<<32);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h0;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb1ef32821c3a52cd1f1f6ca711cd054d6acd0d49a90f8b4a676cd079f006a690b5e8a424c8c888d6fa269e4917138fe03b1b19ff33bcb5c6bd73fa82b194731f069a7d501963e62adb0b3d3afd699b50bb35aed86b7b7fdb72a7a41f108c5d8866b5;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h494c053c17450f1cbba078d3147f2271f8f6c0725e1ff36655728649827a4e334577a93a2732df93e52397523d182c8c38a25c2a717c610c35d9ffe2d950cb1729e36f9d2c7a2af86ee8548c60f4faf76f05d975adce892c607436cef36bae9cc666;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf7d8ae7784ccf35c4fdccf1a78d40db1b666f3bc1300c0aecae36870caf25df143d9e9066337ab0c1ed0118b88703d75778d3d235f46f343d741f9064079b8f7a8908b81ecb84ca204acb739a77b729fedb3b81c0e4a813233d23d6f3aacb74779ee;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h425c5b776562c328aa97538b44b5a1a808c8ad64182741491aaed92bb5d34ec65558e19043068cef6de2583bce45eb7054cd9c817f06e3846c01324ed07eb2b8fe8f6ee7eba496b9c10e2833f2276ad846cc7cf71254d790debb669575afd51e74a0;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc26c4a6122fef7682e266d974dab99f5ae247b52168a5f913442076044d608400ec4dd05d57f9a06aece6c367612af92e5206be1638d21ad5c1682587a1a784afdc92ccb7913d37264e01d4aa78570724bd1951b91fc0a5859ddd56027747eab42b2;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h28d3420435b2446c189f6c7dd176153fd1e8bba42c123782ed2843276a78da3ed250113dd8115d24022bd8a34b98facdb2d2c0473f586e9afb825bbe3e8bba33eb06671f9652f732bbd3c79562991556d6ae5c01520f6844526603c642630988d723;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h18f0801b56f9e7ff150df25d47fa8463523991134baa46ae7b43b56ba871a5cf32bba729d941377628d001d5e176aba37d8e7cf416e8136e22011d505a4160751d83306471815c4147fe7c921b8f88fc10947386e0603f373772c417cb6efe91c08;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd59bde863baa025ae366aaf6a46de01d79847c1957e60c6b12077a1bcc35b2230ef154a9899cd8ce22da2a267ddab69d9aac69d3c76c3e18207534d5df92951d789d8d7fb32bbb2ae3613eed593e6342f7af811c956af60ce62d0deed639d0562b62;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf22e7fd7ea3f533182f856df4a77871db953a812c7143bdf056f66ca11c09325787c3a72faa26b8109facabfadbd44d1980d8afadf313fce51e288bff53d3365436da668a00c087ac29f3568c969b3e8595342f7de8d633245eb326321c2a70cd1d6;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc400f7bcde0c9fdef51cfa4bf68acbd73ef8066c12164fb0f3c7ae0995e8119aa7759faa588bf83fac7c8f3c4a2d3536adf8b94c4f194feda4029017ee41cd7be0a00f084d58d579211c2b9bf41fa8ae78e3c06f5542d23c5e86496090e20ff4eedb;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'haa2ca4cc8e7119f8ca5e7897c6f7cf7b353d87ed1c0ba1f20f8d588c4e546c0d44a26209498e92fabc26075fc1ad2394f21ef82dbbdc782ba46cf72682f88780ba29639538452e4136ee97bf8d33a4de741249f244bd51380bd4a2f2231c4fc96d7c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h87917a42c0a96853417f4f4165a0ec247dda0a2cf0748ee5888c67ea90d9d039ed5d7f4cbf4bddbea52dd3d00ecd97b71cae76a7cdda23d08e3a0c17e6d37be8f5565f246d8dcdae9800b88c094d0510788ac3b76fe514719299a2ab699b22f03a2e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6fd83606df65d9c1e40b16352ce3f4042b996eaafb6775a552c4ff13b600e86d12d25d680db12c24cb7f3cfe865135da4e3d016bb90750bca138cb09cc374ff77372b231da3057392119b1fbdb989afcc58ed836f8437b3f8915699c6399c02afeb0;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5cc11013232971cc3a2216ad5912e975c980f3f98e0f2c7796d438ef521f282561105765dcf55fa1f8c6db70d0d26de8268df05afd7229c8138111db7525125c67b458f5e46e3fbd938bee36782f18da9f8cdbe7794bee49c2644c3b28df644577e8;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1ea3b93d9f64a54fcd1ceac1b88b421b933985e02f11aced39df540c62a5f52faa4e12fd935d545fadf29df967302e6bcda4b5a10a6c6fa1b9e8f6957c6c06582e9c4010f01a3aae0feaa3e042d132b6a9c7a99adc642f0ccafbdd5433fded0062cc;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb1bc4bc3f5e71e680541ae34372b8a517d0b551b05939e3695b43c61cf62c6f6c412de46726720d81cb00720346727ea00b047d1722007a15c20421940fcec34c14a910bfba8913ded73b224a706e8fb2abd6a01c5f576f3518fdd7e2075aa13c908;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h39ff24a13991d70520ed91b39a7081be61be5d94b8c074452e0a3aa05ba54bef29b2507746a110d65d1a57612f7bd1c080acc1947331954fbc73b9fe75dab0be26cad8c5b1e3cb08eae33c1800191d151699a59e255e9ecc17f2c6da5cbd0f44a9d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'heab267943cfcd9e9ac23cb7409d49e7b0f82ce8fb19805455417944e6005cbbc16d7ba478a1a44814f58cf15b3a712ba10511e60c571179db4bb2dfc5a59f30e42c1f8fba9e1deed6ee499e34bad0b8026d74205be2cbd5d6f2db08eb59b8563996;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he053bbb4dd32251c82b0eb070700bc8a77eff0ebdf846dc4d74fcc8d1967c31de26ada1a34fcf878b0e3089804a5e1eb6050f5ecf542faecfc42a0763bec256adea9bb114e3cfbf253313ad0d6fd9595e5347c661af889d1700aa25227c9c338bf3a;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd7890450244d5c932583fab98f1dd01be79e2062f03d107df85ee2ccd5725e56536bf2808bac520bf07519c57c251112cbeb9fc3374697e752d7fb4479bed6d33121820bef3b69da3681dafe438959db17455776aa244e175eb75b6840418b5de98c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha8efade31d81b0c54eb83da5313db0a3b4a2cefebd45b6e2e366a22554c938aef68afc2d88820eefd0d996150b8c9d490f93380c465b553be030face77ce1b7c95d3e1c090628b8a661ac78b0e8277277b605b788d4a24b1f5441b8efbee68888a3e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd424a481a0e3e90f6ccbfe70ce05a3c37b703c9b479543fd1b2fff2d8759461b5d8aea39af0a779314d911281d887b457531cc68bf849d8391a9b2f94252a06b9f76a4a7e6dd42953f739441a05d7415029ca32b1510e3b446766ac4fb64c483c488;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc88566b0a0494f6eb09a2aa26431c53091766b7d03c24cd8735bee69f7623408af33bd5114d22536a8a1fcf573b05577b8d7d8aa160d3396bdf402b8e105bfb257531ae1c85aba662df76249e433f563e545c8fc4b7d352e7ff7c5197d572ca84f6c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h306f5a6412f48dfc06022df06d4ae6284ce2e267b2b9e1ddd99d7aef1c4c2192581074619c0666593cb0a25454f7f24eba27ffb632eaf631120dc1a78ca4c557922712cf704c6fd0e428b336934c0cf0ca4ee70fae6f5cbd4dcbf145738b01a0e36e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he77e1da51de68a7d6df256ccd079cf306ca94ec6cdb9770ca91c7831f542eeb7085a01119fa8c7c97a816a92a5f1ddafb09b38f45879c7af47dc3541643ab4a2f9ac23eec67a600880c7736dd51f78a46e3410793a07d72a859fa2a9c758e0dc826d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf927ae931f517a2801147773b890eea374f67e1fceb4ad31e6a70ca6d2003ddb43a58526db3ee03828ced3c26da1e27adf77695fc10c78eacdd12a7733912a9e22c93add7759c8c98a446b4f72867db0906eb6844c10a2e62ec20c4683eff8ac4f40;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h22e412a812d53cf0d827f615f53c4f9d17e808e273e0393bd42cd074dd36811cf63bfedf1bd7d6ae3021e212f972a875e8315a4322216ffb5698a66a529c81619fe86e762df638730060772cc4e516d1f7977837e8ab8cb301203fdb92156d746d36;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb3a6edba7e9d14318d9ad1a7e8eee56014e171fd01e499014f1f78072faa7f9973964fabcd35d2cf37ed67e322c74e44f657c0eaf2a37a8ecf18450e86dbd98747b08366869d81d8c8c714069b5ccfbee1e2e0574a07fdb453a0ddc51b5679fe715;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb9300ce876dd6e171f896471964a3017ac8c6d00f06bc157786b897184f09a06277811266130f44276c48a6c5dc727839332bc419dac9685093b4b2418c1979cf86dde117f98111290baaab3c49b7018126d53df89a866a200261f0b78f39c233cf7;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf86e8f2c6a78c02e7359289a3e59e15c4b884b44400c1756ca3d639d02fdebbbc59ebc2fc912cdb3968771184151bb05d7dae45bb31b7c7b240785ecff181faf499c8cea4010bf80adaa90019e73bee0fd04d60ae667056a201c9d98424572dc44d2;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7de09ea67305bc19192aecd41fd83783231d70894f3fd47f144b61b0ff559b71bab46043609cfec6e45723f993f34c285137c8388e44b21b258d71869d3f192ea7d403f79a26200cd3aa0e3402570ccacc0e83a642bfff680bf72dcdae2bdb59049f;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1a33e67b21f12d930555e1a4f9ae8318404d6179b26eea9de0cea6050eb769511cada9fda6ca1f4837ddfb6e19986e2b6e5fd302f58d7404404d209863a1c24212384acada92628c53d161d8d47f70ba14a213f56faee81201658e6a7695cf51bae1;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc81d2c46c091e0c908ebd3847b57f5ba94984a7716911316557d5172a4c03aad850bc18f2a2a595d83487033a1c193ec3cc9ec7c0f5165f833f0ab3672ecb9fd1d732a192f4a3a1c08159154c0347ba2548f4348700d424f9e2926efbceda07fae38;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8439ccc3a18ac97b097c7c3e56172531a18652071c322d19783097a2c1e6a83132467c5e948c4c9b4d083f1d8d1c5ac5b9236214da1ead3fb44a55f92f4349edae118d457e7221c3d3eda3ea6c8f7c4ace1c964d37e013a05f1f4a72a0fc82584f0a;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5ecdf796e507729be1aa77ab017e88dc0a3a814fd9add8795e3e4153a7e4c1442c21189ac4cb7ba83cf7b210c76c32ab6348391d529f48087df32b09570259ecdfaab825fa396348360615f634ea3eab27070630aae5c3f92481192d1c1edadfe587;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha19e48f5291d9202ad91430f9d31864e6a372f11f67e16693511d6084648f7ffa416b4be2978c725cb4b475e51638141b05c6a53de10afd2fd02923af9f496639dd972060f8153a2bf7d307d84ddc64c26dd4f02669061a9d332aa7a062c6048eeb9;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h66844e09df58721bfdc7c0ab4eee571a17a9b1dccd28765d2681e8eea9c63df5461cbe7411e835b0d0276d61077bdeb3b57495f9f51f27d63ed999fbbe6a5a72dc34ff4ed3c250b8e47dd6aa8efd36fad87a12924ad2fffa3e865361bb63402e2949;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc7ca79b225d0be86766d7cd984d558c6f340bf483086bb61efffb32c3c0d3b81fa94a8d3b9e1faa771a332f08f06a8fc3bbbd61ed0f0d578e44c50b517c2ed941115c69d767ecddda5b2135960d5becc87ac7cbe3a302153be5483380ebe506dedfe;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h663f18f0f9e887afe121b01cef1b326aaa1557b2e98b813ab00a15a5bf92b1c8d0faf05fcae757fe4b5003301ab724f655d8e47e7e359e9b76807c2ea9164f8d7972e4ec7c4c2e8f5423e315b4eeee72f8081c7c9d56258f5958ba7b079c4923dd3d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hefe81e70684209bb97acbe90cf0766db4d8d74e6a9dc3eb343c1ef7c94721c3f1eb3e891dd36cecab93f46f7752fff12ea67522bb772beeb3940ec6d1331442f0d77b5ea975035a600e8cb5905d74d352bdba480d89ebe2dc0033c4cff07bc25a239;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h465346f216a9ba3eca805965ce48aeaeac37b9e7cf5e88fb6061cc6c0786df376b41423cba7cb8b0dfcd71184e42f8e45a3079e40236c09b5b180f4d3629ddb7e2f705ddffaf3390a28b25b2a170b2e95ed7850410a8c143699f138016b6d7228837;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hac894b37438718c3f2f0a2a5a948610a880c7565bf87f309452691e6c314dbd43ecad726f7f1dda0ffc5c7002abb312b02a1539cef920bd227f6d5f11dc2ab367071d7022fdd5863fa8872453ef7ce7d9e971b303a7a2ec817b6cccb2ae53091eab1;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc116bd1f5e77f45aaac56e7081b4f6836e3a39f3d719fbe667c54271862088c56e8fac4de86e29a82f4727bce253121849c2f422a3dcf593fdeef8a285b520a9ea69bfa2b89e9ef1b21ddffb1bd1102f50f1333a60ff0b42d1b7faac1195195dec67;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1942b78869792cf495140f842f0f0ce5ca189800d6a0f8c2ebc37f7abf61c24effa9261c6eb289bad35b4d2be9048040de794c23fffad23d5e8778048598289fb429a20ca0f8f01af25d40d6bcd3d36a966135f96e0ceb31e94ae9a3d6d221d40d5d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h974a552108399d66e94feb9c62729b6e5574168a088dfe9eb5bd9ad6bb0cd7a9fb652dd08fbc8c21564ef6aba4893ece152be81325ee074edab457df3e107fb4cb23e752041100a8a639f2b64bf03d2b6746705143fcc1c78a550951f8a5913361f0;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdd672d253e0fbabf6a1b54cfbb0a69602515973431dbf985e8404ef53a657c6e760f2be027f02c843cc5dac73781c962b93378f539ad1c2cb5684a5cae8781cd0c0cc53e4fcbc1cda1f9e72ed82bcb5ef4c44fb4da739cd5c4d419e38dccaf813d7b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h937f6407bb85bfb6fcfa44c6d99551d5814c5a834a6b2d894565e38acd2072e940c341557f4740e6eed73131b25d47ae6271a07aeb605c164db72a61df4d0aa26bf37d98605b21b6f831539cfd285339a056976c63007be4f3e707ddcb3c907f601e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h713eb34e0beec2e6be57fe671fa3d006573245143b4aa8db741b881dbc1c20f6b88ee07d922450805c1610ba59cef9ebd03e08dac2e56aa4c4c6758bac9751918bb0a2673854093b3d69c19d54473362dff4e8931fd7614946a46b06769c215b3e13;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd0c79786b3d36709a1644a53560a366cb947402cc40487535310502c185fa5d661853738d587b7264749321356a2fc7c947fb2c54eaf01d90783c66ee9aef68cf63602f57f752e91ec616b934e2856e346ab5de9c5886f6ccbbd8551b52ff94a0bfd;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3d7800c31ec654632650317dddcc7666cb0641fbd30130b80af7ad308c19438532c21378c2dd2a556202e8e81a6cf09a55548db6419d4bfd553e8b535f7e69f8ee2730ea08f5fc19f7d5fe71254961ec038cf9638cdc511fcd80da61563fec0dc843;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd11535cf4d472b0c7f52425407e701f24fed196ffa07c57f294d963dc278762a1b3049bda4fd419a0db6470f6d936382a9d46c580269c42edfc0a1af69095f6acf313a1db325759f44034bf6f3973271eed2578d3c9b5abe81fbdf153e2d17a6fd8b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9d6d24aa5a18f03256df31c98254dcb32c82067c7a3f6e2aaa4db9d64408058f2786d7544a338dc9595197c811bff8a47afe3714ab88c4f078423d4ca01eb44b5a9108ce22f6d21d1802dafaf764bf435b6e8f77c17df78b6201c4ba683b93cb9841;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc37a4926c7b9d4163dc283cc2b5f74db6a5eb81706df09bdcd510d029cfafb120d6695106b96820500ecdf6692bf3dd52e1749a0fba03c4cf3b4ee85fa359305221761aee7a0438427b304d28cbdd8892984f7a1474638fe3f5a9104973ccbda445f;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8817ef949ddf49f05abc4555d6554a95c733ca6aa78d77979e906d34e49d7bf0858f79c4f8b7e06c2264ba74aabe7b1cb6ee92bd5cf21efd1783d59530c12c6c659103e1b8f8bd16fafb2108976a6e93b9a1aabc02b62f6de33e9d19c1f577fa4fa7;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5d02a19de963f71e9226b8386b4c9c68eeb7d6c93bd2a9448dc3b072b4add4832a8b9ef835273b1168f4f9738ad9c96114e782cae87ced17750c430267b10cf1c31f889b51c0da614ef7bf5bed323d62ce108f032f861484a039319dd03c4e25e062;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6f325c606d6782749026d18dd5ebebf0326553bf689816bdb35ec59bd90224e84ca00f96aad13de262584767d0759bd5c0a5c77ec5e4ba22f7f90f9b8d93c7ec047d4489d33c2931027eab6070704797cc212333d9c7079ec411a2884472f9db6f4;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3a9ebb061a2a27cf7bf45d3f94ca30c37797138cf62e38e3717a2fbb90e7976e9a0a799220df3a86b6e04c3bd85fd2a4c588b492f3144aa32fd71127247691ab8fa786e28cf46d7f6fbf2069c2f43aab5648504e10fccfdf19c069aef619e8ea0269;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4e8b85b7651b9e5cad5f6f2251af7c0c18c2f90b5b31288b41f39bff2b977590c0df96bba4617fe6be1b95b23a2f5b1e4d5ad7605a0157803adf2cb699122481f5093ddbab936b7ec09fa117cd5bde370811ea5543fc46043518a2aa30767db8e67d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1d85f0fd2cfa31016113a20f13a834f54f8e3cc8d76cb6bebbb2107f9b0ac7a43fe2884654fb7209f7d35ac0d3d2384506838cbdc13f3ec5877f420fb75baaf347a19a019f00c9a46131ddeefd00832c71671dc2a002c9dac2a696760d0bfb14272;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h408c885cf821b0f7fdcce6af37fc706a6139d9b3862125d5634e6f87d02a3a2fcd96d18119d0bf0c25bc1b346496bea3139c6274e0e7e998ae8d467924ac0f1754daf3496d9ebfb23b8429d108271c1d658fc9233b8f573cebb226266b16ca17d54f;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h409530308a55dda3be2b687b497e7a8b5dd2e57e513533127afd85d65eac745669f93652575de1e80f3c84637e64f7c1e5b56ce2781e9f15b56a3eaaa461c38259b1eca37776116db909d168a275a3d7a9834c439de050f5228112ffef249c058c38;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc5ad0d924ccb667e35cf213bda3efcdaac8b361eea5fbb619ced46cc3cb5adfac4bd1cdda3d0e4f337a2d7201a04a997850c470285a08f2a0c8907e17a5000f55aa72f922742918199843b9b9c4091980b0d7001bc902e65b344fc1d05fab0a9663e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdc66070e9d692ded9ea07cc2a98fde541e97a051e2b0a5dbbe087dc58823a9eee54d6e95e170284612b083e39c8e638e479d2a4b890ff5577f249c488e1728c6515e8e1923f4afd939acdc06de810eacc0cc59f1d52863af960ad5619f53d119a71;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3c56ed2c5731e2dc72898c11dcf23d52d622f9cf3453b20f27bd789ada1845a9ae6b056d25d66920aeec407b8c3eaed0a4c2045bf715a8fcf18a151fb89bcfa7d261efc699730717cd4a2c49f156a40154db44a40e7e79f18ee44148c612e13db8fc;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h31dc9f0696599e88c63931242ea30454bf17ad33a1ebacbb99fb5c530855eaee133b0b34dbed6bc48c5d50d6278844b92b511efbe45b2e95fa3c9073e13fbf28fe79b8105f093ff9c5a1229a6b62b55dab6c665d4f64760d29d96bf788fa395e9e46;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfa53e1919f93ea3a1ea4645d1351d87ede6b036f09209f130247c8fca044e423923552e4feae7940c151016c46d1da01166c677d934eab2b24f9c00f35763a78269467cf5319530524ed575d9952a821bfa1740eb2f198cfaf9bde8c8fe3a86deadf;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1226cdcdd1ebc4db339a90772bc510346ed954a313b1e127f763394ac8e46498394c0a59ae49e3c48c2c673e3928d040173464046228b286f880d54ba13db53cb6f492b4b19e100fcb192140404ed938251220e87b8b049cfa25566e8af0729faefb;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2ee754a60244a9ac31e3d1f3abf7c5dbfdcbe63596fb9abdaae4d3d57b3c148a83353b638f2fbfe97a07421fae67d05961bd486f16d2df9978e61b7e8e4f4ad31dbcd69c5f30e4f762e3175d131694aebd0d4581d6e112777b67561df8d376ca8541;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf1be7f929349fc4041e248bbf94a78f74413ded2be260ab372d99989f30d6e3b63a75d90775e12b89f5d75e3dba7472763ed9a8c8c01c51cb6c2ad0fe3df077c7d46b25d032c35550edc71faac1028e63a672959f28636d84f3373c0b5fa53af3a11;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h10d92ba0147d23ddc6f7988c43904b255f5e8e53947220340ca99162cf6cc15058fdafcdcd03355e5a92b3f233ff0c640ba6d731843a01a34e7589cd3d5b80dad82c1ac2ab878ca0c55678cee66d8f80b945fde719b43d5d0dbdc97f566a60427f28;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7b926e6dd1a674331c72688e434ccac44fbc479a75ea23d9266121f437cd20c5750533fa340946782472ebad3134c9d576ee837cf6bd2860b020207746d6730eacbfd11b795f56d47523ed81a1f657fd752e90ba9a8623cfa1698a845a5bd3158f7;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h516b747c7751e8388f0cbcf6c5c956732e5ac8480146e30602ba9f8b1f22676686cd6221436d16a65df6eaca911140b6d1b4ba297ff7d2f1487a1f64aed9487d5bd5e706dcb7b046aa86f35c117e5bfa299c7d45b0da6bb3bf77684ac17074117d96;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2cf67a4c44bd3cd3b2b4f477e20df07fcd3f707dda774043a32b04445d4c7d70aab2919d3c3be8f4a80db2e4750096b5c1c49684947e520b4c084d38decbd844846a1d68c7b9f6671fcf24038ca27bc209e71988431803aa8a63de429c2ba73daf8a;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hddc51424122388467919121d9e2ec859aabeda93cc4ed84496b3e411b61e18faec24baba212974969bf5bb50b12dcd19b47f00f8bfffd207d6236f1ec2b0ada5fca92f08e65689715a9ff59314f1e5ca950aa55ee41d256300b98fc410c4a2145b12;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hee71735ab202a8099562f0552c5626a1699004fb06c1a087cea5d9994f2cf25eea7f1aa1765e851fd0009af3ba1a17019cb9f01d97e4588f68dcced2f66b5e3b235c624470caefbfa6efa32913d424539851e5f4a2137f09aaba169a53da6346348;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h41fd558f03a771eb38f32edacc37beff41c67a39aced14593e7211dcc46e8a71e851459635793529d84b87863acac907902daee2c9a9b3a9cc01c01b479597fca83432cd6b6e5b67152ba0d079fd4b71c0d8fb61e187dd2b07178973fdefaff7f17f;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hebbdc3aa8c3251350eeb957eb58dd93ed357a9dd01eeec0136c10051953ae62e206d19dd096c3db617cd67a7f3ead76c1d07c8ff8e94641aa9817dc33b56539981372ef6ad23e29c4ba4c1a3f42f61e427713a7ea86e03fc46606e6fc16aa00e9b2f;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbaab7b8fee291e6f2e700240c6d550f46ab1fb49f5f40b9a6804b57e01905a6cc4687f938f84c43ced2ea748c8537cc4eb059d8b822fd1cdcfec7e0e4c7936b9ba826c28b4c5bf5a4fa3a73e91a3f4385978c71c9403a1b30848cb50b44f8acd0a83;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h52cb87ab8bb9c055646c19ce623ec3683780607e60bb7ea157fe66f82d57946e753e81b112793837e912971fa93ce829fdeaa596165e1218bed6bb57436ca9a4c8a8b303790e6d854c9e0b99217af9723efca58fe00ff5a4f35e46b3dcc53ccdc843;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h32ca8c2bfa11a05c9fc4e0f9d0ecedd54decfab3d2b3009eefbd9af6bd1d8ce66b8e9a2fc997d0d2b666fc62049614c91c894601dab488268e9eb6914282a7441dac03f3db886730ad9dc90f782b35e85afe1112c55cebddf9b31e0920782d214f03;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8d9503a738c1dab2bc1c77cdaf7ef1323832179c55e40f43dfee610a07912e4c74a4b78f630b6fffada42c33f158a264040f1cce6d99d0f99497d19aeda2104ba0c7e3213f08a4f1929c6b4842dd029988756fa003789a5cc1d33cfa9aa0e474ca4a;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h819d1a4947226981a6076054373906472fc099e13901579d2635f79aabbdde07d75a10ff333b47bf7ae74a118bec3a3ed26d7cb009ab34c4b8170ae4312e9b2e73c805e45505e3e5716d40415b69b20b21ca8f4ee5855e4b60f35e1baad4bce539b6;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he87bf9a23403c412f9ddbbc46becf7474da61d13bf2830ecb7f215ca4d2f335d02f7db4aa2ae26624572400130cfb0d80d20a8d07a0bf217f796df9059236911d1e8963bb751734e6c201386e9998438903c26f548246bddb0533d0fa5b794c8e077;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd8373e1fe5ce802fa271106dd98698617011b19d7e408769b84e0f97946dae127d79e5906ffba8390ca8bf5ed83482827a6373b4443948fd3ac160d67650ac00e9351ed2402c895b4bc167e9fa97bb893f2672e162709e52244eabb5619a83e19c9f;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5ab4b41b90455694eee1bc18419e7afe20524be0ace7f0227ae570a55505a0670347d322e042e40cbbe02370ab3006abc89484e9126a9867fc494cd316b023f707217663bbf0966bbf118aa68e776164ce015578525f0976f61013cfd58884617f94;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb39b8305e2518008efae7f4e666b4b80d9552f77f6a0c2d13533c42edb47792a7cf025904bb3b0bed1e97d2ca360b2a3a98b061f55a3949524d7e08326a802e4fce87141ce68e58095217b9619af310cff7394bb2f9a72b776ecb15ed99efbf1ac9e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2aed5c2b442d6bcad473a394130bdcf96f65e91f0794f31fb9c55e6e0ee2d862e84dbbab79a521dff7e241ee4a9bad050e36a0a87b2138cb440c3eeb56e98a02e7d1bb599764cc5d5ba2233d63614c2a3589c45df35df5d945b2b55a9392ae6783fc;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h26955a72b2eab3e87d94f341c7a99355f29835515554aff414c0f6c16c394518257d6af06c37345b5d8d78f9dd4b69577367e83647761236b5b4334591aeaf1a57ad9ce6db3a877dde44dc76654e7c1f1902c2fe9e88f083b3593993bb8ee352a5d4;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2ab7601f8acdb1787f8735af8f41523f1d940e4a2d9489a23952729bf2d781fcc6e3d61ff4381f268f5ceaa98a5383383ce38680027313633bce65d50f937eb5503a49d9729171668cc2262515f02bc624250653d2d1c1be6b2d52af8b35afc6fd5;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha568aac5615402bdb01e638f2edefaba99737440323c8fe02c52e0b383cd3963f20b57791dea43c333139740d5225ea45a7fa4c3b2d52efe31a0cfe9aaa759f109469628d54deea3f8f6491a873951df2b23c20491540f958badf5068826b2339251;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h30027d1378635c14a6e5af3cf7f55939053090003e1f3a0d52b26ba88dbebb4fb5a4cf25be54e0b31c0992f21eb420aa0112503d42a8a889a1cac244fa7ebce0dbec8720b0fa19e041db4ca2df4cad6ea5a07334838e546e952e0cb6f87f3f40d0ad;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6db60704642d4ad6b65525d4001f3f72bfa44de8da60f0bef9d1df21a19b472558bd2b473afca1ad0dd5dcd547faae85ce947291bd8666b06655842993c8a60ce702e771dd5d787e7f4b431fea74e6a273af8baa3f452674e754d227a3eaa6984c70;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7667be6b9fa4535a8831d1adbcfb5810feda2cdf17ea91c5b4291893b5d938228d2fe9f96588baa95fce19d8e856ee2637dbf8888d8599845e39de13856e7d504ee69537d67267c5bb66677d943e657e83789795df7a0904328b80563c9e264c9ca6;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9053c85807174ede65578cecd6bf00cb120061a0a6cc16c5c5846973e9e853b61c27befa79ed5e51dcba9136d9f8936489b9d5257c5320a0e2397e3e68d7d6009eb4a3c07616309cd27987a5419768aeaf68c8d6f52379075f95b48cc669a93022e0;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h618cb7519ebf0c9db7488ba2bbc96621d6a1d8ffec5a68df3a203244119e40d8b663266e658545eedd5933248697f64e6d5ce622e0979ae441ad16b7fe4e6fdbd98d0f3b0f0d7cd2e72e46c969fdfd3b72c0427e384ccb3bb9a241cd76ba62b05bc9;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he417bd9b507bf26b2cba8cf2e5f28317521594f43dc9494274a9671283e0b173d477e3bfd6788635f181fd253e8055702f4d2697c0252d3a529461e2b20244f8194ac1abb689834730abaeb8c9043ab7156c1cbe8c98cd91cf58b19013c0bba40835;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6302c128decac03896bd028fbdc6c534f05573fca55f4652afaad7c27502465bac5476ec197f21a36a7821ad62957b3007ce74a2d9c42e0dc28c70e83f8d9b2cc72cd3677c30d8db613ea232673ad3e2b6feab3d04eaeb44501c904a818e40abb6e9;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h57ba8b5070b1d133f57a05450d2f3e4d17d0e00805dfc815f0351e5762223f9956dbd7193b84b639fe85412c9fe6d042247396c1610a562033e1d68cc84821e0159a4b6833529e18f492736f46b85f2e080984fa3eab3dfa4603c9c4638419ce1439;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3d53259f4a365d945de3d5b8f865798777afd8bab6348be26fe94240fb07910e15ef891d0ea63dc8c7aab3e292d9401292c85f2dddc6e122fc8f1f76ca8c96bb498c1221c1e65320e7b2949f9a807a19c3f7b886c2709a10b96b5d87d68e2009c3a7;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4bda4ef9dbf098333dc276bf1041eb3d3b3643a3eebb2bdebf785b49e72518525419151ba13a0e71b6aef81cf8a9874ac28225286309c9b0002a1e281d65d9f58e98249ce6ad3f8dd78352dbfa1131884944cd65d0aac35105897ba2d459c48ed2e4;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1fb666d0916d6a122cb39c1f41da0d3fde99c2d57c4bfd3ccb6e720f84564172750d5c93337b48f5000aea1fccb17401fbbc975c4c357933a4425ee333505e6c458c4e9608e95816694809eac360e0ab29e340de077e58dd1887b31c4a7bad64efb8;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5995131abf2d235e710664b08b5acf969a669fd4721f57c936701b6256954505ca0091c1218b3c446cd9af747f58ad38896f894e4e22f5f9a52478ef81791d0f21b6affcfe8d57ce896a31935a62ab9848c8e0cf9d51da1204ddc5be1a3968857d2e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf0e322b9dac2087fda6ae9da6f75706a94a1fb54fefd6545c693452b3d20d975099d2fcbdb2bbc1e91a7c31620c0aa6dae994329860bd77d9ea47f49dd3d9242ef84b6b5eb742823ed65837cd5fb93d5d58d392fd57dd2bfb17a9ffbccfb4bdf453c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h58bf88eafd76d0bedecaeea8bf01b00532038ca56190341b19c5f6dd1d4f09ae0379f76e4e56d017858f78d7f7fd4a9b9e8a44336478f78d7a450b53afed4e7ef75bd6c1471919ca873f40ee109812d7b368d84c95a0ad1817590ca697f015e04744;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5ba63e044e86b349b841dde1e5391fcf99a25bafd20bf3f8c8da1a1102d624f0d13d3764d14fd11bfe095e66cf2dad07bb591c675f1f0a941a21d9b6b530f3e7f541a139d5fc4b20b148d1e10478bbe890a920da4a5a0ff6c3dfac44de5348d1bd5e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hcd30a71af786759bc64e193185d139f3de456cbd3e3247eba9578daaba60913bf3805a5bb8b21dfd3d5292ad763439818a1a6cf0f17fa58fc79b00c445e1cae350a366ebd8db8eeca17493b0403fbe82b17ce620d25959193128f33c51ba06131236;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h563ed1762b90dd0e224844e32b9e90bb5c6999805544f6a2fbc5e526442755933cfe0963dd9525b958777e20df15d5f984102fc675528ab756ebd050f54cfb961fbb120757a5c87baab2c04e3528ce38d4de6e98da3f15f3a692d21c47f2e65438c2;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha07758f14328b575be233897657d606a9539c2545c60b442bdd4c9ed7853eb808eb916d83c1cf27cc51c18ea528b9186564be3b015f5d763b28327946ba1b0ce9b800e360482f273f249524ec18053a8ef8bde012057218931da0913aa9560bbea3a;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h620ddc357007ded4384b69b63de3f1e7916c62cf702e87156470cf30c2df99b743330ef003d851173e8ac0c4ca6f0ed3c1b8409c001ece7fe74a57f757a9e5cf2b82fe5881b905bdb279196693e023e60da7649aefc2f9f579d46d727360b79ccea0;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h52baee762ea410df4bd8c2817963afd47ba222ea9aeb178cad9cfba9039e27a62d0866a4f244a3d91b3e6a94620b32f078f715a1e769578d59c13e345a2391c6c5a8260bbbe2d2690871f17dfc93e0ed92e430b2ea38ec54d67dc4dfa323e61a3a52;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h442a21a5c06279d5f266938048b41ee393bf51535839b6a85c94ff6942fdae9445a70295641f1d27d1fc8d8355002b1e08b91940c60d73c90e6e7283dfe94a33affa4dcc01c17fb08f552860a6f8fb6d225e4300fb4b249969ca61fa55aa9aa2fa1b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5c6e2c2bbe957413b458b79ca6cd55278ecf17b5ce70b82eb6623f9c455003184b1667d8d887cdf67946b4dbf04398b0426907acdc6c0dde4c9666bda0d7c83fd2eeaed2eacddfb636fe027c7043add2552f36202efb34341e5a1b8e7af878d3a46e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc28a09afbba413e9e8541b4b1a46a911f941496ead648f328ad2586726906e19cd38b34328c312954f5c0becb01b40c2949086e04c298f499ad02206d866a98fff20d4e46fa0b700e506157e5ac66bdf184d02e455169d56b80d43e9b549e164e3d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb908b48c474dd2ee214ac3107650d0c3e372adad40d187b33654cc2c18a5a6cd33a2bd2f3c94fa9230c9ffe979a412ec1d29ad2e4c33843cd09ea09b14c969c5cbd93d8987f299f3cc2dcb5acf8cffd55aa2cf31c74fb0b99e1607ca07f5329a1107;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h294ebfd77f2824254e57af2a78d3c01387499e2ffb54a0a9c7ca70bbeedc06372acbc900c7bcdb4a0911a9bc8927fcffc21d1429ad3f7145bf751edfcbc885d54a4a56539ce7d2dc33bb50d6722df7cbc6a2c79930c00e3c9486dd93d7d79533fae8;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4e05e6faacbdd65b87865f3eab9440a76524ab441db7146f23840390d9036b508649114329cc5f012f17eba6d3d1775478192e0e34c1b6fa87003050c5865de7fbf4b402ac1e15f33973164619367dbe203c71eab775cbe39fbe4bebcb945fb9c339;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h77ac659e1d78cc7cbeabb62a58f172958ccf27024b931c77341f591c09ae83dba554583381e050d7660c346d3d9e8cf8b76e3893881effd091325f40d8d55b62c9531f9c60bede929e3582d54ece72cd9bc272113ea3315c478613ebe027c643871b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7c3bd3691ed865d6dac2955ee6609098c1d36cb28c9e25f08a8b871bd8c241bc32d050dbe000929dcda00a6728d41a33cb8dbc209c0c1b7f700bfd4fad1d1ce423eeaa34b421949771ff8b3629ec5d76c8377c415c989f9cc248c954e4d896bf2de8;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd64ebc008cd08bb7d03dd49f1ad8a90dc5d54ff986688dd3b6511a5b87722cb9b76864cdd8c2e13eec28fe5e4c67705529135cdd3696616f263426abaedcd5b8a829ed3bd13b1ba1674559406e082015e503e8b4d7449fc6c5d3a11444e34f038803;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hed35d118af366dd603a9cada7279b5b36e4fdad8813591a4bb0a636c13d5440bad9d1bb2d552dabb976d98be0c95e0de7ec2a2ffbd0e995e2e6097f80b98cf6fc656cfa95a78fe53313d22ba1c201f66ffc0b486babe8d74b9769593f5296af8e75;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9b66968425a71055058cc4c324f1430998b0cb838831c2ec110ca07dda1390c5a67b1216b8c7dd5f81709882d82dde19a2f3bdaafa6b7c2f51d5ed7c4775a4d2cbcbbceb33df3b7faeeb5db4ae166cf98c7493d8469d644c61030235cfbd10a6650d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h118782987a4f7aa97f69ec686a23284c676fb14f4ed7013163ac3f22ed48219871f585831655f3e3c2db8a658427017c2fe843a7b650e17b9ecd31089e2fc0be68115c7209036e81f21d1cd6ad4ac62ff718f6cfda6aacc1286ac14a955226b7903e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1c5a1b0a6306aeeef2a49412f42efa08bece7123d4174078ba86cb1a9a9829a06fd7d881352b6d81a81dc63abdd95f1babbb215d7a657208009db94b2856f0d4bd57127444815b826acfe7483d2376ddf724cb63813ae2b3abcec7c76fcbfe16697;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb0169f31ce3d79dd45c43448d6b23548614f3d623aebd828980498535a8258d18ed6b052129dca2088a0316bebe9266d9d497b9adbaf1a74d2255cf620871c4179d33322aef85d96f552d3a6fb7ed538eb5ba8697281cdca21ffff4f24ea4e8b5d82;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h75ab5c782075e2e75df6aa248d6c787d6c8ca5b9f774e9ac6bcdc64bdb50168b55538cb1e394bcdc1f7cb6f15de047ba2efcc4505788398137085396470ab2f1a1b3fe8b9b0ffdfec5378ab6cbc47a17489d7e61af1225583656c2580bb5154b815;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7f78a26e6586ab229c18bb85c8b4c8ae876db750e638daccabe47cf79d6817e72c6187154263ce1f42aa00c03861de1b6a5bea7bbb7ef17ef019517f36a49791ae706d31b369f4dee7a27564bb41aaed33429dd9117595ca58cb1e42244e6a61b124;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5f2ab818ece6165314523818b5057a7c0a9a6ff0f9d874dcaa3c1189cd275e3470a69dab291984e16db377b2567cc707e3849433563f54f05fa7ae76f7e7707a1b221b0a0ef34756f0ec3a4f569793d5d5a0c67f3623cc8b7664937003fbebc40a04;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb3ae28511fcdc67bf2ed208473e8eeb75dc00959c5d99e517aa0a0fbc8e086a37ae7a5d301ba12a7c7ce41f0021dcc4eb1270480af9c9986964e0b348423e78171c570205b7ce3a4a09cc616a6f76954be8b31abe8af3143289c036722597c016fd1;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc68f16846cc0bddc8dc926aeb1993e0a56183d4c7433ab8d9cb29588c271f20f69e96be671169ae2c353b7692a079e16552b043100322c8cb707d4f5bbc1b61ddfc0409b87e7e9c8dd3b1d514c1afa32a1cce0633daa1697dd9f034d585725f45186;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h357ddcb8f0d69079debaa09c442e43b6441348d96a41e320ceefd6caa2addeaab2b2919f9ef84ade948157690c2d00fe898d406ebff1f226e88bff97d48eb17a6b6a75420acaca4db211fbe02242ac96a7a53ac69968b3a69806d5c57658bfa9b7b3;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h898e8c7e39097c61d5c338a53649f33b1086f526bbbe2f39917b82d9c2ad4be7088f8fce6c3dfac881dc9642312bf4b59bf8af061fd0139cb2f7cbd19c3ca5c574bfa4725664f4298a8917ef4ca59a65e6cd0b24f4ab56158ef08be4878bf2a57ed9;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6caaf5959a264d4aeb9821d33339200c8d751fc09ad32b2eb11802bccc427c47cdeee574b8fe33b34bdb5d96ff74e49f73db5ff470fe6e6d9e4590e081c4e92d936044d43916ad4a0dc8b8e3d041b723a9e736f4064fb88fe7d584d519ab0f43007e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hffcfa6ee605036443c8173bfd0ef93c942469f6f2d38f4971494461e8c46796f4ae4b41d4aedb173c68b690d8fd5cb287ef317e12b2adeb0d9ecdc2378401d35e25b3312f872203bd160b22cc8da7834c97c06d939c8bd461d3ecdc805962657f631;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4f5a6158badd983d072bea815cd630e1a249a9cc24aa885e63e3ed759c17cfbafb913da046c9c0dd1fd57e94da2f7a088d9029440eca48ed19e95dfd3f91439e4859ed503e8217a68ef5b2e39fc21a358fecf78dbf939e3750fc0882b18b892f90e0;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he1d63d963e2c6b2a7e7806d2784037b9ea0c649481d38ad7aa5d1f4fa12dba5220f035f139c4ee6bb6c4311038460370260d2d75be70ccd416b2a1a8e0793dbd1d0242043aae55b5201beb103a2fcb2b8e76d869554eca2ae4bf578e75c25e06fae5;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3a26c6efc00d9ba39297bfa035ac5f5a47c49b5a303245b69a908254a2341d30836ff1c70c62da998efe58a1ae7acd54c0d0315a7688c896052de1b4851fb8d2120ede0193c993f00d58d8edb1897ebc6271920ba6b27c7228efb5ccdda23ba6d1e4;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h958ea0ffb2f380e5c67cc58ce401e2d31896a3467585e64827c2aee4a89dc921e371f5c9a8f50e4c757e4aab0c20e1c9b6569fb20ee217a43c6b5e3e90a01b753ef3c2dc954f4ca09f823d74b3bca536ed43625ad67a6cd3cd7a658c1e80664c1651;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h40e7fac56241c9fcc1c1536fca77dea5fcf4c91269a8f88dcbcdd1b465fd794f6c0fdb911087cb5088fd33d35ade81597c5e2ed78c0bfddbd08eef85e4426016bf44ce38247cb84ccd78947af9c156fe079e0a9a4d024cb35aabaec0cafef6a7929a;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdfefcc08d6dd3f5c477ba4d57f84ef99b8cf230b330b526c9a9d38abece3e27bade94f13c8a1585b4455373f546f1f81735862d6aeead4609465dc83e886f60515b55c200457c1f579212257b8c31336a3f9ed6b2b8050bb7c03c75f897f1ff7552d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he5e16f01ef3b207ac3bd201bf79b9e3f63b93f59d897a88fd792be2adac29b0c07d5bde6d7e748095d824cbe880d10fc486c5216dc4a6f3ac6fd0416d59bda93962778a7ad572a955a1a2e7354f5d409114a766a7754210f33a41a0ab4e646ddbeaf;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5da6af294c6ae101ac2a16fbd88e74ff68ef32f644d968eb2fa62f300474620d27cc4ad05c6495078f445ec7572e5bbbfc8f7fe02e4dc0d376a7d0b57675e3ad407a98f9ec0dab0b71b1cba4c8669fada65a36d4b023671a6f986b1687434ab06303;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4c95b825ac7c7039f937e205608fbf573d72a6cdc5511dc3ee2591962d846fd8e765411458887f0ffcc2c7dddbaace7408d2a42bf6180f3f0686532ce1a993b523ff31386ea3d27e01a4990fb5189e37ca113fcd2d7de6bd9c3c893d1e8173c9563;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2b33a39436e66e358ce54a12d1713714912e3228c822f88e426494d316444464ce2dcddb213e75a41d87e124d023551b32deefccf9649e19fd2db96e25052c97a03c4ca7a2d1bf362da7cb203934b90f2456ee8e933a3cf72d0091a184b11dbd30cf;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he435ae4542f4187e2d29a4b5b39f6ae57d90cdce56e92113e7ca4141da193e4ea725b1b2d6d3a4812fd11d1cfedb760e4a8adf8e131acd1b80544b66f96653454f148a601f5550f864f92831c15b8de398b5bfffef3f07ebefca3070dc699eec2069;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbd47afe87937dd7cd114171ae8e829969bfa79b9a071cf82ecf3dcf30c5e006763771b83781ba8970a7d2644d0ef4bfd7a98c7868e1f3f65f7a618ec2416d7455d732ccf9bf840fcbd400f9db553aa3422661951f570a899972286122b0f6901fc0a;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h53b2b5dc0abc85572f73128b035094e0d02eb74f92cd4e98cee4cd768f2156df598f63c40fb435ebcfdfddbd639943077da10bb210e0d4324033a81097f50b41100362f8c1d56a15084421fe76484967b3f0060cf0e8698903a81db51081d16f3137;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbc42e664cf65cbd7455c2ef8f2388e25693bb7d4ad1fe103907088301f3ce0370cc67d9f0548779cba0365ea54efed316998c8a98d3434743ea46e5c5df6ed7a2e793762d7bf6bc6eeeecf4d505038b7513626dd526552dac32e1c6d0012600eecb0;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h60dc505053526828609c14ed5e5a4219cee52192ef3fd2d03337803b67684b338418e285358be6c20366f0f0ed14d18771f6fea803bdf430e670bf1a4d6ac78488188423010f2574fde5b22fe19a9a26f2117b95d59235960e98a2a02a59c2f41dda;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2d5e9fd50440b6961c9b6ebd571a604835fe98ffde47ab70cfb28886a334c8ab2ff383d804b1df2531557bbc645ce69b7dcbfec17bca328a997597ed9878a15024d29d48131b9d12091ebc85c11df3e1bc1daec8bdf7588e7276c2a82902a09b19cb;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf070045a46a61fcbfcae5fb90f36f47ca07167b21c56df7a3d76df84a7a0daed7732ec70e7dce0addb5f7b86a6958e3bd3267247d69b1929500be542a91667dce86f7677af383e73d2b2996eda3ed4202489bae1d5627dec553fe7ddf2b525929ad7;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h407f7b966f02b192bd68c41e0feb705ec1c8be3f4279b50f958150889a7fafba3ce85d27fe56e10ae72e0e0b58554f38e175a70f35ddb752757e8be3166451f0048090d136a4fe0930357dc8f446d148d798119a3dd8f179d18fa3860132edf9e945;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6679d276e0b71ec439da4f0cba39f6430e45daa411a4278ab972b1e07b78ff7af7b12b25d024e49cc9f2569d6eb0f1877ddad4b7ef75805915407fe079df46977565ed688a7617fcb2e98302fa4028e42f4607eba79eebc1652b2b25870a98283762;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbb508189a0518beeff79b7cd6d531ca76bbc50fb9276462a792c3a899b239737f14a04700683364d66b0f0e52e5a362c6a987aafa9119c0333e2d099ed1156f8df64ddd08858ede9050284e3a66cf16ff8789d6f6ed1f5076e647eabaeebbdd6b71b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc7b2dfb2c2a368fee9b14207108b0b148dcc81e69aa94ee11cb0dacb5bbec2a54b7560885af70363bc6ed519506159f6a002db8fd8382cabb67bfb030711adeb9bf6dec230d9f8c181ef8253a20faff7f63358e329876ae45745f118909dbbd1e0b3;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h93babacde2281c27f3ee7870a631689606536864e90c7f8e4684c8b93373d4369b6eae596b84182019c64e6a765bee028b1515d9944e61fd6d4983dff92c420a325a62bf13336491d8b8f380c7bf6e03a55f1c5b2a689625a4f5412adb8dfa47a13d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h726470f5c3040050e35f9fa6f8be1b623ba9b747de95e4c058741c603bb220784801a079b389ef5bc8c064ebc9b2966729afeed842e55b23595bb8d6749346171221370765ae7e73d32ad71a0aa5d76ba021f8f13f7684ad0e5c1cd27780d907caca;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'heab3b8c71e5a01cf6f4d176ee6dc7a95391cdb81c966c62fdf99dbfc71df62eb9c1f9123b698aef88e1d8bec6477de0fa6029b6866c41973306428381845bc08f075a13f4eaca5a9e86ae05f47f26adbf56de6f9f041889633b201e6f89c472e2304;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7fcc8d44effb4d9a57a44b6cd32d361e51370abdd719c2c7258000a4353573db0e6cb9e9c3b061bb7f1f6c2f759ff1d1b8ae81972ee2d0d9ba3aea532f56fc074008261d15682081d5e9d969ab4195c9b19de777739e249fb3e2699522481fce58bb;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8398b5e0a2d3cf2b8828b57604a326408015b2f3ba5d4588803e22781e8b1bff770a71af7005b20ef3b114ff01f55504dfa5a2f34f1438ac1a3d2f18392f0206e7abac5ba82cc4563911ab3d9bbe610fa269cfc9faeb227893ff057e0a2de9dea1b2;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha3144759e7ef9baf4efa0a600f7c3fd63866bda0936a1da0e0ce25ab89c265de148cbe30369bbfbf0e18701a797c497676b8058716a92dc4de4a45a4bcba1a7b71c096ee6f08e6255d60c1ea4bd87bcfd5df6caa9abc0679a5d4b9e30b2f7912d72;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h33f791cf13ba80268017476bb8535918ed54f31595fe6b604da3a2fbb03c9ec94372f2973e37762158017f5de400c637c9d109e662b2fb5ed68841fc1e919a20282ce193ef1f089277cbb33714f2e45c7387670cd07ce1c60055e36210a4d4985d52;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbd3fc0ba3b4a232a477c072ebfa6b0f69fcb50d4f35ceca1e2c1919e33dd9a663afa0d6b977c182c1271dcf6b39e8ffef6faf17062ce1a58b3c228dda802ad76649cf13475d4b1c6b1caebea3e6f99c34362a653db6f01a63fd92ad904b96821ac71;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h833741670bab98f8129e5f42201ad0e1d10862f0e7283ba1a3117ba86cd333b4ae72860403749a5537b598ccefbc2f2a28c5131043ad84a70401004bd643479788c9f0ac86a932d0cb98ec99e7cdaa21129bd6994576d071a4d18fca638a1d02660d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h62b704d2ee6d61909ee9a2504a9520f8967192033ef931435b755b5443d6d151a0fec279b95f427d1a48214f5bb0fb018a4a326596a513554f37193b47fc74754d5a9fb786b147be662e83e818f666889eb6d412a52eeb6d13012f57c5b37b37646d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h84bf98c8b5f650e6822357ccc56c224cbf12b2d8f2a9dc83cf0ce4152d9ef5beef0c017e834477f75dbc9befe58408ece996ec5a6a750624af8058ffda434ed79b64951b8f47e163e121e30470621b7ec271633f37f5804b709a28790a6317adc68d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h327449b6b5111099c50f953491e71ea1391978b99e9d1c3b38201259e723086c4a4c3bcd729743046dac28cf40139addb246078596e16e9963d8f96de13bb4dabe8f64a5738cede7323e069df1340cd1ff2ca62789148491aab70061a12d938ef7f6;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2691208f601c13732da2ac5bb2cab436bb211a42ea2bce7e392ed432ee53f5ca83c8ba619c9b1331ab1547f532a67cc2bb6f065aa5d707931d27b2015d245f30208309dd19e7bb5e647930060af828281e6a4b61987ed11ab0e1b9eb33fdbf535a59;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4d8c0379997aac80d98efecaa11500c9a44dce1c67c8b04cb5a3fff4d6735008e9c3fcb784cc1c3e6e030264d6bff00efad4122effb8a95fc6e61e7be3da830c3673a4dd4a9249e41f149acdfb2ba28da73c5e116f6646ee71932aad8a5b4918bb8a;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha8a20fa41584600fb97d1adeae470bee089f09795de6e409acf8a2efa29eeae6bd7e0b1bc86a29eb31939561535724da20ecb144e0f3d7f5863f8d8a45ed6e64ddf4334f9d7f92c9507e7830256c6566c08efb3818fda0a6f4c89c98bbfd49440625;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h857679d8cd43f7b4d5d04afff530d72116ec6ad3867f8fc597d1883ca7799d017ad2b6ab645544ae11053390cec14bd7b4e47ddd62fad21a3e57ea07f2940d05bd807e2fd67352db54bc71fc25d326b9da1a2a3249126afa1309f6768b97c32a923e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h76e3595bf753333fb30127a0aa845b4f86f8eae58ebb1d1543c6376b614d235ce27342b0ef6542bdea42fb5de6c75f87fda991be00bf4b45768cc8a79671c626fe44a3fac5be606ddc48b89488afec0eb90b04439f9620272eba1d8a7592a893060;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1e9b1e9a1db4f519f4510b6387370e98d11fdf9a0233a7f5dbdecf2fd596a4d83f4b5e2cd180eba5b679be54377833425667569046e801295d8f6f14e84b7c2582c73ccdbbd0756a84b2c7d7e2654c57cf31ef19257ae7c8d01a8e7eb9f44869365;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd746b169fd789558cc8feccf3410740bec49d58f0a12c8da01cd4410a6cdab51ecdc10ac6f495258132343b40e8a9adfa3331a3aa8d4814a7b408f4b5b6bfd8304eb49a509651d078d9d0f3d344a10f55a446974f3b7698fb2c5bfd27c999bf3cc85;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2aa25cb7f62ed5c02aa11d6a7d61fab1859a76046d5cbeffb61b21ce78ec59e37921c37cb72afdfe5c3d5bd99e6a222ef30bf3af179ed72c70ef357799b332fe300110a7ecf0c6adb6d1583b8e4ae041e600b92fa2be41e5c790a9409276f370e634;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7cc18ed292e783a26fa7811f27bee976eb34dfda90164fcb3ae694a35661542f433e0016ed7c76e443ca829e8cba3d2a7f843cbb9d2141a440c6e25335032ae4a13a883aaccea0a767f5722eb43750da3fa8ad637669deeeb8b5a720380ffb22be07;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h16d20307eda3e68a58d97f36e04801af42dafac71d9da014f4bbd1328dd17f552d53d091f19f2299eca1398d464ad26dcd172be363520e8fbeb20ae745814e6f2db3ef931bb1f87aab37426c3b17852475d6da772cc6ad0c0e1a8f2cf9e658a25ae2;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h62a95e477002abdd24e6bc0bad24c53bd0e1c50b20b0306cbdc96657e8371a5251c799a0ddc5169b21d7adfd26728c32cb59a7f649c3013682eb14b339385404c1ade2e6eaabfc9ac2c09f80264a8f424950243a0edb1fb57118be17f7fa23cc0b8c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbff5d3ad5843192300d6f5d089d0e9b353cff36b956a04ada1c22ad16438d2746dcf8f96fbcaac41298d0ae5a1c6d5208171f82f268cfdf735a6aa26277dfec158e74c153986ae00db9e699f57d4f70c3807503d7c861b43d3e139ad68841eb56da8;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h753f38e41d04068c1345ec5c9d6f9b3efd6db8ee4fe4af7bef29c0e306b141deb1e71533c791cbde2ba27d99a0b3ba7dfb1060bfa8b9eab1299e1eb22f6b8ff2acbe48dd9363553252bf14590c4d83829ca9b4b7880d6011c46680426f89db36d2cb;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9117f7b88224fac5fddb7eebcf64d0f4d1e92402fa6d0da6f00d1acf78150fdd40a18c7765a23b1d1c452ad466ef7847685d06e00f5dc2976204c48a9d13bedc2b5a70bff3ee6dcc4ac229e29ff5d94cf69ae53fc5bea9516229e084988f7338248e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbd1f7bc338f6a05c8d4b5aba0d6066145fff521e15dcf9ecc234b105767caef4efe5dbe3f05ccdcd4e47dba87a0d78fc334ee9f5e13af7023f7e33767cf9b252cef9a5acf9d9acc1af871f48e8c98d8c438f8243036545d416685aaec5e45b5f2fc0;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h422fb5293605fdd03ccf6135bd39e4e7369f7a1b0a563abca9e3272b26903ce2c413cb289e7a009668c3251deb5842772ba1f014a04e3b83ec7de1dd79f006861e7a8b4c1c8c5ba7e5331822199cbe6b591dd21463a57f8a137986ff849088969b07;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha1bba811771e97df96bd8e8bab8fcd1a4babe47aa41bc0e0257d485f9327330a21abbf033aa200964ee420be91d0c437e54ec11de93ebd909c273373bcae9a269087543e103ebd14faebfc7504496d66b432bab0e9efb9d83f395945878be5562645;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h21ba4a33366471b1946649b6e1adef829f326e77f612ca3df496a456549f2df4d047227df1b28b00b5399a5c571e8215dd986a973ee696ffadeb685ed25fa8c3741a9fe55ef210bffa41912d3fce41e054cef3f1e4799cb1a66be609669d89012a7b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdd144f40450c039130e1bc9bf2bd31007b68fba45799ceeadb7984724a294204b4349b60f3d8f12667a57d8219a63e0a7f9f850fdf6a9a5f2336570daecb6203db85cdeeed3a009fab77bfaee06a7dbe8f5dd0bf0eaf32a5e5902fb79195029d7763;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6fa960ee5c196338b534836da92ac2e592182dc8bb53619ec54fb17a47669cf043b195c463341d59e501538f3f3c4b821310f1bee46835e92417606bd6fe6b3cf1bae45ab8f1e1c2cff0c836bed02ae22657f9cac0ffc59f6470ac104dc58b16b3b9;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd033296c6e500357b58cadfe8bf3a0c5ecc74a7243ace751ce23636a530653220e7d9fe64668fe4a9eca01154368007699f22aefde8dc0d1e80ce837b7f2e90c8f5ed217f4f019f6670c7b3bcc98d9546f6f2ade78978e46c8c0d9aeb9a4c40dc6fe;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h513d846548ae062b6fc68ad72734db1193d5543c287cef652713604000116d98610bb4db7eea9312c3fce2c0cf81959c2e4ec600dcbf080d1726a27907aa66f5596bbce40168a39b5263d2d28fbdd1fe46ae77f46e2d92914c2004e8620d212afe9b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4fb1a50b21d7a0170742edac74288953c29df700eddd6a27ef1f8c79f236a88a31cda0b0ce1889ce5c7b3edf24afc29cd9f5fed8b26d0b02de241f278dab272b047abeb9ae5a0a2c6c1ba6e301e89a19fd320aad67392ceb0a8f90027c1959299011;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf8d6ac8a327835fce9096216bdcdaa7c6903bfc9855d3779d40d3e27e7ff3b41adafb51d073b1f3747934444ba69a460791a3c01a5627235d9e81dcee2b442f69c8b80e934b520e4d098e8d3209c271308d4b9c74aeccac72e59e9b2b6626627c0b2;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5cd05cc39b0cc2849875968809da0d2cb020fc969084aaaccb4ca457d13bb25507e28d07cd418ee24500f5230892bde79eb0c069bf155b9ec82256ae23109a10e64669c4260797a9534ea1ed279e3f9779e1f49eaf34b38bb02ecc704c4bcd0d82e3;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6f0ba3d6b7e103247d6c5e558bdd188c8d6c8f51975000e374411eb16a19c333031154c122420e8f5140841bf3fdbe4ac04f289bb78c8edf146c4561ad314561c74fdef0786ad7da0c18a645a07c3a6389614e900c3b711b283ce12a055617dc552c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3519d98ea7a089a7f2047a7c01ac10026ecb7aa4ce3b26d4cacf943d57e3a878e14fac234c683071585c985c2af73b4b60c67d0b02f9774b1c6edd55f1d20e4ec48caf93deae416af494f9e4f5690f1f6c3042cfce9885be17b74b3109c0bf93e033;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb6cef309e5fe31922626d3fc7ab60bd484e5be808dda8d3e11f84c0498a49f9091d84d0b7b5547f880856cf0d330649894856a203c957c10b1a168d2c30abf31d0f18b4f717947340c128a5a07cc669e659d7cac786267093932f52d87316b68f5b5;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h79e0077ea32dc1abf99c9a59643180a7e5426ce99665effeb19a35f5ba3981ab0f9dd110408ee550b2e05908fa3ad1119f968ea39974800726f8e8fd3a87ce203ccb5e81caeacf5e8260bc16547226e51030c70f33e552357ec5d3d3eeae8fe8c72e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6c75674c356213818e7d3573aca28ebf670d26025da5cfbf37b7fc244082972275342adf83b2856c29092815fca5e7e3e883ca59aa7db1aa0813f688ae8148e03cc9b6605cba81e390e780acc48d02623403317032d095d7c75575d90567fadab45;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd81b33babca45ef29ce2c4d7aad46d66035cfe098fd89c4c132489f6c0b03de57d2829009b216a6ed42444c2d74cb8be657c53558a11454cb82b52a3454cb321b4368bbed15a13b34d6aaac247c6cc5eb6bcacc5c8e2dffdc249a6fe77e87afbdeb5;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha1ef11a2ef784e054e1b174ae20f4ad577ff733d0ce68659fcac50d83af8f7af86696876e06812b2797b9e8bec5b09570c5d19ab25f980f844364445b0b8710a2bfa4ba8f4b21b4b8721c4318edc6a58d83620fb6890149b2e9e6c9eeb78f329c510;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h19d87aaaa94483f659752465e6cfa74cb6c557cb8a4832d1379ad532a8a72a102526b5407861865421758e4aec188125c39c4a521065c922faffb23b4938c34d28354c2ec9eb4ced264bf1d359ce45eaf1bcc10ce3e5444524fa7e8757f6df50269e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he1957bc6bddf1c71b25cb2b6f1ea4f1b30bd75c04a7c841a249a43ebcfeac85db169bba66de95514b9fbaeaa4d280694b8bc63536c27431c7434814b0450d0e4f8cc31cf5d0d7225c726628b76e702321382f7079e705ffdf74b346f24e2c538c4a7;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h469380a17d240bd2e3449478b6afb100af5982d52282c7a3a9839b9d6b6cb8340d6826a7f503edd14f190bf8092c38f4f181345c3c0a946be0d9d2fdf53c7d339f53d947d2670aee74e830058a3fa405095fea7563072346487a026f077d7cf3633f;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8b5aaa46146c0254ebb302862cb330ff2fac45e4060f0b5e6df657eeab4814c31b7f37f98d6f73feb6487cb0c63a7cf56b0985d6fb509be4ec06c7cf217571d49fe83dd37a5b0a2337deceb484f861d73ba15aeb6e8ede15b715881df633e70a03ec;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9967d1449cf0727284515950f8ce1b39c8f6d072f75c799f3f314e798b5ed1bc0f3724a20bdeb7a8e2b23f46883d51d346d81ddf9723f36c9385f7525305bc6e04ad2f23d2b993973b56d764f64b473c742d125e0771283fb1165f3f5b9a81943135;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9f359905a41c23f557e8243c7991281f8acd47743efd30329fbddd57fd134ff6e58ef2e8c23c3ed8a8836f22d35139f66114b4cd2458294dacd96bd5f728e7d2b8cde009a48411c20d020aa450e9e309abfeaaf873eef49b6799a30b4b61cd6e3131;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfdceaacc0eaac321a768f76dc34f5df4abb6554d364f60122d14dec02e04ba67d434a7e99d1efbe40d8604ba926e93988a6feeb8258ddaddfd343b53dc27c666b53284ebf76b9f24d53609e162ed96cfca65b7a4b3d52d69570a825acc679bedd538;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hadb8f643608aec671c557e60622eca9f7ea78ff5fdeba317d8ba3ebe1150dab80b2eab7572d317bb702e3de0e7ffb69f3b4e9109805d2138cd2e36e165c82277a1a4a22e1ec613c405dbd862dc0159b6723c7b75f0116099af2f27a452a3eeb3e40b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h45a22d8bce944a904c24bb2af2a27c0b1149a03b49c88eb2c9dfcda7792143f1937823602459ab1f63c16578e1320531d4ef7235372f7338c2be91032261d1e8aa473d07af891e00a1fc3c4e749ca57feed4b4c827b4e358b8fa24657c1a81f78217;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h61e7a52f397224343e0b0609259f39d72755100d74b41dc486fd0fb83c47344afa87041872f8b7451f5ff10f1af7af41942fd6ade1c79fe171cfba9e27fc6ce2fd2480c7509996b25ec179ac43845ced89d82395739b65d7930b98a1826fe8536e60;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3cac65704274436bf133cf24e9bf1674c63b97cb8b25d734a539d6f1e98cd541835cd546e54fa3533d27e8134f3a1cfa13e012c32ac10605ce674614a167665ab85dd8b90330c6fbe893e8c8c397af54c3fe7ab1f6de7604e708dc78e0d5e7319523;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6842be30cf07eb06811b8cf8ddd415cf9eecab44d27b38cfd9b5d33efba567fe240828d5cf85ba13ecd9627a20eca60b004956c7f89eabfebec0e1f623c0d7f8355a91bac4623bb218513ea67fae65e6f7e197b68fab1eef96f3837e8f59fd9c476b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7ee0829fccf9c0c52efb98b9d6801c7d1d735bab37f0c68723caa5801350ec595a702c06bfe5253617aa8c82b115b9e606559ceeb844565d826dc19a74ba5b99bb49d23a8bb8f1428291d486436ca7522fcb7bf16a8c4d496154d8c46cc1b0e04e8a;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4b4229451612d572e3463f36190a10b9332b5e7df1a51e501844cd4ac6065a5a5c8617b9218e2089beaaa553ff21cc221724a353db0aaecc6adb06b533d7158256d1641101a57d66b65542894f412d356e04c28d75bab5cad93de915d63896c3cae6;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6a1f41d8f5b51f2988eb98d16c4c24a1947c9b1fc9bff5613a485027cb2c9c6ee16021241db1eedd39f3083400b4ec00ee41e883975bf5081cc960f4155b1cc81b375d153fe29b1e88a238545fb9a764ac4e84c64be93c14deded8f54534d9507276;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h68e6a2e2ae660607a86e85478db8bc6d83fce3eb230a9a4590dd76664ef5b4e1b2524b22346f32df73c737ac32dbf53daa3233a44049ada2e8f0246ead1e925685074ade42d1cf240a25cd99084353d82154e488154af467751cd4117a7ae3ae19d3;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6fb74a58a763d1530760080724589a1758a57b29ff20440bb67296016186d6eb866d9e240083f6c653b11d808a52974ff0ce04f0741d499e85a9f1b8d9a7e3da98268825502fe25518fe1013cbbc852922ea7470cb57e4ff80222e9acc16893ab853;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h15e69a3b2f029ad7b367629ecbcea162f2150c917140bd4e7c554f05595c8bf42f09e1aa848a9c45b67dcf0e5309a69ea7541fb3b8d721238085cc90df88a57150d74feb58edc15adc4591a6db983be8906a95e632be78bd6b1fc95dfbbe4fb6f3ce;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfb6bcac9b03088f83383cde9806540f51173bcf4d84efef2b56803c4b802493b9cd24c51b3293029923cb8773303ede662b081f36c76812e3d6c6691cb999d4605da00b93a232bb4b288736fd4b8f104766c393feb4e60ce88cfc04d16fb296952a9;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h49da600da219df265b8652d903e029986e94faae0b9845e13ebb4432a42f39bb4e013e4a29347d46c36b49036e4d5df2e4f92f6f56a7b2c00352a63cb1682a76115d696c4ce6fc36a6ce3320a7d0008e169ab89e149431d739e55643828c63924247;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8861e634d49235983427aacaa411db103fa28db2c0a1e32367ca26ae5a729aea6f2d09cca30c68a2df82590fc5bcba10cd99439501047ecc29504f300429a729608db94885fbe8473f5ce079c0e1d42a35c33d6f2662f105899347fc677d267ea2de;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'haa739a5d0ee595c9458ec4e1de4db65bf73682cc41531d346acf3cba3d1dcb345a70e49178cbe29690e9f174b5f6b726c77daafc536b3867d7505b45ff0aa21b9f9b4e52323176a48f8e07b8c50df7a877016cea2c2094b4c9f0c7bd1a23fb79f3a6;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd32056f260994704637559b30220a44e4e6fd4edae74046b9ac0a71273a7d1f2e530e85c1bbf609b54182598a0dee529ef231acc74e9a58c65951fe157ff5f3f7d35dfc2868acdfd7014a7c5d30706794a8aa22bbd2b51e6aa41ed0f456299e10b31;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hebcb1b996af475818e1a6d9d38be6ca95d1cc5c3457155686f732d78c49cd57db79af699a727175876fd32a612a8dc6ec905cd23d832d59af8c052af3fcaba840fde05cc77003f751705951b7debc779dfdce32a449f090ecffdf8e73c0e4f017165;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha75b05c596551cbe2a61ca68f9f347f8a032195e2890a80a2d4cf6a0e5529047da0b85da12b9768dd050458e8656b744341a9e1aa24c4716cda13d9bdbf474a09f778844a30763aca32cbfe8e55bfe7fae6f856697af6ed18db85fbf3467e4aca4b3;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc75a99d957a249182b5b223daac11b7b4cefdfebf4ddf34b321b82a8a1c819891c8594dfb22185dd26cba4460069de545ef11d0b5ea8ba5f79b6f52c8262d2c7476e671eacf93dbba665d6c428bb485edce0a6e700eb643ebe418ea15a35d17fde1e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hafd0ddce8e34ff3a88fe48ac9c5d1b11572e76079184b28ec0d3381079cbc1acd995f17449ec992c5055518ed2c9247466a87e5a784f2af4d477bae23fe8c14cd9326db76fdea0c140f7b96da1d52f6bf035dae4b3281e41a9dfaeca1fe015163c1;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5c97be4df13387fc099309ea1f8c6b54ecc6167f1883082137643f28973a51a45a887cea45fa33ad582b2bd3dd5fa9b3658777c012cbbe52da8c7ea91e74514f78a97f82dbd54ebd4b0e5eb3cdbf491a9333312cb4a840d460513934233c9fbe1bf6;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2fd18c428037da962853b510f8dc8184ade1bdeb3a953f244ab91b6b9a73a5e95bba141c4ce04fb571c22553c1b1b0af3e57f61dbb95e35c7306c5635651552a7598c033295ec31ac2aedecb3a8439b5dca289bb6640cf58abb9854516f72b94854e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2959e49916f0bd48d64aa45538c11ff008e63ea8fced368f751df69cf78d8174a8593f17853eed730b5a7e59157949a67248e01d587ebfcdd3e2c96ed5b55f3251e909083dec7d27b5d67fac862ac7443e6ae626cbc81d44d189e6fdebb2b292d707;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd56dc6313e627ae8ecba0205fc3d52ac4bca4b94fb43e37f72d4da76938cc5219199139d283fa499a903aec5511ba59974a5cf2ac871dcf8ee7ffd0dfdf4c6df42aec855658b698c0a885344bd9ca933887ee531bdbcf6bfddf647096f0e3daf9129;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h70c8f362df4932e33785679b342403a1bb5d371a225e5b4db562a37c0133e7dcec74a8cca3e724d3d3175243bf9d1dc7265ca174d9e76894ecb7056d972e13994d46d60ce6ba743dd014c6ed6e19622133d813cbe6147cf346570eefed50e000264d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h638d36c8d08d2a3b750fea3337f73214736543dad6d90062c80752d506021d3f11cd51d58cd87dfe28cb4a894d6e5de81837b63f2d5f8a2b569812fc318251a5090b2c9e6b8e981a231ee6437e1ca36c8f5a2c9b1cd3879787e84b0b59d116c70878;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h890ffe44a39ef7b08fe17364f6c2b1d5fbf493e86ca52449099e475488617a837f69d91390be0a17572708acfbb5c26a10b1c3041748f4d90c620dc32e37115cddf391a500012e6472025efbef74d6c65a9c053f64919e3bd4d5fb4129962b40b9e4;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3616934a506e9dca7be15693748cfe412c68f280fb1434234dd6b3474c0b238ebe4e53f18f8db483f08c7dcfffb8e6d3d37aba4db8553d18f29174baf9c3263615b67ee6ebbd2940650c888db84f3daa1e0f60ecd9791988017eb3b5f281ed04cc2a;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he0d410352102fb8cb59e11c7c7b0101648a585e8515bd3f56c6fbf9c0b8186553a5fd924db61b83b5c86283785c5009be972acb787c67c760da16a2a3ed69aabd13bac2822b50098daf8b07093ca07ca453392cd50b9b828e3de3a20b59c54bd1210;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf690afccf75751d0dcfaa9cc0f215b20781daf2c38333b663dcc0fe900bd4d70be3bf0018e8c1de844e681f91e7f46012230453a1319b58f5f31ad9ffbda1d267acc3481ae343ed99c8b3d23db89f44ee0b8272a32312bd2d73d9fbacaae2f956e95;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7deeaf4cd4cbbc4437f8f9be5472640470c3dbdd8391d95836f5d712ea8c0305fed7e2525495a565f262dd13d18bf35880678f95bc5b79e0370ed667878570b6a33c7964abcdfdf80548e827be89534173889c245f6d4866a22265b80c48f431de05;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h283edbc6d602adde68a7eb2d165f399e9b664fba34668f49bde848bb2d47d0ccdb9c19b2eb073ff8f41ae08e9361817a8cdce78a747f1c8a122ffd49b446445877320c75332543e0b63fc6f40b1bb1c915d0828edcf2f7657ee18a5c482f7d784429;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h946342746727106bcbb66be3233b7bf0f26b3942bdd430d2ed691c78813c3c618238af40fdd392470a77a6b51d0755f2d4b00025a47827173e96cf32239c908982d775566ba27449d1bb70ab132737261a6011b32aaf757137ae149cb7026f2896e0;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hcfcc126ee187af027757658b4d3d42cb9b779e147044ba8dd118ff5e63be44b5e93248caebf7348a7ab8b7dfa027e5a4d7cfd74bf4c0e88e325c000cff32b6d9436118bd518651f1346ddc34e3a34c679d1407ab3949936c751207efb20c7456914b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb16b7bb9aa1e43e8fbad3fe9bb5ce2f4c1e9f018cc3bdf021f0a7f070024a10176d4147766c3b0b4e2e98d8cfef2a296e7a7a8727679968f8ec0266170adeeb7e5242650a998dbd34d338ca761abb1d7044b9b22daaeeacb32b79b44310653e49890;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he6ee77b1429b1bf391ed510b2a659636435b9609a829516f0694b732c1057ffa38caf0a068928200ad6511fa45eb7590d5cb679e0f3b63fe59ff9d4e06927f7dc9b1a3b535e97a09d6bc939d8582382f989ba7cec6aba5e1a82573d5d9986d29de33;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8d6b7f5dcf1c20b88fb85296e79c66170f07cbd6d7d38930caf81332c58c61d513384fe39546ba28e27243d4f601989b44ec829291966d5c9f045e7fa0d6794007ed62a03a1318a017530297ebcba0aa77ae3031f3544714605423bc0d1971655c1a;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7e0219c7e5006203de4319586ecdc404ebde794c2a5353a220b3d28cc524ae6c1534cad0563fc3a4be4fa3166aac061765b6c2a7745c7c702900b5e933bb4320d871443c1e7bb68ded28793eea73aba127b3a72ec6b699a4b2629897b8c680f7f4a0;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h88508922cd2f5fb45090c60da444b56c2dc551b8257b10e30923f887e2bd7f4dcd274498593807bffceb6080c9f39bcf864e225bbeec768e4c0e37bcffc39a56e5ebf6e31325613427e5d24c873fca9329d5f48c09df25ac7418785dde92513acd60;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he3002b43e721bab187bf9f80a637f8bdeb5d6691bfb07d9da0886cc6a8238cc3c02c234fd4d10054903b3eaa0bae3fc471548d6b028d1ca9ca52e4810fa8ce38ad166d5fb827326881ef995426e2faed29fe056f706ab477678aa0d972e7f7916d51;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc86809ec5bb99600813db830c03bda2e584c21b82d67536f011cb750adbc43ebca87ed5ad0b2db19697b4f3df704b2cea34320f7e761b975720ba7c473c4d88619daaf6b7a9af6b1ae6c170c64c0ba6b8dc3a611972d58e70385c946bd9ff5ae30da;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc50b8019dff2a015530a907a38af2b8bfefdd63683a52296f6038a4ac97be8ad38b97b33bde40e4181755d642c890c0dbc221694e9861a323536898184c3f800f146f653b81b8613858c9b951457bcaf8a30ad2580548bc4fca287fc571889055758;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb58d6eeb3ebfde6c7dda991079ec4746546a5f79521a30b079a8b4cf6f2b6b3d7771b8fe3c58806aa27401588bd037289e81f56e935d01a521013b0a7ffd2a5e030f0b3adb8aa498a639fae34bd4e95833caa29c34fd8b1ae91a6f926a11b1df2b24;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6790474b4b85be447c42e7982be841531cf19960b336a4cd19cc8224545284aff20d799157be14d0492baf9884ce135a7ec798608f3d8c459f4bbb3a3a468a0bc6574da6e07b4c68a1c9f9ca4d5957a7d90d5b6f771ae7350a397216658193a06325;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hafb1f1152c3ea7823d1ecb46d0df531e689d5ee53c1a5bfd3da41f344aaca9aec8c76e29214499fa0271b918d81c69c9a0378fc91db8d0a4bbcfb55bc50b543d90704181c86e80028f6fe39ac76892dba94c36b56f76bdc1321933694e47d1203806;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfa000cdb4402ec726768cbf90e4427be04f3c02cd57216784f426d9e10c2736567f013f736b3bc933a745eca01ed08c98ee417f4bc675bff7542e5582e63713045c49de2de01aece48f3ab9c74a2807b270d708b1ea245609581f6504e8cd1199802;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'had11788e5e3b6e052380b0021c617d6b110052582238a546cbdb3c26aa6682baf7574014fdf880c1d2cac4a3c26853ebc6500614aa653c6adf40d35ed5d432d0193613a6384ae72f1f0da2c5a4cbda184e1241b4c8c8963b753be55e381ae9bef00d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hcc14ffd137f80245358c4cb892230a85383c7afa484d27fc610b83912df101280588c1164cfb843086d3a1663959db07db51239d0c1b6ec1198cfae06fac2c90e923f7dadf405f198c1e3ef56739a77e76c8ad937b85c8c303c09bfd8b3914ba3211;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7c73c1f090fcc9bb0c5496c7c1641c034a42df70246074db196d85cd97d25e00a894a53f6962e804637843bf689b38f6149c118955a270dcb16bc44be6964fdf80f8f55524c6d5406a3a4cfad15003df6c943336713b5ca2e74b2fb89e54614b9b08;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he080efd1d12e89b4b549b10c12a78d4dfd4f111f8f83655344ab8215da77d00518914858e0e571ca2545a291f647a83f7f198f53dd4c4e9879636efb8bba4f0e6cb8cdf3b2bbac31dbf0317b642d61c092e0296c266db379d186043193cff630011c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h36773d200322616cd3cdf42141a2550c74d58ad6a6d28262cc8d5caeb41070874ad9cf42aaa04f98f5a2d1bf72f46c27dfca1743a66e91835e605d8e5dbfa4500494d3e3f6d7cb2dd3a80c8a1cbea1c0eebe114ea15e9eae12e7a0ba95ca892b0445;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h58bb4aa998229571e05bbcf1f0e7f5f90a9486ee7675945bd33e804dfb203af1a7099f71bba188c2ca979e2cfacc5de52292db2e857a61fe14c9041e411f0bf4228e918f99f4444cd07068296702b71c709ed1ac1ca53c3b9ddd03bfd5a48d605301;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h319eb7fc3e43e63f8430ba73bfda9f9afffa885696acaab79f3f428c039ab58422cb32005940a74b43f307b0c9b8c36290ff34506631a7e30d27e0757f5f1932f932d27a2d61fc33b005d3411f68920b06e54791e4cea977ca03dba7c87b08ca849e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb7d39e1f8bfc1e7f678572490010a6d386fccf52ee5fd3b2528bd42ba2787dbc8dd19f7223afb26902df8011fcbac2ec532da99d641924ed2e23bed52ee98906e7669ff7f64c9c91f191128d9522915d342ade67a58eded470b6f3728a5463a580df;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6d8befb565cb7ea6daa16461d6def5c4052d962b28241821ed545dec87222f26e35022e912adf1e962ebc903ad597596af61b35997f383087e18d67886d8a0f464d5a3308c4c83aec0f8a571f823a3f0c75d711ac23435e4341f71669805809e68e6;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hed7bcbb31e78c66d496f59ffb86cd6736ff8af5f3aa409e8192b03dc8047dbe40d51d006ede77d3c13962bc54e5dd444a68b76ca8843dd9c3f585bd03e7dae07e09e5e38df3e4e5369b901b24fecb0b00bff2a4c3740d3d7449d309360797781cf85;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h420ab81369d1cefc29558d2ddb8f81f333ace39541361635f961189fcc6fcc849533cef8c5d0a759f5fc37ed9eb00c0e46ed4f797ae9d0864409cd5a8213ce659bb772ae044f6b9ebbdd7b090b83f3eac3604649f816511a3cc89d55cd25a6d4a986;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb37b35ba81e8a4b7dfccd740de78ea42b1cf5e0b4acad25e2d677779d0f7013ef1cc34af24902e0554a6080ede3d06c7fc4fba9324419df7be0b972a085ecd2d5a64d7926a4bacf5aacfd514faeaccf84a4064afe307e2783a353a47d123e23f1893;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h968a2f56b441ad33aa0fff40e858a22bbca6badfa212275dc3defe416054db135fe1cce219dd9a91417b877a80a8b2d6c0b9bd3dff58ba4dd71fc24ed99926089112f16451a268e6adaa45bfa0dd863162fe9fbcee8289efb319e37bce29d7ad0e6f;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'haffb8b5728aa1d9b5ac19a784c0d0760c56db6f822fa5b79fbe052223a964d2ab1e79820cb685f9fc0098d6db53097c4499dac79de1757739baca0e8f0092d22a9e5def580248ffb8c9de01ac90d0c86d57d915d0955dc204d8767ddb6cd24af15db;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he2cec669af205fb0194e978cf55296e7e0a477a0cb67212eae2d2e9ff47fa698de8c76c167f3d53929b9a5e8aa9830eb876b7577ebae361189bd6f93436a069e0577fce49bb5c71615beb109659b98654cdee2f23245f025396c5cff9d0bf69c0edb;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha9c3d8a4bfc88cb072daf84b819dcb113a0cdd955bcf9facdb5df04e5ef09af99f6d11ed8d8efd56ea32080319953959601811e5de70ed61b375fe46e7baf23aca565402b695c04059c9b9cc60e41d2339acfa79350241a64fbafb357d7b140ce7c7;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3e8af259190b22012e3a044b3f7ccf1c51e814310b32ad7e9fb0256475774ff507627ae6dc311ce599097545fed0d096c7b074b287f665779363c26c5ca2b2a1b7d0421374bf0827b5a38c720aaf885bd0e47213e9e8cdfc594999644b3eaf5b5e61;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb9973ec24720c25eafd9546efbd18d158c07d34903460be4df94a1308a713a9eda61118bcf38f7ad3f09d757aaa249aaa95edde0e8a1dd7bc01829cd25e768df841efc6a0366de44d3b1aa047ba77c700a75fa32b097fb259ac6edf3659ea615f474;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h184ec456eb41270e7d26e2f10610f845eaf1e9cb912db1e3c004e5f39c8ec0e99da5f0ca88749f3e5f5a7969d5d10a2ffa307c5229d98eb890c0365a2a9b60a467724eb8c339125bce3de8ecbea3d115bb5b12cdaabc12af881b4c141e2f88512514;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'haa044c3a4c180ff4eb95468ec16737bce1f041758b512b8b83f03c4fdce547a5afd60779231dbddddf8508cdc192375858dec06e2ed67f0b79c678188dcb3f21aee20b2b8e1b4430ee1541a3daeeed4c2cc569fac8cf7252a832d808948acdfb02b9;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8223ffb41af7349817ca24761abe01e8a86acd421f596c6189881f5b2afab4c6244ae3e3563a77cb0e5b4838cbe5a19462681da02a82ede5b5d5de42b5a4f96878b0ea9cfdcc690893052ecccd26248ccd53eca88434df641f7958aca802f63c1e1d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfbc2ef56792d387b49107cae1ee489380a43e5dcb3865223702e84d2a63518678464b5ec4b17059fbb0073b5893c42ebcd27464e534e206a72e0b9dedc5703a30d56a2c65901d456270f3e0053fba9a694aa8a14565fb37707ab8268bc32b95258ce;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4ae95787c0bacf2d6c1c32da6f3ebad7a800b12661ee62cfb67f9a99b28c9f2602e6ac040f46af828063710f7d60dee6fab95ea288643a50badabd07d1beba30421e63ffa4dcc54b9bb68bf29d55c5642157aa1e8aec71ad17f224331ae4f466ed53;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h74aa674cc9086aae39d8bcf52a096fa8138451d0be9f7a1af55045f5f23d3d6e26f173a3fa1b46f21dbcd4d5405ea7142c5015b62e85ab2456a585a9a6f80c448f4671ab308c7e9092a08ddd67889888eecd4299cdcd900ffa60a9e7890cb831aef9;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha6662f6216d98c76b5f4ab829f5fd390e2c071af150e7961812d5163abfffca3c9aaeaacdd1af37b932b1280baf6ef86797357816ac1b51223fe8c9aacee608a4a79040825ccd2f7e39815f96072eaedadab5a0448e296e98d71ba7d4c0b0dce6c92;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5dcda3427116cb4cd49d0e8943f79d7e92881bed08e1903792880976a77d66434d741f5b3c7cc3e4181d5036c46593e190ca9bc8dfba801e49929a8002c6f5f16bb1f276e24506951bcc02501d5f8a92b312f6b59f40b7e01116110fcfca356eaf1a;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4751104bb72ffb74da5b23c2416dd1f0991b22bcace956967b192708a2d90e9bd3f51299b14ce2e56a4ffb7d9c2a1e6e2ad03323c6ea9a3bfd101ebc8da6c9edb88b4880544aade69c64cbe3783acf5c83e1ff3953ee8df7cd6ac4296e07252c0868;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1a81d6b1adeaf1dcffd5980283df2601f262ccc3fd3259291af5d06e3c8b323ffc9dfc23b207318778bf9ed8bb2c6b8ee85f8a5969b0c32d620cbd6975fced5f06002f58a1b66136cdeac0c30c7551caa2ca17141a930c036954807c0e58bbda4703;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1d7903ae080bb15ea5ea7ef30ab43576916986360def347ec5c89f5450026a9e2f0bfbd5df1a8c95f378ecac3b10edc3b280fe84b1773f14d0eabb680ea42e7aa80111b9de6cdff5effb3207379e698240f7f3447ba563097774641a1f6f58572cf1;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h250aca86ee530a9246c80028bda136747085dc4ba1812281f2501fb765a96e02401413eabe3e8f359033bf585f81d68e8a548dbcbb0e39fa2aaf30ebdee59d48f8402cc73e249d0669bfb2cae9b499434ae570601b16f0fdb3c80d47d900206ebb52;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h30307e45887c98fc9fe6bf595b71e178cf8674a7af87d85bf62f0e503c761e291b1ea939c1d82759596a39a9ae72d45573b832a0bdba62a1de54f4ce6b8d8ab75472bf187829e5500592065b61f45c3b457b63069d006e7e548f65ed22f39b036899;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc08b2b13107323c4cc4f3f7fc327ff61fb0d6b8142345d487a746c8e482c85d9be9e3d7ef78de8d32f57482aaf3ffb9d6450af1a1cc7c21d51148de46ef48597b9839d094b1ee2ab47ff23b14891efceae1187fa13bc1b6bd567c4669a4148b1e4c1;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1def7567ce9424284a13e6bb5ae1e276dd61c2df5233e31d82a46f24c4f9317171f680a8aceeded8994b3ad01b252e8cdb1f8eedb338f4a702b9b936bb0956fbe661b65eb40d302b3715f1edca7fd2343e2ac45e7db512108fa7505d6d9a623dd2b5;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hedee9f497225f99fc0ea4c28cf6646a05c2624dcc133efb939cdec1cfbcb3aa3b760e95036d81655bbd161304c84a5841ebc54523a183bbba1ca4b978be0cdd3845eab5712d10e40f8cb9a30272790082780304b3553d0566270a3d14d80ba498bec;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'had71a0ff2de0bcbe18d6e79e48a7dde157f3843fa5b4b08e8ffe6bb21b65bf3b0e50fd3a37afc32b30a9f51a22888c87b51f76803bdf2d7c89c5c2c484f7002267ad45ce3590e53a17e375900553d6354415e566d3ddea013d3e795e67e125bbc980;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbb6a053fa5b1a64bb4df93a05e87b001d0a19210c70b334469753f710d3efab103b99f8af84ff0e918fee400e57e9dc6ec834fb1d2eeebbb9d37e9138e33548bf63b331cae8bcc5e727504fd8877fcfe65ea1cfeb215912d6097ebe42d49cda64236;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6e397c51dfe84204c1a1b02844b9d0658201cd5606ed0f74a6944b204f6d028add79fc17459cc39f3474ca69849f60b3b2232b21a0e5ea00cef6c73dddf7f3a57744d32cea4463c250cbaf429bd8382e5088f6f0a47f89a7db3db3709db38922a160;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2dd22aeb6deb71a9f331e88630dc28d1496493567490b601527d3bc5d4efb25e0ce9947746ba7c710d02185243005e1625860edf7fa08c17ea67594b2861e9159d53a20adcb770a0d0ff1f1fde9469a37a34cc2a8caac9c2585ce11eef7d7149b95;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4cdc8cd9f9fb5b50bdd460c74f307d1a8df21110736044b85ef2338be0a005203fbb236bbb5ca91405639e01bc4842b0950a92992d865ff58adeb70f294e11be4b4416d2c75ddd7403b6567b827f3a7da2413c9d30db9a205eb555d1253123820cdc;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he2bbf56434b7be913508a63752146c09de6b53521f743189c875891f63f7a25037b8188badca2676fb9a345ceea1cc75106eccfcf1011238ac6a16a72f93615d473810f94d66f2312a51dfe4aa9e3e3e177cea24411968f090897db70b90ea58b1de;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'haba07fc427df28dcf7e85c713f366a48452814ccfaf088e09e0f9d1042332683f157d08372318d7708def198af7ff12472f54214ba947f90f1a284b44f510a2840fad24db303e2fafe955d993498932343cf4142da738ed0649d9402db303a97add8;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbfc0b4da2023009dcc6878a5dff3ef937fd830ea04155a3132b14b700345852b02359a7f3b83e2d75235e466a1e422dee0dab1b09afc58e3fb65cedca82cd8d0aeb67995bab496e52f8db7d2adbb42d220d80c959efe53403a52703bbcea0adb871c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1e84945b47084cc75050d13ffa4d784e36becb6af1ff53a4e5c47797c2bf783fa8650e095c9d5b8b26a0e3ff31fe82db8a44b1e061adfd2c920c7850723672e29fb0444d023e1bef48c0ad05cdbfc69f7a4d71a8d2b374975a9c0cb1c3649857378f;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2598047551960e085669ea79a8b2156729ebe313489d6335efc42e4dddc07a83d0d20eab6662eb6177781d5bda25d2fb90c60367f564e3f4ea9aeaeca0e3a01715e6eaa302f4b5143324872c16ecb81291625b5ac7adff71457b05f7628f84825fc1;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hddd2656870848023aaf0e65a89df2f546bf5ba8cd999e9204e4b16d2d85d3c6c4d063d5b37c03e5a8079759c43d6f7b9505518739fa2b1e9a7f9a2b8e40574dfcbecf45ac9b85ea5991f78c5f55601dd56259e0d842e643ffa2cf030a3dc8f878185;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9158633dff274c88e71dca4adb999999da5842a72c0ee0672c2598c48665289977a70c0aede165b3feef190a743281b983eaf0db6cab313d469861b125a11278f3aff287d087a1c209cc8124b5df1252bcabe5a37832b406ef928f47e385ce30058f;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb275c0cffefde590705c2847144a839ef15ade6a051036b6b182461e3844680108a6d9c38daad3d77163b8c20fa00d07288f855db7370a40755f1fe6e882fc9a16a66f32d26762e16a8d27fa7ce9fb2fa4e6fa27738c3e2de4d904ad08b98e4ef13b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfd72c59ffa10149bfefbd21d46b83f33d11d3ce3840df904ecba2e7f12d118e1b0d99e756e92f2607e8c9a423143417926595a8fbc7e4f38d07c56bdc8ba9443b1bb799dbbada3f1ac3832c17699480af0d621a6157593845250160a8d4d66a7cac5;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc0ba6954bfb836d750f964f3122039aa6fe941390667acebd8340dc249747029c10b453c7c16d8d88d7de51718b831b70cb417aa74a519492e93e683d4d7bfb2d24271e3741938c81735746312c8747229c3cf12eaede979ae9c7db5ea495362550d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6772e3e53f5dad2fc99aa29e337f0d63c336ce10675f9a7f7f3a1672a1d7bb2378c36208458c24c96cdb3724f48b22ed86544a5cfc9b0f6aaf4c2a3e9ed4fb4325923fb743e0afebda62aa2932d76a0db50facc02ccef0bbb02cf3d57f78d41714c1;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h820329418a2fba874f86dd6b6dcc25a43fbf9c0b78d6ba7fd5a72a54bfd2a4782d4cc614cf7c7f25baf607687a4cbd62f2b53028ad91bd54be9a9eb447ee9adfaba852e17f69963027295ef959fa940e0c88f69e0c4c847f41a05b9967e24770e610;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h33e6fd29e0a1073074dcf6daa516b5792a077cdf8f2ef7ac133074141843daf7f6befac93a2c964d685481a974108a6515573286e7b5419ea00f0d1b776f78bae4111c8ef479e76d8ffff19467bc1e3e4a4b966e32713c715ccfcea5f241ade4e997;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc51e4cc3719c13b699db8c51573a28732e95bcc84abbe83167ccd2de1f15d001ca40d12a653b14e3e624a2badd14f1b4571698bb74e2d78a8e073924ef2b31a988773099593a1aab5de3eec248e817ae0d00a0a950f56b2e9a458772b8edb642e6c9;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfcbd960584d6f123763206b108ee8f94a3fef6fe52d48d3e4ff624472233f0c37dce79e45a27b1b968d96fc82ec5043f2725a2932b21037451cba0cab852369d30daa58acf4ac23ef3a167b1924bb806b0fa2e14590c716c0deb54b5489f1f07f78c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h88fc6e77e3c11262a2c9b8cb092f51878361766ca8cdd7d4b14767f78d067247ff953c90b486230617fd4507d520a4118bcafe81285e85270297840699e272c5dd6e8e28a9ea202faf1ef215d6488eb88329238b38464589c4c09980bbb6bf983fa4;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8c581e4c60f2ec88dd7ebd157402356a7edcf9a9e104dd7f5697d011b830279009484d8c0fcfe9c5f0b90280f31ee53e687c1173ca9e38d7c6e9cb68758498155cbc98850a7f8cf8f9379a43f38908bc13df72c55bfa2d6eacf77b2a32105fda3e09;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hab2b6580e2fe170a2b9fdd8aeb9f6b8436258b7726beb01bd301de2f036d72284fc9a72e03f5152f416ac88431038f340b12afdafd3b6a9e10c2f90c6be6574ee6ca384faa3ef88e09913af4dd204a322779798ab669f20019429d6f322c0147a99a;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h30b15a05626cecdefa779fff5003f36d7915b2bf55214d97b073e3ba1f728517ce0f89e49d3a2306f21c72fff97aaa6024edc0efb934a22298140396123ea698b83bcc9a30ed7cdf9a997cf28bf24f67fc1af993db6167467ea5d800558ac116c05e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8479bfddd4cc1aea43ed88ad3688f31f2c1421d59d152e4249ebe34ac67452d034453177f1f23b08fc0aaa8281776edc55e0189498f953a3681def9646aa7e5545a0d7be8a7d9ffaeb611c0fd8f07cd150eb6e16ca44906c456849c352556a97c733;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he024e6faa7329b5ff5950ccf2ac6458da1ef4b15a69892bf237ea8ed4e4f7f59fc703b930144d66afc8991f42035860bd4e1181edcd9bb2129071304d4f71d179dfb321141095011d7152325f0f3ffa91b0c6d396a780aafbbd47379a2185b1fa283;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8e390643fc0162b8c29bbb015038791f3f0de05561d8d35a84df854feb770421adc4613c7bd4f16308c3689dd7068516d685e7eae6ca1bd5e7f699e962f880d68a415078083ea4037b30828a511675531fd8e99d8893d19c64a3cb1ee397bc6aa14e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha1f88e4d976abdcea1f153170e0119c458f2e35c0fd01edd05aaf8dd9c2c99ebf963828a2949e0697ec4f676915293835b06a18b7a1c713e84027ea9541aa926490120144e389e778d4784f65ae6c792b3922e96d69919f2d25d55c857840ff20371;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h516b3959f7dc59b10fa97dfd1264b807119d689ea5177a481002e02eb83749de9502407666ed1c3b5f20c87abcccd611b832b0ccdb1c06b0e15ad5e19f8de0b52ca2817e7466c9af6a685e17b16849858070263609b5f0887097f3eaa0dfaddbe776;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h62ecb5224531bcc627b27e92c95048f8dfabefaf78bd11d235d5a4e9e0197ea679e7de82bd1f2d70e1f0ff3d078078672867447196167aeb386ad5c843c2422532226bad119f1727d7aa05a2b8cbb180fcd74b86d3f419cf377ee5758ecf84fcbb38;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5037a9ea3724e347a277e3295268e64fc1e4e8139efe8d7cb0f86288611f5379b083d28e14e90f3d786c8f86bbd31da8f889152218c09f6829487292cd071f9f40d6658b6a2388b3119d2cd5233a190f0736d861ae7f5a547837c047a97c804535df;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdb0c47ab2e99eb0d529c991b60ce81a89ed7e1c47d42260ad1a80fa1223d85c74f95acac68ac8eaf17ff2d0bd1dd94f20c079ce275d51b67e0710eb7b9101e3ec9ca4bdc7cd7cd2cab97ae8c1413a2399827ad38bdfe9b4eed670b0723b223d285b0;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc9dbaccd291a4c1891a9e2aa30bf84195889e7c40c97b036c1d90cfe4a94bc549d9fb4c16a6604707b98bf9ee90f3a6cf21f6f444ab930da69d0a3c0f58f6156f61684287673095b2c4cc8713cc1353f08002b467b5d88e1a19cd7a6b3e3cc97ee3c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h48158137dc60c6ac209cff71e95bbcaae0d7016ee9f4f91e485d6b99a51671e71e79d273700fe15582788a448592651e7925ba2bdf1e95d3752b3924b3c09421f4403a2afc5d180b50a33290db062f1c8348e5e9a3287dfeab459226e66f5bc18fb9;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1c03ed070d8a90e8a8d811d0da5dc1585523192d529e96807139f04eef9a8adf0ab0f1d6934ef986244c8691468bfda530f3f9157acc94e073de1eb662a6108e9fdfeca8d1097a32fc9c5a3743c81ecfb011d34e474a12e755b7ef157ed7f44b5ca2;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1f49dffb652f9286b035858129c676ab4a254428044a18f2383166baf06fb56f0713688d3c3f8209eae37584bd3de99c1c9a415aa7f03fe1bc43804929ceaa54fcd133dc16324c23a7eafe14a876a50e80430df83a2043012b7679973a018377e381;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1530fed7ce0e5b79101885756c38d4c8f1c53a8699700357071e023228f998831c6b5731c7fa18d00ccd29b0e952abd4d727ead2e74415d998455d1d43319272b1e1bc78224f78b98663ba2cd36b3d3cfc8f1fc63c0984b62e05a12a9504464a8c3;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h34cc81978d6da0a3c616296d89ad668ca7a2a6ea863b08b5d08ef54df90610471c3b91ac19f00a153edc8bc8dd696aff60cfcad22a57c1c546e8b48deabd3730408a4964a842ab6b1181f01cd98474331eb0724545c589a415a52de2ca0ffd20cae;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1cd9ad5ef70ab03595fccc4ae0c037f6a880bbee92fed77065f8ba1f8c8b54efbe9a5f3e8ea6beaf343a23e05dc033fb2d93ceb435507c5d039a138291fde3f9beba8209a21a85277ba664d6667cd5392788f1bd87a79d9c027fd786e1ae8ee4fe56;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h226df4909dbd98abfaa11fb049c5d368183f1e601b101f3e1746b9bec55ead00322bcdbdecff93f83025925623e53fcdd0833b4ae3d457840ad67f5335faf951f525dea6a6d05713e39dca43e6235335a43a844fcc9004b4979859d93e47b6b7d870;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h15b737c92bcd9fde358197d394791621c62a18645e3eff9479e675e588e31fdaf07decae711f02638dba3f9d9b155145c9d7b5b096b2bf59d971ad8efc7d1f92c137c773325ce348794dfdbcb1edaee04860a15b796c54f67adcdec2276543bc2da4;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9dde114135b5bba5c73914431e28e5df6f72422e955119b0dc81b547ced68ad24c6fc59f147bd88e5cb4950a69761de8387acd5e5fba53dc60c483f80f257682da50b03f1c377da406846bc474b149f867d6bec6ef0dff7fdebcd068f4bd5ad94215;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'had92367685d20eebffd53d9cb462b0b7316ee94e512bdf762c352a196d9a9cee401a2149b02a1eec67fd79ea096e29678590a632d5d9779e6a6de0e73c07462d5c37cda827b09422dfeb193699b910fb51bbb5667601d02a8b0dd94ca1a1b429f299;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6c133747185b9e03e45695606f6d1c165e8198e37a1625a6fca52723a8a48a5e94169f38eddcaaa8ac3c7b04771fa495271c5e201ab7af9bf3dccf9d5eb99eefda9d21cd229e2ee6980a8d625cde0db2be209ab285a40c8e17d8a210127e11383381;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdbcb28b648307e7b0ffbc1ddae606d3a90462afd6c0699e75c74d5b4350c3a01d5a15e077f7bffcf21aa5ad138be4d234ed55ebca5b70f681880094736afa716b333e5e7248c0ab8134b7f18fb9571a583795368dbefa0f66ede612df5f7a020bf83;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h98660231b657369c0b4727880e8f60fc6a2347a5f381ad6b82f33ab2180a4039c4a37a95f49af2080f2ff6c00205190ddad8a79d49afa99e7f45985b59e950d60dd045cc1afb55975dfc871da7b7d9eb234d903c5295dc1925aaa07b8b879eea4bf;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb374d0e32675026b2085a306a471497f03e67afc17b43621eb8925666046d8035314d9d304fbf42058f3af379b0b528bb61be5b268f0ead778b8484f641c34751aef1c50102d80de962fc6e5ca014a47ab888885cb231f7a5484fe85288db56be059;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h98619c3192ae39eb2ff39f205cc1e4d70e131c2b7f90c2f7a25aa849686a8c723a78b64fea60d1ddf8fe767f92fc45819fa090638b2a60ad0924583f708dacb545c20db24a58cc8c226f00967667fd35519064f614486d3eb71561155bc56e3bcdc2;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf45a35d6ad64aa49cc8d0b936f26442417859742950fc82404108301c514fc6c8a55583f0db8191c848c768b277478d1dbe21bce4d3ca0568628ace6678f34af20c2e05894f8e5a8e12117b837d29f0a3d94b6da2f1d04f1149e93c0636b90abca53;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'haea6f3162c21c6448173852e0cdb96cbf66b20e20eda412d4df04bf4118ceabd9d3c052245b3fa8e84b1e0b5d44c848759e432c8385440aabc53efb68711a8ac0998eaedbaf75d3f7c30d7a250239ef771944aa8befc9e6229b8f4efec0f0fea2a65;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h15319b29ebeb11ed93141120b0df18797a79d2acbc1f33dddb6d991f6b4979fe56164b3a12e10cebabf55a015dce1afb99d638d37e1e3cb4adefde9ff17e04ab355bc84d23050583966e47632ad4d0eff291371675626eefb911f429230703c51b87;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3671e382da35982968381bb85be98039fdc378b47866709476032a46c313eb1f57380d46aa4f6859ccda216ad20e52d09d5d4277ec6307a5a5a36a0e3ab94d4bc711238f6fcce55eccff77f5154a5fc05e8fb3e708058bbc2a577836ea47757c5828;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7c29ec82a38107cfd0720ab8577395214d5bc2a966c3cc78a2ca630d86534ef0f625dd20d5fda2731c1d1bb7099814736035cb299d7ae479e84a27ac60fbfc8c080e8077d1f01d35e64891232a258727a10bfa63543e0062daae52543a7e882a5ff7;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7e235aab1a7ba38f24d23a4ad0506863964adba377e635f19af0ab0a6e86b7135f0b7535a643fef3d27544bc7e9323fb95fc0407c1c3465c942b5b29ecb28e476210d403a28bc3f2353637f7dc586d9315a703eca29ef99087722481d1f07af8ef19;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd777084e1191a0092decc55c957377f8ab0f7bae3aa34b0a2dce7f6be74963483b66af6e7447af46cdaad584a9207a795561cf63813d835152bd17448609810aeed032227d99b250fc7366418f2779978b38e23058374b7fae72c3de9152c6660c4a;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hee6444793270b3c489a515f2c741beede1b978ea907fc3af4a302bf5798b85ca899240adb88735c83e2ca5b9d6d2d5d2626585a78296e844f8c7b4bcb908f70a65b223042dabcba4fd525e5b4c6dd0700adbd15af330b7ffb164c9081601f030a25e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8b366c0d60f7055a6508b5f173efe54ebe2a9164c131d16bc200c6da145a07a99ec24e4e6a0a6cc4ff11f0f1b40299bd6bc200880f4d1bf7d32be289de16c28120b84260487970dee4be22fe3047ae9efc7cbaf991fc234f2d273893801ec75316eb;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6720f0e9df204e50f084da1d1ac167799edab22ec7b43ef54008523736dbd70f6298984434b8120918f8750ec77dd092907d15e0e6d0f3280ce4564ecf8dcec43a316a38a930c5b05f68491df6d2b8efa0086e01c07af4d871400e5719ce43add683;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he643e9b269893ee6bafca92c993892a3b1038b322e68a1021132b9e12492a5f221fe3fc8f06cb351b05f89b6799e558318f6ce556d4cd91b20586850884c514a3553946bbdd01b3097e8430a660130e4b468375d7109ca5da472c0160367c28cd532;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h32c695ca7efaee60c1f7285df08b309c5f22f0b904a1525acf0739fa80c11135f6050077fc28976d71ddcfc0233385676becd8f0f1c074f3f1466fb6f132fded4b61393da6215bb8352ac7278342382daa592d21869cd377b4d1662d70bb4b1a366e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd7cbc9e2c83cd3278c0e68417d5e05196cff34f24b2f5a7833c6ad2a78c99ca1a274babc822ecf1ebe6dea4f6928603516f741df1e7bfcaa9af334d6153686f54019328e33ee4ccd590524ea440670f1414a6d500a7fc06dd03c787e838c20a07d0d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbd8a4f5b3c217bbf2ebd96810efeda7f1dbef2a24b4c38ec913e06b4d74d8e7ee5e28afce981d0a36309a66ab04c6a882d0f7f9ffec20dbe0949bad2a5a9992ec9047af2e9d4ead8fbe07586fd3abfa20ffe7751dad1c12cffd92e1482bed038027;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9ef8105dd9849ebbbde85dc1d1aa653818a10b78749e99cdfeb8f49cc7ebfbfdfe0bc20a1f7e8ce2934698b725b8e3aa2c07931457e4e939f3705033e5a331e29f97538a351005f053cda52ca868941144b1149f701bf31de451b2348915569810d5;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3240d5acda4525ea11f7eb043c3f7c52bbe1734b4f6c0a824c3123d5df8547093e363fc82971f645ce569da8aab9d4ae06e814f2afd041f778c2da23596c94a00027055b6e8b01c3de943194b191986fc19cebbe8273fec03c6550256608c9913253;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5738dbfbd350072147c5647e353bcc560b4b1068e8fc3d367fd1e060b08c1a80bca953096bacc0a3504d51d7e3ced5203bb2d8d96525f730cf3a299862820e1bb869ecf69b867ec90360fb2d6f1bad80925978c8a9d55a8ecf2940258296432a631e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb8868842aead1d3116c18cab4d3a5a28b22f5af64228cc61835eb0ec44db4334894c9922eab7acd7051f384002d81f33e325242513eceaafa52be8020f2ffeafd3dc315ebcc029cb6200023be73bfc3ab1c56a831c4c86bc5e5ffb2abe7ab01a5bb6;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he22f723d859ed43921355d104c290a28f531e67e264281a542b4a3ed275157a8e4a422776a541dd5b0b6f89acd7ceb94065a4e0d995e8c980d4a0098b354e7a22735835adb70e875821a1a9a5db87e7e01ec6ba576474bf3697adf721342eaec8ad5;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfda3602725e7a2524be11b41af354fb2c95c8e2ffd076becda03c04b1cbf059b4fc19b555ddaba487856cfd38427b7157b9d9364569236c2d98e714be4c058771f9cfe38ec8d1f3af039e3179f7aabf3a2577aee4802940e481170a666138cf4fd20;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha977b0179aa724435fcf19e98b4e0daafd10d2017043428a5de4e9fbc23bba1ddddbb59171dc4c78203efff6046a43d436945959a0ce3636edb2775fad06f23d5640137e71e5647f8a4c6e436cfdb2ee0eb0a844e9063ad4c743e547122368b4974c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2f94fcfb9c80a517d6acfbf34fe8b4c2ed7c5cedb0f8542306a38665eab917c4da334901b6d3d1e38227bfb8b889f0e3d574a32195ec790e84dbf57f93c34ae99602fb5a9272ba13eba9e144e4e5b5fb0629b1eeb9e3ff9d3178fd02213882987d8c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7b5af7a26b10fe79ece170ae7caa1c79f19badd6d8ce5b6348bf512fb089001fb46fab5dc9bf7bcf8282cba2db8950de0b3bc95ab47576847665791244e618f9841adb368951e7cc36081c06f6e9e1dbe62d817cc74d11021a32cc34fad9f3d86a6;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hede7b6a016da22a114a88ef765bce62068cef5f51cd7164bd6be81fd13bea0f3577011e1f934adb79411a76f5d8302b2aa58225c3ded4a7bb305eb4df72e61bd0525ed8c293ae1cedb1c1d8c4924357cd5e649fdb1c0118e1cd7e4b43bbc8bf37874;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha5a829df76b05992aeda65a22942ed60f6e2a16d75f0b578cbd486b189f523f2d12bd62bbbbf1ec5de734bccf36d0db92b9141d699f65291af3d4d167b89ca427d500b0ec9a1591e05039db1b6b7931a176d2525532a30f1b9c17d80b48a738e0bf3;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf91c4474cb390a189426c5d8460addc86b521e6307eba5d13f6fecc418d4d0a2828f96c384a96ee4f24ff0a26f95974ffb72dfc39ae2ccd1b2b1fe45a3f5cd2bffff042382edf4b54e000c6981f05ef4f2688f3afebd3e68a2b939b8c5a301dc51db;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hcc713bf0b18955802b6a7dd0b9da7ae626f493fb3d94bad27e9b59c3451edd1039a9a7f30829bd3bece1b2c90c3201222a2cc64d9274e5ed21b1a126da80e1f3d9850522785fb8d0c2a9e19934b862cd259514d13fd9cdb38c48e992d0d340a09ca4;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h85daaf7a7d71853febfe3f5007f51b2943e297f0e10b45322f128250049c153a0d6015d80de8921d4d893c20458e32f2c372b6d2812612d9371d40fcc3d2018e3f3b7dc6cc9b6793357eaec197efdf30dff457fb8677d881d5b940d63d0ec78c70ea;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hcc8f7f925c27d73b6e2bac7d0895f425f35c763c287cd94624ff0a0afa7e1e040b2f3c2f90c1d5969edcd730d208b71b5e5a553771a9a24a1da6b7491a1907c5100036b2f198c2a45bf8bd06cbb62d66fb7754907a0811c218e1d8041216600b38c5;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2e14381ae67de03a151aa2af1e7be9d3711135cea054bed559195f624072445d1aa570a3d6fbafc5405258e52597c4f3dce379312fae3250bf1c0c07abf338a12dd0712a0b29ae781274b7a48791a39932cad110b2e047355216c387968a93238d57;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'haef78a66a907d02e2bffe860329db9055f1f12a2006c2357496741885ca81f17da9195383570503db39133c3b039ea72cacddb116e8504cdcb48f99c5d35e40a63d5a0ef3cc14c8d92f7dad87ac5a40cb3234d61754141cbcaab917fe48aa44a5a55;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h59f4e3d66f7a5c7ffec221e79ba29a636528155a22e5aa278c0361b140132fd7d1f5f63f13553dbedd6d003a47388561a0dcfdf6b9285a2df7b646687100b57efeb807e6352cf5380771819a35118b451be93c6b46ce0c9b09541a39c71ed4b310b4;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1f4ef2d187c9446f64247800b0db47babb28327722385c02be74483f028710f257c588ee1a844866322a17f5e69ad16f774232a8bf4af1a3aade21914b125b91646da34f91f872799f591bedcac098e43183d9f275394f8558d10460fd95e7d41c6e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdd5a0193d4954ed5297af4552a7f5fd5f5e9f63355af19ccb94083b68ece27025e665adf39d2092e4359d7806fb559a6cd65fffd866e68e79d446757b62726f73ced2dbdddd8970faab30a595a4710dae8f46db2ad268d609e93d8ea0eac2b7b1a2e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3f87e88d8a3fe48ad2439546ad419c39f05bdea87f4017be00fb51fbdcb1b842afd78554860f6d4fa3fcd154585a5592bd711fcb72279f52a8c587cf11279ee15142e6ba29bfa95191c5ff819e4c4d9d41b769ad47d6a6de5d3a1da310450b84db88;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h107f8ac7cdbc74bd7a75791954b712e66d98efaf0de4c19f38d5a18df59b3350d4f904a47e1fda0395996d57c931336d91d49c9f452904395ab75af172806c8df3a503bf04ac7e50565b76432c6fdef43b947389919bb0b1cec3d89a8a522d36d5b1;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbbfab224ea2b459b3204afdd077f018086c0782bbb72c9ae10b684699eb33a31c29da5c4699810cf2df43ac83875858c1259a0470359a3c5f6e64b281326c7ac8698136debf619a8ae1a00aec338245b962533d2da6f6e388e8573f5bec3a9657c84;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf294b7aa2459cccc8d176073a7286d20220d23de392184ce4a60e86637b175867a2877e3b6baa153589f2fcf8aa01798aab95cb4233a45c4a4a5889a95b7b1c293bddb71728fd043f825ab8e662b0fe9c5ba2023218346b565916c5e755b357fffde;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5a2270d81281a3be037c0faf00453a366c34736c40001f28fb338cc282e5fe5202439883911736a695c116880b935e90987eb65b4282fc6edea196261664a6afbdb3e8ffd74005158f4329fb4d663cd06195158b88035012b148182b37924178e639;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf48ecae1346ec5d80b94780b2caa809cea5859a19ae41e6d18599cace2a72c9d103956f732d5586a426f2262f6091d101f58a0bd8981e356d143cb4f15ee6c505e8daa73e8d35a813e6f9f3016bd966d672d91bfa6a7c75030ee8c3908c503291aea;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4d698e1f4b80a84a257826c9c5ff9e824dbe5e42368ebe9e74483503fd4c7f8ae50b9a533cef738da8a0696c6aeb384df22e344d9ea34350df5c7189a4cac02d1f1681e0cb80f22fb8e28ebda8b075a81a93d037f3abf1b05d862705deedb50992ad;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf8592c97dd4e261ec6c98c89cef7848f55ec78c6c9bacbc54c1b75775bffb7a5cea8a261204876135206d091980d0cf29c99b6ad72ffbd9688edb2dff4bacafcd5904427123ce2ee1141886a6dc857f29daa4100e9bfe7af248b0ba18aa0214cf0da;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2c01fa4abb55ceccb6d3f786b02aa040453a0d5f2e281abbdb98df4c48c6aa574f465e12317d0035f8ee89445219d3f52cb786964704924f504cd5a7265c2765691dc8b7daeb5c240b45b213459b7b9eb6873c9b73302538026a1cf0fe29766877e5;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb37048ccbdff7cabced8e8165854b07d12f2292ad9f584b3be142a6d4afe036a24a2265715f6c41d74fde51aa5b809ff8bef183ca7ee5ca180415482f0e842de948bf5c8e558f8b91aeb04fc3e904a5ff533176c83e68a1d3b9fb132d65baa5573f0;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb659c1c5f7b1324082b7d61671e40a34be81bcb7b461c58032ca20733d4c546ab92225f7f5231aca0918152c20c3f823b705a00117e239f1747d8ea29342c0d0cf93031bb035ed114400f4e175afef570a83d85947cedb71a300198544b1df67cdaa;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb82be7b0560d71ea05e47d31b5af3b297e94b0378ba4211a14d6f85815f078a9605299a9578a97673d19113850e1492d97f8a4e102bf03506d0339077bb6cdd3038c0019392e20b07d6c02086b780ba4e9548631a83ce4485cddc8c25a37b737bb3d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc82d710ff7725b35cdbc6eaf3509e41f0ff1f3725c4ca29e72fa6a7023594d6f334d7bdccf1ef6719b4e655d78b4ce335debb768d79e8b96ee3e0cf3ec0a9279fc916ab8ef914790b90062bb45f66c1d91956f1b450fa6d9d0a21829cc892a80459c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hcdceba20ab319e9093c19ec38628840a335333f4bb7ff6847f78bb758f941d0878ab64a92dfc055dffc48b27059360e14511641b117d84d06fd9d04599edd4655faba8e157f4022e2bcb20be5919b7bc9dd74313c8c5f1568478a8b11bb1d93db76c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h26af538d4b15f5f4100fc462e293e63d46a494e50c2c175c7d8e732773538bdd72ecfd54fb7ae16a78865a3eee6331288fa1b86e0173ed4fe42b3c7cb7227a4adf6a6e48b5b191e13c4de7b072b037be88e71de401aedb15f14ffa8af2090f6817af;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he7933061f53993f94931eec1fbb4ee4dd26a9b80a015d69c8a47990fe03d5d5cb07401285e810e923178af77f9081e913505fda41fff1f3614e6017587fa3a99a837c3d03cc4ec027e545b4fc9812d27d8b929cd673bb04c775306df62bd20e70244;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha208e0558945b715bdb7b334dcbcdd54e79343412fcd64f1374cbd2415452e67b4f0bf62aa375982ca40cccf87f6af2b8a824ad1c30f021b11084b78c0fb5aa4fc643249c8e7278a267ff3c5b9e6589e848be6b6ac27a5150b1b935adc3d99d61e51;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5fac35023d6f2895ba9b4aab452227f44041b35f08d46ab3558ab402b7cc53577a7f0f2e89cadd32f3ce3409549659aea46c8b6640434e4c73f775950d10486eeb984f51a63fdde98e9fdc8edee6a53d92c6fd2489a6c784ea40e309939c61c3876a;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd30b05888138ef20ace52ae0d27b4b8af665ed5e6276890c07e2a46ebacba8fb8d4dece48c4d1b3f1fdd629b8016c5d32bf04b2f875a9682a0095385149575ac56faea1318445752f141acc13d409c2ac7f17bde4c511d90060a0e4ae50ad3c5738a;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h55f83672b570153e3f429e38e2acf1e0904ada1306b20d98059b44f04d11f10aee95f70d136200dd6762f091cde7469ccff9095f2069050347c05e87191090e3816182f296748d68a99c44d9d08ef1b88e44d484f20604f1a4520ebc9f5f59c95254;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h448a9779c9936f68a2f37b4506bc549163f53f44aaa2351b147c1e99d7d17ae828480349459354a7e5c04be9df1171b2ca6426e751f4101bf78a6671d008c7186b10f9754db0d112158477cf3b244129d67b0df3b076f9ab420761f547e0bb768e27;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hcb472c7e1e64b7f19d1190bad907811f74e9695803ac0a218b4ff894ab3965956140ba85801cb4f66ab64b968a120d894575888a89b317c7521e5aaf0a110370f73229fc0f9fba42e2212d9c6746f1ce6ce77d4c68394fc4cec21891f859c5b15b48;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4b8352e19c22b4691ceed255672f1aa2a749add785bbfd54a53a8e24ae50ae2285eff8e0766b9b15776a1704f3423ee40b6d1fd72cd920b270d09ca9f760d7a9cd225773431a49d13c8356d91926a1ee3adfc1bce43212977cce4ca9ea5bbca21ca1;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf6e552b5cd75da40857179e360d331700a143f842dc736a2a34fff7a990662929566ae2d9673f234da32c78bd8f6f3aa58b8b04cabaff8c71b3e2c300b14d88db8368dc1735995d1874ccc8c8afef08ef738ec7e1530079786f24155b84129fb1370;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he4cedba6dcef7a0353786f955cb7532388151b043d3efec880e4177f6ec5beba0cd6a96a71cfb2b0493c4d674d8349fcbe17e61e1260d05c77d7a80f6516c734ba2d2ce7ea64f61f59896d894f9eb3ac95e1d8c415a141a5f68ef0a6b0cd7292ca49;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7fd1465cbc6dfef395e5defa133cff69238458f64ca1f6f6139af16ed90001fa1749b944fdff21c641b99cbb98e04fd103bed4f75ab7e682b7aa48bcad0bacf7f0784d6f48239826357e2b6bb4da565ecf8cd9d64af1e0063ee8d3696473c8d935b1;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha8901d8ec2fa2ca8ef997360ea84a949e356786681584b78be1cbce23faf82e831bdcfa74da95ad4fb8bf7f210febbdc598fe2a2cb74225b316a0a098f5a2825fa29b300dcebb72b1e82f41c3fc3db7f59deed7a76e1da33ebd3dc375ef13b0f375c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h699cc51c4b0377462b0eab5011a28f204ad9436437643112ce0baebe6d18b0d0a7cddae079c34b4624afb66fa078a21f5a39a5e0a00278d7bb84287e77f10f99d7e52d54bd8aaf3f2191587e3c29d58910c4cca26b3eb5d77b287d45985417dc5654;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4998ae2af492a87fb3f839a252984b95ecc3fdd5ba3d53b6d1a1298f65d5609cb014d8fbe38b27eb838efb099cdf7bae26271eec6d68500294c1264258a7c883a936eb3635939e1b9cbf8ac4e8d92da0cd3172d5975c363ae3a6d7368c36c6dc5fe8;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb708d95cf086e11e4a407a215df59c1301959618379e4e33af09e73f45bdc264cee74cc528a6c3169ad8fb41d789f24361c9344d70c047b77cfac68a9dffb06731dada7c0c204b3b7f45525c0c9f4df2ffcabc39afc6ef0c5e293ad150897bc86fa;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hee6aca9231179ca550bcbda59497a51e165854d70c3c3bf7f08d89308bfc3cf4f1ecd59091d2364f29038d25410885abe38cd179093eac572bf3d34608dae1533d8863021b060746d2449ed0cb8d3344e6b474099af34fa3eb2f6061f5342eba3abe;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7a07b03c5c27be04a156371838a5cf263aa43382d336ccb4f8749bc8462647ce414fa4edd7051fd519603ca85e6f48acaa620f508bece9d9a20b94347cadaa4470a99e230dc37b67eb434400283f9caf5125d52cdcb4a168aaab0d5112ddcd3a4a89;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3356f6a8a0e02000445f05b47d0cf3872456bae0f99d37601e3c3556097f51c057e498518cfb9de1ffc22e0bf97c1602e2455af8e982468819f6a155eb7ce7669e7b951dd9b9ad5c3cc32beae24b149cdbcfec444e4c04340c228d6f95cd68fba634;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hec1c700b86145d9ffb5ae46cf595575850f0c637ccb16853f0ad1a9d232a5011f67171b42556e38a9aac906ed6a0d28bb953940bcc77354f622ddced3c414dca52a3e25b8250b33c182f09762d32a2fb5114534ab5cffe6d21d3a9b2ed724c93c72;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6e60751a879f3adc8dfa4ccc60235d24229964942333dfcccf89b052f2f6b6e041560bc4b2fa8496fce21a285c03ed1183b54ca58e9fd45c981fff4f078457f6153738b1b92031fe9d18138c28dc3a74fa834fbed69b9e15189b3c17f6de490e47a9;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h43b7b4650ccd16a16ff1e0ae9982e30ae2a877314be025b1276cbf368e5860d75539e605410810dfc3f780c65ae44ef2380824e0453d8e5f4c7415427cf3c80ef8aef7adf190a87140e14a4d7bb09ed51c1ffb844da186cfcf1b11be557cf99d81d0;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc73f8839a6275ca060fd47aa375457921d647f640a81b5236c3c676b6e22efd750a04f7790e97e7d524be4663f23b85a9844c81630004430ba2f20f4b268e84d352b77134f124f5ca37e39d98f15c0ff3b972d3e0521cd343e713591dc2e4d8a7fe8;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf8ce29f5caa227cbf1422a978c131724006757fea84eeed429ca5eac9d81ae86ebf8527e4ba7beeb94d4677e3021f86fede3a316e04f8526f3e6322c541f6285e91ba2f5c3c15a6dd01296d4477eb90854baa57181f82a7a378a2a87d3784c6732c8;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4b8b5cd307a86fc83817dbd551ef706c33b90a322cb7f45e241a3f9d3093c408f786b6e70d58205a937887cb949723e3c646fb4555d9e5c0313435e0b85055e254e56e98ad462f5173d06aad0492334ca05698071c4b1f4fea4cdabf1f913bba20b8;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6983402b01d0a7691d6e0fa8c0d5f6db63a0b2afc10092eee5ab2417660dd8d3087b0f38861ab7e97d2e13a1404fd5549f344bf91731229bc4c990688d6f8c0d639f179827f9047968b6622cc6f4e9ffc8e0c985ab773eefbd0c5e25586c18fe1c03;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'had464bbfafa3c152005b2280010eb6e3036ca356d859ddf857c7f55edff0ecfcc9719161f4fde7e114754392ad24e74865699c5d4752f8c2cdaf3d797c3386bec59f4c3eef24dede8a5af8f2fedd33598b2ab45713340f8b3be8a5bd2ec68c74895c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd7fb5de9fed1b7ab179930d3b8a6208c93ab2ffd8b2e245e6c25cb0d2481f67e7a60c20fc7b4c08bcbccaf14414a8ddb0bd4e53ecdbe5d9156680e60c834185ae75f9d5964ff1d7731055de89cfae8ea8481b4efbe4603a1a52e2685a4e897e6ee9e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h47a1d605a47d785819906b6659229934fe805de0582c7140e0d9078d581f1908e0a28e276783a0e195d806e0d126505f05a0dd5c3b92276d6f9aaf34212c4c34a411fb80118e13ba0ee68102cbea7e1b78540aefba1fc293ccc1f115a3aad189f9f6;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h65f5f12fd7ff77fa0eef584e5ed9beec63a31c9dd29a0c61ead95e6921e4b41fd3458b344c49dabf486c37830c664f0961c36fcfb03bb49d7e0ee26238db4fd5bf4722b1c9e3106dd99654f590664e49504780a7d590bced8ed7f9d85a059245ab25;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h77c9bafcc69263cc37d4fc6a3153a704dc4be629c955afd2fa60e93cad07b68b3389bdb248f7d978123cfe2a2d1c74903681f7576fbf6ad2d3e29336f94f6a57f758091e87fdc868e8a45094ad626c3892d82fed7166ff1717a178e8c54cfd933ac2;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf583184c6c04a2b4413769fbaabb1f8ce5330c46a26b7e7e2596f209d1de99ffcc7df2dd53523e912258ba3728e3d654fe9352aa53ad793e93620adf09024f3301a377d8d2a67ade8110bf2c195386de1a3ceadae6a0016871bac33fd992345156fa;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2ab7a3c49a3132b206bd53799e5b3bea8bf7b1080f22829df99948a3afddac7e0de684071d2709ddf176590e04e3d63986f4c2c5b2de7dfbae6f5c9b416aecc9e67e65624a6966bcfc3c3b3f7ee65f8be57d792172f7d44599242c6889ca96b80f4;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h52de789a0978b62a92fd7e2d8439a971a6049e8626b9a42201330374c42982e81a35a925c20ba7d5282ddb8096af17547056441c5d58fc9f6acf42dc6c3246d881289ccff0d364b96b365629881da02427280e2d99505a1a1a55e65208caf67d9c24;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hecfda658260eb1d5c5884609485a6f36c2eaed84a5ded12e71a8cfa690af342f1375c8f7b103788db69cb055ff18a29291e7d1d3cc7ad4cc8cf036bc6fbbc169fb534312e93d294a7962b7d642ca9febb7653b49517eb9950b17f49894ea55736d7d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4e9944d3d9f267b10141b2e13fe768c4d5b65e396a4676ba70d1733c041f83558261e340091a160e47bb5f0165b1d355dfbc7e2c4505e0657dfe0f26f8d3bbd3b60e7cff4a5f7330d454f55b3b57b189e9c0f13d1aaa1140dffb828e82ed155d5fc;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8cbc45f5d455d90078f7a64b67b86c4da2b4c69ce58d584915b4375ab34f6fdc1b28f4dcd281966ab689c132cd466831d11c1be0f1518be2fa03c3411f27e0dce32d959e7ec23432890dbdfa7094c4a0f5cd02e8dabf8be2dd861a273d4943fe6605;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb7fea9b9ae48547ee818fe81cd62a1e907b38a5f460bfdbb58647ddb2be93fb1e21e1269d31b1bd6e22b252f4f650d6a82d30b97bce77ccfcece67388e3409934bc55c61ab9e50db365e20b559e3087625ff499a1895ef05ea3f4b9f8eb36e34c295;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha1a896ba0e3548c658c1368a52ceed1812056065932d5089dd6f729c313c9a8d444da064a3152c0a170cfaaae46117dbc1a12141a453d0f56adc8900def99f1f8dad4f98c8cd5026cafef318b7a223b75a06b72f496dcf7bd227b6a395c15230b930;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2319a133535919bd3d9019f50e89d63fbc1e2b042d37dcefa1f218f746dd2e1b32d82684fff40dc22b05a22cdc6fd359a13c60247cf3d9ab502dfd3f29d41ffe1ef3087091d6ace224155601c6737718a4b5e3d8839695c19cfbd5410139cd0a6dd0;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he012cf991f5ac3577111fe910e994167cfeb214a485d5c6032ef108112482f4804c2b972a08ad4e35b4ea9be909e34528a1f1afa98684c7d5bd9cd26cb92ee356e2457437eebf5c414eb00c2c4188b19d240df10f403323f673c3c1ce31c65246365;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h280744a1cd27bbec9c56819e56fdcaa19ad1a814eda12a3bd8d070aa9036cd3d17d5b66b2230aa8e52885b3b21fad611ae70f19400e86f3c7bfe4b05dc6e859433a7620fc0f11334f1837067c4695440245ab3b4030a00868fb678ca7a900f146fa0;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hccacab80e7001e937d63d03a5c31024aa2cd23e748a94a803fbb90b9caf951062c02adf44dd6d76455bff99d8adcc9646ed52327c6f0915496d7e29d053aefe35e7f36568be06f2ddfca87e3c7202b42afcbad5ee01e3b452bb624b62ad1db535872;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8f0a754ac8e4149539f74c006c11000522b10bc76e3ce55ddf93a8e977bee2569df8c6d3355a03cd8efd39fbbb5260309e5ab2fe3d2d459770b376332b3a49b297219cf86aabc123686b00c8a25f9b05710d248005c847380b7e772d002b751f1f1d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha0e04dc4dbf0e5a7d852b6a2fc5b82bbc62e8a34d3bc1256a38f96d6858517f48a652daec158a8d20514c88020136ba68a1f8e04e719a7c003d6f07a786ce974babe1ae15e80c3f3e52e502a9e7d3402a018f961cbb3d505dc707d2c6231116af13c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h57b8d94241f4add09f4c7ba91fd2a31e9457e7e0fc28958ee3cc99dc25e6394d8d4b79f6b653610f30c84d8b6cbff79d75fc5c1cab985bdeed5a3344fbac33a366ef5bdf5e884c3b368d7f4b1879e0090e950df2c6317dc16980629d86d9d77c4c5a;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h557a4be4d1f16e26778a1d118296f4bc40791a5af42a6553b136e5a486b64b5e9abc8e31e1d00b69abd7ee721b173e2b56f6f1479b7ba4ba68aa935535aaf209d7552023264a3b95ce40fb8cc60260e93b4e9f8bee1bb1d61fd66299cc43323d9070;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbda5eaf96c3118dc23309513913088653831ff72790d37b9d3f921c91713ab7c71489cec857b48f2b663b829bdf0e3ccdb920654cb9a04ba3d80b8094eb5b83384390c8c86ffcbc3ef804c11335325723d6de27c6c121dd245b9b6afdb10776bf003;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h95216f54287e00bb39ae2e16b46c7e1d9b39cad443af3419143fa807a0dee92f8822d15a0af31b7e14e382a1ca3b265de77772bda598022642af900e00c94523684f1bce9278f0f3a42d305e029313cb2f2dc3d49d33d077eedb7da47bab2c0f385d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h53f1ef06ab2b07471a87b394f7ac19f4513cb6119b862e09dc8b967e3728530b230096be4fc58aae6f611d0af3c0f30a5e2198b38e5950824f875d3922e9dc2bdaee2ac7214b365636605865f44e1f88d33f59445afc29f4ff88d36c9c61474d9abe;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hda89de5849a5ccfe23bbb64377222918e31a0715f5bb9c509ae9615606bee6debd392ec2b1d2ae88485d72ae8d4e8792cb515b71359cb04cca18f8eb7838b8b05f7623c21c724e570d679b25dd38b51801c8468ab29861d06ade01685974b04a2aaa;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h91d74ddb5236308fb59f745e713641ed6598058897fe35bdc5c5c6b9ffd7abce63b7b01aeb18705d6e20357a9424947191edca06104fa81807d2729c6acc67e1ae5d346c6743e92f8be4068ba3b2678fe631208d51661cd3f3e43bd9a93564cdff1;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h70b3fa36736015f77fcdafcfa6b10ff217e1265e0a5e59a28a5b8566145709ff5525b3bef5d3995a4f4ec5ef85bd5b9c6da67a47d4b1e391471c7932915873aea16cf846fc723c9602cd3d8871651aa8181ab203d61510a082806b09b1e2ecb4b813;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3ea1fb11baf376672d36418bb17cf2fec2eb8447618e33c39fbd961c680606f441ba7675d2c12b8eb472b8b27661071f31ed3583a8e1fffe75059a086bfb4a35552afaf89d9dd254ec1d24f6a02a4e3f2e17ced892db7db6de1c674744f5f421a77a;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h496a5867fefbeb54546e95a9e4763504078118ef52428d955bb3d9ae209a54ca96592bba0e01614b15cc3b1f9bbd8f38d594abd5d312035addfb464d118952fc34b442814773fcf37d09ddfdcaee0add7b544506b388f4820b31e671cc1685ea6b24;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdebd4566c22c0906a6a4f2fa5656420d4d8312f437d8b1a498e4a30e9e8f5f2b3f1c0c2487876fee75eba2f7803a0e9bdd578be0bd6e4c3d99bfd0587381fc7992cd10e205fcf32460617e92e299452c1ff0bdb0b38760aa3f9d031c04cdde2674ee;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h14ff1a5d6756d75408096af9eef5d9d4827f64478ca4c9659b33034c3634eae11f54a20705cb8d8f33853f7d6ddde814b35e022c4dbf6f621e8e05bd24aaf87c4168d8f430619c36484d02a046aac79ce6a5be5210198471423053d9c5fde6531586;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4151bf1454fdb9663934def2f25ba5cc7e59a35fbce4b06c56fdd04027e7647234d1e7215f4ed0ca85144e8095ccc49b446b94037b95ee2a56c1bd0784c303823b27dfd80fd808b8fd39487f25b1a963d68d7186c840eff578b9e1286358fb80311c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h47ceefaf36c38ff0f4b0b6bf0930036bda83a399515e77be5be136dc037a66de656250e2c524956ce3f4f5b2d134d015216f0283bd495ea4f0bc0561317edefff3a4ec8879c5cf5a83b601b6011ce083673800a525f67a1943314f26adedec9aee13;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hedb40484d4846a98bdc389a89b2879b0669788edc4bdeaac3f8be22db2f67a518bfbe2f21f0f9ef3a4311b5b03a62446f3eabd989755ef8fa9ac529f7ea45e02cb0d1c041b9a66549dc345792f15dc8e434f511e84c00b99870e349a8399ad35dc95;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9ae5e96b08f8650fc1a8e895dcb55e590795382cac023842bae8d0d69e6fe3a553dd88f40a59d75328915eeac81eaae3c8ff3a348eb4ac32852aef3c8b2c1f3c4740298a9607809cec6cdef373a4e75a236594431bdfacda0cc3c25947284401406a;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8cbe4d0cf07b4063ecf534e3cd94cdaf1b99e4da33b8ad56816355f55b7965b461ef12272f967f6c51f828b63c8870a53e81614478df64cf31e3dd3d91d0c16f24bc7392b3ac353718a0ea75e445767ad2f9bebfb2fdf42ec2fa35590f4ed6325de7;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hda3fad26208ab41d5539365dd193ccdaad13903c3726852c067e058a0bff0ddf9b5585ff1cf5b3f707bfe6997cb3f0118d74fdbb80c0e382d54ae16693c47c7f1e25554bc7306f15cb2fceaf2a40879d3ceaa47153d3684bb0091b39e41c62649152;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h755ca9e9bd68ccdbdfc54ffa1c189d9a9be5cad7438022f42bbe1241ea4f18b82c6046279d4f32343e89f5e8283ed50b0e1a1aef3cef0ad7e76b70da7df3c5287ec4173da426b52600031fc60c04e4ecac7c5ad6b24611c3f4d9a744b596467b26dd;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h98363ac9feb18397cea4a7b819f2a013c6ec1cdddc3c5e740535f86e65c2dd3cc18abf1daaab329e2fccf149ee725511b3d59be79d00cc28b77815d338bcafb1f2b59977a279b01909727bb3baefb4994bdae34adec80a9390038024e38b63dbe923;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h463632b9f7df899914ba6e5bddc5bd2f503388961781e8d61402fcf6e027e9fc4542e55b870eeec0e588abfd13df98355e9525ba47ca7840e8a97fe04520e3bff70fa4140ce0d366b54c258221d115d5eebea90bc492d9123972b454150b854e286a;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc0adf01c61a05e5f5ed6bd34ab4008e559bc8ee08c2486a9671f3844cba3ea383a3407d43dac4c00d0f6388db5f3f668759ae0a89fe0f4d635b7e1a6705adf77a353d15e1b817f1892fb45776d59b6b25b776e1c627dd287aa0bbc7f07f4d57be24d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h37df5b209f79ee4cc8984e93ee7bf37abb4b42333aa0aad31f61275bb81c3c989641b0471c455a13572986621a237147cd7c47215d77e887c86a6e166e2f307a51a558895b3b833add1a42e65917cbf83df77a4292fcdd28aa39392d9e2a5be2f8a4;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6cbe6e37dcb8d8eb5a20abcd3cc58734f04163d71e8729c580b8fe6c5300fa9eaa0fd5dcf4291c64ccf606b8c55a282fa97d76564cbc6642b7cdb7a678d596cf8988520fa9f3c6d060308cf01228cfcabe26f8257cbb7d90356b715d337cf88aa19c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdbdaeb711402935e4f314847402cba910888a93041f3293b2b7d4c8b69a42afdf69b4d525f8deee9662915a631ee0e6b48efb2f84aa17121c30d02bddf99cf0616cac3a6a824d95bfa58b3a9a4bcf5b63b27b600edb85131722c3fee1d97e1fb06aa;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hcc8fe1311f554ab951fd04dbd1129c6d41a5fedc7bd1f720bb269414a646fc0a7c37b22125a81dbc07730ee36f14a31bde6a3d5d10fce47a45b2c0d3fdf2aea1efc98d752404b180e30238e1f9c93aba634c724e3d5a47ae1c58c7a037d04562fecb;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h401f0b20080841f42ccf62c4c35681307a6a0193055fea5de08e76352d3d91c48f7af1d6a19c36a60e47d6033ef58e6a2851e54620e232cb1734fe6137f1df1eba2f822c06510f1f02631b4d94f65ad5a1b3bdd0ad7815fea03256ea9f172804f101;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2ffe5b7014d2e0c95309530e2566b622ed756161945a502e8af52cad6ee555945ce7b38d9cb36c7693463bc934bea68d4f1e46591ac6cd192127d3c09208b811b0673b7390bdfd4b131a2cc7db9275b3b10e6fb0214977d4d60a92caef64d7161293;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3082b93e7f9adb35ebd48709a5dbbb7de65805e418b0e5f6e0fe87c11f1f858b1ba6ad1e3c16ce598bf854307a15981bfd9dff9a7994e77a624f5fee3372c495d61246f0a05a35992e098e051bc6c7feb8c849e52f36ff2c073fff50285d8be47fe7;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfa511c03aab618980d376432c3f124182edb2749c24660e99bfc0061c5cf9e0667cbc4b9932cc03ef2b065b3c3d76a5583c6aa4ca83571ab989c58f963ab47155d51d8dc891efa203fc36c93944d5f622a1b38a24a4ad02b612690e0bf02176c6e46;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'heca2bf3ef014b6ed9786414118200597591fa85270d7bac5fceda8f51fbc6e5bde730c6c28cddf6a28018477e0046a2d0879d27b510166eaeeb38c2211b6e89b0bb75006596cfa94019a51f23431bba394944ab6e69298b2f8c1e18fbd1b549dc60c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hcc5f3f4fd2322060239d357cd30dc3f99b502cffd0118f136cd610da010ed7e05bebddfc628d6ceb10662a6f32b660e39611f8201bcbc845cfb563d6bf5d89b0e4b7a9b40470ffdef71d28c9286254f9b808c94da225089cc65c0f691ec5b806e7db;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h12b85acd928080613f9e399b78d0ece688e49ba6e7d0269a2cbaf06c38a0121ebabc61bdcf46ef2afc87aeabbc4fc13e1c67846a8ec87b0cbed75858316ee53554a16c18abbcdbfb81092e2959009342971b0a09b7e5497a1b6ab76a7dc0b205f33;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'haeb20a8b0816be4a83e19b97baa64c17a9be334c54a43c3915b8f092f13030c32cb8196b27bed4ca05e4f81472e50ff1cb0a5c99cc6397dc008d560d4298adc1e642db5cbce2654e7355c54bfc812274ae88cf3f1f907e4b8a626cce5b27269ec446;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h698753ae783b7a2753ddb69710a10fbdaf2c743c16d2e2aff13f47653a4a1fcb9bbe68752f9f0a21a8d73c3ba748a63ae541bc7cd6266588d29911b17342a3b0c41667c8bd73418dabf785e2cc5627b4f43b69166e6ba2a069a2a2d253ecf6452aae;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h47e8f4f3b2143d3fa96a0797996949f60ac16e685424fc1149537fd69dc0cc432e05ebc4e4f0c1ef6957eda3158d2d285dd62195ac15aa7018de6fb372bd20d60a7b348965237aa125b514c0af2ac3650a36c28fe7905633c690cc0ff66a615c80ef;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf758c157d6b686cec0dc0d7204ab61e27bd4225389159fa1310d06cfa231c9dbfa242d25eb442da3aeb8187b4d72d8b7dee38ffb672b2c01d988db2b994e6d566bcdae404c39e9ad54f7a431302bdf6f251ad20bd016d8549338835314e02fe84f47;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h633d7eb5b62e00321a538fa5ee573cbf5182ce8576b328b601bd36a65ef24a06cff71b86c1c5cfdf9cd4672ef578cd257774caed0022ed40b9d83abd8bc33d041bf2aac486237731bf0cc1b58c37bb99bd1f56ecd37d5bbc5a352341f5de3376f800;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h43a78837c02209b4b3d24384c0a4f0e34721bf26c9f9d150ca66426968a903b237b594800bf06497271073c40202b693ab5ed17802faad2bbff90af4611741939062d463893cbf9dd464f974a959b4942d70763a5f4867be62c23dd1f55e781e0261;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h36ab89ad134348aedade4800ee588c9f3d2c07e0a9d4a96d8f2635a3bb5769d29603720e21ef40b1a77c26712eda1f427a9c781a2607b7bafbbba74ec8e4f40df03b86881c9f0c380f5ab07c9b378f80c4a2377e7eb48af6ea06619d8b8a37cf4a40;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h477abdfe3b75b31b88b5fa9188a554bb2bf4fbfd7d0cd1e008f278b61b13120d52d877d6704c6e957b66a364e3b13ab2c21902eeabb75f8f219f4d1d2e1f8bdce120c175a4b87161c53497a21aeff2995944e546d86582161503bfe6473827f27f3;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha8e3cfe4a0cd895fa77ac0e84a87a0518aea07bc69decb99bf25f6146195f6a138f1cc86a658a3b0af1385b7de6c6d50b0c0e86d0473cacc1330612f0144c4ea7a3e22e7d8c162d376d8521f86ebcb0a8062fb54d9051c4ed7014347eb9b6b2ea090;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6482c0d74552996364ac4152933e99ca2febf3cd2bd93d8d91a25e1cb063954f319b0516661e823944ceacf3ed442276ea4ee8270ebb16319b7475087347ec8d0930bdc3c8e64849fddc50978b4668b6afb710dc54029ae6997229280a1d68b90f35;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdf4cb4e0d0fd300794edf982fd483d6b0f4ac0f2fd2a24d24afcc897a5869816aba4911ee6ce309b220ff6687c1743d79aadccbd5ea96449f9e1656cc2b6056ebe6d6839786e58881fd498d27e4ed960dba1d070834eae2701a4de2c690476dba098;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h425f2d2074a6db9e90063c9db6b2d1a28d6c9fa47cbf3ac53257eead21d406c04bbda9b5f86c40d5949c17aa61fb44bf3bff60cfa42ae8f1b645ad0e4db4871d75d912b2f0111a91e7e84d7d4c3f1d2b4d2c7aafd9c4ade8d004f26bcbe5e20428d3;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hefd21c626139ffe8f43a95620285cf150fbb7aa05cba4623150fee8834ef9b741a09428165af935594ae77de174b56700a2f4fe67cb0c486523ebdc8e50eef9140b21d7d23faf7c1ad6e3c29985bcfed40cec8029d764f4a9d8f04b2ef47745b37c0;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h75cf7605120c431946db4d5dbf57be2352a19f8ff3a8c8f5e3c92869edf2709d8cce6daa476a46859da1f907f94a3bf9058fd7fc475ae5642b25a33153c452cd9d262d3baf8440d913b7f71712c73e90e9d90367c1b0385d1fb2915075c6b1b91c25;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h837e43c0d4ed3f23e99186d55226b81f6d57e0eab01824257db33b7188e85496e98164214c6df1dea5c45950a8698d267a98021b4ccfd6016ed308003bd58a6a0d7a0a142cd918d843b8455c62e80479f8dfb51ba6b02691d256590c721ccd0e40ed;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h46e10aa64ff90d348ad716f0a4268496eb668adcfefa2277754b3092cf68c8f1603c2d8d56cef8571a467bbd7c241ccb496401330e5634d9053871bbb9d9aef786e88fe4874ee332fafb4b1170bf425426e293d774c33daa816ad48cc7a77e2ea9df;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h37b15a458459a041f525cc2748063863f6b578610666fd47f167b42859f727688569233f5e31d466e97768b540316e7be4a7833e243aed6c24e9f52673d2c10ee04519c8f7f2b2e7f3ecc228f9d61e24658f2acc0e3b8d7aa5da418a5a8c4c22be04;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8c1f38d6322fbd6b4ea5ea3da182699f300d43d8abed7c66cfe6a57648d3ebb66fffdb4e4821f73496e501a56621e8410847ec0289b1e1e0be41ca95167d9091439fffc027e096d11863849249b6513255640a08e22d135f7f135ddd24f482c6ea1e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd372ca8e83ca0d89dfe6996def3128e3466dd9e43b1273ed93003037bf615733edb78450170d6845a5b27c6179c3f78b0ca94bde84f24262656f5bd970ef2b602e12f02bd403cd9fcc3f14b0295a7386f33a42276b322dc6ed63ced8c74b12bd19cf;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h326acaff4e7650b4fdf4ae7cb7e9628afe77524cc62a9028b0b43fac1015b6226305a4d2bb2b1eb960dc343e6e7022570f0de4611a9d23da05ace6fed866a33149a9588a71d6b9ebbc3fd72d86f71ea54c1b12cdf61b4c03f86b7f1f58015bac875a;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4ceae7e0d469e7d5cd99b90081a96bd94eb38742e4657d3f41f160897834aeb1da1dc350b9c57da9c4d3094717cb2851e4462db6e7b15336bba13069f64a81912929f06f45ed8221cbe3863f0305c5c91e7e4c9abdc5c252cee78b6487d1926717a6;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3af6d8e368451d7e2e3e6602d0a07fa3bcb40b6ef00a6503a114bb673e7393fa4f874e961e1c0f68f7001aa35d57fced92343a7185b87255a0b5b6c374fc94e26a597b88d259483e0fce856ad1eab88ca498541856effe4d10d9ca5a9e62000db517;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8fd6d5d76c3f2ecf2fe2d3895bb9dd8ee4bebcfc84919df8d184c5995a00d86a8322832f66b76d011ba6a4538de96732e016b1c3e30ef127290227aaa413a2a4fe677e741f68eb8a8b35ef155de948b248b97588a76e795d4b08ee2599d0bce35b60;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h880f2b39e31aa96c9aea64bf8de1286fd595257a5a634bcf94b56dc0240d39371b854e3fc00fdfa3e17f190439cd3f2f1dcccf38111655d8d57bcdc47b80eb3a87be425f8d10cf7ed7e2140980b4747a57d3f7b38d9af275c4d65f4f65f468084be8;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4f15776bbc8caa93224e7ebd5281826cb1494c869cf9c8d44b92c6fd85e76d39d4a88c1579dcb0fe039d223016dabf54bfca59bb4b4f0192ead6efb1fbb7f342bb66bd5fb48cdfbd506cbd63eb3779ebc4624e855a4969957c6b664cd29c0b7ad930;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he43530bd717de147ae3559991d6f5aa6e37cb6a7e18bdc00de697621120087f918a1fd83c1032b45a784ecfbc3a0ccdb97a48723795e132906c7f8229cde15d2548c317640200c94fabb12d6611f32515e0cb56a86902e6ddb0d8ea81dc953b41be5;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2f14e80d1bba10b5ea81efbc4d5301442f65db255ed6299b30966e62d0fe4aaad7937911272ceba6e06fba563002e652a491b46b9006d24ef5b0e76dbd3ab7e2fc6b7a912c0f0c95b0be3a695fb2e2de111a81f80f961d31ec21175981beab1da151;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h31c7b8bc8fdddb858d84135ab8a1baea3051488ead34baa8cf150298aea0b84ec74309acc072e2fe3f16283b3696277f5480b6cfc8b852b067236fd17ce2c27b27c89e9404ef6efdd7892f6ef739802333365604bbd5ad26fa2d95da548204af0411;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hff3a7a7328a9f50218c12ac379543d11a1e01bd03c14f773cb20a27f5fd560cee18bbdde158358c42f88d6aff2baac6d9bb0bfed5bafbc6369fa59bcf97049ba6aa20500bfac251563aaa9118a49351b4e6de7560181f3c13f21cce572f3226bc4c4;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6943b9ec6082e1300a0cc311a2217cb97761a5bfb053568961ebd2f73a04a4e10fe687917a65bcb694f8314b1a2c618c1d4137b68b72a53589058d90826f744c91e86c1a0bb46b820b7527b632b761d5477c567156f0fd6167192fedcbd209dea0b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h90d80383a3d88171e6c6c9ebefa35504cb65aa3f4a1797f861333962c067e97f6a683ad78d5bf69dff3ed66752f0c9496aed62412fe0c56ee762a39d4c8d46921ec1bbc126b10085ff2488ff07c19192bd6ba40361c6494b9c27057f75b10c24f6a2;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4c02b725a1a2cb8aa87a375fb960d9f5b99bea054bc1f91df1f17571d3a60bce386b74eec8ba851322b706332fe6c7b38b2e7c532768c5a52aa9eef93d20aed13af94befa4c13ad0dbb55257793bfab3d7a2f2d09aee56231ab4703de232e32ced2f;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb301f309b5687ff065df1ae89f9a32cceca019af6724d962a09d3720785f27819fc6b28cff691321739649e0ae63bbeb4f3aeac0d0b698fe6c403f95a18262caab07c7bc186ab6d30eeb3667d99e8af1096ff51ee3d799c43f1df441c83689764354;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h62ee8bf102e76934a76196fbedb604bdd02ff393e5713a7587bc3a8e91430855a9a7c286c8848663ae0c432f30321c372e7c3edb411af887b7ebfce5816a77a7cb4d30cb84cc30359c64d80d52eae78816869b7150e61a1ea49553515469a8f53b8f;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdac5a83a579cc44aa8956c65a5882a6b737bc7a7111bdbd6aab54957660a2aa1ae901f98af620d28a32761964b870515716aa9a85fced36210cf35cafad48ad15365adb60a7e2583b08d581cbcd011af24921269131f807d8f1e295979a883efa267;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7a71af24de40b8575e6be42794d5ba443f71741d10ea336b6cd8023344c20068a291def125e5afdd4aa09e4e0e1276bd4aacb73d21da54d4fef3ab750769721fc1d79276464a2b091a8c12f033736c2d893a348ec6c33fe887881635f9dcfb301102;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he0fd775ee2dbe2bddf7e874911e55ab8d04bf6b05e1783e898f8eaea1a486503b8956bc34cefd30e9fdac65087e8543bfa86d36fcd6f010e4ecb434e7d05e26bb5042104de99863040f30010911c29dadce6d8074f659f3af89c410f1406cc3d2495;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3d80714487f64e2e687a4f57d23570b7ba02e8283a1488d19b763ff31140eb705ff358df92cd9ad4fa444ba43c1178961e8afb5233d5615438e4d1e3858034b1275d1613d2c7e2e5b13eb2afdef3588a6005dcc2a5403aa5f3af5e81bf2131d16f9;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb6de28f8fe960e297f60e492e23bbae05fd07a327b82d0af92e432551d4063937f0cb8f1c44a376be2d998b7f15649b325491d0494b5ab858a192ce48ec56ace2c747c47719e69f5676d6c37943e2bb4829f7861fe0467cd50fa0ea6495a28eb6474;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he123dd6bad4f5317f2f3109e055b5f535a6a3e0e2e6819091aad10026be73623615d40c164001860a9d6a8bc140f66515784baf86fc437ec365237ed1ffd09ef4a5949519b33614d9ef00f5dac4e549f2a5559c890ef69e936afbfe2588db70a8ff8;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7afb7eb074313d026a5cd263ee4ab6feb0597a4bf41c61da49d774668475bf73db2dd554e3b35294df3cf2d108d6927ce96679a48d6c2f5b52ea3b74c9f54151d75aeb7e493134df712d1be91a010fdae18c99ffef3b54c43b4db7be11479cefccf4;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb80569ae9f7e82a3c8be6c6d69f2b61a50c47b6ce36a5d9c6f9f253b5fb15118e8c55a58b6842b034cf82962782ba1c2637bfa8856365432ed75754d763291d59e1e84afc5171f4cdac4a8f97863fa5bbde5ed94e715aea836295f8320497d3d9ddb;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hec4c7496dae267444e195263a8efcaf5e99f0a69d7d1b605f20fa3e51dcc7232552d8a75832b1323cf030d4afa5fc8beec8afa56e767f93cd7f2f0eaa7ac0356c12a0acb079e1845479123adef5f1788b7f55d608f529d30a831448595842975d1c6;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9ff48bb0cb8ba3f46dbc9a5550135297fd5942ab972c9230b0a78fa2784efdca3b1e66e55a010f6931a142c4b85b94f125a02da479c74565b5ab8004d531b51923795a46f85365621921980b9f61da29f8e4dd62ba2f5d4d957e4d285ec3d5c6b1cb;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h101e24ef1bc4dc15cd7dff25a7722a1bf93bf815b3a41db5d716b202e52b7f43f1cb800c7aed158864a557951390d08dfac9b23c27aa75f0f9ab783364423174f3a30657c3e140c046db83383c128ab446c787ca4fc9b4e0d489810ef35e3e5b3182;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h105f7459c8bfaf32336e019bb6c108c64c02e153b2c0f3ba78c9624333699ce2000adafc8e9c2e084bf92f5d57f1e45bb7b8955c7347b528ac72ba303f38855fd37b6dfc61cd5b3636ca569b8000b0023d3287bce1bc1b0a7defb1e689431cebb736;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h70f19b88fcf2c79fd7f671929366b1ebfef75dd9f94b10bda93e46c5c9b7a062bdf3ad245dab94ca258bee819710c00e6581d3562b7b63029da1caa9b11d2b297c818781d40758439de61af83fb405eddef9425b01d1b70e7a648dfdc3a94e439813;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9b8c5c5017dfa4294fa130b0e8b154e60e1a198522f49764bf3f3ebe2764065e3a96629dd130b335e4b253ff9c3f5e41821bb825d6fad6f2665092c3118eed9d85cf15102a42fb77785ea5e6b8356b521ea8066d704e94c2ee792d0e6e89a243b514;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8048956e03769cf1360da4467d0cccd7e68b5b3fa5f8d43c106fa8e7e982cc123867fea6814998088471c2e313bcb8ba843ded79a1f28f7005e8448c14b77c6273f1161ae1e94a97a11ae6e3443176962b5be272fd37763cf8e4e8967224cb25f9a3;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd7c59fa745e7e31a2d14637310c4d9a762de6fa830e8fac0a151b4a57f5e70d6af122b592ba27a115ad407871ed05884b4499ab592a04bcba9fd1ec2d3475e0995e37b40ecf945631545a2c74643959946f585e6b1e423ab473e152b43bb5f505746;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h93f1553d502ca26e9c5ccd25fff70e949ef19bcfc8e82c849ce323eaad0e0316e0800b500f7a975bb2d4035d9d7795eb1646534887a74fce5f3d9c383cf3adc96e8b308b4490f25a22535b9bffeda58dadcbc3e3615e521369b89cc0c17f992fe872;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h440695297b5c3b555a13ffc3e4eebe9fe88b8397347714fa55d5662ad779297e6a0ae80531c9eecfb0254289e220ad4b2ee6678b15be168bf55c3311ad703753a8f78d445bc353819220cd19437c7e1429f9f588bd21e7766b98252f9baa10f9e835;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb6305659d3452c86af247117a3bc80a5ca3bb0ac7adf11aef468dd30d6f131b30c5c3e9d4b237dca349edf9f43f7192dce84435df982e9c8141a9694c3519b03b8753b5ba146ff5c71e769956f7ec97e2f7337ec357b6ce463c5d03a652db119b9b4;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h27640db4c655d4c773ffb67daccd3670e0f4f4d6195ec96deb607be4d6e0cbff4f59546f886d69f3bc86cbc698f1a6318ea5457c73999bb5a2f9706cce96084da50e60fb77af90145737813311eec57340982894fd521cc52241992b862609d51c97;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h631e552da52240a792da94f38b1e22be57c6901fba0b8abd94c1a25a342d03bf7e3a8ff6a1bc50bc3094637a8a7ed49c0d742b4ed771babfa65de17d903f28218eefdb68b9abf69ae5d4e30542e589eeea5eca65f3e54db86094be00d7cb4a821249;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h636212857259e4cc203a79b2eb8dbf12e4026407bfb350e62611a6c2cd5d026b40790a24c63403d69a1db46faddd05b02afad8586982d726aa90a7d5900ab42f64351bdce58b0bc403ec7b84fc9786d3985b421ee0018d874ad52e7a9ffd161c9e8d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h12dd57443cb7de996853e4eead166ebeeae104a35c3d348f9228d8f2892bf7f5636cf7aad9f9fb8880d0967302b0be100fa0b25183a7c32b22a60d6354228e895714a7885d69f9c332a7fc25814266c28ff445058a67b205d3b2253920ad3cccabee;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2c991f491bef751823797615171058c5f845400cfd8a7d8b8cb3baeb60a5ce4c531c65d58fcdee4478284d78bec88d9baa4c2b22e000361ff901cd57859a0b3215ee27d68ce798f20ebf7f62a9562f8e6a0d8962e69672c5d657224cfb98aaa7035;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1a49d0fcf6944b2bc1f86177a022954a8b64f7b68a0f97fb791d786066fcf35afbd79a52e2a44de1787c00314893f28845f8a337dc4124e3f685b7f7cd15cbab7e796ab662991ad93987492b70c87c965723fcdfaa1bee991b64fd2acf02bb6bcad;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h38f5f2df27ef01a293650d0eb8adae5ec10cdf5c9f0b7ec795191d4b5f702018c8ac5084c69c2c05602a137cd1d155f34a2702a6a705f133f25afb30f3ada1ffb320a3096159f3ca642e7d67a053a5dd299a2bd617e47d959e6105acca16b5617a1a;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'heeef3b597e3640319415bf1fb0c0615f719972348fd1b27ac00e71d8569a72d88822cf7907d83916c264e5ca4ec09519e65da1bbfdef2fe10f29c6643bc61b3167142629f588203e358ca8a23df4d09493b27ce35228cc236a2cb54b7b969ea8eb46;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h50071ce1842a31089d1b512f6eae0784a474b5d882074dd058b1f104f1cd238071e7d38db7d6eddbcd4298bfebdec0e72fa4759fea63e241f6ecb50acb3732346eb7462cb5f92bb432fd38a45764117b513b2885a62385c084a0a84de7b52afb1e55;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h28c32cc3e5967bf814d75e51a0a6b3eea58cb8251d6490e688efb17aea9ac913b0e1e155f0eebda498ee2d454fd9e70c8326ed49f00e99e404130ab80a97e4c8d23133c8fbddde88983cc25cc000fb5b9f255fd90868a829099fc0bb02ba4e59ec2a;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9eae282ff347ce1fb9d6c9d72d4138b424852ce3c4d778da7c2695badb0f639ac96772fd678a4dfb23656d3c71a103942652c12f6e0e164c53ad46a67408ef5755ab7fcd0acdcf243a8345c28a7671f82e18e0e927e558198eeec3fafa7d0f18ea0d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc5c2fc11fbd6b30b48b977530fffc2d47d2512176f7fc0124a523bb383966eca18119b167abbd98bd6785ba162f06de3be03ea2d9a536c01f81cc355df0cd3d11e198d84abfde5bf00b670a83a0de51801ef4c7734acc23ceec3de7948e2e37c81c5;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1e71e0266c52e72758e1e1361b968794665552e7de599df61472ad709f122974d1cc9a421090d08bc76a7c8dd2514cf5a1c46739f049715b34ba5fddc5fa07bf55624781a4cecd37b8e3cc6b2f5e3d07f12b8e512be0fc1806e30798a1e6f19e2a86;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he5896c56ce9fb927ea2135ca1cfff18b36bf44e081092da8ad0f0eb9082696041f8eeec042a63f59392bcfb1aebb7d2d849ebae398899d9aec8bccde90bb3e66af33b68446055fcaa15211757d4295992debf2aa053a996d9e71f31705c6552e854e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6ebb3362bcd56e474a7de0dd6f08e50d36389779d5c5e98e8931a465751b2bc49a06d7fe4b4e6171d2813f7c9836769a0193fe73f582de00b9bca12275901dbce36577a33974de397d0ad22c71f6f4ff6228504ceda5b0036e98dd9389d693aef19;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h777f1d894da45e5d49d145745b1e40d5e65100b5fe5852f6083e77aa9ad36ff54112c7d97e5f27510fb5c3567e62d0d6dfc7eb7ac3a5667c0684a0e69cc684ae68c016b015d15b532aee7f8481c980c01765c0506bb6325e8b3cb56d57df695a3664;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1e857fe89318261d64daba4a2f5a8d3870154aa724e1ca296500733a0ae25626c359a30edb4e658df2949042340c31aedb501474f01f008be26bf36c1cea0ff83c0ac54fc4da3199c17503d1f530a4a0242cb1f9ff7671223b0c508a46de5557feee;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h749c41caa1ce87f4c364c06ac75ce63fa1ed19f5edb796760ab2882e54f95f7776cd96e68601ef3187f0dec9587735c62b43d0f4a30d6087290542db3c1013d6aff2ba8d3186381f86b671027352b6c25aa0838394cd4f8d7169ad728d97ae0b9590;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb7a91d002e94d05d7d1a83b0b58409a65c9784a3440e97a6da04622afebbfc866e924bab83e884b7a343e4d61d7ae46efbc20f7a952d2cb249db993be8ba1939e9d00dcb6877056b95027f271d5c4fed7417dbc488a95fd8f6096540915664cebec4;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1bd3bbd310a30ccaa312d02b2ad620f84bf15de37b53f79a9296da28241d6a2637be01c085eee0ea7273bfec566fc49dba7f5770cd5ea6a4ff3b7986caf370bfa5fb711e05c2c4443b89b0ffe5264f7262efd6b8e0400e2127d17943ae040c86371;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbc08360b6c9b6b0d437c06f1917ea3188a3e07505061626773560188b1a48072825ace888b29e97e6186d69c9d2d97e3fd40c28b466ed70685f5d67b540503b1adda6944f10f648f73ad7419d4550ddc1972500999f797fec784fb96a5cae762ebbf;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8707a5de99a6b3f60953a34838c8e736831c137afd1f2ee2096cf8a18bc2fad47fd5597a7c154680af37cc1b1142de81f7f89e5d9fee7d2d6d0fc0e3455b5f2887e220312323f682f696e79ee91662a0c8cbe623731b7b83304e8c7a7ba3b1449f73;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5c161e2f35245f53f6d87d11bdf22235d22783316a16f900f73ed7a31cac8cd574bf05cfaadc3674c697dbc1bf324f8b1775a81c9011495a04e2919c6f012aeff67ef2a66daaf82040e6a15edbdf1791557e541cc94e933d36e7f1ec6c386e93d0eb;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6d1f42c6d60051733fce81d235d8bf8402021a3424846a29784bcdf47d6d7d5045b1115e15b66ac1130b0e8eea1dbe2ff67a9e193b3e2599a8df8eeac881e22e3dde17d64268b2731ddc6afc8d9c086bb81e7eb5eb249ff348f0ded6f8d6cc8463be;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfe9ba14887d2405b4a401dff472bb3f806016d4c17d31290aecba4a907f5301ad0bf8bd19cda0ed688035f8e9d1969109c83a04c57f0d5c2a3103c42c6ace39a0bd29e01465407a788ef86b2fa90ccaccff064af688648b2815aab044b5274b9d758;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he51bb35e2f8bf44afb669f1fed51b891e2a2ece3bd5cfafac82f92932819f1cca77cf8c249c975d4c087a712d2326f338ee9601493b7ef3dc311e76eef66430a51a32191b53a08d49ce64170bda4d2f26f9e99eeba63417a58bfc27e6d81f59bb8a8;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h646d420f27dc3586c008f3315d188a5b106384852a496699d15fc7f711abaf9cb9f34d00814edde4f211727c557a5724396374e010521ad36ecbe55185369eecb611e17ce89ac3ffa339c2cb5306c7c9dcd012284fdacf8306990560f20af20a58c6;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hcea35672adb32698e408c61c2654013d5ffade86256f49c0f9018e3696d5720e2ecc0235cd620e249a7b6643099eb7a1c84d203bf06ff969a9b451852858dc4ed17da8bd63b43baf29db4f7b938af6baeff41f53d5941899d4435785cdc872b4b441;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h651c3ff5b76e370869319b9b900c895cfe355d9399dca694443b072bd2518158276c68700937d4a6586f8dcfd05f282110c1fbb6ff4dc01ce962b812bcad0c8c8c6706dd04621d51142cc46f25a5689ce7b65ea94a94f8f10049c5d6811e195feaa4;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h45adcfdb2e76d7c4f8fba7c7be2516642ace7275204cb908e81db6843873761ef7ce7d828dad1a11e1de002056257c2d2d880887ce39c749260237a131c3595851ff2a1e5d3ae3d73e789f2ec4f2de026e4c3d9046bd9bf61639e37a4d5066258536;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1bef58dab89239deec4ee680858b039f9b9e9aa6076aff750d52f050a68c596ae6300e6e535dabe0020f62dcc246ae69169227c1e23d911fd974926c96484615ab58617a35d702ff912976dcb885a5e56d189bb46bba46fe669d380867bc3ebd5fd6;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h39d954cf195bfea35c532e84458cf6a1ac49a87efcce1f7abbf6107e8f826a10e35755d187f42e695a50e044574b9991c55948003f602e03ffddb1612cfa501e0c8aca24c618dfba12b7ccce3c51676b3578d05eea5c1151d741b30d9b42b4124624;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha9eb7a207de81006a4f655ee9b487e94e57fb0042a0fd849d57f58848def718b71e0f3f8b00524c70d80b660c30e6b11f791fe49264f961c49e89a2b960ea39245b1b15df572b35d9a77d2a5f463dfb1a614c0a9a0378ebde8c9edf13df2586772b4;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf66ddd03ed455fe5872edb87f5ab948faf0749ade89002f1f8694065b3d6a4d36d349a78ab890c658944be4212ca8c34232ce27df3b16ed4f3cbc7267b71ca292565e6e5401c78a50ed20c065ef55b5931be377991b72522e6d5eb1bc4250ab255d8;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd39749ea26568e51f5cef3cb6bc4557d02049b3e6d99771b23d603969d1e7317e74e433d21c2aa9b3095fd4aa0c714383663012f0092b9a9407cca70ef54ef63d76e1173b869c0f191271e6e87b6dd7dbfe3893c6a7bf8b9301f16aeb300a1ddbae3;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2d9eeca872bec2bfb171df4beec233dba48e2f9e09d0fa3670ed7d8626fb7da239deb95a962d4000b9ab6d1dad9213a95bc792964f300441a703918c1d97085402e928b2bc0e530614ab3590a3624035a6fc545b39609c596fc5ebd4589057b080d7;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h196c0d42985427d5cb6e93b8fc8c5689cf4556f9fb7973f46a361c72f5f88675d847301b651d352bf9e6fcdea602e07f40f9837c40885455e9f5e135e29ab883daa08a21a07e3b4dd812af3939624fb7d57cf73d96c96dec1f44b95ecd7abfee85a6;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4ba90e5aebecd60f35ed300062395d5216d338baf1710dfcc91c78d38e9301414dc45ab1e3fbd434c021f8c24b49f264109a6191e93a200e6e4e2139c12d89a721ea73ec8886e02e8cd74f8b037ee7129f31c1ed3289b19cd3d3392c0307356d5f3;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h446aee884c6e0717413c75cf65c2b9c2e4ae5064fd030b366704a624a7437f65efc38587463edae1458dc82f84534b2bc5472102180a3db5298bfea64778dd861f0ab560c7abc3de64833348ba090148927b3d05b3db65f0fe1e08c385d594a5ba8e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hddba16cba999390042c867be2c1f7751ad5a1418f8e90decb3d35997de0ad790aa25dd06bb3790d340667bd35b0ed9666e7400f7ca0bace0edc3db25e27a12b579676035ee27e978e50230672a55ef21e0ed271932880847d65d0b8576b123bff1e4;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9f0b0bde960ede268e0c3f41397af02793041cca5a5b2fd17cb23dbdf443d1a9a2b06656fb4675c15027cc62a2bf8673f7eaf8a1afcb04b73f6a90985932e0b3cfc05ad8ce1f5e6906281fdde251af712691d547b3925e8ee53002b9cef2a7ac4724;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7e17aecd5865ecaf1080b7de0b2cd23dde87d1029166132c1a411f05b741ccba5c883c130a840a6f0ff1bb0ee6c4ec3efc8cbf7ffadfc6dc122e1fdd7fcefbaa1d936c22905b58e5b5c3e0ac788c77616d6e9ba77f835e3780335b9d374870b4f756;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf2bfcaec53dc37116fac2998c37d20be870b326edc2f44dd436f0765d6e7334349cd6382a66999989f8ccd26181f5e1b718cec06c6627de389022b48c26e51e13a9b8e7d49385d0710a8b441938a0692b63abf63b84ccef696d837cffe71b85796ca;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5255abeda0ce603aa68800dbbde05c8a44e3658031e574c98568337f039431c4fcf0ae8bada089b1e11d067f7094a4d06485619cdc8a27dc97b3e728dd3230074b25cdebcfec02d8c6a19123cef46a7ba47cedba9c02879f5cb7ff051e16346522cb;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9592a9f42dc080d8af2faa35b5ade6741f47c2b1d8bef0e02f39c4a01b4b5ce744387422b13a703a344dec0bcb1b7f9813f84c6f317b08aabbf6fa9ff479bcc36ae262a0c47e4bfdbca9d238bedbd2eb63866b9649da3f6b17bf3c84301befe0702a;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hcf2f1b8db2e7a156e2cbcc1dc3ad57e369b3a1bed9b6a9917d6fa39e14d20cd199319299800e8e1ab4dd6fac84c09925c62b1fc0eecdf8789b1d483ff837216bcdce150f4d6db8a42dbb602e2652756e88175574c169c0e3325ee8174639a0fd3ced;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4fab97584d37599945c28ffbaefcd1cc547d1730b3116002b6bc6fe467cc71473480f07f1dbb08c6d79f681728f1db062792edf3103c707e820c44c059e2f2723b3beffa01f35602b37cac2753e90727eef6d1887203e0ec20c2f9dd4c4d73167f6f;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8e2e19477a6dc0776485a51db83963c02a8e0f7e7c69780893234907555ac08e63b04a1b419d46a89c329eca6f659d3e78694ecb1524ae36c3b8d31efba3c153c07448b8cd4e8a85a841a7d2edf1adbd96bfdef347f40b497d355c791ce1e232ed3c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h32efdc1a3807f90300c4148a21254fe8bb641f4ea960eb44ebaa52a4740818ac3bb618c73748a8333a99815f34f7485f8a4c176f15b0ec4c2c8d8d18da3b426fc5b5d779f280c62d80600e608d467dbe4c56453745859422edd2d235f7a1ae476529;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf35374db300241474fe92d873e3bb1c7cfb05e762a196aa8d3ea3dd127666c2194c955b79b0a229625a294823ef7ba92bbc79c3b7c1451c707cc5681760dcc089bebf56d21804eb7a8fd4f9d13f9bed4f07c96c6ba00ca9496802cb0d6b1f8b945e7;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb257d0e52c999fe01bc92806569d70fca52f57209782fe5e8ab443329dc55ed7467ee2474a917d6528876aeb0ff8893ae740a371e905f2321deebe19e38612b1d6fd8c40b0aab0f54c2a56822bfcd60be5d3606d389bbbc8dbb767b3fa72a6058798;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5d7c2ad9073ef45fd4e99bac0c0d94380c34b576834d58089d5268043ead7c3fa22c0f16312645e5f739dabf724b55eae9cb4c00702bd21e58a9ac8413b5931df655e1a61771525887f5e32a740abcd1dc635c1eb33f1a9b7e4418a51f23850aecfc;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h11ecbf869914c0fc6b123a7dff705f82d6fc1c4dfde5649ab6aad3dfa1833a720c5ebe8f197d3124c7790c156f96a932e7c49ded0115ddcfbc9bf5f55e6f3b62354d73ea59f15a0a71fe0b21ac1082ba29f6dd9fc369996cc8495c00ea0f963ce4aa;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2586f524b69f49ac7d1a6ce405cfbc4f1b3ce32207006606930bc4256fb6077cc774b3518cd4d176d81bc3d73056fc42a1acc0c10067b582fa19b235c015bf1d0a41871405e179420744002213b03acfe2d8b2d741fb5825bb3346c581cd292e03cc;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfb9793a7cbc7a517bd8c24a7e94f3da98e79ea3baaa4e2ef05f501fb1afd71d2bcb9fc837ecd1894b6b7713d0f69c3e897393780f2a482bccd8a764892fc983e34ecde0be53e0a499877c8b19a460f5158f7538ce03b7638299e620753fec42f0259;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfad63a0cb66e5cbaa226a520e2704336fbf809c6c8f56b1bcf2d2927f9cee48b4f0ce33b2b4e6ac958ae57f03b1fbb9b753bfaaa4e33c9bd1fabbbc4bdbc0790267a4dfab1916a90fa319ad57a314b5ae3c435a8ca1ad77046433c20b19598a9ec4e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1077a3b9e26bc1243f5305f6a324abeeda9c4e3b7654fe26ad71cea4294f1cb529f81f13f010b6247249b96c24bc46e876c4637969048cba783b1c548a953fa0786ee779b1d1f21f6d7e08da18cc447c159362cd20d0243d0980b9aead15aef66bcf;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h601ab7f5dfec2c29598c119ec53e373799deb1fae898efa7e3e5596ba3b5552a15d65adbf67db113508e46223bc3b04d89ff98c23a3bcce905e980182aed34e533c419369814b9931ab39ac429304e0310901232024a82f5c86ad0a4e3f307e0c62d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfb83ff67a07e4ffcffc31c5b38d966df3283701e9143ed6e6ec556b6c5ebe26e50c260f19ee3de8f3a7394cf5c7d42e293b3f9e33e6025d7aa101d28f8f97eb29dbffd7042d2b724ecdef9b95ddb1d38927d652eafe31db1b00677b54d0f294df696;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hcac1d025d72d8658cd8340a99179cb9e9a099c9b4d72b19055e9ea75ca9c4db33d43ec0e0c0494f7e4174e36c867e9fc478e6be3b2837f47244fa8b4c6b4f7e0ba09a646fa0790c3668498c5dd69731ecd10441598b53417efae1eae7f6deaa4587;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hffa5d9058a3ed10eeddeb36fdb61763c7c9ab55cb6e5dfff450ef02fc1c284a82a5e9545d4e9c2a6bee5c1ed956057a84cfa40ffe17927301d2afcb2756cf92ddd48e99e9a9d0400d9b6682e6e1281ea3723ef8aa8947d0db0343ea445a75d65e955;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfcbe3da4a9152ff7e22e0051ad508c2148a1572c00c671bfcec7665a518ff10f6a22b5923b97767dc885005594708d01838efcdb0e2b42d61a8f589d043d3ec3816a68764767b20babce0dfea769022ef3210bd81bcdac6571e8ef6f856d1370bb1f;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h48a3ddc73a5ba1680776c469b2b651f5d7f96635388e4630bcc67ff380dcbd5f92e923303320687d4dbe2c0c8ebf61fa20b79f38c969461e1ab99bf1a8864acd7aede59fc0dc207355f8ea46187c8625036845fd2db669781af209a8f2ccdfe9ddfd;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h45cd3a2f0ef8e1e9cabd8fd19db413bc8082f8abeae10f5159e8e404645ec6d58f9cfccaa55c3365294e8359afffb52a011cd16534bb708e8c9da12d9c0002ce409d0ca3e144c8e5afc8d31d9609dd5f6b39da2d307ace864c7748b19e1d504a2e06;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5af72080f89cce25f7a88eee3bf15d10fc376b221c046f82e813f1ba14ea1ac134d66a1b70dcf3587fa0d35c14737748caf52de59fd65c47cf8fd5efc00ae6a891f74ded871af6fa8f3ab8d4cf14728d812c557e77a710e58e75420502b785d9d48d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h52ff406fdc98535740640b4cea8a2f2e5a8483f5724bfbf67425e0c013edf771fd7c92016c53a856fd33b55dabe8c774e7dde291322e2e9475137f155062ca78f61fbca61c450745a7797dc285555234ae0b9ae880da90ea27f1dc2cc3cf093da7d8;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h96d444d02be8a59cd06dcd30f7c5cd722e875a4b2a83aadd22f86f9054e9c545b7d9b37869483a45c8621cd56c93be7f89244b268b9a9bd4389a522d0d8b38da0d590c9d1cc808c1b47086374052112e59b8a24a1a5b852f109c0dac339ae337de57;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5e6427f880b3952132d536d9b1871e972aa864e1f3345f6f04cdd9f86454bbee20d04b721b83c11b49fef2b983dac3b8a73e63fa22b2b29e9d0080cdefbe9794b141f80811699d3df6af9485abd9b7b38527d58efb1e3d30f027ce64dd88833da329;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h13fb52059c81849d97d503242a19acdd9133c7fdb9d3d4e12dfb0ab3f76f4eea47cc753a8605abda2ec759acd8e1e44ec2d3e7b3a61ce12e6133b24102ef727e9bcf7e71ff67b3bac9d6bf767f7c379f6568c5c7bf4f36b5e67afaf290b16917be0f;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf2d0a493a8dba918d1e849ac9acc50395d191a6af227ab3be62bcf28807f96388be99bb6b394f915c89d1cacce98b3ef8cb16f92ea36a868d6dc040922ff20673668d4c8832bf55a97f3f2f79382f4ac4c01205b43f754560332688f2dc8be872f43;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he81622a5dc7fca33c6d3e03d44f3bed1fa576c9454e546fd830e01488e42ca68d567d2f2d2ff4edb51879ded9333cd57d8a4f3d5c7d55871fc2adecfd7cb977eb37b8783d865336080e1d36427724769c6d8029c117954a030aca9989ad3ac561c89;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he54c18927e3a0cb6dd194daf3cfb8600ae30b4519d7e36033fe0aec02ec9aed133193e947b8b9510b1a2972fa3685a3ee676d0191cccfae2e76494cf1130392a747c0b3f5fd464a51760899adf83ea60c568c5c7edff640ad90696d5f5d80afc20c4;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2696dd8498f618da08ca4a2181d5faaa5267bd0427d45c394a384bf73b71f12a163f8b7b3197c05884a47ea9181982f282703f43207ecee07dce0acd79d1b47e99e8c63f14f6234df9d8aacd696dbe186339c8bfc0d71cb9261a4803c49711a5011b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb93f99ab92dba1e827d5a1b8e256138dbf9a1fb49a4341843c1492e1890dab6e325bd1b06cb84749bf1765fd05f2a63d0ba623f0cd74bb734bfa65047b6d290b05d372d66fc24b814b6b568fed955fa96ebf759767ffaee9e25523d6dd89a5fb72ff;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h47ad70d1b1d07becd007e956c7b3395c302c288c591c32ad50b0568f7889572315f939a07eb788a20b393e9a0eae92e27174676fc94a776a78d6a01c8cf067a9ee8211e326c2915a462f739704222055956917e0f2410b230432ce471a025e117abe;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5cbb4b7e5e570a587f2388a7f5354c08a815159cf7dd4c90c3f088f88e5a6d85f81d88784e08c9fed67f5184d5a7609a0ffc47f19888ae6b61749381957b7fb5a33faf3a59d9d3f1e06e802bd52fc70bddfb74354d5d76e5bc6844967ee06cfbaa47;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7930307713b15d058f007fb86b44259eda9bd19d9b778dde84690d097114ec00e8e17bc2e2015451e0a4f0deb901050e54f7609e0288fda2034a38ecaefc7021aa2bbdac06acc7c721b5d99d8ff6a3ba468b5fc538cacc1d69ab4b226a08f54b2c2e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdd39ddf73664dd394dea401fb77d76dba52c7ba884fe7178c288847da723f051417bc42ba1c94c9c6f75bfd61aa0eacb19e1cbbafaf3960637debc7f283e8a0991b1c215ee8c98ddfe8d7e549fcb44c267d7f6561af89c3087cddaabfeeefd993af5;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3cb0b3d65c383843360de5d9239411b86b5554dd52b0f0c2afc904aa4ece99c324bd3c6d243030d9f826daf26fe87c6402b6eb65dc4663a9e66cf2fae6e2737c0413af6f4c5746c4a777bc29bdaad1efe928b96d518dbcff3f1370cf0fd6b5e4d358;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbe99086f2f0f9dabc832266b6420844a6a92741e9e82f42a1557bdae02a231e12be588ced829e670c0239627509ae45133c53d1453fa75fea790271c74964d14129a4443a8df5ddd5ef8faba73ac38bae9c3ff888f9aa541fd918cde48e295bd920e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha1ee4ef19b04d48c5338116682cb8a67454eb6848ade02eab4f26cc4e3c05bf0863317ea9b74ffaa483afa300ad3be1d41dd66d756fa2fbf7a0c205d424a13eb57180b3eede642df25dfcc88083ed65e8ed1ea353bc249ff85c898fdae690757970d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5685ee44f1718b618bc8120cd95a357ada2a82d082a661462dae637e02a258097b62e709a785ba40cc7254d28894e02bab3b54cd907a03eb0f4a461bae39449815d7774986464e83274054a0fb78619202aa40785a6347eed441d50c93e7ea1ed2fe;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h10df82d9e9521a46093ba3ff8db2d5834f2ae4f19f2f888f5a4e3b978a70cd4459648bd12225a1a3e550464e6cb322ff24ce7f76f4cf2b6686ca7241dcb8272fe38d6a983b318e01697a86eb67933c3f34a0622b0497819fdf5b4c28bac6aebc8209;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6dccbeea24937439d64f884be42eaa9545ee6ead491951fe6b73dd780a43a1479702f30211c4ce5801d6da32e4e1b8149e5de00dfcabb14326f02bf4e123cbc776b38f286f5c750429e0f1765faf4aa7ba0608cce0cc1f12707cfd68b266b10b8629;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he58ea0b48f2cb7abcbca229f2e4fc2e931448d639580541ce8c33282b97097e241608ceeb7a601f1de027ed57cac407f0583a5ad2621a5724d19dcf8a0a2e6fff9dff1ad58140f1f010a842487f272dbae15621c94c138a1ff68e1f94a4fd7b38a31;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdf6ab3922f04783402002cd945e20b3580613d17e6f06e1f5d3f12d68f0ea5c94aa03ea6ecf5f3602aff97de9329aba583e3d84c423d69137a8949372d3c75e2e53f03175454da47c98db229acbabcae5df588cd766c52bf2a67c32cac4848b07539;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd9f33a3c99969b21f9dce1d2af2448aaf98018c2d1966d41b2d5fc6800c48e0adf77f826c259e9be4aa783e0a09b08d07e9fb0409a3a8ad4426c3d5ff428a1a6e817b5a1b28123842d8a5fe42cbce963315b127d25ec7a43f2c32ffa364b23ae2051;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5da7ea6165724e3fd05383b0e9a84360525697c2ce1aa67145094658076bd0eb04db9e07de37e86fab764272d3076a3cd22f4f708e57a85df27dd57461e2aa30260647c1f8669abd906a43a1122a78de44193eb741ffbef3b7324aaad95a9169fba7;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h363ad4b4a27c1cb78947e8734f02709c17d0cb7918c5403f427137cc8db6f5717847571927d4e000b8cf361dd51efebe14f50d550757960965e07447a53cfb403d94726fc6bf17b3d4aa51ecc1e4fc2b0eff4c03fc57179f761da60ff9da92ec0cd8;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h708106e3018d9ae83a736db27a4171469f3d1753ff55619a6682897d499a8ac5d3b70eeb7d7ca204a9690e7aa50e256795211ae93736d272e24d161398ccf888c95b94d6d22d04508f231ae6742c59e72daa153fc5b2f55d994e7e0094ba4a677de5;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb5e50ad0a64542ef104415045755f5ab54fc706926f75cce5e2f0c8a0afcd89567f990515c5aa28b2f005b70c137eff5a058f28ec4d5a3460dd844d73404725ef7fcab8367cb2534dbfe143c460ddb16d2117a21ec5f9bb46eca7f5c6d31a4f26235;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb626ab5405f0647f22a54deb5d8c52c576df0e361bc27e46e3db80f373b47f1f36bf911fde56d625933488598f580aa335e0bf4325cd63a80be2c90a3e3e9ecdff125eb18ad0a6e30f3060039215f25a253cea2f337e9b50df98e681303716ddf6e9;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h71b94018690865a0f7c281af1a54eaeb0ae7459295cbaad9d9ed7728fe1489ea1533403c353c62e7b27453dd1954207c59cd057f352e08e46b56e47d9b58a37b937597a1ef3064493ee38827fb718b2af905f73c1204f57c70fc2f296f9e232fb406;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h96606ee57385b49fb24dcb010a5ed5603887aa8f9ef4764e0cdb9f2fb7c9e30dbb61c954859627476f79d41e160c38975aafcba9c58bb95ac855ada72ee61601cb3a63366860584a9d5dcfbdc48d8cc67945a8ec11f044316a1d59f620c483f051ce;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbca778a6cf02dbee56c3f44ebcea00083de9f74b720aa7de6fa3b8af043180b6d86c0167f0bdb897eb9ccf10a8e3ddd5a0ca1af147de053675d9563aa3460b863bd97a17abe606cdeee0afc5e059200eac8d78270644cb44cab3ff3fe678fbbc961b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha7c10b1b2b976e21afebba9f27a4b3266f220cde039e7f3d4d9e77ec8722dd4469883b1469666adf834e9306324ffe0b63702e1375a924b2bea12b811bb028b713dfae7f6c9c53506cd6e76433f76319cb9d617a89c3eadabe9bf2bc824ad15af1aa;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3fce652fc9d8c6e2505f63d6aa21a658f002d00dd238900a962db1cad4fcce5aa6424dc721ad887c82430c7105896c2677f1b1b3fac41c609ce27fdde0383de0e35ab569290e677ee333dc05b855d2d20baa3cadcbac8ec8545c68ec3c2693d02a9c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h23c32587190bf09d453c3f7b9c17e7206f415e2e6f85b96da8086959e6bdb77aff4f1a7987564917877ae54a936df3d827e6e32b4deb48f960a5d69cc9fa37110ea1c03d25b04c9525673095ae178d0c3649e34660a6b009fc8052c540e6acefa703;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h64efaf01b7036228093af36223d4155dafd3b15bdaac5d1d07afe246dde4dcf1262c883cae43df23c56b15c20c66da376735afa29ac3b1e4dccfe5605567f82348ab7d1234a709dc708c8846017b7ad4520a2410145c0178f18ed0f58e706aac49c5;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he86d3b77c2c72c5337f42c7ff7f36600b2d4bc691cfea581d22e2558495c748bfefc9a50c29528a593b0fefa89be67a2803e24127a1b6b7fab54727b5d3a659025ab8f3ae9f1f33d5751e5cd57b38b5fc03b9f039a2d589b664a8ad12f00977aa895;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h724356442e9bea1c0f813460413963132cae64e252d8e6cddc15608d4e14eb48f12160e8294dfc0b613a2fce0286452fbd2309d43d23003df5fe2bcefce70c0c07914c3b4f6e30e5a6cdf70b24b6ec895ed7418958c4000546715b10a20a008c1acc;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h46742a5f6d5fd0b2da8d524ca884a5e8087afe0d1368856e579b3517c5e5b479c2f342e937b1d801f2b7b01c445a46258920ff27e2ff2e544ee353aaf3a23d906663a1e878115b112e03ee284581567b0a269c272ad488b0ea4239232320f4d6f073;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc6a22d5f96ebedeb1c818e7646233a7302af434cb21ce0f7df957a56216e36c44871ac9e7f5e42e903b341dd951d09e70b2dfd91a8c07ea92841aa77886df71af30b76c2c8ff7e58e7570c70274b70910efbbda6c13cfed0cfe4782611eca457298f;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'heeefa222dee2030b778a300fb353d5c1b289f31175b4589ea87dc7b1f02b1ebbbb56ead490e714c7a97d05c6bce2fd493965e0b481899659a5ef25756afa01c0ad742495eef77d6953c0488192ea405d0ec6f9ee37bb4afc38c6e6949c5635098f47;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h12f929b98aabc51cf3ab12b904b0175a70b365e7395ec1a0aad2251bed8437dbc7983164c39eb71d37f7089ba4bdeed5e8236a5b549639a1c69a9fb3b420beccacf414b4735aef0b366a00d83a93627e8dc18a064bdd4b635d707ba1976530796598;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8df7224eb9f5ac2bff9fcd0d9ec28dd6080273d8e0eb3a2cf1d4a25c51921a154e51eedbc595033b1ef6ea102e64febc5b6d2cc3aa97b0684f93c66f024323ed39410a196b2a27f8e370dac960cedcfc4da820e156105fb89e2c3a35d81e9e5a0229;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdd7d07455f75438b2e750005e5a9af84fd966b9309920d612c4034c4d0f713c3ece7faf10fe9a82b50ce7a2d786217d73f4816a3230c661e451ffe39c9e9e147fe5099ebe666a1b29dfc354787ef23bf813dfe821f018c00d170e6a5c3b89a145743;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbe8829d96da203f2707de0cd73b9c8d0d8f0ef1042da55042714a93238d48fac6a375a4c56e1be1328a5b18f199880863ad51f0a2c6cc30bac1879196c3b17057015dc9b3a41d28199a5e098d4fd762e5722aa3a628f85b1852c423ff18ff41fca72;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9f88d673cfce1996d1f0f5b4d21057846e2bb9a020f466ec58f75760ae027245cec583b4d8118f3300c2d3e1f1556ce418c1887cd4929cbd2075977f488759a2a9d0bb1a3143601e2e8e0931b26e9f244431b1e0f766e00ee212cd2f6ad43ee8d70d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h415af0589e4f76ca03df3b25122147d4f8afcf3a2ac82e3653f603cdfdc9527c86ea2764ee2056935dc53e356e3c3f56187e20d1542690c572fca541a4a744e2213de3b0432c584842bab40d0befbb92a0cc6ee4a0e17c6237b237def1f47c43a6eb;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha648abd78c2fb437111c73a88a438a7dc6cca9dc03fa852edf6ba9c0178c33525649536adbb4c1a5cc8621081b681122a200bfab31f8731b99a898591a6309f867c75dde458712aef610c5c6700f9e8210b8961812db914e3f5c57834c0421153101;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb365c51b8f8ba70e1e9802a285a4ce45476ce29ed375367dee968597654304c799758171486908e697e29f325ba4d0d3fb9db8eccb2e60dd405d9ce129e2dbb1b33a53bb2421a88b4dca01120766a91f42aeae165ae1d394b1e54bf2e457612cda21;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf43505b4c9849f343b4fd54f52772530d6c4e6e44624bd445b165e0d8e3f68d99a4f3414880fff8e16a5061fe4a4bc8185d77be188d6ab5c7a0df2215f6e1274a104300d07339194a7f8872de27c8a682f44319e415e43ac8e97ca90cb894b82b4ac;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2c7a592c585b1b86f14bbb19734ee29e2adcd2489cede6e793e73de6716556cb7df34d80c10dcebd7926cbe05ec7244f57fb36f72f3ac22f12c61c4d6c7db0e6d6f6a11879ac28df4d3e7aae12a745f0a22a9c6e78db2c7678a1c136469edd5ade3c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha9349f79cd3ecdb23ea1ab2f646a318fd05a4b2ae7ffe00859c4ca715fe21b009075f7446224882867e676169b1301baa4dc3e5dc4d90a3dd288400274cfd2be99db40dc3fc2827f3576546ffe7509096cca72622ceb8a63ffb6a837884427a7c130;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'haf52c6f3eb1bf45eaef9e4914f46455a362fc9dc89f34856a3ce5fd94eb959a77d9c49a7068c41534c2b2922cdca77ef35fa4cd5eb11e5626d0c6c290e3e99409ffaaad4bba18e133e9003ddeb9cd050be610e143f9596d4c2e7ae684849f58d5c57;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6f79adebceb7ed4001fca6da7a51ca197688c11525e0373a0c7b5141722b8bb9d256e2a605206a7a084ded0f4c5f6678ea0b9178065a3088bff1a5768597573de7a5be5ac9679d19a2ccd87ed9836ebb4e40195b66012740951734166648856acb2c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h20841f6282de328d300e627f90f88268283705a11baf79bcccdebf706a18d9d03d4bd4bbf8650b102f115be0b244bf1db08bf2c42862b74806dfdffa32e37c9384b012462ee990d45b5ea1870b2587d9f372cc7de018cf2c6a89871a5f5da0c5358b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h780254ede8d62a5ff65a5f86d19b1446d32c603095d4f97871807f408e9ce3fd3235f58460b951a186567915f9b42faa27125de98ca3963bbbbac5b1256073a13f12c32495ea8843817a24ffb8b068f55bf3bceef276739465a8b8550f2e98068b8;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb79874e5d5ab6446df6bb7e152f4c7785d1f7016ba9be89499ad5fe11864a949b988680a957bc5f62ec31c5aeceaab07bf793c6ee9f0ed7f9f602ee51d0f3c5fb9597ec065f47e65e35c307ea091bdc2fb51aac66e4e36a5beea8657ffedc9aa481b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1f53eaba2d5740814e1ead1d5629e98866f0a24a61d15253ee4af8e7869a1053a14816903a235d166eaa103015d8e26c52560002d30987b4a83d19aaeb297540faa950c3ae6cc060a0ce8982e10316af553be4e5ed0e35bf9406160d45c459813ea0;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7c85c9e32b4bb406dc15ce4763feba62e6a85f957efb933457a99c9bd05e0c865a4181fbdc4b9ff584c5c550c42cef84fc0d5af3d6d99a9dccdb2dc8da6252d242afa5ee50551103979bb1b51bf98997bbcdd279850cb69dd9a079c2f25b22222315;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8b4b1b735ec2c5524c1a65d0c21051ffe42a205f8e41b9e26c1fafc865c66d1762014c8aa9a025ab1164e9ed1111dea64574d32d93884da4026bc7c208b5e8beb4744647ae282881852c66ba5c7ed596493962621bedc5b4e03bc7045f04662ae499;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h700cb0d602b75b66876977a2bce6c6a04c8367b66157d9a8d5b414efbeb6d17c219ccae448fcf80f88546f49f63dcf5688705739146316a74e4406ecce1eaa218a44d47bd501de52af1a37bc3437e21e00e6c4061fd8ecbd0ea349435f4194e5bbbd;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1ddcaad594bc4e409e46e72178bbbe193646713550c5a9137f77d3c7ee0e6344a536d41a684d2219b5303928d69676618b595d2940e97566e833584c32976e017c72d7daef4bb89551d11d8556e6332eca1532fe7ab12f672e241546a6d5e6a55779;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc27495d1c9fab47cd2726e422355a253e1e80aa0a0d1bd0158c225f51e8293c5fe252616a7cede9ddceb9494184b4924ce5f210284f8f1598f8ccb9609a78de854635d88357b2b6621ecd572b9ee1e4bbbb2a0f6729fade6586b4856228fe8612f29;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7c59c8b4023e12f9f036accc7b72414df744afa3b486664ddd42357d5a6407b8105a3b5929cb244d820f65a380bcec925328baf169150f117b69bc7473c61158bc3c8b0502aef6ed69f118f164580252e6e9bac3b934181ecb2d0a76123cb86d1285;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hac33a626e499d3566d622fabf9f1c157724f2001a6d71b9c4b9b0326b58cdd2f9c1b9341cabd9654ca91063fcb1ad09cee48c3bcee2addc8be54b7416fd281b24bf5b55d050ba9d529611071f7473479dc89aea9a2988dc0f5031974f294bc829074;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6ab5d578b13525c2b9187b67d4d9381f5c5d7b5cf64f0c66967424c0ae07842053332dbdb4a2cabf2ad7a82fafab98a7b91791d341e1184481fe38edc396db8216d8cc20feb9909bb5057453f2f225a0e02cb176c2982a33e10dd486ac07f560d318;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h55306ec0bb9bd6e594f1277dae866e4659ff0c2bb0c494aecaa9e8ae0cda5e03451f7d809f17962d4a029be89198914c2e8f2b455188a0defefeadfdd77bd08745f548c49da229528967796459cfdd74f82515b334b64d38e95f13e35981d114bdd0;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc8d23d9b4c3ba1ddda27839788fef9e55b3d75d7643b727dce84e2708c5c186962c8c010e0f6c4929a16a45bed872197bbb9d28ac62ef5f33b873d8b20cdfc26aa9e4f9485f8ed431c92e82694c4f37607e34f55e86da925e9aa115cf9283f6fa137;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf2f3e986029b4b19a46ccc969de930afcf9dfb699ea23f0f6088ea708c7f5c9b6475916354e20747d9058428c1153f8a2054ae82d44cedc910f44d64fadf8eafeb5b2f5f79f9f495b5e649815887211b5c31b103f32db4aea69834e661042af19686;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4a209b41fc54b3e442c6d79e3516fcbd1b1a96c68e733e1824c020cc11b310459496a7de7865eb3e449e14a86c24a139bc08ae618a5ea5edfca82dfece99732c57d46dbcd3ab28e765436c500bce9c74c9ccaabaf175bda8d3ca724c5cd1145f6aa7;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h69ab2bb102aa54ee67b752cc4b7d8cee0c9bfb7eb7b29586ad06b2195af92ae14564013b1d4b476b9e08bb199c02ab15da0c2dcac18d8093f8defc60a20a41767f10028a22b0ab5f7ba5255a1a6a4f6a4dffb34d71b956ef1b6f2382981b509767a0;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3fe0d31345abc85347f77e0c811cc5dfff28d3fb2939f6ddbd6773b851ed7598e9ace7a65a1f025e6dc77eec408f7efba5897a58af536bbb7d230132797c18d041b704be4bc6cf8cd0e78b8aabc1dd2717a37f4c0318f4afdfc8790bc515d4ab83ba;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf06b5a871598a6f3c4347c773393ef3f767d31d56013fecd2e672b0d564c5c77c69ef908680e86a778457f3e4fc812e70e68d2c727aea2c1ce16619f7980d4e1f03e1dc70c59a0b8a1c4967edf2f67afc51e9234f4eec2252b8b78f7a18ffa8daa90;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h64bd05801d447a476df111706fb9dba99a5560217f7031f315f53d0e029b346553edd8e5187b90545bb4b4243eddc1fed3277f9f2dc28a56594a583ffd8bb12854c7d6370823f1fc56759495ad804582a73a8f6adbcd230a5f37057ea7abcabc2813;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h31fed1a17660db7c5990d9e958923947cc3a9f87764ce5e1514583fbce878cd874d2b93e7d3eb99d2995403664f700239741b009df9b1e937c6019d06700fb481a552be06820ce5fb0ae4b7b22b8d19682f4ad072b636e0a59a1fb541b6ef4009366;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h66f37c2ce93681fbaf27eea35496bfbf9bb01f0e4e79ce201357d54f662df429ff5022c4b62a896a244c938855203d2a3e750decf001c4cac65703c696807779bc4af0d7350e1b8efc5ee8a677d004ba992f6b79fdc2db216c6947c55ed1ddedcf1e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h474e356ab27c92164afdd7ed2876482d9eff0407e9d9b2becff686da8af12ad646e29a390b0122352b41a2d5417f5c1829ac872fb5d6e40b16d9defc28d22d08ae36b9f8094d25cfa335b2fb2b7837282f27360bf04cd3c8dea5464374e3912c0714;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h44de6db946fcfee0436771597199143e64382817fe41f29174995220147f42ce65a2dbe6d08fd7731a5a471e16836636c0627d7c5122a8545e992fe903b87e6924f19c232f5eed3977f3d282de2610f8be7340a210d11a23f485974b557676f4e49d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4512896dd2335ab7e545ab49b9b2c30106cf158184645477856de1907c89cbe18f7163afa191bfd65216d0fe16c772ea8e29e3b698b2b4f595f7ef75d4711251973a4cdd982b6878624359e997be474c6b379c1fbd8e800ebc36a66d8b564f7c9b0a;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h745815402b4d6264863c3a9eececf0cb391f9f97362eeff0f96eab8932bcb239d4c6f9e2bc1ed5ba68fe11616096c47cbb2d49ddcf27c6dcc5b6ef4bc525a37fe20f6bd255d487f45c273bbd6fb64478289ccd94aea52249215c4f982ca384b0753d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h647202bb9d064c07a67f04e0fa07359e2e4450ec20ed9c90762d56eeee4484ee2cc0bc9361cc643e8449d712059fc4f19818183beae6702b9c0083a923bdd41ff6bb4e3bacb0065c32f4c4616cda74127789deca6fbdb9e54d66094af33f48adb545;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3bb8016479dab04ae1ce36c1c90a605f3cc43b2fff62de5e6931255a8d0547f6ae71bc2ee63a465dee622ec617534d2e2e943726be2a63fbadc7ac46ab97dcf3d365d52db8b9898de6bc1175ca923d4c42783312527d6cb08d1f0eaef326fc129f6a;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2d5cd1205a37397d0e4e8196e03812c7b3fc89e1362830b76131d5afb02d9db6afd3597bd2d41bb6832a328bbc0a8a4d18ac2f4afbab3060ef49243283c324551d9d48e30e61d65d25f936f54af36929262ea8f4c93395de1e19136174842fa630e1;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfc99eaf35bb094f44056fea7e5144fdcaf4f7f8ef32ecdff827273c63f65f067652d3884fd68d9c9bbd7ba10587715ae2a893bc96b1a08c7d0cc802379bbd9a4952ffe9e5ebd3442edecfa4163a29d89050fe83524f8ab26ae6b2325d2919612add0;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2e854b6b8090d47ef2598a130ad4cbc1a4e43abdc9f941215c7fc3a5abf69ce2f7ec975fac4114cca1fba142228d2b5868dea7b0360daa1e6bc94fed3b07e898801aab1a5466a84c1bb67bc24743202268708db21009208566c7352b443da564f266;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1bfe12aaefaefb4f95d8292c9f99ecf2f91b50a7b5eb12a5d0a753e9bb84205ed946aed605dbf8b4c5fb47b77db4290ea0791bc9d6110129ad5b392b0cf8eabec52ed60bd0b33940a21758164b66e87ef4dc04a9a4bd79eae61ceb6fba22c812c081;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2726dc4fae654f81ab5197e91f042414ba5b2eb3cfc90b2e08471f7d98665fbe4e5cf2845cd441fd4c1ccea0102ec5f259cba11393e5b59357bf8a7c2413cc09d67aa4a755f1a87850ca9c00fc067c8b894050a2db790c2bcf363c24fafdc262386e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7835fca8c45b3596a5db3f8b30faeb459f2150345765ff9acf125a69e37194008c11cc54722f2edeed71ef57cc4af3335c6bb10fc35a789142008e7aa01567e2cf70d9b618d2ca5b4ec449856c934fe2625c1edbab812d75c53ebd446b2eafdeaf5;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he89895e9a7139df4016183d6693d32e11bdc62f7627d02b6e46cd5de8ea9511e9862dc2df738c36fa44c2fe42eebe61d1da7a6f841a07f318067a977f9ff5bdc41f1e5e92f3710f8aff9b2cca9a3e545972c92a0829d4ed3a3a123fbf5fd4e63657e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h50f8b91d1acfed13f43129a8c9877c5b2d41cf6296ac7683e01e047d9fe15e1deed8c30df3344164601ca1ad346997e02a0d9fae3c7dee9cf785315c833f4764f9e398d6d0fd4bafbc2117e7840d313f3dc6ec93238c5d9179f64235d80c22142f04;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4fbf4ccae35303434c1f7a173fcee61067ee5092354c822c8524fa6ede485ccb97459ea5c8e0acb0ec6050f2e5a7e0e061b73672ca38b6e42046b268c22333689ea83147f94ca6735f93027cd5735efa45ad7bc1045068a6b4c98f4b140d158fac3b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc4a115512e8646fd9c74fdc4dcbccd7cef7c5ab90eff1304647c46c7691210e30fd6ec3fee49c5f9af6ac7fd5d4ef4ef0f2af21eb3db00ee29571ca5098f6a67fd16706b20f401bb55bdae97b4c7e26033de7206f893a58dd53dd0c60d53a078a1f8;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8ac631361b71ec5e5d346fcb27c541cc6ddb6f8a4261d21c69f66bc2ea7735b60c9b14ac08bb59c4e3f457a9cfc330b893562de140f87d91b86a63c07b2aa0e42120136a22f6192beb3c112534f35e44b8d8fe35b56def8e70b5e4ad4f5cb1372878;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he10cfe0d318d30028fa606bb13ad5f65b2400270b852614460216daef9667f660b8b16a28144aa21d8095bd7cf9ae0c68a213bd95ef73090869528733d58c3b565f03da46da44826c87da19a1d0321063d277c8286aff4eb10c6b4abaa9ceb3c80b4;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h295878e8805fad0213e11a5f4bb955bd2dd1665100f6f974cfd1d392fab8c72c3865b1b590a9215605486cff7ad968fe6ef42a2ce54bf1d427845ff7b027e3edcd205ce6afc3bc8291aaa54917cfd86e3d5d3c83804d2fedc52fe3bea50e35f4cd33;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5a7ce51977cd3fbc7175c72977956c6413c2322ba9a261fba6df07f8c86eb2fea6fc644dfe06f436a6b120ef82ef28db41b709f6f678b65039c902014d5b59955b8dae5b8e4fb7119ec5148e07f61fd7b1baff3bbad8681c0b84e5238b6f2bea0ef6;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb48e4f8e0fdf2af7972056c0ec2aebce3a42139a9765207b4b23cb2392a61eda72255c6ef1954b6c3c22b6b6ac46dcfb1639acf0a7f60b9169bf5d480e44e811dd1fde69d068c132d1c35d30b8cf12c94a46800f4f108a9ddce019ce436073cc8921;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbc6d5a071ce7e6307806ae4d0f41dd96cd8dbc3d9dd532a93398093423f8a7a80e3ce583fec05980eafa089372911f48a0f8e13d18b6740b062e460a8aaa64eec3737fb325c0c45ada4deb92367ae79194b60eea44846687bbb12de9107142e8a701;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2988cc6ae69bff9a4bb6c429f66151c906cb383e640fc5c776414e5fe7073cfb29453b981b515915e79f0d9f598f4a21a06d777d03b1a8812d9c46499ce9c839c1f237c40858dfcfb30aa5792de8691958c0e139a0c68021e66ffee6614fcb20b476;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6528d408491e6823a98053c4620133d87a37902a5ed2bce58ceebce6cddc8633bbb3c04a52d438d0d668403be3c6360a6efc35c068aeebf90cb2acb9d9abda7e0f9da94a5789fab11694c70ec2d21eec6e93da7a3a5af86992f4f843690be79a7ae8;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h50ff2518722fd6bd245f99b8b5f6d03801ffbfd99c20e35294e1023a4b9be27c7f680c809ce4177527d2e5de317482416eb40fa30e4b83dd9d200df591b7a784260fc0e547a60a7408dd0732c76a145ba0ba16f33a98d07df0c0a85bba0d7b900717;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5e960d0215482dbf819c1c5acd634f4efc68dcdca7768887d5a438cdf1c5bece89769ea61f0d8c6d6607fa8e71329b7994c9f691d71a1781792fcdc90f57da3e20b2d50110323e01514975c5b8d14ce4d4e44055eacce57114f961bdbab9f05add60;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7e4e4e6bd5175a9fbd658dd4a76d839ed6feddef13fc289b42dd40d12b890104da4dc556107fa1473bba1e8420898881665551cf25e45c4a2b8e7c9b15dd9920f65b3874916841b31dfa3349a275c0dbb40ea20882fddf0662f40120c3696ab1c3ea;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h85dbe2efe4056f2a2120f9da8b6ce184b79bea44acc311053038edd46a6262e6d99a8bf86d5cc9181d7c90aea741ddc67690297cdaaffdce6a0ebc903afe483f8c6ebfb8aaa76f6b3cf6aa607a38d1e9ddbe6e75e6221ed0221713d80041e684b419;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd95841466c412e5a295e24feb3bbfbbcf33ff3248a929925269f7cee78688b9513fbaaf5dafd419b33666ac0fdef7f44f1c7316e192cdf35a7a88678df45d9077f473894b3307a8fc689d6d007442d7d54cf84bcd6e676d34c9c99ea254507e75156;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfe9e3c0f019217fa3bc5ef7f65ff89f3f3693e330ef326b8bc4dd9da9ba95caadbee7206f2f8d234af56fc9b9a6b995aebe03f81388329d244c0d9fbf430ae3be2c1f95094319e6c0253a160c26eee0003cebfd0337a8353f24929e6ff4c52b30dac;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbdea82d269a5ccad75e545cfe43bdcbd80cbd29f1920872fe5a1a0280e86427d6068f47199d55ff0f1eab5c3421b2eb958b2b0037b9ead69e2415da8707c5dd58f32c1b6b3a6cda02341fc58cf6dd5808fcd442ae085db1fdd99939c8befa187f11f;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1111393cebaa2a68a34ddbe1d08bb881b3b5621baf267b1c4fee6354f12208a02e6686cb5a561c59b22be203583aa1108f66fadabb10f83123c726f503a9c6638f6b395c66a7b0bfa28946499df643abe0c3050c28398901c6b9334f4b5229d1c9ea;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h35d1d1ce25870aeb2cafac9eeebb8142e93354c638ae9dc7a597360cfa8ffbac31e9424716f48526ab4887235f0726cea5cec60764651b6f10fb265c049e98ba9d53b24763dabaa9dde9b09ef1bedeebb76a1f13b5c857c6db7acd32aa0f283ef235;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h992f5da150aab5bb8f5c1a5498028c0f056b6d29a935c312022222fe9c07d4b23a8ea02f714dfe63975f9a40dc2f3d928c05d1ee4535206ceced3e2b28a913c7069d5a12c011ac662ddbff3d1af32c25b38c69d923cd9d54e357b21f51e69781fe7d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6c34c0f0c50c7bfffea2fd4dfbc4c99d297c7ca03bddb6c10c035e487d467ae4eaa966ad2b75c25e7e296e6d9826d2b984156407c2f97ed8b330b3cecaa4bcbac86a4739045aaa9dabc38882860c3dfc32deca0825971af5bcf5fdd332d232488a17;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc076a3c4301f9f5179d93796aacfcf99e99be096ee6d96a988c655f2405609ed7a57171ee6875bf61a9eec3fe07c83413b0f3eab9179a298ac71f74024498fb3c3430d9ea4d7425aef08a72468d47dc02b2a7fff97d347562b03fa9dc191e999ae6b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h504773b6ef040c7307aba2e4ff91564c2bfef06b5cc1d07e218a4f03f4b8e1846f645ee37b42925c42618f7746790b4a475afc60e563be9717a9d9ed3fb26de2ffdd788bbd1f9ff35db6e2a0ab5f8a13c11e04ab36577e6f49a8e3a71ed90e5ddab8;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2938f7600ac42f50e3e2f657558145587dd64cad57d1c7a3bc947f3ffe856649047c864c6ca0baa75ef41fcca4031ae29fcacc52a70511d1f071a7f8d63589fe711d386a2bc7519b145834ccb4ade13be37c49f3381d5ef01487c5a6f372271cb4c3;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h53faf0c2e6bdb41b3ceeed5c4dcd779f0e2a9d5eadefe9bdecef6f9a7dfad9cecf1ce2fff8c382dbc12dc20c46dbcdbb99dadf3e5138aae8522e8e870f65ba6b5306dfcf7741528bea7f2722cac9cd4be4b50b56f6b03da66127c0c2a8f0ba3db296;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd570100e210240054ffe9009a9470cce6c3849f184bfef338d1a0e0bf47fd7c8d30ee6295cc4ee2b04dfe3cd775be9723e55ff7009c6635aac24220290b316b047a2ae47ab8c1ba2caf460a22500c3d6a48424bf92314f9f30f86bcfaa5d48343531;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc4247959bac6deeb10d9d09aef1a5b90197f3fab2b02edbb9f2b5ab7c43a7fb66b82d6c668449f103882cdaeaf88cc89c6803eab7c89c9ab151ca3c4abd27177a6ae2f4fc0cb46727d8a0d558b9d0501b07da91a883b7e3acc8128113baefd477729;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h31110baf20b14ccffc726a12228ba3bfe90e6b3c489dbaa6a8ec99adcc47585e4b165f4a71da42a7eba9486f8c2b76c7e0488842672427638548601bf8d95c30b7fd7961a7472c3d63545dacf56a489765a61c2130bf0ffdeb66ae0392a94200df0e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'haede46ab3ef06f711ef2d4ed1014bc8b1b06ce5c2c6a3db41ed0275ac94704d5c9d07fed3a957f9ef11dc133d4d5a97ca294834fd892efd971417227a4ec385aff77aa02409226a29445e63b25b5e75f7ac45c60aeb2ede1598152c1ddd56d382146;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8549ed92244cb02d3ea4434ac5cc9ff758b19d517501f55a992bdb711e916ce9125b7329d918597eb71a8a2f3156f4c638518e412635dc780f50679ac4c84f09c4f03db8dfcd82588824ee83dd6a7f948fa81ed2d91574df6c3e591744972e2527f2;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h348cf40b7fca54dd6d38829653109c3e0f121566775647b5860699cd2d8ada832b09918b570c37c42dcceea622e45305e4b8c6b295f32b24139885f70ce24f9efdde2ef8fed4035842649569e8888ddec307554109d8ee429dc1977c741aa920b251;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfd59d623f60bdd2355c743718cf288d2d141d60c98db5052d606302e4697f6daaf1815a33e7b9b28842f5137e8a29ebdd16f6a302f7d95aff50ed27d205584e1881b3e896787a3ee086c85253281c90d53d245da89e69f55eb67dcf9fae328f7b279;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9cc066b4df8a0e6f554e79d94f8182b9d818bfad8798586d3f8cdcf723fd7ee129c41df9a44a7ccb52f485f00cccd40cdb3a665e5d5d98c2303b2ce1b5d0b19f2a8d86f8ce0712c4c31d1f8fa11232e9fdba1543a7cfcc910c25209f246e8ecc9802;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he54dd239d567d05f0a62d35eec75b627889838739607a3067357942f4d17da1a6c90b600ebe97bb67a6514828aa3178eb0c66d8074447eae08bf8ebc4d31874e571d5b8eb6a6e1ef79140fa4995588f6b2a75dbf25770f164fe99e66cd7b0e3a26c3;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha4043242f16fddb2a3ff4afd16d05313ba6cbdd1f92f1c4ff34f0f087a4f77d61e288df2ea52f065e6496ada8b63efa0fde7ca00880182d63f8ff8f1e4dfc4d196120c65b530e8b71441e61e58c658edf270e462f8f4cda3d20e262e01ade3664c92;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6392f2b3535412f94440cb76797fa53fc5b64d9335667d71c06d338ca0ed755059c2456ce9c85add53cffdea02161495ccb8874dc6ec0187d2161b7d789a1864633f038de0f9da05e5237a7d8683f4fe9b8ceb774d827e18f2a7adadd1d539e983ad;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb31553a6a8d27eb1ef57a3c8f87bb7a0197a7c5f7862dc9ea846174153a9e36bbbd121b7b8e2d8ab7624d500f887dc1d6aae0d7547f35d2ca0a2587b10ac78104df26e0483ab6bbec49d3cfc22daf380beb18912bde48fc83e67a43cb1363b773558;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hde71ba4228b8d1f5f8549200e04dc537e2f863d4b79ad73904f0b9773aeb4fa46134bd243c7928251bef4bc52db154e8903023030e41d157385e608cc4ef51f67d2460846f7f10aa9e42e9df5a2131dab96f392cec9cc674917c3db78126ff809c9c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h463650009a0633e5b1f52c7ac57f01fa672c1ef7cf5b6533e6c6da1dbb2797e80a6965837cde94328a6a5eaf00c8ae7aedbd9d6ddcf4473b5013490e3fcdb5024f2393b7641b5cb2bb0a69923598bbd0f51ddbc8d688872bb8cbaa0b6f8bdfe5e166;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h56c3db49b0ee6b8ecc5f9f65fa429bb2823609048ea2b068072a6b8db4b5feea435bf97a3828f60f68d99a7fd2c062944417c8381bfe397ff5fc11303825c6eda348ffafd80c0f4ed440443b5656cb6bfbdef10291a8286d786cc62e82f17f001ccf;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9cbbb9c89221f6f8149f20d979e4edade8416837d462e0e4b9e899d5e1b369b6fb9f0842357b17418da14a4d4b35d254c14506aac1d4a1f8ad1cd00e48ee19ce4ee6f4e13ca042e4d47565fc3ddd6c524c358462aae35931147fb981d759e7b4f902;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hda954a355f68c12f5a73b923fe02a6dc1df7d1e16da1d061e6ca31968bcb5426665a556cc4bc81103f679691b1211fd35ee9d9f7cbc06af73883988fc2215c150a9cd8e787740a8b65a89d66f18a56fecb15588acdb16ac3f7f0ffa5dc0d0229207b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h33cac2ae9c2a0dcc66838f081e705d46a6f841b8fe9e67cc85887f8190ba85355fd58cf96c51e51195f7c84c77b28e510e7d9b3626afee8add027b1a7743ead5ad7a52768695222a1a8a61a09a2eb29921d735a9958d34ec0268610522723223835b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he6b7e560c0c13540ebe76850c817fe52a05c8cda1f8ed1c1b3f0cffd6431c8916a5a48acf6de0c26551c7e9fa37c9b8fc36d5aef6f25aea98a647de62a75dc827c548792ed94b20d4117d279a42381740ee8d425279c1a518ec13d35d9b85fdf76b7;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he582dc5869f1c28070252abd45fed8bbafa8ba832d77d2daea3c7f7280d6628f1254cf969985a9b5fe4decb1b34f50b764f99f3fae5c2dc5ed210389a417fbe78ab2db1beb2fc4e86eea8dd3d29ac3aa5171c20b09bd46cb59bbca00495c6bc442eb;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h86b938b40cce1dcbe0ff53a80793567555ce15838b44f2f9918424dae7b9765e99c6bfb461d2707613d8827640be0666f810406183e037cdc45c1660f09a14f7f96b2cce7e5675cbbacacc60a56c970e5d625a6d6ad930db62f054d42ffc4fd71001;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h57b56f5320ecef18b0f718002329427d787549df5faa6ddb1449557817eee6af161d8ce15caebc3ecdd99ce084a8333218542462a2dc224eabc35495db4ebc1ec1cac96329d15b5b52dded9f2035d63f559b1d1a6ae5e7cab3af88c8d32aa0eba824;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h96a96d1f55f4799915df7751399647eed1e9d86000a2bf95e99e0c50a9f017762f6cdaa3480ce88e1045c42af251d9c8f52c5053d9f9e0d314a488a2ddea74725026e578d91d9c059420ae06ef01f4ef839f73f27672dfff173b4ca33f36eec3bf61;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h61059666749635a1b766cf41ca125570b8108f93d07308247cd2333398d095f7c347a365799daec342d0dedce1400516d6874947c2e91814f6700e1a5eead08b81dfa19f669dae8f5c956fa85f92e37a2f9b947d153c433c6b0ea2453a4c81262e5e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9f8762551b5b62038222e55442d2d22a13257090540e6a96f122a9fce6f13cc2c77e0903b5171a8e077865a8f7f654a67dc5cf13db99860dca1b827fd56e8d401ced96db62805753775d6a972fbbc64f1e138989e016b1ac0f9e44bf0ba33b9beb00;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb2335b06cabb06db74d0d17514b5e8cfaa30865d056a959cd0c45c1262899fb0c9ab3d992fca3f6efee8fb3d9a4b59c9090a62f674aba3c10b35df8e62433245105ce8f13e63613c368e5c09dd694f8400977018f273c5daab89bfe318bb3ae7f43d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h95c7e4b8f6d55c675b00c87477c5a4e019fdc91444d2ddc88c5695bdf8d153774d89ee4cd97e6aa3e4ea3889e5538e28c1d09e1e95334735995c8105cb7bd0729216bb4ae38d4efac545c7dfb93802063a5f7ec5ec7680fba91a27b7f8d99a7666aa;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hace9605d949de9613005abfa15fe91d7cff72b1bb53b1b94c2d3114bb53efcc3ea16984412fd757fa8826e7069df19c204a7add90777cfbdeeff9db0b73287cd664c835e945cbac5cf9715e5f906f07410b0f29d820de9801a5f364f92acdc777e74;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5d6129b4229162444b9bcd4f4ba2d3b82a42537838e3fa406d13ddf1989e1df89f7505f1bd33f2a8167c0a865c7d81fd32e3db48c545e94cc6e408adcd91be42b411fbff0a366cb0b6c22d46abe7463b07db04194182be45d9190dbd59da96f6a024;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7423a464695863895a6e2d867f537360a726c340eac342257facd1c414f87f98f1573e7f18dbf8d3bc3f795631ccb76e53267c48514e214d650a1eb1d7ecdefed81783088be066cf728ede335ead230d82b13c2b67f93a99c024f2d816c7dd3d2ef6;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdf57da48ec545e4b24826e508b978f1f2186a9f8a3bd664c1e3a72a923f77670ebda886f085cd1fcd4e2a2efb1f1563454cd784728a0e46f0f98c86316c26827daad202bae0b882c21b2d74be2638a21794efc79425466889d892e2e1ddd26049e47;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5552bc6a36f424c72e93cd5fe481f3eb30513fe1fbf84c380585a0e2c48b3f1c3e4ed9a5cb3909081a476d6061152b163cc5690896e4fe565fbaa6e797675a508adefd524e17001524d171ea033c326c73d0f123b324ae86a53d4f4316192fdb854f;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb931910f1ad2fdd02016227dea457ba53b3dab24465fc87602d41dd64c451c591c08eea1a7d34041fbcfed52393fd33ccbec29342df892a1ba7e41bd2ee9d6bf7d506ea115f2e9eb1f7ae40b3b25b42ac0eac1f28073413f0281cbe7a8af9e99906b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2ea0d4d1b7040f9f519b26048eb21330414e591e147d0a64d8ba64813c6f2fe60e7dbe0e5bc805c6f148d5abaa4e65954f70b3770ee4863d81610be078093c22809f8cbc0f55ee8a368e8e4c44bb3e215232a268af501e0294a55b0e9ca3503839c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb6ebdb04406a8e7a784e8de6c1e6fa4ffa64a78c40ab10bc0033ca3bc2df742b3cc1e6c9cc4cf3e626f21f0326a64c44a54b48afdd8f0767a87feb079de5bc553006a0d6cfdb8a4405101cc3c0b28bb03fa4647e2339d1a837c94a949672f80e3270;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h28f573dc4c4c90050b7c8e5e6a2973ba688da2718be13e83a15cc3e196421e2bf6d3f995208a5c31d646e199e143d8522bcc1ff9369440e5fd9b5d1c478574482f6c658a6f8e8dd4db6bd77bb679a54ef4d6d00a216624c40f5764a9c9d7709ae8ac;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6e16a00644f87cbe234a9caf985b473d37641ff1eb496ff640f82fcbf59ed6c44fa02bbc9ca047031d72e3b99626218ddcf0f541e57bfb4ea654e5edca3ae3650901048a19a9652aa869c1f12ecb45451bdb1d0e90622a25e9422975d46b8779c922;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h166db422b5343f691317373565b54ba474638bee733d94444c7f13cec1ba0cecfa653b8f2cd8c260c437b7dc674fcf2eb04c503d5827458d0bdf8417e8ba89c0c0ed987cf3531ba27c1e827ee089c22b0b1b4ee0f9b0c69c9f3f3e6cc1a4cb8c0cf0;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hae570ec48a5dbb3c4828921b99c1261c16c28e97963e258f3f4c72b95df576fbfb5f7154a916978e3937a9348a00ceadbf34aa4b37becd8c61014f75a6c261adac8cb6e39001abacd21eee0a2f13841c59802783321522fffce4f94d011c906abe98;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha142be85fc8977e7d09d04ae02d2fc4ebde3f747dccd81d389e74a5c693c2d372870cf3a3ad56847c6f05ceb7ce844fa2cf929731f6035182ffa1cce093235d7559daa48c1ab993620f50007e7235eaa5b8ce8d4d127484de4508d6ff93d65ee5ee;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf249b7316d79c5ddcffec49cb612fb757375344f0f6121eb96c7ae8da12428cd09e3709858173fc7bdffd1e06b4b40392efa51967d41b1a4b2749cb0ba437ce6e1e4dfc19bb6c2ef2fc367b5b7f3a5369af0e91545bf9498741c572527a312fd02e2;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h62e2455b2a8503dd2f0c60553cb807c2c56fbb1a425425aa9c0a0125dc85adf8d83364713d6eb29cf175826795727204993356fcd05355b2e29eb1d8c82f0dd390045c38cc9892f228c79107b800a10c046896efad2b8950f209cb53f7fe8d5faf1;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h23b950bc83c8220b2c0dae104f53aba604ce39518ddee9b66cf5c3fe311d943d6f9f4b8bdeb0af89f119e35cbc9c4af64c1d0a3edd192436e759aefa97bc4c7870b91d8397087952a5e643c9b48c85a557dfe46cad93391c68d67184d2e1f5007e38;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h426b2ea1815e17de7fb88a3d05dc84d7353337335ef2c23ecf2c0e210fed5ab742fbad82b2ba29476efbe7475af216dea1fb8c82bf9849e3848adc0474f9939a8c3dc3bd4392a5d3956ac418bc078becba28e4c311f736ee541f7057ea0150ca5a1f;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1392286de467a561faca2a448879310f5416934d42572ea266a95d4f6f794a15eac63adf536835d6a81b1decf181a53851616fa421359f05dcc0ce418e0006f8c917dd312a544cceab9d826dfe5cdf67aa621c80b2df58440d9a922038c7c9aa37fd;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2e351d0810a76dae2273b8ea4f03866f6c2d8d2402d6357d9161cc9fc39bd4f4012d39e6a4e96d31ee32ab53fd2d990ce24abe73fbeddc347cf69c47e06256e0204687be1098630595ff8e92ec244e8a7e1208d5d179dd23428961fbeb62b1bd6570;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h83202e069d38c5b67ae3d5eff8b06e141a2c4684d5aee4454122d07eeb86b3852b770921ef9bb295ba0a371020aff24172eb438b95151b8c7215303cc2fda9556b0c3b6c14669f9a3da667edcb97cdfe5227fdcf8c69ca9f7f2f7c1f0f5ea6a4ffba;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc1f4ec14610635b8ccdcb47afbb880be9efecc4db7b46f5ec936f3cd91d2dcee8c0af13858de8685185080f02f11d5cb487a846301f7d6a5ebfd535f5ea3111e369a0700ba2d8e7361c2dc51c8fe03703120af0f8adb88b54d43cc62d68b690ad5bc;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdd9937c13627b769beb4294311a5c3edee0c93bb4856fd28c4a32b5f7cd72ab04177e086a73bcfb2fa3dc878dae5ab489f18190762fd983241da0b82682b3581a954623a63e35687dd9ec95d8f62ea5e8c64077c9e513c0db581a3b9ff72dd157249;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h439a1a1d8de72ea1ded22f05be09e6e23aa0fc8cb2ea07d9f36a85f0d28fc048a85b4c1cd61a380de32513ffb81adac2db95ae1830e082b61550802d6a2194f4085d17d9b6202fe0c70fd24d0930131571ff1bae4535519951b8a28b1d52123d99bf;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbe4b9737ffa8c3bbb69c97e8a6ee0dde71965a04b00d1612cf04a1d45930d3dd2907dd0f6b5bebb2a19cfbbd5ec39ea82da82e062e3b3c19002f5efbbe4b36d2877ddc69df05f50dcf005ff0ab52edb39f00491176c296b7210a287c0e942bfeb4f3;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3eecca6fc97ed4a82abcc16f2a742d4145890b3a9bfdebf67e99bf2f1161fc80c3d73eae5cbd61a75a40dd0bcd9e3af52f33aa3f27300a206668ef5f00b4f62b1a9af7ea19d41baccb3f9f76650e0fc5101e193e83ef50b6cd03b7b42d27a37d24f;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8d4074024c786aae08366292f77d047abbd2cf94d7e70d8a6a1e21dea85e765094fd70bfd446cdb798262b679c3192d1b1e11d5756c1c23f8f81f780ab9340cb08a72364c0aa49a827e3b8b3e59b5b394980a77c6d78fa01cc01ba13a8974f9694a;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h575c537621e18a3b05790913b6fb58f64f3a70a94ac488d50116a4ffd46265525821b7b235b19490ae6e28aa0870191c2d9a7525c6593d9457b5bbb1ccb88f3666edd167d676cd693a6cca70862ebb57ce6260620665d8d6cbab97e376cd8faf9f83;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3772348f334a21d9dd02f3ddaec39b9cc265eec0a99821401d7456f213d5dc02fd9544be6156cf4f8a88665f550298056ce959eca715d74ccb6227a59eb1105f64d25216cd33a4458073bc9f111623019d4971cc161504e37397059b683e2a3a2987;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h992b6187188cd815af92c7b25641f843e31f04c8afac19c094d5e165532a38c118d2acad201354cfb3ca1c3b00fa563fcdbf5047805a83b5974b8d9b814ab4126c19495e25fb339a09ccd592fafb2220f984e21e8a28f64a734df9c9436dcceaa8fa;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h27c6c69415ab55becab993dbd3184685c8cf3ad8420c90c97b2a6c5d700439d571294df225f3b74089328287d0277a45d4093d2edcd9647c73b977ba9c9341e40a25ef8ec308437a5dab09047535516e1ea6f7839680da6445b2610072da2166b43e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8505f900b997c29673e50216caec7e0804e0ecc6f6faf56a5994dd2f29128c51d97292b60d66bb2f5fb493d7029a618c3841f5526932d77aea41e43001f881054db259bfb69804871dd44f61d07b3e2fb4a97c061a3cf1d341cd4bc62e3f25b22b57;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd083d7599b16cd2b06e3b5263cbb8fe5449df5da760ea07021fdfe0eb1505263da427303351609341a926c7cb76fb497b762c663bdb900cf0ba78e675e8dff5de4531c28e84185f915257cfb015d200e3df450bb6264b75b205ba8f5f043ee7c352f;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hed4dadbaf5cb5ebb7401714016a6ae5adcfc07066396cbcebbde8b7b7ce9cb74983bb16d1c3672885855ccc9f71a03b3392cc5b130fe53e49821d72d0af71d89fd2c3b7590f733aab00cb94645b1983c00789bb37b0cfb0e1edb5485eecfdee039fa;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc4b25c19c42a8ec0e192d0476e12fb026e9a6df4cdae25ab3144c7c5dbd42d5e42f100f722e199bcc8e3f6de529d6594023511cffb9624a343886caf888ab02e164b0733cf1135ec47e8b65a6306fe4f84e3e795362e244eb8ea90376199529686f2;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hee4e0120c0fa1d760a10eebff46cddc7e0e8991157924d208ee926e94538c6f554b2af7bee1f402cb96afd8d9d46c6b838a8ef319107ec69fd11ceb98ef7089018bf8c9341df32efb17364166244a3f4826455768060e44610d8367395643378a26f;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9db214004ff4897920bd0a57c4b2440689b8f4f1df18996817b4cd3091d808250853b31c09af9b47d733e36e85ce8edf6369acdf6afae53cf4f89a9c081f4a408ba5fd3933ea5daa38a494dbb2fc36b558ba527fc527b351ffd7533845d69eb92565;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2f03077132a2fd32f9e2eaaf70c814efca0f03956c749b89ff165746f297b82da6d97e5a04c70048460d27d9e7a272f8591bb85b678dbb82d03eff294b34203f568b4011dbe6223fbfb771e4a465dfe8a7a1521b022d6a9fa4e899895a6f2364dd47;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h90e14223aec5c9a121d68fcbfa659ceaea08f98cfee2b6b8bad49b1f0ff43b57d4da29517a900ed1731c5fc0760df2237186a49a70385bd38613dbf061e532e02660b93faaec4a124e85c12be65ed42477a40668394aa5b099a67d1d7fcf0a08a60;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h60abb7d144a64c2b5f5f83bb2ee584278d028a5256625253fb093270608e4aa307678c5d49375751d49298ed080d4018fd4bbd9147c311b49b80ee69112427d38c63221e1dbebc456c04565871182a58d48755caad99362a23c03012b49c0d466fe4;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc81b70b5c97742c998df8715ef92185dbe5b82bb79515b36324636941466ec212e5824f00e91b51dbedfae60beb930d96fd78682867e8ea543754e39308c6876f2b10875904f145ab50c187176e033f4aa8e0c33377cd167e1ec1dcadd701ec58a48;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha9385142e847c4dd01854d657968a62c5e7f0f74ea1c7b6a1556e47b218734b3f8edc784503ff7ddbd0d2583cb77f97b986d1eda36c790b7bf2f68cbfc8ac38025c353a4f90ca76c1cd120ac4533d1278a371293873a3dccd4d5b72cef17e2666e39;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9e281a33b2abfd1a1a14b06479c2d7d322c24ad687e45f40a91384c9cd3037d18f7b318f6def004bb75f77c20562d9d56c47865e312c0a68010d28fa5d452a46df87e5805b61091ce0b426b5f7e0f9a88bed617bad8864fff0b857152407940b3324;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h402c1e23e280033f1758252a6eb7dfaa7d0364045cab292b9849e0538256722e680f6c940f30f62f59ea3d269919feeea72d20142cd5d54f7ba25b3855efb92815f225a5d56e34e4e6b778e38fe2ce899c2d01df2202132c846b3dd710d0a050aaea;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2c4b74ad5f1aa9519fa36c55b959dad2cad3e74c91715fc22287c73f1c750e094fae47343cb3b9cc55e00a5764a2d97abf9e12a4d1cb45fde499552fa42bb7596512804d80630e7d2736dd87f527803ed5d9717185cd657bc5cdec9c6083af1f48b4;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdfca5bd727dcb0419a83d2417dc704edb66fb4056d1014eecc5796bdee91115cc473f6ddf6bb21a836435c1c8218d36af99efa76a73063d38136edd87021329fb4fda17be4d6f72d5bdca1028cb97344e6fec7382513a9effd6305c9f055228137bb;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb93aa5d43789b8b7a25bcdf1be57e90bc879820b065378cb09e87f515303af8efdd935d0b4e5681604d3bbd874f972039f66dd658ea1f5cc7d8a33c14a1ee74a257370cdd9221120455c0ad41831f8d1b1d434a8878d80832c049fa89c5bdd26b58b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h38c66ebd32360c89adf1fe56a1d9267af7d69bb13a75be4098039f0de49d30d0a705c8b1bd85ce655ed412e5273f6b4b959451564f8eeabad2ca5a5ceb12468bc29ec25d98f60bae2e4b4e2e5607f8b96440f8a135c7d9a57b635fae95f3d92b18cc;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he9db9e520b4d2bf80af72b1b5a85ca16e2a5aeb5bc63ee3df80d7be31d0f76cf12917cf0d1a5a8f875aa62594b245851ade84f730061d9f98e131815ce5a09556190fdbedb48aa831b94654393c668eb500ece7e255e486a48144f066ec738ee897a;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd3a68eb4730f33d4837e18e6c869acc4a552a5dac709a0202c8da455a7261684c34960db8b88968a72b21672db314b5cf97d298485ce3ceba6dfda6f0c63577f293829c630cffb00c900dcdd974a0784f2db252f7e1fd56460bf9c33f60b4e10f343;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf77e174ced75f33cad3247c00c908aef8debed1d6a7693e6dc14591ffedc4065399ca04262c16bad40b14251d79fbe196c3fad49357650a8b1281120e79b99c59b6d9028c166ad61f06d1954e72d726d75ce9efbe32c8e37f6d9823a4cf11d5b358a;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9a3221f018f471124c2c3b79f36df2e9ad40ba48dec1c37570ad09d42e259dc2a50e59c28fb5ae208874feb919351e04d0b3e1fe9fd8f70e6905d28dfc37f72a68a83edbfc3a87fdfc7e185eaef2b635a3b2fb68191cb8c9a1a73ca1e68347edad8d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3a62d4279392b7b6c5c3462d8977bf031025a2b4b691728b07be26ed945cdd653b0ae467ea7eac17764b16ab238d27c9318e14c9610c75893d3aface0884aec03a83c780fa652df60c82d369b69debddbf1744bd2fe0d1a0d9539da210d1677e54a2;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h75432278efdbd08fdb81f9c0d5100cdfbd88f287c23cfee0a6cfc97e6e706b2af61aa1df95553b5397ae128e6f098afbfa4c86c3e8be25ca367bc4a5fba8fadd8d7d84b98465da2a5635a65b769ffb69c0d0e7ee72030ebfe28c620bc7b5f2fd1cc4;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5cfdcdc77ebd3d94b21dfc10e7ce3973c24a088d06c747212f461c2cd1c9363f2802b3959427c17b67929e36a105512d1bb88f80314facdbabbdbd2c81dbe16479c9b5839afe5b2a34563fa151ac0dbc414fa60bcddadb4cbcb7dc4d99f9689ce1b0;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he7f158a7c7e1d32e476b9e55ef0f9c6fb754f847ac127ff8f6487668227623ff3723db1a9eeec53f45b5e952bfea367111c74624742c2f8956b4b03fe8a8f0d707ad2ad6938d8b26104ad65885ddf72c0a1e17bd34359b837bafedd7891c5be04b5d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h95871c65c6cd4ef7c5fa060d075f23c56c30f978ddf6c02a350f8754232bf41e686388483353906b56cd4cab795fba0f743dfda9094365a6a6cc307b34c11815f7cdb48e5a530b2e9d3ac485fcbbf9edaa789cc17a99502264426618dee56492ab02;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd58e60b58fb2a922b76974bc9de180c877a3f426d6bdbb655a971da6ed3e4517dd3ef95761191499ef1a196780ac4206e9ef878281f4dd47914b94a39cf1cd20dade14b1770fc7f173bea53eb612bbdbb93cdf330ec7019085e7c29c74c4d8c4f447;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb8591cebaebae7e03dc75f7927d2c43bb1568304962debd720cc2b35052d6eb5df869c2a036b048f04a75d83adfe193a40f3553b7219bd79f2e799d366ac7e44fac06807f60c66e3ac3d5f75b6153e89c911d68dd6968a4a64322dd330f200695a46;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h423b0c8e3f47c4964be24793154f6c82d3dda2fbc681ae98a4217263eb018813e58c557b9e60027d14d6fc901951329c7d6a81ab71600b24df71dca43050f1a097f7c1b0f64ea84c9a1e22826098b643123512a7baed27dc51b8e49ee7dedae7da35;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3fc660223dcea00fad3c555eab9e0bee358b8f3e83df357b2bc4c91936bad0feb51affa0cf0387443c80b50a612c9787695e67b3c2e245eb2d752538120c678c2a8c154e9df4016e8dfcad9d5ccd1db446c5dd7fd804f22c30ee2aa3c2a6b61ccb71;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9dca537ba7f02eeadefc68fb1df44a2608e284b81c7e81f8c60226d525ee0c5a7f60f8f234d2be77a4e9e2248474777a1b695f3a39dc6d6c3c0a5a5165416442acb7ba2ab434b750250971d1c798ae56890659b1adf9e5f8e462460b14ab86c54b32;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h430e38285fa55f8ebe7b4a8ba6622d3b31339ce765715e0eb3b8cbbe79a06e464a1d3200bf6c969fac0bb9552a0e60bd5a15189383a50ae4925f5284e97b62b39d1688185221358dfe3b8b2c4f64358e9e59a63a278a3783ffa67acff9ea0453ba0c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc891d250c40fd1ce0a013c1d1932dc8a8710b0334e7eeec0a1bf2ccae8513894788bcb01808971966bdaa072bc086505d6f0de0bd43b6ce672ca6b801f4acc52bcaddd80be7c0791436e4ef4a86290cedb2f550a07e53a8250f7fd2606000f30f93f;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1416b402ea1087c15f101e6f6a986ae50cfd166cb1369f0265c886cf08c4789378de0b0441c793ad441d117d94d7e434b4826e03eea47d3d494aab469562bd289c1063eb159069151f0e08c24a0da00a91a0191ddb9506ca191e58a0df8fcc27ceea;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h83f966ab7e14acb9086f916ac9d002418e82198ef5d9923192165b6d5d3663ed9a72552ac89c11022aeabb6c4a3f90e361e5d86d09357651427d61c99c1a11b8ddcc98ac0c57fb4115dd4372890a3f37e963b8d4361a69137094bed0c46335e5b397;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6b5e658c8b7d81f1531e6a003186b6eeae0d0a0f146ac6867a09661021522c2048acea48b2dc52f450031dae57fc97a5e8a175f2b0e2423e137de843a6d05fb77af2da555bdcc3549f18b61cacaf9546e08187b6696070221d315bd7d43fd0bc429a;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6c7524c734a14e3a58f82e28f28a67aadf7ba43415fe2e559488e4d793f26d89b78636ed2e8c28e3b810b5bb5117e5d93cc77e328f6040d1cccaafc05d087f1934efd50c96edcb40a7f73fd8d2b85cb91603e6fc98fd449ca26ee068afb8dca3655b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6cac33223647ae91cc8b8d1e045d00290d4df13293019e28110a770febffc096d6bbe772b7f829f33739a7a28807840d8883949f8a8574301a5449bea57c9850d6a27330385e132119b25ec7247019c5b235f1c6302e087254e4113e0e524350c7c8;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h65d0dee2d1ac2ef1763530e4e182e313741cab8b7f519399cc3ada139034886fb397624906f40a712fb79646883fdd9f380ac98b6e0ed19a5e0886f1206fdaa9d31182ca5b97573deac3aeebf4b51f497e3bf3bbbc191d2e8f6f99bc358240afcbe3;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h896fa4670010e69f9f5b5a77b1deaa99b1c62e3c750954c7fcb4affaf07d992d11400bc49af90de6358ddf93745c5d41f807ef6fb83f93fc4c44be2d3ea757e620db008cbc25a65c720caf31c684eafbf6546f3391284a35e0e2e1e49268c90910c7;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1141bd0bc749a9ca67b92ea52eaf48f696308b94880aa47df0508bdb6d5e0712acce8524bb1c5a979b41db2e33bd8a9fa4b23634b5695541b955d238b717ea728cf0670b5704c97de5b7e84ac99fddf2cbf7c222aabd12ab3f5a80c05079c5be6bdf;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h751f0ceac98b32ca0e8651a8c4e6b3a6b7365f195ec173e6e8e83e48428a08aacaa880d7ad1fb58c5ea7a65733f7ce3bf5b1a6a2b5370035a87ad8f8dbe38494d99fa074cd91df084ad1ed5e11849734ff0eacd14592875c6e5311fd91eef7bce3b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8ec7c1664c5217b97129c22787165ebeb7c2544c484e3b4ad5dde3fb85b16a72b25983f35e4c82def0448972d9b3f7087816a73ddda83c0d0ffd591d533db1736fe32e3921c6b5586949fa34f2d8b5a057838660fc7a2414831d3c844b349716fa58;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h32410a2cb29f9063a655fd1383b3d4518a05aabb4336d5cd45859f9212093fdb73603d57eee0f77c80b374d9f8a623b06b410bfdf165c0fb22ca7ddd363510ba3d6d1937db6b61691d1fe42dea8f4e3db91a1e9a9bb4792d8d1c98e9ac2957da1b41;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6beb7562cc72292cdf6483d6a773dded68934b04751cb6c46ab09691bd625183c5d86ee88aaa3182b84edb38006c267870cc2118a5e9351a6c2aa97a8e115aea62df498efbb326ed5046df03c45dd359d9a107e6388244b6eb567f0e4efa0e246aea;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h349deeadb09d97d0cf045d5223e497d051b4448c4ddbc26f635cb9cef735f3e7ec75b0b682aa3c100cd9ecb53fc5a080d8d9a01dff50572c0c5b6fb715ee323255f77fccbe5a12ce29a5c3dda8f8e4aeb87d63ac89ea11a148097ebc493be894946b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3f489f914de117b6eb764953962da1161936c8d60696bd09a2c5f899d679968f6f279e7618a5ae640c7deecfbb1d081b53e4f10516390ab45cf0db5292a9f4242ab9b877a18d1c14072c4caa4e4103e7c2be60765a53dbd0506b221a9abfe85cfd95;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h61b2c2e2f73788c3b5791e1022934ffa57707d4eabf4c7716111a6f05b3db39ddc5f52a6d8d26d16e57360b2be113de4125230ff08f6dccd6d9d738e27c3c51d9c326101e0ed1a297f50ac2da4b4bd84ba9067c79b7662f500e28bcd28d9a971e7fe;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1f46bc4791a47791bc38f49ee44e5ff2ba32acedadba5ba0c44b708e7d5e9666b87cdc594f83622a4c100f46e105365d1328fba651f0402f58ea17ab6d73ba7f30642d5ee02c291983f3adc2063fb3b13b6223c215aefb50d1fce2faad27d648c369;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3f27085e6ae27fc08e86d9773a97ae02b59ecb4a80abac8b155beb2dab366a24b3d0e0521e1cc13ed67b538bd0c939b6e31f2de3a8f7da321095129d9531bc10d9df899c72c61181438f127850cc3bd5285a46ba2a2d95c904c14b897a95dd382955;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9eadbf531829fe3e0ddc14fb661f35a3427bee35ce4eb7c7e619aeeac50e1527a66f344f1157c6b22a69bebdb82960f2784322e0779076228eba4b30566764baee3e4bd15188e778d8d652f155fcffb8725c15e07521eafcdf36ed8ab0ac5ec03f26;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc859f9d44234a14727f4e0d191582b1ea16930d133dad85c6dd3696dfae721c16be7c68f658011ce9971cf8b168049fdd1e4843f572703ae920298da982654ddc87de4ed819f325da00bdebdefe1589dd11d84e95f41175092e7dfeadf1e666f8cf4;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc24fd4879c751c0057d339619b6ed4d929ef978daba8dca810c52c9c834691a3c9bc8f87d117b0995f59800fb9464ed9308dcbaf35df4a2eff304d510dacc3d24a4e36617f9732c3d83dbad75c34cce8782f8ce069454dc0a35568561f9c6effdde9;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4d2216e9ac0ba7b66154d454fb468181df300a9b6cb3e769aeee96cdfd4317f24e13721fa27cc803a32a3c575131ab7db7e5b921863d248a4694f9e5cf5bbf4eb1fe6e3b03d78766ca5f1f463e10c3564df8af97d3d7462c5bcc738d7ed35c6e92c2;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha8a17832eaf705fc8ff57bdb20b93c626f53f33c4c74045e1e0ecff1a11fc16bf2910524ece19048014f062838b3d00606c33b526e480d8476d271b149aad99cbfd9802b9f776c636ffc7a693eaef51ddf010ebfdb0bfefde7d59f767f5ea7e5d549;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb36ac3f7d1d836d94c2444a02237f6e95ae8c11cfe457a733bf20be46cce3788193306371c1f11e8d7c26088d884e81f72077b85790bc1afd6d0d189b176efa6641517eaf81a6ed90afaed60b1300881bb851a05393a9de8a7e0886c8c2f8f4c952d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5aa1a29e2d587ceefe126665b06711a4c23b10dbe66545947834758daead454487ecf1eb66ba8369b662bb93a61c78782fc90b06b0eb62d0f5b93d1388ecdc7f559b8788e1c1e943dc89e34d0807089b957ac1b669d68118a6d422b8f6ee6a29f650;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb067698773097252f1bd82d4e2c1c8d2b3c926792b0d39a98573f0b3d975c5b8911de66e5e38158ceef9d89cb5d0d8ae25e5d9c014777440609c37a59d27a02ef2745dbc620e2ce541adfe0e158ffa2d9f44e0b4b6d19a718b813f52b0c7af542c0f;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h28eed9da284339f8b1418677e1f693a2eb828aa07cb07200cd46afe05de10ffa977db59ce1d8632681aa40613f511a491833bbf355463161853421b195485f3cadaf06d9f4e8479eb18a2d5c7302223044e884e9d7d4915aec068c03aacbda63bde7;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h569044c4a57a45fcd980ddde59526e6411408f11108e976884b32c553af1ba9e37187398da63fe7b788c109c466ac5b97cd3eb70ca4159139b01426a48b8810a5b17ac61de502056ea35e42c7ecbd9fccb450734824cfbb8d15c61974728be98c1c9;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb56f844fa0f8a2b8f8a62f2b328641aa8ee01026c83c439407f34dc6883997f69a2a5357383a834a69c7cb380fd9d34475b8d2fa1abdbe99c346bba294652d434b8200b20a9d08381051580909e6769a555117aaf4886a82bae6bd5447c0a93ddb92;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9cca8aafa098b28104eb80771054f7de2401b4688a20f4f159afde027b092ae9fd930fc613be1fc82197be1524a52abe3c26ed35f88f063ee19401d5939abf79a07e5ab9433f9c4a23f3ce60b617980cfc423e1d43e93e17dc5130932ae8d46debaa;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7c895c5431e34f4ac67b34e90693c6bb7ac56b6d9c2e2cc93487d677374247575933910f320a0a8a31804ef6f7f78b62214e311f8315329429aa9c13172b70ffb4ae7a824cae6579d73ce34a963efdc0685ac2ad6458824068948d78400c7881128f;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7232cfb940f23fe89873483b5fe1f05415734d1dbc8e66ed4e71a5d64febfdd8eea8f2049cdb3f33897e7d5ffbcf570c15443129ee642e80bc3f3fbb8d241e63a2ec0bbc502f2ad179583283d3b9b341014db7f481df86d1e09213cfec2cd876b8b8;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3f9127bb9f32bd462f0f3188e944ed8cc6f71a5e51c283188b9c20240824800cf2b1f1fba33d379c14cf13f785f1294fa7a8c13ca56eabef02307cfb64db72dc6a8434379394d63df806fddc35e32930b8aaa3bffd42d043718509b4b5a9160ab1de;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h50901ed67db45611fadc9685383551dec242b7bc4c9f67b8871f014a67161e001909c09c277a904c4b4f585f34bae66075fa2aae91a413a786fb6dc49b68e4a26755911731edc185768294165793f60d8abb896da3924a9719fccd31b9a6668f6e66;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2407c7823d58e221fa50e1b2a65f81daa72f05fc8c7b8940eae2a33d0f7a4748881a8268f95d3d717d6937a12cd6213ee8f6f68e1cf6c74e13c1752736c857e489474c49c2f550d63de0a319280b8ea37a1d4cabb2ef4da83bec66d04fbb434235a1;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h413229b08bd7efe39de372d0d5c05ddef231767700ad6629c8b147e6853ef01d04302c78eb7e12fe20d498b9dad417b9d59fd4b9c7381b0f5f1fcdb874e0c36f352edeade69868d81ef4135e0a0b60415a44ca69921671817266fb9022f8e850e857;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2645204f2b1ccf8de0c11256ab44dc4ef6a4e6cf007f816e4d9c5bb1becd8a01cf47edec7a7a9404ea0b26d2f4fdb241c0e2d77fd5ec3a62f6b0b40664c7d02e7db042ea2142c084101e703c602abc297ddbb25af665e86af19262c92071059b2c4;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9da2af53412d2900ed78d816084af16fba7ea9b0311ec9ae5b4b481dc0b384800e94285f55947c50c0213166df7f5707708f68936241c464f706d87c7222a259acfa47901def8793069ea4563544d7350cf1bfaa086acd6fda30b56ea2f463767161;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4d28501e16e3ca14a0052bcf7f1a919e19506e91db81bcbfc6ad7f96a76efc6d422ddd66172882b250e6e9cd4ec985a9fb9f23bd97b627d3ab27d1795bdfee88fdf0d6a5e7313ac2ff1db72bb2c921f1408bd8cd20bb20b9a44e45054ff857460957;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hce4ff742473322d8f77fbdf538037fb76c71c3923fde22a6b90ae95151e0738a4ed8a3070b984fee6a51a9efdee0c625a1deb6f01b50c4b9145c0c69d3948c69e4d0bd54ee668a2fe7c97a4775ee6314031e74e377d8cf5f892df4b8d540067fbd2a;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hae98af9ff22c3e4c8b51017530ff578c9de39531b5b760f4c3e9164695e3c54973c77a764e2b775cfa2acd2ecc201c0433fd9507200e850feba5205d5fef123856eeb527c990f1c7e9b4bb18e24c45d2f51071bc006b2bdce22532b1d81684ea1c64;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5336631a7025f542e84bdc578e47d677fbda6c71abd902633b07d54e48063ab9969fc7347c8bd01dbc2a72d23a46199ff085d1175a1f4b1aff31507b9153e70a394d92013c218b32149c8c8602f4a9dda8163e5f46b8aae2f530aff7b3274499c962;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2458c57f0aa4a1c7286145c6ffafd21d2ad801c0756fa3f288bf9d4a0c50b9f98caef28c09ffc27ea2d09935d7394856e1d7c86dea764dc4b1681c5393ec714e4bf00a6cf9069508bdbd365d33989f77740cceacd62d3669a74022f3bf5deb687521;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h31e43e241cce9be1c2cf1bf3f6773784bdedff7668b3635959554d33d14b9697e663a6133042c3aa091d4fe2c338b721fe5569c97fa8e929c461ed93d9e7086a038032c9a9633548eb08af5308223f4c7d0a2bb8002a1a71e7c4670c3e62cf984d58;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc8ac6057ac71444bc30668dc01ba5f8829b6bd6ea601253338b08fc47cddbfd031efb9815b2a1c5efc59801665e29f2dfb5492fe6fdd8cc6ada430b5c5b8cea8c33d2b41379f7b0106952fa3b06388ff711ce2eb5a7b8c80cc2365c4e40ce80e1cbe;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h10a623bfc25e4545035016418267cad217dda086b218d984dfd8d9805f883823ea057d805dfb985bab5d59a8eabc4b143f6844fd3726649170885ad35bf0fee30fe3949ba8cb7f3c878a39b249c9ff9cc7630b4e5f745aa2d0fbdf6118f46acaa1ce;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9d0b80b96d34f3950e6f3047278c4578d21d438b66857ee9a135ee4afc257a281d48e8d9adccdfaec1d113316cc2bb11f561447fa226a385e023c726e5c9ad8aadba7351e3f5e69358b1486970bafa366b97edcecc37cf2d233bcd891d74de5157ca;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hcc9de6a4cdcd8efa25568e2e2422eb1507a538904947a1fa49be1714caee9686d1e89b942e7c234a008722cea99a98176c942c9150f57948dfdd39729e4c8506ea92e0240ffe7eddc2c7fd1acb7618e26e2aecb719308691d0587f1c4fe0b82a15f2;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he7d733dcbf2a413db75ffad9d5329a87b7ee7ac27f31655a241e74c12af966ddc40be38c6cb221e35c3c4092ea5d4705514538e61e76fd321b96a025969e4548d2cf2a69120d32d071f650dab3b770688d50658c7e391d25594653e4646d798e250d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h500f72ce553633be074d48e9c21063224545175ca5b144221e08fd67d9e1acc85ce056ba9290eeee44f3ee20bd8c73fc1b64964a2d1edaf3770259195d5e8ac73d7db35932ae09ebb2354ad3292b92cae8097dbbd2211f0dc1bf27093bd32478d858;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h433019f0e021078f64fd734e14e95f2b3db8d1b165b505e10fc27d08bd365e17e767dc7d6e68241be1a1e4491e2ba564313cb854c4fbd6a9ff4e0d80c6374c8e13be11ae3ca158e52323bb284b50325ba3760d90f77893cdb92bd672bbfbf76b3716;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1303bd0fa31a40ea136b8e6150e5590d68a811adc84caa4e9c8a8f3586bdf2598ec2a3b9281844bd9a4cdb8dfb2b35bc8567664186c5aaa86e3c65502c0c60224172624298f5fcbf63cd24bbfd8eba037d8e299c6ec0fb1638389e743f0c62ced256;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd06e2a581aca49ec8434733fc2c380683a12f18ee44b96a444cde6d7f9cb2be378afb642f8a01c97f666ac013bdbc78fb054365c7f09079816f08a38b4004fd1a5e79c60b50b5d115798a24de44c71d5b1895e7288c32c08df57b5dbab18e360bb53;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5c80cfce1c3111529630b81a0009b58c3e421ede784d81f5457dca40eeb411a8c19c889e02fe90191fd4c2476e9b0e6439e16c078c6423ae310ff8e92fe330990da55518368a8be67bdbf0b0f81dbf7cb0c824da1fd4e6e5bc3a537f29f14755d94d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h37e2618aeb02aa83b9ae990db4d63f691a7470005043a811a0c7571dd9db89ade68a80643691da389977c6034fad562d608d03dbc2c6e9a80f3fcb450474a0033bf6d48d434855db6626176cca16f647915d7a6b8b6c59542b1d2235ee41bbc8001b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6a306853d964f186bd3b1d4eb65899076185a784f7f1e1f01fa28461aaa68e5f2e156e27f5965bc692af19d92b330cd712e3a9bd85cfec0e31ec92a79d1f22394c2c6e7ed22420594576b5768f3e3fbd37452f258460cb14aabd1de4d03ee92f52b3;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h79948b037e8dd3775cd99db8fa6620b53426024a01c3f8f469946e1bd13c986ffeb0cd270248ad4c03df57338f1c9853d2a268f0ecfce28f5b77ba864badd004faafe9b667e6b4124d17d4173950c4b66a52701984307f8a6650c9d6c45440b66108;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h99d2388c7d24b1972cf29d5840871fae21d3fa2d20c7e0cd2a3ad78065ff604f54f721cc3061938affbd1ba5c4f2ffc42ad8c9a7e236d769fa31dd6f4daa1a0ff164929718a703f141e30ef167bebb76db970aada848cc067b0d9b6e46cf4cd275df;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc44b2ac5ee8a976684a9820c328b5cb90864266994ee4508195e5a4ef62243fcd44a984b251d1aa9da9a79c4d0d6e10d49ecc0cc314dad5ba64220cd90b5f9327e1e15670b965d70a96b53eed4f2afb12f42afde0f58efda2cbce6b64a0331d0d68d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1114fc7945577e73e85b0eb0d9f0344982485e70fe6ae005553600e010e3df0e8c173d74a403849557a9c9d94706c57c59eecea27dc3167c622343e7edad785b00fe2061887bd3021a4570f042b58b899d750df853a381712be83c88030720431c6d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3245b9815c7c7ce21d81a53e494f936eb03ba07d198d1cbc993db0d40b80773bc87236314693ee769c901922358405101f112d8417fd18e58e6a7d9600eeba5dcfae6241c959009730cd27f40da6efa360ebb68034c076fbae15f4c43d8131b9ab75;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc07adc84869439a7495df6f6dbe10d748d146102dd1cd206c2f772f1b6e9a6e38bd888b6fd774a20c92a99bc1bcd4fb10c17984c229751be24b38199548841f7922f7f815f59f8aac2a13f85891acbbfc8772780f524f41c6444b6f2c35ae58b3a65;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4d64f5abe38b1fd3664ef9c06e7c946ccb873e19d304e96a1fa5eda47eb5207d1d819d1d050a774db64114cd71e6ecf1b4b951d0ba0b432697d13d4ee322c79b6dbd0edcfccae13dc167840ccd9482716d937b6915e377321bb024415a16579588e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha022be8eb45b38014150f4b01424fde841ffa40ca9922c9b56a3e85755bd60bd1df7a0ca117bc637808c14976207204ab064323b16b1dc03b13c0c148adb9a71b362bada20b40eb854c1a4b0c156fb55765ae372c198851529a31503c715cf360eb1;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha6c6aa7695dbf996f173ac6f159b75c620b826244194ca048732dea38eb6a08602d6d7f389e68d1c72ae9bd9c843229747491bed878f32bf63ec6e2b2c85f9a2144dcc48f1591a5875420facaed2268ab45cf179881e96590750124cfeb01a1ea52;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8300354db9136b370b37bc13a5c02ac85cf1f357679a3019a42b21eb2d1c22c83edef5314769a200df1cead1a19a20d98ba96a30df0c487178b5a18884e0a260f253027ac75699437da74a87044792299d865eb96d93e7ec1d0fa0749791b41f998b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h987a40a5e157b068ac1619dec8e539ae360e495469a0d484fd2ee0576ab5189d21529ea73b995c9ee0cfe52325665ab8fc43c89214332cc68598651bc2256aaaa7238b49002d5492069116d459fc7a8c6f831259a7a0489b1996afe642110745536a;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hee9f8c19d50b6d64406947c7e99589c1645ec23a29657dbb11fd2a68e3770773a88c738cc9d12102794c29301ec72e11f0780ef9d81c55c6147f7d95bb13af64e29394f5240196b9b03d547c4593fca4e4961d0594c8d4d695779bb8c3c6e450c5cf;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4f176e7e3642bf635299e704e31f53cc980e9b07525f76f3e163a3909f716fa8325737a9b431322d1a6b86da18679dfe7e8d644ecbc1151796fc108cdf045576e0bffa60a04fb5609a55f345eaf8b2e324151d9b7966ca62929266ac9655c9e39981;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h966a1d5ad850de3119d88ddcb50da861bf7f3352f6ce581bb95f52fd15ab17dfc0a4ac2ee8cf8df779abadbef1a370b8e02077102db3654d6626357b8a63a27308ca74836d1b805570c799bd1f486cd6156f6971938e741725e19ab4071c602153c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h884ea48255df379a8f50a4305816eb94205b9c37f6a558ceb8c88ae749ca32871bc275c874ef3153c4a0260d00eedc57b4fdbcf5b9e0c4f2051d7c31a1e043ca4c9fe7f8d829174f81f45decacef2de0558a16fb896760fc5031d63270a25096602e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hce815cc1613e939e30e443003f027f0964d9895db340b76297f26b972012bf9b8ce160b0c01ce2ec6a864609823982e35abe2b56c356d107766c7b1e52b8eeb37b0f04a47030f46bcd2e4583374ac11e8cb61c8bec349b355c9f4c089819a371f54e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdf853704689d306ae8ea206d7b05af91858db002766c6a539c5cbbb281aa234d2a9176ff2fd483a2e4f37db3474ad857a49cac1cf2e0c91d8a7a43febd7cb1c63caba376378a124f5e57e9ba218b82e4582fe7e42f4ddbb4fc69d04b9b2d0654693c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h39a622928e1c8698b5117e8cab733f7ca021f1929ef8d6b5f37193f656a9d1b25eb91d64834c1498c06da0d9f7a48012a97b1c381e4a7fbbc8b249dd4464b16755ef62ed447a05557782b9fa7f9e8cafc29b379528bd01908d3fbb21bc33c2258aa9;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h139d65a276278d40eeb0edd6011bfdb2066bcf6776b82f7dd62d874e0114f70fb4c8d08a4950b9e78c64b7b5d9e64f0780b8d5b91d43ca7fa244020871f7cba3ec5132ef0559dcd959d93f1c5854ed3c4ac540307c17a8a0361d7e41de8f0e4df30f;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h61e163bb3f08abce2d70af848b0aeaeba671835a9becdc5caa1223b294d4ef8d5315b717b4e3b01675a631367c63273326680a85b5cfeb793bc69d66f69f5fcf29d9b8de397263731352962cc91c99b7db01b0b11ac3cfa84bff57dca557b0f3b5ed;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6d843d5391355c5eceaad6a3034742c473ece305eab8717ece8def2d9dcb73abdc564e55f8cfa1cbb6473852c7c7269d237e37889a1d42332e3bb03001bce77602a24151a270b37d745d36f65390201c2c0c419835296ad333a0fed9c74cf48c814f;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hcf73407d9bc27596a5377cdf3331121212f442e016dbcba03512371285a7118c40ba199712a7b5dd831c0ca8c2128fd0194570dc26309f0ed6403d77be271780d286f14c449cd9298cfde5d315cb84b1c36953d5d4e16e2b5c8fb3ee53fcfa9c80b7;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h51471a7e3cb1500226041dd5ff00a6ac8c2c895a6ed4af076f6ca87948857ba8a0d45a313b827d098fe7163d9d7c29ce2b9f6a2cf42b3d61266befe073a14bf0f8f019320f1e35573299bad0a2ad597e9dafb79a86024bd619a8461d0df45a6b7b6a;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hab5ec29a7667ed795039f33734a3ed65c74d01db542471889a19214faaecbcaf613079d26d76fe5a4fbfa4c35f283c3cd747fc48cb916553d63f4df0b0d78969f44099868e2b2026880c9ed576440ee08005c6a06f79f2f5f2f3452dd03a52f38577;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h203b5cf94300035f310101d6e5a9cea64f710492625ba286878eefaabc260e689a5669b685905814b8d56d2341c2f3ac90e1a015690df7cfbe8a11cd891468f32f343d06e6e8bb62aa258e07510c3afdf31fda955943f995535c132c961d840fae6c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8eb7efa1f3c709aa71477ed66196ce2f0d03d1664c940ebba326817dcc015f191ad29aa2f995ca655db1108cad9a1b3e0e6178f8d314a31b79628cde2c7c77fdb447277fd1a6db75ee1716fc1560a84f99631538b81b0cd16258cfdab09cb6383b0e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8d8c9e08e30cf8b65a549e021879628a16100608096f9ce4eef872c19dc71e451989a439037b0536e2b2d70c03d7ac9204a66af3002f20b72eb0725ea31748dc7b3b1dac052e46b5de0d5b38f54fac3035621a2f7cfa1087d1c17587616e2bdff10d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4d7fb9cdf4a72b26ce16994e4ffeb920d63a63e0f7fad04ea987ee4c821af68ec65d1513918e84737ea7ed2db41dae75de40af3f1fa8d9225dadd43569c31db4e0c5879b16a6f1107690971c6c56e6345edb9aefc229340224616ba4c1a4a80336d8;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf230e12af5cf673e59c91680e59f6663e53ea553c47fedecbe435360bde2d1f9c5b75aaf69b384e4867bb5fd4ed6d2845bf2c348c94832b7cbbdb2bc4dc90e67284cff3bba79011cb00af418d8f999509104f2b998da5b7c8efc48f6a29988735f66;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb1a7b66dde2848195a29b6c58b1e7a93b11471dc28aa50560603d75964057216936412180854c3f6f12a7e9a233f90c8b3c63f1b6c059cda821e337910ad9c8a53d55725f4a19eb52120b43e5c9ab196eb67cac4fc88abec9d03990449e1ca4b36d4;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbe355cfd2fad19604dbce80ff1c35f99e4000793080d27ce29807be45a584234bc11e6920d39897a57ab50999fa9bbf5d2a2b68f896acfa78d272fd77f728cc1c9adf6d78c77d5013dcec703f8d87e9a9ecc4d28bc7bbde0bea24e638a9a00f7f88e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb0571c033ea888e64704dc5be72e98de2deb2bcefbcf0f31269728508fc364f9bc0e84c539329bd45ad3aac84e8fdf44ed6c907749443196151f26b0bcdbcf3768dca26e78691619f5457b1980b61fd71f9a52726913abfc44d8dffc3c337b455e54;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he5169172561c1de2e5744c52d2e53b210df2efc5f218f056e722b13929786893eb4c0b5b4672c4ace4da1908b4c8404e11c04a7e4c1f321da76c11beece15f8bf245b9b0772e916c2182e55558100d837c821cf45ff5b35026c9f6380d9850129a3a;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3d5f65c15c63e136176689aa85b1733cd6bed93d473273a07df5322cbcbbc8edebda37f4bc163445c303a7d4ee7d29be7e43d7d2a30e577eb65326ccbcf051978890c81ac13e17ae6a1e91507cbbbb9af63cc95760b5b1d53e691c9466562c0fe383;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc9b70b2c525242dd1f67329df7fc10a52240ddb4ced784fd0e6aea688b400cd4e5509113adbbaca26678dfa541d558ff1e2aee543039a785f05faed85d39e430ec1a6ed1d85ea5a69ff735bae1ec637aa4e334cf9fa1c83289b03430dc486b580bb2;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hcc13f997d209e5e35b2ce5a39361a0a066e9886623ac6e12e4646d87c014ee0858d3b2a1c56d3e5c41e799ab465e398f196bd002268e8217a238bae315f080b3ed0a177210cc745cd14df9f4eef7a4a5d660395ecb91124cabbd32cc91527bfc2e99;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf3b3f2d190972f37ad827c0f118a48d78adb2ccdffedf858256d077e8af847d0543800e463c19b5b22e1370a3321bff8ad34d534b3fe773d91f42e9bd289e3496190fd0e1fd557ae429c6fc87d6a39302494d6297b4c2f05e94d3920e51bac43032c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5e778224a60c17e7134547eb6bc68c5ed9b37a7c52b58342f414b7a719dfcde8fc917828e0d1cdec400b7825838dfdae44ae862a20049e7eaab43928813f3ad74f54ce879a1369c5b53348d60f5dbd0cbdbda5a38ade1c0edb1f3d39a58e0f25a77a;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd09f98e08c374b2e7392f65b0db8b953783f6e002761efa621f89445a5e259f4d035ef827695b06d14b7a8350850437d86372461c6eb5b22bf10ba3af4535f80e036f13c1e6e70587433dd2414861271cb9c0e70e6f83689c06baba555c14118d13f;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb597c1146d6658287d24c83108bd5fab908844296ce2a18d90bfaef16664ef5e3f815072566fc06a382e6116889ed62fbbcd2bf0c299dbc3856ec0828be12fdd6b61f5a35030afcd5a886d99a8b1b7e9eb4912efd3eb5e486605c972da488bc679c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8499b323cb166de28c6c90547300c3be9718138f8dc3085f129763a02789ccc8b5c4d9027c8480bcfba2a62ee025e46cbf81e15b07cd791ac5383f22aa607a825451d0b4be30b5608a02bc13070ff68c04e98a75e3c25c55d194370cb5d97a276765;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5dcc6de98dae7744ca81d1c07fe4776430bc021c9fa7fca3605fb1f6bfbf21d49bacad140366a8ad51e129dabf30a79270c1c64e2af7c7803f932c75dbe2657fd04737ff11772b819c563789df91343d2358d7ca49a2511583fcac2a025605b599ed;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3ffb6cf6db8a898f897272f5400c1fe9903cfbf1b1d19d2b5ada6fde8ce53714ecab83722be13a635289341bf01c7b93575ea14e3dcb7ff9ded28c49e012bd0a88ba23514cab9cc1cf8bd3da7926adfa64b19e0f25216823f870b5e05b0cf3ce9d8a;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h34425cc5762825f3db065ed5cdeb631442f3246ab427bdef8a0492f30d66bc359f777244b2c51767b673fc53189c97238802cc9871d474f7d192d29dc4567ef4264d345cd8e0830948a7cd9542714f171d1bb73f628b9e197a00e1e5cd36af44bdb3;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h45c3cabbaca8cbfe346b156b2849215eb1f012f7c67e7705f60b7c801237f56e6bfe17586dea744bbf2ff0ed24c384321df4e258d33ed5412732c999cf0d599cdc04c6bcec5ad04d929e7983a9040f8f120f65455cff4ae0624f8b4411eedf6dfa05;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5b5d87cff9b9d5a20885d65fa6f90016e248b3dbcfd8f68efb258bcc016611c6041dfd610b9e9fe69de8fbdcc6c53b70c2cdac49912e27b24c7a26877466a0bcbd9375e5380e7f4af6402005d774d572b5d8b2b56281eb05ba560ed1448e59188b63;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1bd6def75e01d6f6a4b1a7c0b8c10a20815678d3be838ce8ed7d73d0a2fddf99b3ef6e331069d268d32242491e16e3af53a563525e3bbc8b62d1deda5bdeb384c5dbb91fb09d4d7a328b3b1fd8f6ee88cda2b4fa8eb03cd13f41c24630003278fcf7;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7ff6af7f42aae654645c2814dd54d0c1af5cd3e6cb203d1cbaaeba418647c605039c787ae26a8fae8cef61c1f02b683ffdc0e7686005ee39426b878bb05c83168d6cd42bc18b1ebebc3c7012c2d938cdd21d5ec1524cb9f9bfc959bd5c3dd2f301fc;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h47a7b2422a5854af5ac2ce7adac59ef0fbd8afb274b666496f895373b30f8aa624a0b936cfaf5af379a2960683d5ce398e37fb61114b8d3098ca7d6a8d36e8ad767bd82d0438d371d911bca88a06a265db5ca58c0d10d1cbd8c030aafb434538d12b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5b1ef4feb191b8307037231bf37dc5a550c173e66490a3f97f94dadf4723ee773271a47c18c5c10b7fd9fb317944fb24dbce53e7c8f92bb7a61371bac323998134d2d3976e68edc245238411b45aa7938cd483954d4a7bb88ab2c36c389b4f19c0a0;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5f2d21661a5e3e4cb9fc8aec06cbd5635d8b8bbfebbb4d0c126f49716604aaca07328c9bfc6c44b3713c1a6b369a0fa8be1740373d1dd8998c0c50ddf6a566f0776b95fbd71e2ea19e6ec784d84048f96f8ba31a42e15b642d16c025048bf6bba2d8;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h720365f25179151410b68f460b3c4baf03232a27d59dd720e5ad9b5a051a90eecfde2713896ed330e675cb47656e549efd7ddc59bd58dfe3f97ef993e7d9b03695e32a2fef4643e593b3c489f1bf9944e60e1629a855b34342ffc2ed6f21d61e4ed6;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h301a38f03bc42e73bd663710bdccca452fd4e2e355e747d41fa26a9b77b95a7904cfab1eb5055341a63ac96b9c043868b243945b558656d6e7c42baef49181a72c8d7e9b2f4e5f1a7b3359d83814fc4e6de09802d5ff7d831b298e33579fac577b3e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd03688c7490edb90f536adfd5177b7290d9808fcc6ac85f3474547c660436c4fa23c442f0a0663fbe601176957568e52cbab24a4c12a73629a2b43813b3874d10d4380613e91131cc68f0475541f379f40c60931f54119db2060abee2c63dade7679;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9713869876236611a4108051979bfaae9357c266326f298178a971427d817c2c128d94e4d2f7a1f37f1bb6ab2eb241bcbd5ae75f974fbd9f039cef585f04e4cf32ba52c07c77534d71e34a10b7b94354023aa2dcaae33beba335352a7a67e19a6a71;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hcf40f4c66cd3708c4f4cd05fe2d4c9d11127913eaf53dd47a5e242ff277a68918379195b306f9351d2eb2e09c00508f458eac623f6276456ec6c1aa491f400b7301e1dbcd5ae1e9afc512f8090eac0b8cc73c3e8315275a1a68ad1b1276a272104c2;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc4ae27a27026f1483d660f0785c24ff8ae75bf8fcbf4d94185073dc7ec7204959cc5481a6cef3d5d22b50f3fe31e1e8b66392f210aef3fcb58920a3b0cb1c75c747df6e18810349a089aa3473e7302b2a762ba5b2666555864dbcba88da32ccc8a67;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h51be7ab1bc24bba3e497128e7525e17588b92235decd096795babdcf8ba66580a3b864fff37f66538d5e0f869366fab9db858ab1af7a7fdfb97de7e8a556cafbdba7590f8b2bdb7fb1df7bffeb274d52d006eef9889d5ebdfefe091f75ea9fe8fcab;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h254c11e9ce19082ca731184f1f2f4dcb47f1bcbe69fe024818077ad8cd903b3bdcccebbc5abc16255fe7e2ecaf3dd807e6a4648f18c4f06815ef2171a8069f3206049cbe046773f853e0d3025067e35b9256e94acfcda2735e346cd8eb9241558b98;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h592f467f9c2c31e15a8c24abf23efab9752fd6c79227f4e1f141d9126de10fe368c66a9d93272576c99bdcf7f3550448b018065ef7c41f60dd495d059062987c1823d0ab5d1d323951029a55aadf8ac0db9cc8c8601ffb74cf1a5fd207055dba8a8e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he319ff0acf811c88059949a599ddeeb6c2d0b7baf562787945c5117b45c8c2ddbc6e7a180d5be22651779cf71dcad1230405454a58b0c2862b75fd9543b0ca45215c21d79d0c186585b13de336d4d0f61b24cd8317232eb2148af443dd8b7443ab5c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hcf66c89203d6666eece6682030ed2d820e7cd696d40e8fbd0c186e7c9c81a0422b5099d2373016442cc5f6781bab96052f0a1270e8a92efa75a6d70c78b554d40037f0d8f384d3860524a55e750fe24914c36332fd9bb5c09763faf998fb5f957d85;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h69b3e6754ed7a363fae2d50ce2b72ee9c94296d26751ffe0a318946c4f52fb609195ee1959ef2eeb4364982f0589194d0604a010767296de7804bc1ce45c31b356f2603a7997f9ef30725e6b4e6752e54de4c2b9f7c8e47d9f5b197b0b11b2c42b43;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he09ac0bc42b2ae9c356a1fe5aa0d20e2d52ba790475f2642371ef07e10781b8427aa28f9cfdd5804ba432deb545fff9aef81cfe8d88fe9197cdb173b4ac1c3a02c420ad2bfb75c7887ce530f48c0338930c879c5dde2c0f2e09b6c0e4d92f42866b9;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he028888e9e45000a761039f00b9caf4e9d9778fc3498dca10e065cbd9e85f4ec61ea0425c8d406eaf47b0b4739964352ff5fe926eb5e1422d74a53df58f081c7f4063cdf96777fd995c5f34ab8809ad9bc18a950c494ac2584726c51ce210320eb50;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'habc6de08f4c7e9c3dab201336ce5ed2ac047f161d4a0938c66cbf563ff14bfcae6d93aa642423e56170dad16a9d6fdc8bb599f318391ba522e80e1214904cf7851108ffb59b02995d1c3a03b43390ff01ea273b8713c65b214b26ea0d5a5b8fa14f;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2100382b2968019afdee5783c456f17e9a03b8110a99f5145a59295d24910a246414913b328514429763a88f27a35b233879c9d2f1c026d544709c2fd7afd2ef4c37ab249adbfcdbd7e3012df7777b4cc6c6a09d65c7453cae7c163a4c394b490c98;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hccc3e69d93ceb0b256d5800bc7abba415a8d7b8a6702b525009b6b1f7543b59d0d3b86942f54f62813a52a15d2fb6436ad50ca0b114565beff5eabd2fab7cb83b00e108c3c56ce2e9fa3a3d8c4eada672709158d0a62f4567b49e63b294b999c4e39;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4d04a5706c75b7632f8b04b8120e53af5d310f23491c9ef9fe95d4c1ad1fe0f8253dc53e14068889649d4f96420de5dce1f745248cc5282d81e9386d98d041d8c25cbc0d56665acd6a8dfc8436444325db7ed349c866c5ca923779faa041b5fe0b73;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdce201d05d9f6be47eb43205b70bfb2cd6e845f49bdc72857d7f2bf345ae9a46fa0e3695ba77d3f0f7b7230ecec9f6f3c83c45f144d90ca739e245a895599846ec203157ec7c7dadeef40ae03db08dc6af14327b1092bbe6bf8a73e227a49774653a;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2073030960745c0816de57e40f0859ce41bbd049d967c2548b74fa74c52dd83707475f24ca646c37c6139541bad913d80d95d15fe0fb471cdca05ee4405943429a1c624dfec263724806793c272394cee80dc1b08865f5ab2f876db291170b7c8f10;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he745c61bd235dbdc40256bea4a2c50ab2e50008ee5f0b1f55fe4fc966a239872da1b3eabfc15bbd89e88098438db6b56972a6e25ed9804eb85db00c5dc9c8154c70be374fb67749c25d4d73d9f7d29e2b804fc6c5726671304879310b11a55044037;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h36f77b68aa5f27079172a74f92a77243044bcb8212ebc5214753b1c9a69b1b005e179d1f4dc59f8b08f9c77e69db478ac0584c8cd62f1e668f538e015d79a7558666b4331f15b9b5e3f29f03cefa376e9a0ce4c2c348f804a66a7626ba92ef0d0a9f;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfa04742e426144dfe3639c5033fc9c24ce08ede4837834f0e552c6bd9fe5d7c9663e5c212c93d83d9c30252ed5735a8ccc590cca6ea930718ecd1bb1365975268e505ba56f34bd91c2cf12b9e3f43fa5f14404e0f81a7bcfa4448bae6650c60b17dd;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he91e8195eb4fd1623b26740f822c08c18a47d5379598d9ea4afb3b93fe16354127002ac2c0a65110294eb5d3f22e41a09900787a81c3f2fd094f63291f413ef7ae23438904605af87f00bda52b894b73182bd8494cf1d3e90d203d5599ef05b75ed8;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he6d918e0ddbfc910d35787d08373940d80ef65f619f4f873447f1d521556c95483b9d78f8afef84ce9785237af0cfa0c26c92aa9fd5bc393a4aefe9fc871f828d09dcdb94caeb7c43ef38b486293ad1fb3304ea6f02a46b6fa9b823708813672b557;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h832862316c1ad6075eda244bf38fab7caefcf57ab3775afa239f8d1743d12a7cd760ebd9c6b1d37222928bb8881c15e01d1708ff3ef59ecd4f9f8952596a2e1dbcdfc970f659a1eb88ac1458704d5b520843469d876ca8001232f8353aaa068e6d3;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h12f33732aa940d9fc27c15c0b728b46e4b06f73218c0e560851e767d779a0b6f4751f7cbb1ad92b55a97302f0da9f6ae41e55df43a99f3441e8a95c66c4347e0bb6ebc8788913b238e404b2c5a61dd2e6d7dce769056bc400cafc227b8d2940c8ed7;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6c17061646aba9db01827b44dea61163fc05fd872847c5743d75ec8db2b51828ea9f58bf6fd9a506dfd86b3230ea7cd1e672766588e47b8596384b2a697d1a44fe05573e91cec2e1e4b32ec7f4e345c3cea7dcc764c0db00297e2c6971c9f7cb2522;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc2d1fb223f5c936c808b702f9d9fa737673310a1354a963f0e8cf873ffc9bdceb33d55044cc708b941018e60afb0ec96b3298f7d89b1a2f2631fc88fe90a85c881d61afeb9a7bcf90fc7d5b76a657b3c7bb0b4cd1e1aca0ad3179ee1f68e1b6e9fe8;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'had5b80e68166b9c60f8a39366e9e3e9609ad94c4b33e1d5ae51fd87774392bf17e45e5144410b1584dc173cf3bc9d5288ad695c433cd91aebc67edec8356f478c16e74259581f8c435d6253fcbbf83fab039350d9b1f5be187b54307410767494302;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8ddd73dee00d689ee8aea9e2419cf1ad5e2e4c08b3e223c4b1c669ef476351875fe51d91ab948a879dc72d0f0f3b2220488101d4e13e7457f2da57ed0da3b1a1b27402ac0050453853b644b73747bc1bf7f641fe305bc4a1f29e3bd50b2460a8b0fd;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4f953e207e5741a182e96cff075cbfc73dd5939eb8ec4e2abf1c1b75a6fd478a971af3f251687562b55f6dd0f3dbab811346939a4265bc94a1692dc567462cb178ce87385a4d53f716b2da7b817168e7b891186f14f15b18de61ef14f19d7586da62;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h97232069afc9cbaa9da5a040be281340221bf311672762e157c10c8ee99f69b5d87644cfe1ffdfb3a24105f4f3fd99f075a2b5e5bb5a701269881ff008af87d3a781ed5d53334a70c7828104446dedde7d9751f33274aa860f9980d678e0e23fc773;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h180c5c2d19e8e087d8b25d3490a2d0fb64fb997ab03251071d9ebbc2885f7b54b09dd6181c75860b284a150af20c623b0b010c9ff431d4b82f133c0c9460dbfabac510fd3a66c95ef2f6e66f691d9f8357e00a50d7e1ad3409abe5a51681791b5a79;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc95a951009c9741d23530c375effc41188c588d1ea3218193afe9081cdbcf6879a242bb61055436852948cfd01ef38b4286bbed6d1bfc63f501246bfba68aaa543d30426f0b7d8c05d3b30c29a333b39a2efbc38282f4c9976a4a954bac1f7cb1d0e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfc2d3c343044cd1c3365424f24635d04b91bf9e49c1182bfd88c21ef93f26c678f6187759db933f0732d87c8a97dfaabffd99c714fda090377c40dca85cae8d2e9051b7984f0103834cd07b142de0805a86986713d3db0298f2e3df9942ed74d6de;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h45b8bc3533d25df7f655bd76c72f4e6a0a0a88336e2c05c01110a805d8420fa7b93f14a4c5c0e8fbb21231ca1fe6492483c0fb47a90dbb8819c6f88afd8f9edd7a3c52ed6121ebbe433031f4eb31ecfce4641adf9399c930b1847c4fc009a19a190f;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9b331b01652456c4a5199cbc356ff1f0853afc7d1f85724502c4257481457029fe8939363bd615e9d03e17fff6bd5f876ae08ee9628f902f86fdd34f6cd6eb81990361dad9ec17033c71357d77b0da02886162fcbfb3ff6b33bb001501d04efef999;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h11133807eb9f3ef5f9502c86eaf6a9e0cce123e8291403b044d050315ca78857de090664afd5c7e0979bc3519aca1c8b1ffb3187d7bc3aaacd441dad84292c5b71e58a0203dd126df75b3b82bfd3df1fe95436a3a75e2859782dbc4ca5ceb8bf3646;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha9f9730cea805e0ed70a418e00534f2ed2e1fcf7fdd696fab61b9be10df88afa192de20e5e7c6377202a35ccbdf994a79027c6d4414638392f90d4c9879f3bfd192294b4b850bee32075c225ca7e28e0f32be696c294060a1c924de0eb932afa10e0;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb51eb7cba6d085f8130fd70c310f8c4cb9b3ac0899c3ce894c190d51b97f8125fdcaba66ef676bc4c11fdd6eef7c386cbf33c0bf02c167b2a8045d32e97a55640acf203a2076af2fc21e6eb8ea9494259a1740c068938847c9fd5ff3d117e00d29aa;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7dbd0dd7a89ff0585c1a00d25c9c4c621ea0a8eed60307cb233f3c08de84b6ed746c21d36a0e706b8f4c40ee66633a4e8cf3c5d99d44cc9f15181eba338bfb2b1232c4b592ee80e214711d8c415b57149eb7583e6fb58e52494500541bbbc4397b66;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h788826f21ec0945f9f2c89775786a8300ea814003b770db4df02cd9f48bccf1f0f8c7d199ba270d3ef5de306f374b66003a6c9b0af2bf4d3140ad2d642402f261e4f7e49f57d65d4e734748330063e8840025cd7db6b3977de72a94e540367155c1b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h80cda401009ef576680f044826247ef150edc02f2076e293cc696f2e7dd6743287ebd85d845ee8d08570536c73483cb4cb0f843744103b9257e9d3844fc0fcfd2363db4824240832196fbbbce3720dfd3a13e0e13538ca292d7e070f3309499e9f06;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf77ea242a466a28e51f092e280d9c79503bb8ecfb387211375c4e9baa5af3faa82984607842a489645f42ba7c092427cdd21e519a9dcb1fbfc3794be2064cfd582995eb0376ffe3b35908c49f44408967b8ba79ebc6628af544464b45b172cfee035;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb07f864e1229fc62907801dd2684de755a344bd3425b90f7402637a5b4d1fca32e2c96872c75416345b07e5e407fe65f183ca249b9e878072bea803ce6cc2bb389516ea38257cf3a00c8552272c1632489ec970e66f04e7fdefc27c9a8d1a3f0af3d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5de7539348f5a71a167b8d44513934ff0dfb28fc51bc908e854f8a1e844902b2cd1a8df7f31413a3ee410a3d3f3f77b3216c85dbddcfb282ab32866170529c6045c455c86a51a215a8c45047f4ace5c57d14ee36f9ab1bb68685b3258f1dcab0df9d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h92a965ec14f623f1cdcdfebe1ada36560b2a909c07b79065acb176ed617cfec6004dca0f0028740468eb5f61cf4eb88dccb1013960446febd16104b0293164df56c5da405f86364dadcadff253e21f6024017b6053867386dd302b0a1f102a4639a2;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h85592380ea3d81aed07e67560373fdff3216ce524588db6abb159f018659f355ff61d33214872b0884a6ad4526b609d336998b168d702d245d6014dc8ad88ad6d94339131a1853a21f50a3924fd64ec063c5b90110390c1360f6f8111fbc9f9734d5;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h613d559f68c77b62d1d5cba12c4ad5d9ec0a2fe33f6d465b6450f1d989d44a8d6301e249c449398709e765239b3bdc5371551062cf53aadf28907d241e5b90e5b2a921fc75c8f99b54272dd24f2bc3ef3e526589707b7cae4d6de1126786910b381b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hee626ab213b349343573c624eb459a8cafaafd69baacf5f9dc672f841935a16d7becc31075612af48027c7ec3c11cc4417bc2fc2249c0f297aa1e70aa70a10702e5cfc3ddd284902d47ac661da3c630ffbf58662ea613daf5c61ef63a63edb75e2f9;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5ab719033991d877be99e7e7ab1912693fe25f587c97173e4d22139ce8b0d951c1c0dc11f922e4958a0ce024882fec75eb18c376537672a89db4fe3ad9f40498c7ae7a21286b7dbfb33e45479274b4c2605f2d58c1b4f35645447b2cff16d0f1bfc2;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb5282333527face4ec2d367fed90a5913b41e19879c69f11c7b34b12ea902747464bed663b432c4952c95ed5e07ae09be392f472763d181d473a70328c6110acc81f01c837994a4c7b6f112f271e4fe90b79f6b6ea8c217b8a61443037ca4963c099;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'had1fb09382f61a22e3e75b6c7d7c7c10e29fdc578fac7cced1a4e178acd874aafc6da8d167df7b9fdb8beb69cb62b57e159dc444c2961f9f22d11862df9eb2ff1eb5b02913338d48da167c20253c82a3468b71dc9978dd83b62997b3264aeddedaee;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1391041b070b2073ad2952be95eec16c6765cece188dc9b3bc1076ed7e1285030a4b0c39079e42f367e3dbfb28e0334710379037a1d92dd5f9b9fc41092e92c868609cbe6720ca774050c40e588d6e4a3eb842925870a87408863de95adeab8d3b57;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3dfec3e56ad42fede7a7b05a04ebad3c3bba0064ac17e0cc070c73b247b75d011119afa0fd4494a73dbbf883de7b3c17654d3273433a411404a2e2fb6cd504e8fce1739cfa16001fcf13937e87c9e801291fd50044b42c7cae675449b4e790344263;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3a12d0cf65a6224f63d0fe3e061396bb2196e14e131adf5fc7d8b0a75e2f529218105e073c44859203fbdfd00421a45a2149ac4e411baab46ae0bc4ac2605841147aee7cfed1e0ca8acda1ac7e6b3292a4ffdce23ee2741003b5421637b6133b618f;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h64d44a067dd1aa80effe2a6b04cf05a9d790584c92791a1a06a5c3b90f540a2507cd4f7e68339a79e85976d2be84eee84c7a84b0f194e4f7ed9ede54b2e63e1164e2ecd849b49b1ad64c50c531bb28fc1a6d9f54d29ce0169682ed93dd054c020d7a;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hda73be7b4fbff0bc54e9f7f5b3f5265934a97b4bd09290448a592f48eb06f921caa2f81b6306de1d8516301d2b79436605d629f8fc3b9391001f58dbf5af16cc18c87e47940e0e0e029b340b6e3c00d4528fa0133883af7ad5b97ee4357d054a607d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7049a2e1761a0f84be74742854fc953e40b823861735de43d0763ac4236d094f2c197eec2d042c33b234f85224f71cd42ca1f63f46493bd5566ef22001366202ac02a9e8459ee3d2c5f9500da5f73040f82895edd01a182322272775ea32c4d3cd85;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hcf027b3a73aff367caeac08b1f27c1c027804582818cd903ab4b07f63c53183c8969eefd98c5a197c50d19c75dd56b6058db7d44204d4739b33c549bdcef512347fc31c65ebc193085fd17072af99c1c8dcb1ee4178553403687f0c896893f0f37e6;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbbd45ebee41a96b3e29bc84815aa0334e5593cd58e0bf9761e73e7a9f288132439d2f86209cd2461b7ea05b78e34937d01cc771a4d2e738f6559ae949dd696278932dd7254431cf3eba917b8a07f7fd818b13c7cf07874b78ed1d6f09e7d7e270a60;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h573bd7104751da9b91b5738c8125c93a4753a656c17d3ca8035729f2764cfec2e131ea4a550efa8ba6a42e8c48b2944d246757aa5cf878e82f8bef23c336c1453ce99961e5bedfe68462a255577f58567e8f108582bae5662ca1ffc9ef21e3304212;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha7336aae575a04fa19dd6ce7a892e7fa3584a0f100f6f6b6e9439c91af462d6efe36c5f10e4284b4d7d95911e97a75eae94f831e01cbed6386b161a24798257ed15eb009d3b6261389b53718d29bd3b01c1644aae8b98e83700054ede4ed59ade217;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9b173f880e68c5dde425d92b9dbdb2cf60a0baaa11ce908f87167d2a96fc8ec95431be0afba9b8b4b9a810a1427c46e80b06b9fd961431ab71d7d18bb2743fc210997e15648b87d928a0c9e7d3a63138c14c7b788c1928e55bda8f1fb06047415ddf;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbcf4e7b7c403f4b1a93f1eb4cc2869d2839432aabfeef26c35e1c5d9fab6383c7c26d2d1d30d3022208a4a25bf3cceadf83d160029992274376cdb4bae9c3420df68d3b3c6190f1eb928869248ec6ed60cfde191b4af136434e9f96187f68b37705;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha5e310fd9ca463e4b0c73415b325f09cc440f280827ba195decf4bff26c2690c1bc2084d10c117d504ff6a77f2c681e5ba93a1cfeb351b07b93910c97a3ccecd10a973e305039bb6bfc7135fbe5d0c6ecea9f0f72d1fc2140a7986434036ee47279a;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3ecf0850cddecbb906216cee7d0140e9130d174f7b73e3baba7b003e9b0e8ecf7b028d8e7e43ef08048db893575c308dca37e37d76b4d486ece1f7a498d3294cb2d24d58ade6671b20afb86f3ae7b61f73bf087ffd1c84b8b1347c47a448bc9f4541;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9ba3232defe6d2b39a338592829796b7adec1d5f2b745fa9a6c67a60cebae737c89c07dc3a081d19a134cc85ee8988f3bdded395b1fdba2fe54cc1dcd8358646e5716a2c9dba9280a3dd38f6147d472bcfb51619fe182a869222c5b4e3f03bc4f87b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he8b797c50b55dd21835edecb3ea6d6a970c724a8e112366730a72e32bb21743349ed969fdb298ff856a236dda823f2aa7643a28d974425954f052fcf6e0a3f1eb8f38301003b541668872fde5a7eb467cdecf02f9632cb8a46ca9232f971416f7b92;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h40658448b04baac6f9ebf4060ed0cd5b361e085f6a83a39893757d83a45b24f5158423d05b7c86e9aff6b46fe3ae6976deed1da203bd7d9c0eab4dd20013243fafdcd567ab271f525c5d2ca3c9718d2d1d5171eb5667d691eec6c6e88d9b87812e5c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'habb457ec3ccb200806c676cf70fc351b7a2821e6f6f46f2279765f6a02434e5ba2cd1659b7e7a2efa3830d2911938f335303e6c8856aa0210dd9f6c2d7725a0cd5b3044541eae8fd66795a3fc7134f24a16d651e177b69b2cb8971107a6900a1534f;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8396eb558e5bbf15d5358005063152e03d17a26c838b9f8f8e91ceddae73e3edefac838377d82b92cc6be86facf3430751a03eb321517444b32bdd29a5c0659163713d6f295a39c902a8eb6ef8f637b8b302adbaf764a4e3953b0e601768a2b5aae0;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4cc0946838542ef4daeaf8446dd7be35b1cb0cf57cf21d7ff007797b09a0e79808fc4082f573a615d71e43667eb28cc10fc3188d7faba9252ee16a8a036c167f6a3d2dde36f85e59f6464d7ecf0c7b7f00399fb2398f4c316280d9a54e63b20982ff;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9d8daebfd967b4726223e1b41ef88b44c2ee0a7b496b59602f4d5452026df1a555b48198c04fa5a2252a1b4719ce5cb9272167e9d06422e4bde3dadc4e0bf8dad49f9c6c61969ae148f0322b2c04633c80f77a0e8260ce6deb12552b48970a6a2e30;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd4e4f31f80c1674e55557dabec83bd11c4b4699088d383b7bb37ffe81ed136f8a91107adf59ecb8969155c6111ac9976aeede03459a9c2cc751011e31f3faddfd860210545e149fc5b9b3830284053d4d6ae6bcb94d1c9f1b4d5a7a5a471798a6e7a;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he56f6215404cb21acdc0071dd5f50d415c6eafa7a42715b4db0b28a16d9b9bb368ce69b28de05a51337d51902c0463ac4641371af8be30a2b3ef67958c5efed1c3e79e80b7d6ef64a43906d633ff762aa1e648e5ddf80c35ad40d3df4da97f2a8e1b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6fea88e5f6d6a3cc0cf55b595844bf682993b95153cb7b786bc4689213f037bfb1f1791a4b238f8b6fdaff8b5cd5d72fc83756b73cf9552af90e6c3150f4214c04cc6ff8af1c6c0a41acacdf5415f4fe66565489b551ea8906cf4553b062ba1a3bb5;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2f6b8f474987e40454ff04905058a2bd5ea03b465f14e768923cfcc4fcec6fea167cf69c26867f2d6cf2fa7f50585fe9a1181eaa8a3ee85cae7daf433aadfecee5414140923423ae2346101598e38490c9d0d4b349eff90f45d95326336e193e838f;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9765afd853642bd040c86603daa85b25e442b49a30faf4c1175757c01276772d5e437bd4d47c51b384a66806e721ff41972864af0c59a48feefe049e2a6305615137be0b8731eb9efda8515f219a209a4ab46b35de2e1bb2ae4576f4539f777d7fc9;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he54ec54433fef4241dad212b90c20a10526c881821d7b818ba90e9d31c8950f318112f79f142727b4745922006af1a9a881e85197b21b6be87fcd8f4fdc79297fecf34f8100f1a0def58f64f8e53885cdc45cdf666626fa68ae912d944eb52827674;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he11b8d6faa25f5a29c1199067a4163e463a821d970b95cc5965d3444dea17b56f8248679cb31c19f3425203739e8ee10ab7caea02986dcf096999bc14c98623c4e49b94978064ebb3188c39a144e83e4964ed3b588c77a2bdf6fe11898d36082815e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h17b45d7bb8e0b88e702242ea8852f689192489f0d193ed82940d1b1f54981b8a8fc9643e15781d002bb23547929d380c5fe9f030841a8232a6c38a8f6cbcc28a417d9417328d6a40f1efa8ab03bc8c99d675d3d6ebe18fde92d534a32d31b634d9d0;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb9ae9c332e4795a8cafd7db38c8513dd24b67ef036b5bdc3cead990e7f7bda7d01ac1eda44b14c3805f4d4600b553b8bf4effb031a48b3b51015c32bf812a36f1f9643a392139c3493f9c59eebb5a810b56a83a4b0306d38e8dbe5b72d54c9ddaa15;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hadd62681caed09ff18b6dee0a015f2745b541705407b7584a5b6ccadc136a42c2c5eff5f8c10e63af6997259acef98c1a3051a5b254d2f2df530fef6e566cf716da26ee7fd3fb69a91646d9667b771345e1b9954b17bdb7c4077003c9256fca674a1;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3960ca3dd2069a3bfe40f25a0a731c274c68ca410dd3908720f5a1bf0c92a68bf5f4f8d4db989091b274ae288f9daf6f08310fe840c06f8081f767474cf3ee381a84d326349d6ed925adef07be2c324127117d9888cb7561067d53e4891c385a9571;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd968db806fdac2b9e20558c95211dfc55ef9bbe3b0e09ce4c625646eb7b79182ec62b400adb83f441d350c6848f041af67e8536994a8070b195c29354b3336d3833d9daa73b1c43f401162e9762f0730adadd672952c17c5d24b15ed9ce90c7ac201;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h317fa288513544e1d00e8103f28e204f28b61400c320d96e5c7fb7c27f7f9f8e6c69a58a7d84a1184c20095ec143a7ad7794fd8404cd07f33b08b2caf13e3f70e0b544cdf76d43d717d1c68b123b033594fc14a15947041aff126a7ef9f01c4e1bf3;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha12bc4c8c03048cccbbe66f93b91066acd4de3655f1adb97c22f19d3ed9ee0374eb135c50bd0d44524e7bda56aca71d42128840087dc1e68ea5ae579d2d5848cc9bf451306bad73e1b4bb2855d42ddb2c942bb4b054bba8cb235c5a2e4427ac9e589;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he3bb9a77746f490dcbbcd8f6794dae5f41ca15e056d19ba2aa451dd2f0289a3f50f5b4fde513b06327f372372d65d909edcbd4f341bdbdc3cc1f4b4b78cf1c1b049ce42b6cf20c36dd106ff44203bd36d15e1d2d97345f2809aff08aeb1fd4a3b870;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha806f74b179fea0b9ad56f54b418b465e6427e9aad47c8ac6f503ee28adaeafd08b7f403c689cb1bc35ab33d2a596de8cb1514c019a13de3eebec834dd25f29ad30034cf86952924f2586dc5017f490d952e2e869ea2abaea048b8a5c8b9c28f2520;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbef5653383dad1499d639266d3c9ca16e4261caf1b36952e672264029fb486a2646f92ffcfce02c55c37155e04447f7c63f53d9cc1fcf10dd47b99698d0f9eba55387d5ea9b361e7b1ee4e79d399b3cd458eaaaf4b6cde35fa6484d8c413cd1c35a8;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h920b9474efa8f7355a333858eecca1b3080f5603124f2a63a0721b4cae31c0ad349615c0b9f94e72ae454e6ba5793be7d61470361203a1d0e652465d8b6342724fab9b2365d62ec5818001b0f58924cbd1ab2b43ae341668f42cbb803b6e08e1824f;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h84e12a94def03ea301bed99baaac6aba3ac17bc1e61239ce5379c72c0f7f6a182a852cdd3fb3c8e660d4fc0bdc2cd10dc64f8627d8085369fe0b2279753a82576c03eb5960f9e65ebe6d6372f129dc67f6c6bd23fdd2cc13dec5b6dc6fdce7702386;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8100947826f38075ce5b9ba0e3ce46147c3c3e6ecba2be5da0827b745a64a5e4dc190535c1bc90a14ecaf21a630f5854323ce73164cb57350bb86c74e5641c08fdb0b196aca83b5e2bdb881c94835927aea86a068628513f4344110f6c86f0e39d82;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6990445191f6a615aee78bbdce14ac133984245c3fe050ba2d14d13cbe76dd18a40455ef2256b6d4ed1fd20e6165c35dee7ddb4d8544b39cf5d491a138330a61558e5920cde87fa863656f2719e6701e7bb9726610a159237a3aa2fce46f26a2b1f8;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5cd937aaf27f67fa209f2b71e826711648367a0f52abf24f987d088a338f098bd374c72933e82ddce4577e561883cb67e45bd5a5cb7ba1cab2dcd119c6dd22326aa88838c74ca06327e5df4fa05482d557695de4d400b52196630423d7233f338d1a;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8936028b8d4a57a8e9b03f700f3ca960909ea30b40318135cc94eead358e018806ca95801f0a5d781f597925ef422dd71c189231c6213a61a49782e074e1e98e13bedb33e8f164885bed836b214047871c6da3fe6b998f295ecbefecdd566a4ac361;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2025c0a0e529494b7d5e1cb9923a22c9d43dd9e226d27e809ec595dd4d514ba9014cef158846880a4bd5e65a9ef783c988305a00c350aeb0911eaf527a8b3f344881842f82dd72f585858b0d5d4266e0456a53f415e5f5e9916be065e3e204f6c229;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd63c4ffbc7da66d1a84e1132ea521f30aeae08446ffb52c72e2b7acc46a595cc94b52f10d5e85ba5d1b549cc919e813793c58fe2a426a0088372c64807e217fbcc48b96456c7a63419050d8ac32a82882f5034de0a07a593621448bc74fae0de8ea7;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h11c3c275433ac3554d25941b2b31b42cfaf1e92cce8e95088d30ee1aad4015423486655a590e4cf9c9244e3b39b8c5ce3332e6a9d4816de5106ad3f78c9794c3cfbd85bd432f9f28022e4d2983fef1d11e7617e0fb7bf4db1b267bc48fc8146652c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc7dd67682f5e73fa6ed7d94c5be912f63696c7abc912108be8903fa164aeb5bb1ebb2e9d6c33a48de31255c9d63678669c308fb25b4b4297c7c1273ae2ee86f4dabbb7996393e89098c92b62a05c3ce1f136d86a97d711ca4d96e7b6af7278dd7cba;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he968dbf9a2f0971014c2d933485c38ee81e9e75e1a37c7929e52ccdbe916de9bb71149fd3cb6c5b8f4f9f3d6f5d47fa036d34b4c552790a951319ab97d115e710e53e4eb4d08e0a9ad6cf6554e93ab436dab8c64004bf3eaeba45dde73eccabdb428;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8f85317947e0cb6a15cb44c0f8d98c1df21278a0da9a1a569c6e6f78009fc508196c4b7e2fa3b2b660b0a9bd826ca1ab06b8c091eb80dad6f06a91c741b9f25732de1105b43768b1f433b0dc2a2d6810a9570196d98d969f29b61ff92e1bf676a45b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h42c872676db49c94a2c85438624a6f04c95f1604f5a8b7b4156d8bd3183cf1c92c7ce0cfe11eb4974839cb0fd842f436fc43923680f2ce3a354f89f49ca46f1f36cccdd153a5c6cb30ce9722a344c628ec0bb5b85611a94a27c988e8e567a89dbf8f;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf3d3871c118dd142b78ac0cec7729d49dad1c4bb024485d6be6ea58fee079c32f2dc2d8ad7f5af90820eac5336667323674a1ef0c0486cc2949e5a7452f2f0fb37be86968b786044e973c55118ff6fe91bc02cc32cd77de17950d76d4b120cf52134;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he2120da44f69aced570c060cba47c3681798ca91f08fe7a25bb59897a9e3f090e64b3e2e4f3fe76617bb581c0f43402c25c6b88dc48c1f033e1e38faaec888022f529730cf1f73a20d744a7763bd4f482b715150f1a78c363bff4bbe94c2290dc90e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7db8ab48514198bb65eff7b8f62cf3302e32e1d1a178b002b0383381dcdd57db9410b24b9fa7deccb5932dabc78249771646f52b93ce95a3238263f572db10b4695fcef94d25e9f5f98f46a9ac1243fc2cae2f9f959dfdc6900953e8338b792dcc83;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfceca2e87708fecbe478491753acfa3e75083e887b7a5b48bc5c3deea081858d9fd367737a82c5ff411fe1705ac4b0692ccd2ee0de3d7c570e718ea67d66099c04e42fe13b7aea2950e8e5963e518481de0b1c4858948782ed0b7d3e39e4bc0a0bb8;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hda41e26590586a4dd8922ce9922908da11bd0fa9065f488732a34706b205acbe3df26c58cb9b740f3b2c5b01e558d203e9a4cb118ee90e9e06076435e3543709a3130c84db225d005aa3ddbdb4653e0d2830cb36689e17e21bd2558ba854f86e2e74;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h466db04b738b9e28278ac79792360e1cbd1918fe5c6004ed9838e1cd17a9645cd14f90bcc9dae088359efcf44dedc73ff783c162769fe9a4132e299b7adea508097956548e3688b3dc20abf7231052ac1696df4862a4f647c1c123dd909008f1add1;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h758eeebd759116c0c9a3b8deccdf9522f1b00d0b5a9bd0995ffadf342fb797ed2be81216db069ab5ab2c7030c08de154b2064f1081aaf990ddbe4eed97c5c3d448e57e1bf9451a97e95e710b47b6af2f364cfdf375b0a800430264714d7259e36bf3;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h222ee6e0119aad4ed18cf42402fe7afa2f682a592646b91d094f0b0312313384f017cb1df035fe7b2e108be59d574ef6df455a77892f9d8ae0e7783126d545f2ee2d4d0d7890570c0e734ffdd3d6b0ab7a36733e00f2ec65d5f132440e79ad682dac;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf812b7716387e18414221799754cb0a9a69a8b12285f93ff8be0db3e40d9699687c909405378655cf76e073fe52d5decb8904c11bffaf64a03cc550a9fc5d0bee6706306364c16e31d635d92102147be86f9997d4d4addf56a0c853d325496ea6d24;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8d59826e518e3b89aa4d0b346820989f0971ebee3e460f72b5fb14197bf5a02554ccb83e9b7d16147d1f05b5e50a1efc050ef8718229656ba5b04a5df98ccc70f0b96c9e8b3fd41d15de417282b22d207036d4c84acef68fa57224c747d8b22e4a4f;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb55ffe3e352cf9859557dcb9bf21e0d2485e813952965ab581387bab44745f5da616cdfc97d3f666eb04e643fb615d4e03079f6783ee813e6978cd6a6f2fe72ac511b4ff3de7337ae71c73b82743ce7f526ac0e6d358a17aae1c6e55192091727846;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd762feca9144937eab952fdebfbbd011246e29de0569382d23981ebe223606a61d7beb365b339ac3421503baf0ff9331a5937cc87cfb0085e2b39da7da8bdfc7a7b49607523bb90ed12246b6b9e048e80f089bdd60a54af775c35b00061aed977d1a;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h83bdb0abe0c4aaaa1879d658f9f50a73555e84d7fee1f3173e98e4839a36a9beecb1d979c8f9ed88402bfa46e10637556d9f80c2cac5a9a986a4b59024df3f65ef31896d08a00200a48dd6aea90a2a0651c60471d77b8d55fbb5c437794535e66127;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6f4aed34ee6176331dfe6d44faf92fddca5769c4daa8cf0d89ca3e8ab3ad33322944f64b47747af5333f8459f48d83b111ce26cf319c1ddf9188b651618590396ef476263da85d2f1bc744d079a46fec13e1a7d42e44769806d8fe3a318825c22aa8;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8c792dda506c9cc1c2a53689ff791dc24d3e47ae53a9ea27d624d56e133e5ca4aab5ea03d5b75c003ec4c84637ae332a258c1efa68ffaa96e4670f161d5188dcd5e2fb3ecefa7089dd954d8a81dc487dbf2e69ac79264477954e5fdd2de330e355a2;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4ce123452f6a4b8a07ea3dda713baf7ab0162b4a865939242fa8e4e9e76b3ebade6578c121dfd4b9581ff744f0cf1aed4f894d4864e210eac07a33486ca49c32df1ed7c4ed9333af674b00bcf750d6a37752b14d0beb7598cf313ff9d2e3195570d5;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h111ffeca390b10c198ca40ddbc11e73af64f103f7dd6dee969ae4d86ec299f3e2e32bbac6651598e151d70cfb781e987886d994ba5730df45a6cf9e7318f94757ed9c9c5ddab09bfd18428a2c3149dc106e058b80d97e957fd128c1cb832fbf7f6c3;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7db0fbe7e1e9c49a23f04a607f012000eedea9f2dfbd0ff6b4813cb465f2eb85170564bc112c9d01d77e57f5ee8da67fd9c907956a01aff8688b14d4229a115f16b093da1409fffaa0516f710f0225c9097e9fad0c982f4ed47e67c9168745a3f1e3;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hebd065c9a8b0bb09631151844a974424784dbac265981b696b862eb9a2ee1012c84ace92f85dd88ae195f0a4c29969a37bb6659a03f751a368cba288ad1743e9fa8f882167fb43929402bdf1370513637fe8a27e026785d76c1948e6b88b5962a67f;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h99e351346c55dd38230f46b7072f0b66a84e773d19fc26ce3fc2d83fcc8515593d893b6e9b57fb121585de3c7467731b508f4752baba991b7eeb846cd85b82a578ee0b29321e5db57baa5bd96137cd1d213693cc15c7b0382b9450f4e5a5ad46c593;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7447ced52b6c1c91cecaa5be2af0f85e0ac6ff11a3d99583fd7aabe746fa508dbe30a7a2733f4e95db811bedb9e3b6cc9262881612f572fd8e2c0c74b4b4e7b2ad5b79687eb8257c0e233e29384e50be6aed6cc35868318690fcdb6f323a658b4b02;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4248ab2a3dcd50fcc9672ee570553a8b9be0f17dc29af1e06876311a4ac7d9ec292c7f5d33b7d6ec1ca76c6f90d0c5b30f420576d6f615c5ef7dbafd12c5965050cd31ad90c08baa58eac2d1239e5b792180256ede84beaf1e11517110f44aaa8a57;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8e648b5e1189c4151df3d028b26acae7062d925923fcc33c9680e5c3675a520775ce160f6ede0472568cb842621e6009f30ba7e0cbef93e9975c4db2e95f7bc5f7c0660ce652be1e879d7ff4757165b6f4084669f2f61c1130dd60a6edd2700e6de0;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1fb72e48c7b28791640d59302bd858be6d021d896873e7260760fcaffdf99463cc32960de5c8961d7a414bb487e42959975d0e83a67d1c97545091d784f7959234f74a0e8acba581bc59d479b5f21275feba4afff851ad0868921ddb89ca1d2aa631;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbe32ea03806f4c2a99caa6aebc2f19bc5b0c343eeefe86d24f9e7286810b3ef144614a1f336d52848a39da49c58030232f7c9fecf63bf76a96d57c13341beef47f1977d54e7e2fab1e24e43904c6e39c0a4b6150062fb65a3b9be1cd9eba8f0fe01;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc2b87481975009f96999add1fb2b82a83406cf011640b98ba70674b347e59744a8360d35f269709d86c0c7ccffeba69173d99272462b769a636024baff507f94808a34cafc290326b45ce3fd2469e76e35741543fd8fac5df28fa23172c0ade12966;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hde687af4b8138cc3f4c6d854748296563505a60496975e13c603d29675ed318d4024a87e577cb243470f9c7d39ac9e04f139b8a4c8d109195534797ec574745f7b7f9c08c10901309b9b4573e327f3afa3dc283b5c3de974da942fce42635faaa199;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'haa904197c4d1943fc01604cb41a86c943fb4cbb176ed93c81078d09fe6dc3d1a4574696eea8c130ebbd111952bb5d23889302c7af4e4adac01ebe3a178f4d5a4341d207f9c53ac4b21a752a155857a176f473af275c4bccf468ca89e5ed13fd68421;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h322fdcdf1bfc284f15621bc7a5fe716d93c28d2c9cb5cff33bc9b298da91cdac68a41982fb5b6d055f043c85deb3d3a9c62b51d936b6a09d852fec3d81b7055a48eab40e7a2d75c7d7f4958dbeb0c48d84b538117a5b54f238b79aff2be6118311d8;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h111adc4f9bfe944f073be3c8b5c22e5108f7127a2fa4437d153dda52ecf6a375a740a26e09d9f40614d790009e32704d101dcda7bd781e2d32f552f3a785b3ee6bfec1597d49488af583072fb47efd57bec053047d742af6c0b7f23976a0fd98e969;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb9d26712cec45f12dbaa88e395f1891c51bc14882237df452b076f2283a60a42d3dcb08e31e55d60d7ba206cd690c9a6da5b44fd99cc9e27fc791c48608193d9f894c5d477aa1da942a9da34600f39e89d82e0b3374f77378445c4e10d493b9cbb51;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he5065b37b27964e2c14253dd153fafd438be7ff1c59e0c36e0d114d2bc899ca93be485080e78218fb9f2fa193509bdb0e4385a351a379b8a3b44828339a2a47547a69e7a3916a7833abeb1c5882b89c3191fb9564b6047309992e9b333f4746f0d12;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h66a326c47f0eb828dde3c9a2347e8a5e374a78115c1931a2095fd95c66169e21402bd07285c3bc2fd2fbc02b0307d9056b8f6f5d96edd2047bff46e1803d3b93b987014c4bc4e114ad17db57231351796a8021e897374b511047c9a06612c73c8717;
        #1
        $finish();
    end
endmodule
