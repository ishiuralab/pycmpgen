module testbench();
    reg [9:0] src0;
    reg [9:0] src1;
    reg [9:0] src2;
    reg [9:0] src3;
    reg [9:0] src4;
    reg [9:0] src5;
    reg [9:0] src6;
    reg [9:0] src7;
    reg [9:0] src8;
    reg [9:0] src9;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [13:0] srcsum;
    wire [13:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9])<<9);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h0;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfffffffffffffffffffffffff;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2599511db2090a783d77a8422;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3ac99deeef1c3a604cf969e6d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc18eea0351fa8ffdd1c7a54c0;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1a0aa476f45af56b2efc59b99;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf2be02180442fe1e1988c1784;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc370ee12b20f7c10e05c35acf;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7593b738e0cb1c91994f24f4;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4b993c8bdca1b8da1ab8cf406;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbe0cbaa13e0c08f998a7dd9f9;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h46dfad2b5835d192d524d4db1;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4ee11b442bc36f87c9fa983e5;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc58e8f194746fb9750862098a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4fe7b268c3b634097876602f0;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h78b3fa15769f3dc63ca28a586;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1e966b887f20848ef94dc71de;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7899c151ce12392aa4e18834a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hcb07d3778e90db7d1cd07b013;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5322f6630dfba5b37158994ff;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5f9b856f478b1a7bbfecf479c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7d13a8209201d1a1c7bee5c32;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hde528e053ef33aec0bef155ef;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h329b4d648ee21e440e2e3a637;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf28cda9f52df3d43fd147f008;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbdb7a50dbfb73b9ab8140732b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2ba089cb2524ff20c47e77539;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h29332af8159669b130b18fc1f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h62b4a2c0554929639a5b0f6ca;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h476e4a749afcdf57dd5dc6ae8;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h79c453173e432e779e30f1aca;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h82a888fc71535fb8285be4ad7;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5e489b47797a407ef79089bba;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hce0dadabe5fbb1d124b30b345;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h82e2caf0c51a48e37224a7541;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9e8048ed1bec4e547a9ff762d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb67bf6179c4d6880ebd468cda;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1ad707a2f26224cbbf81d7d38;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5e19c16e29a95f6d806deb225;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd0506f61ba16cdcb49a546c28;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hcbc6874aae6dd29977c28df2d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he508356b8f032afc3672788e1;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he54edd65138f036587d23945f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd20bb6413f927408f5006155b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfc6ed6ae1ee2c129671e371e3;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4a7f33e80838029644d9cbb1f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h411a47aec3e476de899a83937;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h73482d0f1c1a15736185bce10;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb745aaa0c4e367550409a6cf8;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfed17b8ec978ed27198ca78a0;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfa162b9328ca569f818ae75ed;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7f80fa46e315a833bea12fac4;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha8a4a79ac25533bc39b8bd32a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1ca5ad52f88f810a020fdad64;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h470688231ac32fb3af16515c4;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf4a37ad6839fd8d8190f3e7d3;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hcac7fccd387af0679d5459da6;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h67f2da0fd57eae85edbb81614;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h940fc00e3625f6ee593c12392;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h423457c90e1a34c2fba97b924;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5072cc533164a5c470fc675f6;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfd47a04eb6e21538b27fd191;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5aa80d623df90bc8cd5f1b474;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h97e854b7004a888beeb81f60a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha3055b515b58c797bebc8a021;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hab15c6a8f944c16c90506c971;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7477f559c4634065dae7160cc;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb87a862b7d78e9906ee0a7589;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc8e1d0041b5d6d4e025293934;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha688ee84f074aabae5d3196c7;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd70766fb0e63e1079e0c67e29;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he57a78bc54b9e1502ddf230a9;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdd13e891df1dcf9b712145bd2;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he0303bf8f4dbe6bc43d77f404;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2c464413122689b4642d51ca1;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf0500b1a8e9ad713211d450c9;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h794aabfc62fae0a21808a9397;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5edef5b01b469943668c87da7;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h851c805666a0686ba1dda8d49;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6e5448f48d50f35d6c606b54c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2e59abd8f613c9542f1308739;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hda90d745651a29bddcd82683e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4bcb6ea779173fd11ad2659a6;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7b05d66f846cc665f9610e5d4;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h74a973d5d6d34153ad9efe568;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf28d101c0e8d93ef256bfa727;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc6d0c5d49dc130a1127f8136f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'habccd80a4b93c129d1b97700e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h52973be0e9bd63026e2eb5745;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2dfe86128b487667ec19e1345;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3bd7fa1b33b46a60366a879ea;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdd855e6f9760521a0a2111166;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfe6da23a17f39762ccd84b91a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdbcca165aa9ff05a9e974bd12;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h21ceb4dbc7869909d6cc544be;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h41d630cbe72da7161d0efcfdc;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb32fc52ca86ce2da81ca225d5;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he7374187ff063524e0827a5d0;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h28c52c35b5cce295500beb8b2;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha67aaf95e228a7f19c2df8a77;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h360e89409b638886c4d6d19f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h76c6b83816b755c803b70bf2e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc5fc74ca21a940711778bc6d3;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he0b50426b598b23370f88786e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h22709f859144d7584fcc80339;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8e17ada3d2e91e8cb534c89d7;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1b81487cff6f132ff553da230;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfa334bf2528bad22b4edf8587;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdefdb2e89e2f1027143b0fba5;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h946f34f7bfb70920066dd21f8;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb0bf38c31bd2117a142f71654;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h956034ff1e7c63e12a8cddd85;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha2ed5ab89e09aa8f556ddc399;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4419ea4dc9d9f6c453af8940e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h84c3654b98a941aabea6d8dda;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha25822483449461c9fbf4c945;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb0d93fd929bba0f1e6c6877c1;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h41d057b23e20ba82852a99e8d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc3d7db2f9a124976e86126d5f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbfd6cc60f1d067027ce1885c3;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfd8fc0afff883ac3f9f7540a5;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h89f92e91465749cbae0f4cead;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdd2f38ab355152a486588c36c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6d7760362baa71e1b11549946;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h650bccb3f64e2ec345abd085f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha0a0c0a654e33a0db435cb5b5;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7aa164cb7db3eff7cab9a6d3b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha560a8ee07c8b78ec52176bda;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6a87bd52092d1d92198bc6db4;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h26de6eb4196ed37ea0ca77935;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h758f53a1624d13568811199a2;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc881d54ff70911e52b699cb0e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4b6660275799dd5feed0532af;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'haa401c6d13ff2b6ee6e3af2c6;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdd4b8a01e245e4b0fbc4b02d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5a7bb4516295d13a53c0ee82;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7492998e09a8acbc7e64a6a00;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc36cc96dca10ef90757546b9c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8220e21242c485c9fafbf5438;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb53b12504d587bd36377caba6;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hcee6690214c955eb5cd35a522;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdcdfcb89d5ff7b4cb6dfd2f99;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb96c23f30272be832f16a4830;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h26d4ce683f77c26703c0a8188;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he2e4be1c8cbb29f2feffe6b4a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3d72c7737227e975c60bdf2ad;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h39d12ada1bbac7924e4af62d3;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2c920676f10256a207f0bf8ea;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1547fe477d5a0b0244a87b046;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h10ec99aded206424731661cea;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6f8ef8e23255661351f1781;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb0f5a8cca6d7ebdde198154eb;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h49fb946fb7ea39cc7e11fcd1a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5ec6a00e78f9029437ad17849;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3d29bf6a8bd13a60218fa6def;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5b7a38b30f6933783741c8a87;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he4b40adac37f57af80a55eff3;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h19fa7bcec2e7e3739bf777431;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf0733b43ef4ef989d5e5403df;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h295fc37813909dbe7919b2014;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6163ece0e0ad86cfb780bc233;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdfed8165221e98cec3dbdc1cf;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7b24ec9f43e5f15e591f6d1ae;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h73f9a2178ffbe82b105b961cf;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hcfec7105f4fffb91bd7e935cb;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd79d09bc27e0a0555346d30ec;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdd5fc566a5e4d6d5d3f85f421;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha694acf9938e89c682991c6ac;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h35977291056e87b68b70be616;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h32c24c1d6f13bada9da99a22e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9313181594f167519b2df6e6b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'had0380de37d7812353cf38cce;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h17c3069198bdc350f3696bf8c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he13e7e5422952e6d5847f76a9;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf7f6418e1de9dd53d65b2f999;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hca372c7c6f6fc7069938284ab;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h82226a137d5177055a03ad283;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h424b27711f385696ac296e7f8;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hcdd3ade6f1e1d11274a37d26a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5a6cfe16c8c4d34e021373be3;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfafd3e345f6a59a68b99b2df0;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2dd8f7bed7e437e750a624841;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbcfd4889ce1f8b49ede923dcb;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3890b04d492adc428045d2512;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc371c103d71f25ee7c53bf238;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h32acf9dc23cc30a53b4442d1b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8cff14933dd172210fdca6374;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1f168591999df84148c328ea8;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha62959e51e570a93054cc1c14;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hccffc2f64c4d9ca0dc2e90536;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5c25cff680273ae131812508a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h51f27f98712e4557a07f59032;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbc22d8423f3b85879e6e64e4e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4330bc2c0b9f0fae8dc523ad7;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf398dbe3be7cae2706cfb4c6a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h72a900995db6b0336f0605c48;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc12c0dc03b9947defd6a3a72d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h46b903b76f4f2266e89ea30d3;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd4a69e55debe7811db4f2d508;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hccb9d43c0ddd8004f14fbe4fa;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5501a39b65ce15fa35bd492fd;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd31900864ae80e211f5d12686;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb84bc048f4cc83477f006404b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd8e3436eb51c667a528498201;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8165ee68c5f0b198f30d51c6c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h974ce23a9efecb7e8c2dcd6fa;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd9bb881807a4dd86287e7bb92;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3dec91a7a0e9adfee542980a9;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7655d913bb7b3154d6b43051a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h13049fabd59023922d5c76f89;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5dda829e3b806e9757abc5a8c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he5b0ede6ce9aa1a68a0a9ae2c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc3c085bf59ae43d182168f6c0;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h820d1898a2662d6f027efe118;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h75ac6b4c9bbc9474afa00885a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha427e18a89f93a94b7ca2f28a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc82076649118c1ace0c7cc5f9;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9a373c47f97c1cc1343c92f4f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hab67b068d6969145422fc5fcf;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2a9f573649c312a646bfe98a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h60ec755a1bdfe7fe19d153c76;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3cc6361ec3f769f793d987cfb;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h36b337bc7c1aeb8fde13195dd;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h259185a5c52226c030e93dbde;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h61ad8c53fc546539b049959fd;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf3f377ca08190e467681c009f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5cdc19c63cc9454e97f4ebf38;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9cc99e193915618a72a3ad1d6;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1d045a99959d8cbf81a2ed901;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8306312a89731075b3d9c193b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc9f3f72059eabcca3b7ea5144;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha2ae9bd78276d4f7963283820;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h23a1026b178a762ee2efc908a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbdb4562e515a7fb5ae82f654e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8780c98fa4d9b41fed36ed5c5;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h25e935c1d684e917b94b4efbb;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8e5a149c5f29fe4f3ca5938c3;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3484cd930ea035dc231c6e23c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h68531b0cee5a0e2edd23f3d1e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2c740c41a76174f4eeec42a6c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h39f9e820ad7fae9886efd5a1a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h214fbb187adcb04348d3a794f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he6a9e942104feefc5529a0959;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdba17e1886714e7cb35f38a62;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc3f9dc75f037877dbecce533a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h977446f38b7fc6a92983e3870;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h403e7fc5164a824a95192adfd;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf60bfdd2beab5915227795b10;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h770998e2b2200d01f9525de55;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc88258433f4dd49daad16993b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfcbd60198d1deaba2252fed8f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he99032fd11859dbb9f02a7d6a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h37b5fc8f5913f6a1259c1c69;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h82c7e5eae9e2ca8ae59fdd81e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h432f5e65fc1c3783b435c4167;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hcbf5160eb6616d17fc6afc2d8;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc934c84e28fd77147ba5018c1;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2b5f5eacbe1a2da077ad930af;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5091b28ad51509a54208266f1;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd7833d9d245b79a92e71e9627;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8d988e6a5fb8a211b55122033;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc790444947cf8ec4387587d2;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9c2201fc0c9252e65140e571f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h25bb8ec5e7f2d65ebbc6e0e9;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb56ae003606e9460974a2ebc7;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he1c65fdf6e480cb5cb31cad0d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h989f4519e49e791a5ba1a1f06;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h893a770a499e96b8f99a879bc;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9fc33c4a602d17e8f47875422;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h55468e2d1c73d3a9454f0c8e1;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbdd50f052b14012d5b4362b3c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8fcfcfc512549890f9279c23;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he296f7d656d2113cbd94304ed;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbb42af8dff2bb4ba6eeb28bf6;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hcaf94aff5e9eb012310ac96ce;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h63967e4ab3e2883d5c4a50b13;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h20661c2723b5e5cd942049db;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h80f6399a9ff5cfc570297f229;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h72b38452589218e0868e225e4;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h90bfff35d6aabc755e4630ae8;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf83cd7712bcbef074e4201a01;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hae44c65ad4ce2964a452dfda9;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h399fb6dbe492a21751d4c24fa;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7aa18cb7b6f2564539f62929e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'heb633de45fe358a627126ee3e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbd181ef4a29a5f81771c14105;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h172f7134112c7cb61a75f50de;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he12a93a0b66880efdd562b75f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3cbb15dcc0202c206a32b42d2;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h32a6b5a2fa304d63b863bc424;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h788de1e69f55df93c28cdc1e3;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h11453fa5f6800978acb27345d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7aac78da7938028c430ae087d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd42f63491f8dc6a6e3fabdf16;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb4a561b7a34cf5dada6272656;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h75004c237a9f442638256ec3;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha6f952873fc60f442ca43d43e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9f4275dac53ff77fae42d9619;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hba8e846c54049f9da12741df8;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfb5b0d3804e6e02a591ddbb5b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6d2a430db127b355106718124;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8b469122581f83e2e62371fb4;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha5c73db2e4e84e1a0f81e91d5;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h594f66665ed1b28be4a7701d6;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc8e811774e60b040afebd4c0d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h91c5e2ef7650992444e8b79a0;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h24da798e62513ba2468e1bcf3;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h55529358f8d32339b92dfd0f2;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd8592ea6dba9fe3d0a726e982;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h11cb56ff767ac11d712e37ee2;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h57b83c8fb199ddbfe46612de5;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'habe6ba41777f978645447a53e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1d62c7d39f95bab59640faad2;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h34891e71f0c60785c72f8c2a8;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7147c8954cbd5f98605047733;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc3f01c0be21ec281546f66621;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h750b037ea0f55f3491b1b750a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha57ff1a8ff3bfaccbf9f4c4fd;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9b8b0d18b2b745583ab753168;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he482467584706c226a7a1be7e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9b0c49a27344f30af132198df;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha864f9f4b10415fdec6340352;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8c7ba48e5fb190e852564ed09;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h901e90e06f819adc85c596eb2;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h12a5f72e12c2d996b2ddd500c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h44a293fbe15e3eff2127f2e02;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hcdb7fa74b00202b9c9b45be78;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he8f701102b4a49c5a7ea5404c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7eb95fe937bf10fab667308ae;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1290b520a54eb1df462598638;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h23462b1039a27cc643bf525f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9f1526ec70d0ad6a44c9783b5;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h875996df79433e97b85bcd5bf;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5459e9deb003678270274b48b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h19c57f2d3a6f09f03d5389e4;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h93d2da791ba063525549141dc;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he71e0d50bcef17f977f2abc8a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h31af356cc1518d98cdeacc02a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbe5670610d2af6eddc886ce35;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3fea1a886aaa49881563c5707;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6f060dce1ee557128e4daccaa;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8eb166c7a1657c10763259351;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1bce160a86880e788dc961c5c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf2c307b281f8cf1670cdaf29e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h494ee8ac3844bb10887789cdf;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5dbf15bbbeb7803b5fc144cb1;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbc4afab18aa8cd348e29d2956;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3b28fa040d8d7ad066ef0de64;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd8770e44987dd85afa796762f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h70c20f320b010fc53cd6659ad;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h558fcfcf6b3e7dad11c60d9a5;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc91153da4b19827f6ccde1ebe;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7cd243d49da20f9954158890b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9d9fdced8bb27d42dc6f00a62;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h78503c69cacd58a445ce116e7;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc75390f594698ed5e31cfbf7;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h436949b530e5926e74d5fa4d9;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h93670e14346fddbe2007f12d8;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdd16e4facc54f6b0e627c7914;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha425f811db5611c8e38dc667d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6177d13a1acf6d8f2917dc6a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc75c99837579a126896a11b65;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8d7d9b7d9a7c3828a57c6ff0e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2e128f194a8fd8014dfac9821;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha8209c135bd9fcd5b8d1b40a9;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h37119230e81d78a0021876b26;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1258d1c5769654711012939f8;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h158989e146f7bb2c43704489f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h32fd701e0a0f356705a0cc657;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h89009f029b748a6dd18085213;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hddb27694cccd7903c09b258d9;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdde5c29cf132e2ed30deea621;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9dceab52f4638a7c8e38d5a75;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf55fbd6fd937e3628885ba32d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7e2e56dca5c84f0532c035d97;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd2698d92a2cdb144dfaf085c2;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h753b7d2c87d8313b899180059;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb282dc1b5442566ef2c091b63;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h72a33b58f13c549c1fbbfe917;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3e51ddbb6cd98cfd68e1bfb48;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he2bad8af4f0bcac6d3a52c6ad;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2ac8830250d0da0e751b63eb;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h715fd4b088e58bb2c7bb1d9d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h49c34caeb03e453ced2a2767a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc771c9ae261aa65f5784d9cbe;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h55d5b0ceb0d40b81dd408e365;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h921da8afc07362e298c2fd6b8;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb390ab37669ee702544921e8d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbb51c2fa0e86e1ef002e9c14a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4eed997bcb6ba8f7ce5a068d1;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9f0e955336bb13f4c22342fb6;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5fd494810cd86223a98cfff21;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h460f9903db4bbad5f63982e00;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbe9b32f2df69acfa2b83c148e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9057adf9ab1225c2fc385cb80;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1579b1b60393345a74a543a91;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfd0978a87aa0bcf67e6c308ae;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hda61c1ef69f72ffac684c6801;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h516e920677d79c3ac3a142ecd;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3200208a475beb9f8a4daea6e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd03547b6ada742143f87373d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd8d0a9e4edc246e285d8ce676;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h60424722ee6420cd3bcf8f43e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc46200ca39d78241aca7182b6;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8fa4db7f12991f264315709a3;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hac2cf809fbe0a91368edba2ae;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h66e9b7876380cb200a07b9177;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h59c2e7d731321fd1066b972bd;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf6639a88e30831e7d4241becc;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h14705511ed245756eeb3294bc;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8057537823318768c55edfca5;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h74bdd35fd6cef922f2383ae34;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h725fe533dbe4a8df7194ff7fc;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h702317d314703cddad900c417;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4672a5f657e8dcbe1f5a07db4;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8c59c6647043b173d4b405d6e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3d7203282a556115fb285e6fe;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h354364ad13ed40b044d6c9a6d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h514ee0dd9a8a8051d779cb1a1;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3c1effac596d3abc675e6bf99;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h16e6eba46238ae381c86e36d3;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'heebd0da3feba6faec3c7e7772;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha1e8bd778cbfe60f9f41a6b95;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5a34c3c1d06a4e53af8f36263;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h270b93cb437dd34aafec1a7ad;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc9217485eb7b4b2da3f8e268a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h33f606b59383e21f77d12b619;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h39101410cb1d31689755c40a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h35fccd3005945efa9dd3f5e44;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3760b67f5d15ae5de754e2abf;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h61f6eb48fc1ad29258f93d4ae;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6eb23619f2a46daa3dea73ca4;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfac56054c88c385efb54f3f7c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hcad239bebcfd4d7ce5c095b2f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he7400287e41e85bb0605cbfdf;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9af9bf04cdb2dff6f9d77355;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h530349648208c92322c9d7e2d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd8df1cd0b91437fd4c6a8130f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5e074d827b44bea80f5110f2c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h32f4857d198d407f23afad4c6;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h764748999742b71e1dae8914d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h14d941fb1ada143bbf6a13ecb;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hec9a4172e7a79ff56d0b6fd13;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h810e0c32fdf11b3ac9c5ef5ea;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h630745b0e24eab85a9df14ce3;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h63a05a220470a6d063f8ae9d3;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h189901b7621dcab7d8bf4ec58;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h160061c6760f10d7796ac8b54;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb85e4f412de66f858ab81ca8a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf9b0c1217a388c5adc326a933;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h240a1a228b005bb0eda00612d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h210beb35bf59ef5879f566bf8;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he92b34413c9c878883890851d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc643020c256239064f5e742b7;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfa08cb2a91f5513651afa4914;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hef6275e16cce2295faf9c65f3;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'haa5925c9c359ad558b5e5695b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2e90d60255ba682d088638561;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he3c073fb49cdc1733becd525;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha7ec723ce48e1298ed4d6051d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3b6b2c47ea583b09cdecc2d9d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hec3a018c7445b6388b548de3;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8b01ca2e611a9ba3fb327b3b9;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8a912b1a114241fc56f6bd422;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7277fdd196d5c9e6812e7aba2;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8df1674444fd96ebf0e09113f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9fa8887d254bea7b2a8004244;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6e5fbd776399460cdaea2faf8;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc5be186be298201ce5bb4406e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6d59cf00c07539dab6e9dc35d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hafe732dc4f95b38b25fe8f80c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hddac41c4bb34795e70c946517;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha881084c85ee6c73412f5ad20;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8ff64cbd37363c8b6ec02f3b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbee4ee297f214c79686060f14;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9ddb29abca93a36c2a117dbfc;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc1124b5aae11747bcca07d017;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hee730f5337a723f24ddea2f23;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h29e3872904ebe79ecd6e1a290;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h923b39fe4897b0d7bb09d10e1;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he470ee99519d2286a06d32166;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbb9765357083c5e255d7602ee;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4ab367d2fa3610241f6142ec2;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h273186320a9f7a0c0be062bbf;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb3ad605a5769910a59388eb3e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h431d3cba3e30af7c7ac6b8d22;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h814954da79e56378052734514;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hcfa395b08f9ba453726c78ab4;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h70c049661d5c61c83e32db27f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6a1b31d1aa34466586ae3ee99;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3ab38aa2684aecd01a1ce83b4;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd5894abcb25c93ed3e5e39310;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h76d68cd50dfb33a20f38fbfcf;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf76deba00870e1e656230353d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc9e8a4eca4ab02b1591743f58;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfc34faa9601c625db7367837c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf25ff390aa5cae9e64cf5e5c3;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hef8bdc56705734a2265219cd9;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h54f5cd30af0b24b44a89f769c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h38ef3e6499f199d7f4aa41103;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfcbf1625891df3f54a58c6c54;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hff3d25bc86c47e0334361eac5;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf64114a52f0039d58d85ba8be;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h95933d709662e6bebce1bb2d3;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h53cf8d828ca1ef5776a0b082a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8e0d261f41524ad711f90ebea;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hed9b35a27568df8c0ed073f4f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h670fa021776653a95f389722;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h449345f3c5886272bc0841fc;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h30759be0da71306f4cc81d8e2;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h51e5cf63840c16d2ba66f1e95;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb4dd46b8be6c1c1fee397aa0d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h197f3107eca1052d0686a892c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h29101b73addaa2b35b09e7748;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h827ccca85a42f905dfad821f7;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h644e72d648a2c5aa3a76c0a9f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha1c2a1eb8627ca23485344e7;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb6b6aff7a5a10cde8d5c5f85b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h579a97e40375d09cbb13f93c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf50f54a317b93b6ed6cd46036;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h16479370b8a69a457d66e761f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'haa3e61b58f6ee808e71db18ae;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h618188d01709b9b17e70b890e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb2d4b3d4a251798a6bc63da3;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4e018de81d28b6cd63838e157;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he1739a9a0e63389765e52986e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc1c4eae81e6872605ef6ed0ab;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3a2e3335c32129570b81b6f76;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h41c3bdccefc9b85576401b04f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc46af10632c5fbae176c9358a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2adaca278def485b84ddd670;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5ebfdf2669fad1ad1da409edf;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he7044c9438bf70b1d17b8d8a7;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf83c20c80f686c1e6adccbad9;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb9f9f9e7a960dc83f2f5084a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hab56ac5f8f6ccf66c775b6545;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h800071b6e374fff54e922286c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2e09b5050fcb8d53e859a9042;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h22ac4d3f701b5c07066bd4d42;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1a459a13a2f394d94c0ed2478;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h67cc190061a085d8f77fe7b97;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb240cbe124552184010f0ad62;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he1e7b5f0475f2c88e22155502;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h89ffd27c62cdbdb2caf84a699;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8fb0ca1a7e52efedad3526d67;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5e1dab66d84e473b61965617a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7a5d86046a5ad000946f6d879;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd049cb3fb53afbb8c1995bbd1;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc8687250249fb421987ec5b7;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h208fd02549e583eb03d07a56b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7eb6596b09803f10afcba83f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h48da8a41d2ad1a0f81f36b7b6;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf02774792e8c3266bbad1eda9;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hacc469ba9f957fa3a12ad7399;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha1a1985736f2cd24d5a9bab78;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd6caa107198799b8d5f2678c6;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha20fe2b76eb5888760a6b80a6;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h13b6ae5eca0027f74f7f27a15;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h90e214f70e22a212e68dad5a3;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3f13a8fe7065581bb008e5b55;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf68ceb04aa0729cd38d069cd1;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdf071bfb2613d643c1bc97f5d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb626bb883d89480b9f276f27b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he6ff5dce2d5f7c08266bb389;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbcdcb62bc52e9b036910770f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hddb421c8be7ea728013a9ae9;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h56aa672d2b412c47862d63ba8;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb40788ff8cd441feb0cea7163;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he517a185ab12e51c4cf45292f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h730695dc69880c888789f9c14;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hac242253d9060809ddf3e8666;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h333222f0e41fa7983f8fbf210;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbd7e9586e73d5e2c443eed63f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h372463e6b3c315170fe4b1a2;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he699cf7ed987e0f0d46c8bbfd;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7cbd3cb8994c89e19099d4b67;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7fa80ec61edfae618d3f44c60;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2fff571b21216bc9c886b4f7e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'heff12976f08ffe5b68f481c7c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he1a509498ec16d478c0a08c9;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h99b081de87d863fcd4d8e2341;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2a49e383065b91548bdc2bf4f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h957c3c730fb3705ae266b2448;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9107076f3b307a4e5cdd277e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h257e0e1f5e812a1d6fe15009e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5438c522519b5779248af12d4;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h36dcf5f4dcbb71669fde65297;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3163dc7b65ee88587529f920d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h94b51eb4120aad42b4c657908;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbe0cccb82650912773383bd71;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2ad971ae346ca542916038060;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h18a481e0451c3bfc233f37a2;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4a0bb704c7c1d7e888de78130;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb3d67809f86ebbd760d969365;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2295ec7f2cc111c44f775063e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h68f154fb45ed460f1d87129d2;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he48a42f85ceebb228e38788c1;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha8f47bc7ec6cee70c364facad;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7f8246f00542323855e6c0cc9;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h17a5627ecf2259f50b3d9f6c1;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7474c3dbac97325ca4cace2fe;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbbc8c82416032b4fadcfcb760;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6708c2ee31a3298ad296c54bf;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h42452cb49f9cd59717521a47b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7e6f2772aecb4680f75de78c7;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd74f703b7f42dec47c06a830a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfacb0be35f95bb738a090dc09;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfd50c5ca0b4922480904372b4;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha1fd06f50b73a2a5ed9fd57c1;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h91ea8e2974b83cfef76ae6bec;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h320789dccf26f5f13273d4402;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hcc935bd385e0fa38bf74ad85;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he927df37e641b65d1eba3b888;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h65966fe003c9d70c231d56d8d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd13e3b259bc84934445bab14c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc8e6cfc5c11902cdc0fc6d046;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h583ba0c62c19e34a9fc1a95d3;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hcf44b6fa23d2e50a64e072170;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc54a6b1cb35ec97b3bd6bceb3;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h21d6d5c1d44027cb64a3c9f3b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'habe13c06bb185c538f561479;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf748972a1c55fce92b296ec98;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8d861596c1591df917040969a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbef53b4480c7c7b232d9e6414;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc3db0006dbea07cfba6b2167;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hcb0b2a168a58b0feacbe24a34;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h661cf83e41c6b5b5aef8df157;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5520e3a724ab6779841957844;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfcfb9bc7c1c5317e858000e66;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc0342d03b20f356d42db823f8;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd0534fbd1f3da1ff002354334;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb8db55f7ac897cb0e01f60a69;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdc25efb1da0e2d9cd3314284a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha5848ecabbce121ba0dd41e0d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4fba86d4fa582ddd566649d01;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hce69961780a65c32d144a8e4f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8098544ae16278bd8cebe69b3;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h38c777716a2292b9a76e4e92b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf21eb75f040e58d16624e87ec;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd1a96e38eb3e8632d2d0d4a8a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha6425f7d973a5731c8e13528a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hebd9f716990fa39dca8925f3c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdfd468ffd96468d8e064da33f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h705fafe84a1afc1684d96174d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8cdfd7786591d5f89dcafd66a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1f93d952a54537dc50cb8ef48;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h93bd0b04d3122e292b1c65585;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h59cac83899e95e3cee6786b80;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb1158d3a0fc51deeaab646f59;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6bd02276568f6085d44067eff;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6ac447d2aae799637934fcdb0;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha5dd8b736564ebeacd42d1ffb;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3e7f71359b6f08a2d562a6495;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hccc354e49a13fa13d8f38b341;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8c006e502e960678c3b9492d6;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd01af3bb950674dc4e1d913d1;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc3e06b1101d7026fbc86ae61b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2907936a2c75f68728476bef4;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h87ac47a029d2f495e4b9b644f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha319bd75fad3bea4f22745cbc;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8fcc7683c49d0cefbc62b3a38;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb0d3055b36d213891e1a8d399;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbb00861a9d9eabdc80ce53804;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hccb60b99dd1d2d3340df181aa;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h321229b40dd9b665496aa0255;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h939afa1fd35a1805d451dc11;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h38c716a9b0248030ac7bac933;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9fa2333f99e33f3d6085ef5c2;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h98ddbcc08184797b0088ee40c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbfae6219e7d9a486d5410009b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h21b8877ae0a4cb2707d02371d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h907dca48800fde300ad7cfbe9;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3d29e195f6762ab41b99204f5;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6b89c63093c4c9b760a3fa67a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbfdf6eb1c30ea923831d01470;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h84ca81db2cdfaec75871d69d2;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbe903a2102dc1601b64804207;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h13c221cba685cd874af032253;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8ce887d2b01dd3d841d6bbd8c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9e782da47a1f29ed854240936;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc992011dc47e0ec8df0854f32;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hcf9d1329396a927ed7284ffc;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h91c009fd2d68ae2c2277f5e1b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8ba692c4c4cc2467eadbf6b04;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf7372d3a962c3f47eb8e246ca;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6505cb74cf918fa5b9f57bfd4;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h799a594ec05b23d30e1ec58f0;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hda28acb0bdfcf24d1f8854da1;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he880ee8ceaffec0c87c09d214;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he6023a38069212b11b0289a18;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he94a860d403d9ed4a9eb7be0f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h20b8104180410dab86c75c13a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4eb2d8f0b528d421c061dcce7;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h428cf70cf20667f0c1035d39c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb85f9b6e1bad2ef77b9a6b0e5;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf083a37fcb853548e10912efb;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3b90623cbf054e6399c738ae2;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbca08e1452ae94a4bd16c6f7c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3982699171b132e86fb0cfb9a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h115b5cb7ffc8d380a5e40968c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3b3fd93103746c7a5131c1575;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf5252fc79f4de5b7410a5a287;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd04ea972e2d54b0b3c0da07da;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he414ad4de8c563925aca721d8;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6c19657e5c5dfc3ce60a98a2e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2204b6d30a2b4c8a9594360be;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6cd1888dcba8b114d387d104b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6d66b0268febeb1fca6d84865;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9b1ec459f3c8edb908f10beb8;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd16b855d3b551d4df0aebb60c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1e933471613d75e90b18191;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb87837b0348bebb03569e93;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha1155bcd8413ff290e1054f3a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h342522971e4c020be3aa5d3be;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdef0c8ea9a35a29ce30356e04;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8c75294d7e7f033fa7fd3f4c3;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hcc8202e25d9ee0b841a633a8f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h85041ee271dbbc8a354b4136f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h95b2972acc132359d0f7d9ac3;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1ee00a2773262e4f00550c3a4;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdf18a6f8a5cad68e504e84c9d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9adb534f2ebb82baa373e10d5;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9e6f23b6b378014d2ef12cd53;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h760ef23aadf87fe6860e1835;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbc28c07df25bc19c36495a97a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h82f9e638677e728552490560e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h32fc908af02f956f801b1e379;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc0b478b8282162ddd079f4898;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hadeb4031197e67e82d6c2df8f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h25228c5daf66488cbae0943be;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3dc2dc91498900deac4815683;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3da48004cad9662799e5412d0;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h290c2dad3b7dba193a796670b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2a2909e4b1f1f8b9713c76402;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9f67629a1419aa8a06775fe09;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hadf8fc91bf69c642229d5e88c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5de4405adab81e41974a70ae9;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8e8283674d282755a3d2d3540;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1965c951f1223eb9cade010fd;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h57372a5f8d0c8272d4b191177;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h60299ababecf176ed7a35992a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h42b2cf8e56e86ffcdf4ab51ac;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'haec110c73322d74047256967c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h20b9f2d29e93cc5fc4aa7149b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hcdf26048bc6d9302e553a2501;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h803b5d4121fdf3b241330cf84;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6031151f5f59d407dc7e9444b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb5809f7792d316d1a62b4e9f9;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hff071a8105019758bb1a0f6f1;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2b969eafa0c53761e0fe2155b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h67d39a71f7e6717a58af0efb3;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he7105fa010176a9e423918e06;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h68aa589315c3d45a267f1114f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfce014f175922b850ef66e313;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha837b1bcf04f7fe00d471cc80;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'habdc1890e5a4f089e9b665e5c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd79e48bb26ecb8f9d65c74e08;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hecf30dc6c76618fe544558acc;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h62c5fd4ec2c79d019ff2ecae7;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hee8333c81bc4e42fcb2353b3c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8ffaaed1d101dbb423900694e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h93cb256c0ae0a3377e79d96c9;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h958a52a6baacfa51d886cba63;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf65f070dbf880ea8441c2fb3e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h69949abc6e12165be523ec319;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h518e5fcd2fde5641f51f34ec9;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc14ac851d60d01df162944d27;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfe042612d8160716a8b3c3e56;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h887708a154367ee9bb294868e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc5f46ddc43f4a16b9492ea48f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4d9a57827764e67ab655f8e3b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h797fa5f4853b516e04b64bae;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfbd7d507ec42febc7a1757ced;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha1689a35fac43f88f6dfe7e7;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5528b25b97f5643175ce97d22;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8f67ad1876571974b465c7bbd;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he00d8df500e27eda332b9e60d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc0b6a49a69a0e66cfb316dff7;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc4e2e4f4c8673f4c412385026;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hac8ae48e4a6aff0ab45335b7a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'heafbdd431225280d0b952d4f2;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h35b3bc904e9479b6d1136501f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3d889cf59818f0367b31afaca;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf3ab3e8f6d9056493df7b0a32;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4269576f366f3b1f9fa917f50;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdf5e2c8abc3a44df890f613e1;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9c0fc0ce6c3f5eb7288649f84;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5548cb9a217c2ac066162f772;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6825422d472ec64cc5588f159;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha17fa5ed5bc67a936ae019046;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc919532d8847c22bd945f5ef6;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h60621b1ba87fe1491bf2c49c0;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha1ed0d0683c41f348ade6f4f7;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfe465165373f47c5cad85e59e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he838f9eee4c4e3aa173ea2026;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfab043c2630fd7b8c2ab0def2;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd918afe7bea565369b02531ca;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2b8c42cd2fd5e158950b585c3;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb4f0dca9c93c0e93800919d5;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8af973f15a7945647398fbb20;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf055166e467b469551c3eb46a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5fc4e712022cac09f9a81e501;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc4530562879271e9e319a4b5e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hcab9c44216498a574720c7b81;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hcae3fbd23f31d8389a5984ecf;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3cca6cc63b84fb97029ff51c5;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h655a27c47b0012b77da7881a8;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf1116ebd357061b054886bb8c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3ac214faf77a0ea23a6025416;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h823e8265eeb7e0bef8cfec3d9;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h45b6ebf569d9d30a4f888ed83;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9f84463bcf57bc8eb170f0a9e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h609f1e0476f5136950100a95c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3c3fb908183c35dbc317eb4a0;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha9ae88645ab7539538f144bc8;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h23783a66b4da52ea75e4afab7;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he125805af7009af29aebeeaa0;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb0defd579e813ef9c0d240fc2;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha0938627fa849e218613902a9;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6ee88d8c6c8f4a745ed51c713;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he653b34bc743ebc78de0b20d4;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9d32028e4f9b2b44732e747b9;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hafe83d5f6760cda33496d38ed;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8aef6de23d7b7c8e32f0a9ae5;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he7f521a7af6fca3018a7b3268;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb36683dfc4969c90fe6a87a51;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2ee4aa37ae088fd4092fb4b5e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9e2383b934764c867fba30b2;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfae24138648d61dc6441f234c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he7c8541dc1685802653213dad;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb5dfec8d488294ac777433bf0;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3c3cc5c66cf75699c518a3939;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h325cb17704452652fc179e3fb;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h83e9e6ca155bf8098605e7735;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6496819e0d35716f0471ea6e6;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9267547cdced8e2f0dfe4d11e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb27449d3e12acb56b4e140319;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb5c5c153fcc50c1c8c58f6eed;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8a159e7848f99e0e0642bce5e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc57e1f62936ffd7ea3c699d91;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h377265dea40e3a39c44a5c30f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h916306f90e8ec87f66bf98722;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1c5cfca3aa7d9919073761ddd;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1d64d6ad46bca7220de9c27a1;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8c0cd46e442827af524265c18;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h692befb23fb669fa47e1c47a7;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7e29e760574382c00baf3deed;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hef35bd5b8e3df8447c6e32a2f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h438028b0d544e5bb02d42f2f0;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8ad98ac0081438afc3007157d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4206928245d6a6e3a4528935;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h556c5286cea3150f27023a198;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h12e4c8aba53377ba190b12585;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h62d20662dfe05a54a446dc772;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h96f1dcd6cc1646674e1046a6c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd5cced7d8bb719aff9106c756;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9628abf1783290c7b29638462;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h132d05433b62894dac9fcff58;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h75fe1806aad4c0f9891f51678;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfd9839ba02f18968d54fb9d37;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2ff1d7d13bc3731f1d97d102;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8e39caf7358785d56b3ade7e5;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9f62a3ff4e30e77e6e2103da2;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7315106b212612d299e2a800e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5e4fffeb2892e4b8f7c83a47d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he655de3aeae393748524e0c63;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6ec0aece3e1289c94cab42ba9;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hceefcf993406950bed78d7e92;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h27b5cbc80ffc56d611f7e962b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hcd782ec3e78bd32a49fa9c5ab;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfd4b585b3eb5b46d36ea15407;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h22b4c62d755d371488bcda748;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1aedf14a3624aa3cdbb362656;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4e6c9572af36c52938ced769;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1453381925469291538648dd3;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h25086c088f115f29c4c57c6fa;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf3a8f7c4320e0980a5b61bfc9;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3fe2bd00eeb5b8914665e8ee5;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5f3d5e03f71093954ca0c6b1;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h503cb9138f00c4cc13f4aa8fe;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h491937a4aa4a1e2553a76e24a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2819e986a509d7ac9523caef9;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4f0558bb46c976d16d49c847d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h858fd92d845b13b73cc85f1b6;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h34f848dcb91a8cf845153aaae;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8f2090e6090578ffe6a1e7e3e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6b27459b5b1554610401135cd;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc03231e81b3f81679d8a6317b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7d1a12a8d67ea42fad9f03b46;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd0bd7f7016eb1f8b8eaa8a8df;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he342ff5b2ee55fcddd7328854;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1a3d7fe7467b0deb3cd9f9cbc;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd3dbd5975533a1bac6fb3b8e3;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1f7a429033f3847beaad7605d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbd808d9d7cfbefd48b6dc5af7;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h220ca7e2efe4b7c4036a20988;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hde2b6dc7fdee7ea7c5bbd9849;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc3d3aa5f5665bb663d43d0eb7;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h725434a77bf472c889cfc8d8d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h32709f05d96591561290f49b9;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb203006fd6a2798f4f2aea0a5;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3c1c5302679ae238716ab8699;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd8eaeed75370de96a354e2461;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h52edc5691cdecab630300b4b3;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha3b0657925f4b7df3526e7e72;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6bcdaeafe9813eb5eaa1977d4;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc205e1a296e7c164614e1b1ca;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5ce388da63757edc8e52cdcd7;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb3196fc469d7c1ece4adced47;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8eaa6bb16a1f33f74861ca2b0;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc1635c15d22076a5ca5403645;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9bce2faad5fd21c92285436d7;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h32faa94baef1ad5ef46b26d79;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2fdd3ac9a12858eac4b440bf1;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h75b04305762578022b129eb64;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hab5f8e4dde542aacc719417e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2d048ec34c850f59f71976e84;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3a64653e334bcca0c2e320cde;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb042c1560a172c9da477e3650;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h80e646586d39bd8b4644408d7;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he33ddf9509a3d2a1a6ccfc08e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h65d8d3923a06e2c6559bc0de0;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h786ca5784175c8d8fc11afa2d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf0fcdc9a5874996aa810cdbec;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1d312ed37ca562d55e5a4a4b9;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5c3f0db684f5dcb2fa9f8ad56;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha5cd755183f7271752cea4d05;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9a5029823b4e63106974a9e9c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf104f93a79d091404eb02edda;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he538edd3f95933530765af99f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h633ba0d6d5ff20fd24192b9d5;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he1cd14e2f44e31448a8ddb368;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h50546cb9e02ebc91eceac3198;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he1e95cbbadc184681fbd46f2b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he8a44a544d8aa2d0de2bdfbfe;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1a84dd4dbe4d0b373defc0e42;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6dd074ba4700b1e6c240fc555;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha511e06abc8b9438487296692;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd46acfcbfeb575b381af6e718;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3eadce55ca5b15a1964242c0a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h95d3497657b7d6f9741c68c35;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hed54df50d04c29f8b234e6112;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha60b42eaf91c2deb1cdba6d97;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1c983c6ac5b87aec4df58643d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h18eced58ad49694bb12cdffc9;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he0f934fb20c096113e699f11d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbeb89255e9c372ab012808661;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h220be79de05181cb67b38a816;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h981d12d13e134f05ddbddb0a6;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf57651318d3f9aad786351e50;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf9d100ccdaa123160c6de750b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he22c176f3ccafdfda97bd5078;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3bc949eeeb783f4456cdeaffd;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha39c746aeee100a9a7210395a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3ce1e2116e92e132743c02559;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hcbeec03c0401fa1e6bb653c64;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1565207fcac568f50a74a025e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h98d569062d986f6af03a44b3;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'heae10bd66887d3f041f253a2b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h67da9e0fab19c0bc6e59b8c38;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd15dd39a4b01f4b9927c9c287;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5e6c33a5aad5e9bf06c764d6c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfe82a2b2d7764121b93f3631c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h39b95bc94a1be58b958f13c03;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h735fcc063c03592237f5cbfa;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7d8c12f4093e3f06569295b16;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7e002a5ffdd98fc97b871e9ee;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8d3f9eeaa547f4307c9acad68;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5d3bd8e48180f65b7e69e7574;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6ea49f891ec7ce08d487420a4;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf71e4ef93a52c215eff5fddc2;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h72bd3e63afd89ee5cebd72d45;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4ed6fe251eba5b8ec0b73d994;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9c343d82796e470a8eada01b9;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h27f13980427421970397e03c6;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7c0f2cfc57ba9888f0664d0c2;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h35138a550e057add8c4301cb;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5f0f18aa90294e8d6627d752;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2d9b939226f16a5633f40459b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h57ff89b0032b04ea7cefa168;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8faf916b8d4e8c5c056cc3eba;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb070f04c890604e7692d55a63;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha492e2bb0a63bc804bf8ed63a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1a5345bac34d8ebb749f2ffdc;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hecbe875d979b10ad31d73cf09;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf83fe2faded7327f988e18882;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hed50b18dbbc3fdd806c722270;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h70836926d981f0591b72e2fc7;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2b6d543c532262fffea24fd68;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf16f0d32126a448a874be9a88;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h25369fb7f2dd5e77e097653e2;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he388c841085ab4edb7e8a3c46;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb25b756611f6d3404e3c55269;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3ac3514fe69f34941da79f01d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hea0d59d3634fe7d1399afc391;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h565a0d85eb974e50db7b4c442;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h250f9fc031aa4ce7944f855d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h893563223e4939e72e78b4ad9;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he724353f0823537ccee7f181f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2f2d3ee0a694c0a3a088fdf31;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9f9f2a4c9a16c7540307f7ee8;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h78f84d7084c8793f3817487d6;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h81f2737445d708f7a4bf6bb9c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h11a71cc3833ad4645bd3ab723;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h720381c8219b8b069e4faacc;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc32c443006265aa4225f48bf3;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc1a8329bf931b2d78888f59b4;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha69883812a01277d8bcb84f3f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1bf496c14016acf760b330beb;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h98f2b942b9828e3ad24a74275;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1180e42c75a0dd91db81e55f6;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8a1455f7a7cc4a7e55471a319;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1dd20f1f6f2b509a11527734b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h71abedda857e1efa9a31ab4d7;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9d2e3d9390e991fdb00188a56;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he0facd4b6dd88b1c4bfa557f8;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1255f839f2427f4eed1f974bb;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hcfe4d53dc0a5827c7fed71a2;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd9dee60218be691b4a438b1bc;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h82692e5ac01c8eb3c51f1635d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h37ba69ac3dbb05002a0c09af3;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfda1ee36f81b3ce16f3b1aa30;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7f31156153e2eeff8eb6866fe;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h62aa6b22789cbfb42507e7bdd;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h534d7da35002077c9796c709c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5e52ef2bd2686ea26f824c188;
        #1
        $finish();
    end
endmodule
