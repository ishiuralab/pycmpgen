module testbench();
    reg [0:0] src0;
    reg [1:0] src1;
    reg [2:0] src2;
    reg [3:0] src3;
    reg [4:0] src4;
    reg [5:0] src5;
    reg [6:0] src6;
    reg [7:0] src7;
    reg [8:0] src8;
    reg [9:0] src9;
    reg [10:0] src10;
    reg [11:0] src11;
    reg [12:0] src12;
    reg [13:0] src13;
    reg [14:0] src14;
    reg [15:0] src15;
    reg [16:0] src16;
    reg [17:0] src17;
    reg [18:0] src18;
    reg [19:0] src19;
    reg [20:0] src20;
    reg [21:0] src21;
    reg [20:0] src22;
    reg [19:0] src23;
    reg [18:0] src24;
    reg [17:0] src25;
    reg [16:0] src26;
    reg [15:0] src27;
    reg [14:0] src28;
    reg [13:0] src29;
    reg [12:0] src30;
    reg [11:0] src31;
    reg [10:0] src32;
    reg [9:0] src33;
    reg [8:0] src34;
    reg [7:0] src35;
    reg [6:0] src36;
    reg [5:0] src37;
    reg [4:0] src38;
    reg [3:0] src39;
    reg [2:0] src40;
    reg [1:0] src41;
    reg [0:0] src42;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [0:0] dst26;
    wire [0:0] dst27;
    wire [0:0] dst28;
    wire [0:0] dst29;
    wire [0:0] dst30;
    wire [0:0] dst31;
    wire [0:0] dst32;
    wire [0:0] dst33;
    wire [0:0] dst34;
    wire [0:0] dst35;
    wire [0:0] dst36;
    wire [0:0] dst37;
    wire [0:0] dst38;
    wire [0:0] dst39;
    wire [0:0] dst40;
    wire [0:0] dst41;
    wire [0:0] dst42;
    wire [0:0] dst43;
    wire [0:0] dst44;
    wire [43:0] srcsum;
    wire [43:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .src31(src31),
        .src32(src32),
        .src33(src33),
        .src34(src34),
        .src35(src35),
        .src36(src36),
        .src37(src37),
        .src38(src38),
        .src39(src39),
        .src40(src40),
        .src41(src41),
        .src42(src42),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25),
        .dst26(dst26),
        .dst27(dst27),
        .dst28(dst28),
        .dst29(dst29),
        .dst30(dst30),
        .dst31(dst31),
        .dst32(dst32),
        .dst33(dst33),
        .dst34(dst34),
        .dst35(dst35),
        .dst36(dst36),
        .dst37(dst37),
        .dst38(dst38),
        .dst39(dst39),
        .dst40(dst40),
        .dst41(dst41),
        .dst42(dst42),
        .dst43(dst43),
        .dst44(dst44));
    assign srcsum = ((src0[0])<<0) + ((src1[0] + src1[1])<<1) + ((src2[0] + src2[1] + src2[2])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15] + src18[16] + src18[17] + src18[18])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13] + src19[14] + src19[15] + src19[16] + src19[17] + src19[18] + src19[19])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6] + src20[7] + src20[8] + src20[9] + src20[10] + src20[11] + src20[12] + src20[13] + src20[14] + src20[15] + src20[16] + src20[17] + src20[18] + src20[19] + src20[20])<<20) + ((src21[0] + src21[1] + src21[2] + src21[3] + src21[4] + src21[5] + src21[6] + src21[7] + src21[8] + src21[9] + src21[10] + src21[11] + src21[12] + src21[13] + src21[14] + src21[15] + src21[16] + src21[17] + src21[18] + src21[19] + src21[20] + src21[21])<<21) + ((src22[0] + src22[1] + src22[2] + src22[3] + src22[4] + src22[5] + src22[6] + src22[7] + src22[8] + src22[9] + src22[10] + src22[11] + src22[12] + src22[13] + src22[14] + src22[15] + src22[16] + src22[17] + src22[18] + src22[19] + src22[20])<<22) + ((src23[0] + src23[1] + src23[2] + src23[3] + src23[4] + src23[5] + src23[6] + src23[7] + src23[8] + src23[9] + src23[10] + src23[11] + src23[12] + src23[13] + src23[14] + src23[15] + src23[16] + src23[17] + src23[18] + src23[19])<<23) + ((src24[0] + src24[1] + src24[2] + src24[3] + src24[4] + src24[5] + src24[6] + src24[7] + src24[8] + src24[9] + src24[10] + src24[11] + src24[12] + src24[13] + src24[14] + src24[15] + src24[16] + src24[17] + src24[18])<<24) + ((src25[0] + src25[1] + src25[2] + src25[3] + src25[4] + src25[5] + src25[6] + src25[7] + src25[8] + src25[9] + src25[10] + src25[11] + src25[12] + src25[13] + src25[14] + src25[15] + src25[16] + src25[17])<<25) + ((src26[0] + src26[1] + src26[2] + src26[3] + src26[4] + src26[5] + src26[6] + src26[7] + src26[8] + src26[9] + src26[10] + src26[11] + src26[12] + src26[13] + src26[14] + src26[15] + src26[16])<<26) + ((src27[0] + src27[1] + src27[2] + src27[3] + src27[4] + src27[5] + src27[6] + src27[7] + src27[8] + src27[9] + src27[10] + src27[11] + src27[12] + src27[13] + src27[14] + src27[15])<<27) + ((src28[0] + src28[1] + src28[2] + src28[3] + src28[4] + src28[5] + src28[6] + src28[7] + src28[8] + src28[9] + src28[10] + src28[11] + src28[12] + src28[13] + src28[14])<<28) + ((src29[0] + src29[1] + src29[2] + src29[3] + src29[4] + src29[5] + src29[6] + src29[7] + src29[8] + src29[9] + src29[10] + src29[11] + src29[12] + src29[13])<<29) + ((src30[0] + src30[1] + src30[2] + src30[3] + src30[4] + src30[5] + src30[6] + src30[7] + src30[8] + src30[9] + src30[10] + src30[11] + src30[12])<<30) + ((src31[0] + src31[1] + src31[2] + src31[3] + src31[4] + src31[5] + src31[6] + src31[7] + src31[8] + src31[9] + src31[10] + src31[11])<<31) + ((src32[0] + src32[1] + src32[2] + src32[3] + src32[4] + src32[5] + src32[6] + src32[7] + src32[8] + src32[9] + src32[10])<<32) + ((src33[0] + src33[1] + src33[2] + src33[3] + src33[4] + src33[5] + src33[6] + src33[7] + src33[8] + src33[9])<<33) + ((src34[0] + src34[1] + src34[2] + src34[3] + src34[4] + src34[5] + src34[6] + src34[7] + src34[8])<<34) + ((src35[0] + src35[1] + src35[2] + src35[3] + src35[4] + src35[5] + src35[6] + src35[7])<<35) + ((src36[0] + src36[1] + src36[2] + src36[3] + src36[4] + src36[5] + src36[6])<<36) + ((src37[0] + src37[1] + src37[2] + src37[3] + src37[4] + src37[5])<<37) + ((src38[0] + src38[1] + src38[2] + src38[3] + src38[4])<<38) + ((src39[0] + src39[1] + src39[2] + src39[3])<<39) + ((src40[0] + src40[1] + src40[2])<<40) + ((src41[0] + src41[1])<<41) + ((src42[0])<<42);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25) + ((dst26[0])<<26) + ((dst27[0])<<27) + ((dst28[0])<<28) + ((dst29[0])<<29) + ((dst30[0])<<30) + ((dst31[0])<<31) + ((dst32[0])<<32) + ((dst33[0])<<33) + ((dst34[0])<<34) + ((dst35[0])<<35) + ((dst36[0])<<36) + ((dst37[0])<<37) + ((dst38[0])<<38) + ((dst39[0])<<39) + ((dst40[0])<<40) + ((dst41[0])<<41) + ((dst42[0])<<42) + ((dst43[0])<<43) + ((dst44[0])<<44);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h0;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9194ab6e7f3103cd6620f8d57dcac6f282ffcc67a2cf221cc377b0ce0bc7c3e9695590a95eac6b75da079e8ef482dd38322740f3a684081fc677e8449;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he935097d93d17ad772421b21d72f9d754125f385736f44b5107920e843cf7b219e388120e3a5749e428f6a7f9c1599ea77418f741192fc3d2be273f63;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2a7dad91a1682932b33d3df74d0a6dd76763a0087a657e5c43d5a0c30e268691eb4f9dfd5e0ddc7138d561c80bc1c9c104781aa1005a9ea17b7319e8e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd5b271b10dd2581a0d670db2f13a12d59a919c356c7b079da0421bfe01264ad2759464dc37399def73f4652f1117e20878a18687222e3de5a77e9b922;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h96a7bcfd91f33685999d0d0b7dce7a5daf2215a0c5a75acac3c7dfb65f31751a59dc89fbd2df765d1c4ccf18873d12cf6db78b4ffb4287d537d936f7c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd0cc6b6682a97b4db5099f80d6ff3b8b546a67298d5e1404fe704d8826031c95e1e803c995343341df52df468f36b1e4231020feab63708fcef482d5d;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf051b82b15c722ab5089c75f85f1c2d837eff29971ef3cbbea7a6c5012a370af53c41288ba33180829eb022ab1cb7ea71f56b7e06c4159972a70ec159;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h696cc0b76e1ae530275d1af439f0ed584eae8b5d83c077ae462fc50901386a825878f9799f5c0c5ea756e209fa6fed0b63bbc55d1366f62b13e781c95;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdada2356b6554cabf5ec702d631e3f1fe23bc1a65d74348d9e05c14251627b71b15b4120a7369936d5ab5d4acf775c4be6a9551b772c30426770c4aa6;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9b1869881fb17587a5f4982d46715274106874631d98e251d192bac38e31006e87f587f6d8c84bad70e622bd38aec9e5cdafbe2dacf9e046cdfbf27c7;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5a3af8230033e5c5211bcb5ac3188c15b31eeebc4fc14cdbb2244a36ba1f6b952c2d6aec0c7125c00c8998a96f42cec1c4b46e741461a1e08a3e80ff1;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5fc262dcc39f7c94b8e0e2b7eaf42b9a22b6993b815ebd655300a5133a0c421750acc649343a44f428c2be7516d36d25e13e0bacd1e63fbd1c017e97;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7a65a2e05265f132719706ac77b7911a4884f1a923b3fe245cc911560d7e316dcec586da90124826a45485aefccf52bb172a9421b69612bfd059205d1;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3e8713af2452f9cf3c4216645e3896751e2d48d9fce5d6eff4224960d879de4ce9ed1b96bc05278226c8200aa9b02a5dd98cfcb6d983658b18cfd05a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h20d3b92086b89c13464f6bb01af962ddca0244ac40730bd0dbf98336f6ff400bc1ceefe6d5a392feb5f3f6c90bee409fb5a4364e3afe84c233c4780d3;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9516863e9a3b22dd58fe65b72ad6e8c72677e4df42ad422661a8aa251199d51fc48c071b601eed699929666f16a47661acea60301112b7482da48a277;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he6cac9f8862493c234adf1ea715c89ce6fceace592662efa75c52244683eac5e4cbc94ebb3f73bb4d766d64370117a4ebe1613ef77c0dc67fe6180faf;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6cdd06962b77af89b532b308a01ed1306cdb933cad43051af7ee66a0f797d5fc08323526b14fa66358318b36dbdb935161a4744c26d0c3a468ffd224f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd922b4dc8d9f543d4ac748df12685ed68bfd7805cf008560e427461982c35569bde5abaada1e285458bbb0fec914373cb0ed3051d6af4e5695811c4;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6c4a81dc1ad0faf27902c05090b6ed90d8930cc1731de1792563556be90ffce4486aaae1bdb9c3c88e5f6c88e363c730539db296563347add52e1ee66;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb5e066e50fa32a467d1ba397eca587d072cefaadd0b55fdd54c69418fabe8b71a701c9f0c29c3720609b6d034356386d8e05abc20530c8a401eed1438;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3dd71d54ff2556d4730649d9e62b96dca47118228b3d16e32ee17df4e84726d2a6a8bcb88ca8ed93a68685e0853509f9fd6e51e3f5f6710337cb2a4fc;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h278ddd2852a09af342f5d1242072bc444168e626a8ab5515536b454e518b187b233f31c8f1de279836ca9151b57c8b3ab75a662786907e49e1954dc0e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h60dabca11461bef78a4796770051d5090b3d5bfc2320c34bea35dda172d4447f6207763dd832b26b20904e390e5236aa937fe733dccda92c3ccc33206;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfa93d19de10a739f40dceaae72e52372e3afa4a356b74df8ba340b62799e7ba546cfc0c83eb81bc92fc68b1770b7ba757344184992d1706490b7a6f41;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha176b9fe6b2e9b62a1ed180b0428cc1f2c0317d618617cefcdebe8563619dfce246226796a7acb82e563a5372b623d612dfb4087dc818fe814cdf76c9;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd86e8affa7f086304474d2387cb8d477fae0a6678f5c73962b903365a4a6320b7660e2533a4f296abdc59c3637ea10a66e19f481f5ae60515ea3d9763;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h20a19fc13a399cca21e923b44be3052d5e05a77f2064ca2c23fbe05d56ea3bf79712ca27dbd84f2a12ff5626be5259eb2420b2bf918b02f825b5b8362;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbbca2b0fae8e8a2ad1bfb1d2274aff2dda986c6fd2461bbd22049a08bf836b95b8c58a381f5be172fb8fdada781ca667b4c7e370baba029eea4a1d92c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h696844e34e5ed3320698440b21af8deb95a2dd507a97a7d0e64bd09880f5528eaeae59d8885fe317bf79fefcbd823c95f6d8eb9710556fd8ea3ab1f7f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h55196ad871bd0f37d63bb1f07e07253d91b4b5c71bf7ea3accfbf9bd10ae88ea9382fa589ac60a7dfd47a7759cdc781b4810a3a83697efe1232cbe6f7;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h650b319418ff9c71128c496827d064c4e61f8e5f6008b9dea4aaaf2d2f5bdb7a2a7958e8e3229f86a927796c577b558af279c0c11e7cc24dc709dd216;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h662465599dfa50f616a53d35c9c8d9446097fb852a1021500cc6b023d6b833a801ceeeb54a397e581ebb21793fb03a239660bb8a0f6338a18d1be88c3;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h37dc7259b7b8649af208dcc3c5f4f92989e42561e4cb4a9466ee654fe7d99712d96b18775e8bc38144e7ba87e106facd6157d092223e63800a63de89f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8e4e6042cd32dd56ce19b12bd116b5beeeb1cbd150946b870ca2e9be24cc3d21a933472c9919e8f678c46648fd990acc37135055b8757809e9e3fa73c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h35aba4e34d27ecb47e333f166151d89fa4f550d3885fefc1013cc43c2fc9d5ffa84bf77df9f7d5fe2470a85e685d5fa96b9c74558c47b7ae625177084;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbb597e7d79950c5275bb2aac4b12865ccab1f5f5bdb48fb8e5627517297fbc21853a3ffd6785ec834e404fee0c1f1dc7691fb59e13196209981b0d061;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he758b85d913e285a724585e57e8e9c2050f0742f0aad1c2db9a2cfefef4b3677bb8c98043cf46f7c10debdbc0097b196bcbc244b15c805bb134413463;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h91c5c0a56d0d2745d9fc73ac5b96e59e2a5afc02e943b2b161db94c0e9ce9ec21f7cc9b08c77dc025f0fa80aa167d438b6b09a7de0dc12040dc835861;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc74723b90fcf46fc6096d0e2c7254159eee33a7e3576e9b6d245f9d0b5d551d268da5137a92376d8b7ae4dc1269f31c1d3abca8393a68b4cb6cd5932f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfca855fce83bd533f52c66a36c53dbe24c1852e4c8f86d68348ea38a3135148ae27cef945c15859d537421c1d262d912f1d7e70471b164edb76bcd6d9;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb0c128f5edd39e5ad0e4cd97a49c0438e356a8e9fea8ecd4f34bbe62fabde5342030cbca7b8573c9de8d050818aba40abadd5ace80d92d3acbce9402d;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h628eb417de27a1ed9d9b626f510f1844495bc6c66e3508e5ef7ab5639a97d0386d45d132082ab51e570e3ae7c866b7109f7e778a8dc7e3b43ce18cec4;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb2131cc1d536a840d95b9e5bbb4172489b0df8aef694a301dd85c72c8b342e172d7db81a0ed3f89311fe6193bfd26e4faad879a1e7d66c7d38c67b740;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1810450928e151748d350242b8d568cb6bba9026583de71c0a7253a512a15e4aa35a279637942c592306df0924013d47a2398548a0ba11ed75e75840d;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3bade7ee2d9d37f793169f6dbc6d6424f222d4e769e2d8d40a86fe5511592496d9acd0ec0b6cf68f3e4a86b3f18b50a215b317540d429b7ba35363d60;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5f53ee6874665833291f68ab050b6b1f6b9d6787aeed87f0fc5511ddc62a156be206cdaea92b820a327968c562ae0d3ce270774bbe2c7d17be9e3f492;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf3d9b2f7853d405d9971560278c8b8c5762aead3693d6af725dd827a8ec673f1ed95c4df99bc12d285b1dde9b6664b01aaaa05f5d2beb3108469f427a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h54db417511d242d60a6a8b1f22346ac41bc3714dc3df47964c6076aa1e864abb6a60a62eb4e52681a7831cfe185c4a5d3bb282dcc004252a7cfc84daa;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h92f468fa4fcc2da0b510e65d8fa6b9b7e927fb710f74135c4f322ef1acd6eeca7fd6cea91dc9aa16ce6a7562e377ed9c9be11ffdf57ee7247a745640a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbca1806ae02f671680221321e2ef73f16454b58fcafdfc6d5063229b4d7095bc26d88be0bb4df707c5777ce57d4677b661d01517d8c89b42a935cc8ba;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h49731fa96496daa62730a380035bf4b63ab41aa6d6f3ce83f415aaf9afdd25ab8a11f688575e905bf42523053e396be8d3bf6b7a67f524ebdab122327;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h82aa8247dd0636dd391ea2ff88b7f4303ce8966496335a458606fd56b57c727e55b962aa279fb173da3355e3ce179d792ea6f854bd62e7ef3d7fed851;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6544d2525d66d6b598ef6b9a1d602955dc5b7612ccae5767ec133f67f4d7cd934d09b487e966b1ad11ae9ab67c8cfbfcbdd323af5d9d0ec05ff5785f0;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h698536ac2f81228a71c2289e0ec71f95ab4728f8024bfb8425989a43b71fe54ce1f70b50872ae98910e7645ab2653a515d348c2b98f99f8f79ea01dfa;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h68410ad566a02680b10e63dad04b1a05ea4a780cb6572b43b9bba8b9300a749f39a3ea65a316757362fad3d8751d9f47c6bb01adffb6d3f6871419ff7;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hebf20403dd8d4061314a015488e4e33db57fa68d79918766e2c9ecb282bfe4d81e7fbb9ec3d2c45e4c01cd3c6aa30c954a888c522f7ccb7b07524b761;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdfa5cc5d0536000e3fc3daebe2a1a1a0c90671435c720d5f2e4274fbaae1d35e6ad3e0343471601b7789ea18fa13e130c45e34cd7fe05baa8a177254d;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h65835b6480da65f2ec20fc9603d1c68949243ef98253b1c1c1c72ce28aad70aa0ed11ec2a375da5154db0b0fe50cd3592568320de481d6a8cda7a0be;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h92af4526aa42498a848a53c1ceb9f84795706ca54cf5cb0a1c73c21379e5acf0cf4aadd40de8c1eaa651db35a70d1e61c889b63e858a09eafc1ad039f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h348fb11cee6e114c7c085e3eb97dc7b1b288da7f22a4d1f00d945e7e24347ef302d62c558558a7533a3dc33c81e7a57d0820ba9e33b019a17d84a79f6;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h667f40f6e33c7db54ee218efe5d0fa444d6f9aaaa1e38be3d3f3ae73aff1607d8619fe405a408b6c0434363e5520896bdae695995b55ce3016f8a19b1;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9aeefef7f2586a1a9029e8f2399427228af646b76e7eafdeb4b97324fcb1130c8204128b61ec3b958f56620c4a106b68d9bce19390c2c99350faa0667;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8f5353b0ea701da6423b1ac5fed9825973915ee08862c8ed16ab98d54bbee3b6f13775bd4223fec3cdca7fcca75532a9413935ddc0eb1ffc87decf47c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3f624f05b9a29aa7295eb77b901390e2cf15fb0ebf7a1573a7fab804e3c25d646877fe61c742256d9b4bbc2017c4d1d28ef2da7ce4a4f462903c2f2d;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h72e82b199d7299c45c26e5e86669d8e4b3835ab3aeb3c03a65bb4dd24b6ba5011a549cd504c9e26cd2a769e366aa98d7a1b1b1f7a03a543654d5749df;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he2a0ac030d4da01cd27ad2f58b4f9afbea2dbc311f44f4da5f9c562e9e4a63c9097c724eca99970c3878ad3d871dc3dd784fa2584a950515b8454d759;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5a0470e77f426ad035bb892095cd772a46529571f71bdfcec32fe8c31ea45797d78e44858c1ee1f80d20173d8be839c452935a5048fb92b603dd3816a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h579ed1740dbfb6d13b3414936f6409b55c158536c8c5e00919c6775f4a9fac2542dc38a3c040bb198b0a5996859d2c5f750ead5c6046b7580ae31853d;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h68e4f85917135fda504d8c6e85e3403c052024b7af9c27d2ef2a2c9dc183ac7405e5f98599a1ea895960589882317b7db6566dfce343364f9d329ab57;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he2f5f2eac1719f79f8c7534a4c94bcc2a9eea75f2bba669fe9d227dea29af0cddbf527a5d3ef8a93b8783d6a89f0a94c957029d8e4df584ae82e203f4;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2610ddf33a68b07ccb8491e6d5ef2daa221d0225a22271e2dec17fd83d0c6b09dc9d5d1eeb5747b11d0f281e3a6cc237944057a71177872531b150e9c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h57d35e96d37beeb4221643c8c4d69046f05e71ffa86d1a144f43fad9017f7229ed3b566b305c4fc7fe236227d855896381d7bdd8e1fe6a8fe51bcfcaf;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb3bf8f436b005f447d8c5c9bc05147c376472608fb198d82c2f6a7a2c3f652bf5b3168aaf51dd7488c7eb2d844f1f842b54a45d86729becabc0b993b4;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h839e9af7fcf8a9ee7d8ae450ce94619bde478194dc26b45c963e836e012edcea49b9d2f5fcb5f5a0756e3202a7c25129751b6b67f090426af8b67934f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6f451d63116d8cc034f44cad7a8ad0626cc71fcc9dc6dcd0bbe33fa4df96352fe113e67c7fdafc508005609a5ec0c372bac95fafd25113a66f497108e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3109332f31efd3032279b7d2e74b7632f75985562386fb2acb2001e20b3e117038c8d89bc86c7d7ce3f9b7f642228238657d11a0125b164627c475db5;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hee4ac82e58560fd91c3ead7a69a37645048ca3775562317591f97976b4a9c33689c6f5fee896cf26765119400ad27a45881e6929788758464c3ed9f08;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h81a2dd9519b27f7ad5fc03ff5c915d41e4520c2459847f4122879c6a6539ae0d838f7b75337c737600023fcbdaf7f8ad2e8699be00ca3aa91cf64f346;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hcc0b2aa53b91e6d3a8118e5344c2373ab2292098f3809ce71ad8161baa7a3bd9de497ceed451d86a1020aba6bc7e98372808da5592cb0f97d0ca2d2ec;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h16810c8fb27b7b76c7c1dcc151bf545649f32ded16f1173c2fc587ff2c63ba1f7ab91c183a15c21bc1455725491d0baa18366beb37e7165ce78c9a798;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf2c50f46e7345c6c3328e55ca33e5a55b524616b075fc32b608c0befd525ea3bc9628b0b493cb313a7bab4d16279765405a0a795ea806d80f343a7b69;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc57445d3eeebbbfc5c820f8749ff71a271137e35ee9c9cbf999085dfd6682748ede2e07d747af3e4436452cbd1a971029da4f51ec879f21c104430e40;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbbc22a7c065814915c33308f729c40f501223c6857a7ae67f24031dce8dc49dfbac19d1a7f0139800b3e9b078743d5414f1fb29dcc72e55a2a99730aa;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h40e52b78e059d5799bd609840accf2b5d1f790ecc6ab22577f06ff600a62b2fac258ba76a5148853d657403d0c55cc8334b07e45157d8005fbbeb26a7;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4f29d8f5680873c961b3c98bbcdefc07844c19ee3ae6ab4cc0efebf94c5f255508c8daf0d36c465ba147504022b8b6cc7cccb36bd6b6301f1f664054a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc8b62a8013ccd219fbd79d672bb9cc2dea69cd42dbab1901c5a283691890430f71c6a43dc437f05a7fb72ad4b42513a4829fdd3cc7191c2947e24e447;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2afe450d5b28cf13b00929f7cd3e6dd398641c92a066bec883d800b329525d2f7a119cebc710e84a3e1d47a038726428632c969c148ec02aa1bb80f45;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3952ef5287109472c2b23bde55bf1af78fceb5836cdb6cd3724cfef5fed87393f8221263f6239427a0e0c53b4d877593b27f941899c5980a2c6e88f10;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha596299f0b5a3e11fc9251e123d7d38949f5fa99d0bbb51866aa60d0b34988166fcd4b68fa36548084ef709bf1f27c351beaef3ad4f9566a2b0fa0984;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h94f52ab1586cda9f2c059185e6e7f9c7cf1fbcbb82461886d33d861e92a029d2c18e53ebae52d80e9d051f97a13ad2a9d5688d357e8af0b091d66e1d2;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha5f0986a48c69ab1633ca2b0a8e57e944cf1d9a03ea1155217607a116a8a050b3b0bab54a1cef03db3f40c0c180329c66d3f1a365a4291f2ba298a5d6;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hee72dba986f93abba6fdfb69a74b5f73499dbf19407af2ab3af29d86b1acc01365e8dae474f9a4c1f10f368ac199498c5acd03682279757a61d9a3b82;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h98cbe590400e08becef6410cc28b9817995a87aa044a7579bd3d1052ba4b2eaab36c20a37488de24fee4e2ea1f3a653bb7537cb0a52cd7281eac737d4;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'heae69888e220c5e6bd24143ce41f281d40d6b26bd4e182fe422ce695dfeda44fcca571307fe7dda7f14c95ba6a9ffd58ef23f7fcb4d8a3c4e7426e8bb;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha61cdad6d669990bd0e6fc17071dfb6339a66ac9a4f62cc8b9f67eeb41f9121411c67501b32a86a0b1c158aecf054f2822e21746ff27276727d9eaabd;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7920a4b7bba6753a581a1e3142ba081907384f7266a90f0f41c4deb85db655abd9b7aa9a7d81b9978c0f4bd3579730e9677a2824043675704fa964cf2;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2b9250afba8363c6a3355775779d7b7513edb3486731bed756ed911c2adaf7412240383c765c58ec20f910e558fc895f7fe71109d8698091b2f7a5cbf;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h767b1615247e90d13ebb6bb3ab91363915392629f4b8c1551e27dccde31b320de8c6aa97cfcb1065df0aa7d6ebf0885554b7d699addf90e7d08f634c3;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha39e2609b776df3d348d963467ad0aa71f6a896db54a236468f7c1dda83fc264005207b9c8bc71c6ad95b0545294af97e7fc989ae4012c6dec7f77f1d;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2616e91f61cb8f368bea8e324223c8449ed5e17e9e15b0a9e58ac0c3c23ec7781ab50b97566b57e3b985b5748593b9488b14064942cae7285b2105822;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3b40b34c066c74a4bde0b6d410882acf25a1906430984bc845b07705ea66097103640c4fcdf12b35e31603b3224fcbd1e9c1191975dc181cc2e9e0c17;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h30091c5dd52de33a47acad91d04d3a97047a0e1e8bce897b51cf92c30ab84aa7c95035ad7dce4e4ecb572c51dd34abbae8cdbe3433772c94a8279733;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd08a04a7a4fd4f805d128e69881bc6885bcbae7c58aad0c0b4ff69e61ee8963cb80b0a045dc8f4f9fbd5b50d41e98896be04549a3d359c6af2d3220f4;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb7992a45c629b764d255a0ebdb9978d90694083ca57bbc326c075020241018fcda7ccdfcad80a269a56546f48e610dbc3004cea08957335d4ec21ac1e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd0204e087e7801387e52cd2cbf02cce13037d6c367d3eeb8e5a8180d2af35ecf49dbb91e1dec6bb207e2ada3f54386c065d61e845a320ee2be5b6f037;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd6508289937c8f04dbfb86beabf7e115b8582412c729056cb879186f1b3e47939ecd41b31ed8542690e240bfdf96f04a35710b628944c4ef296860fc4;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he5fddd6e9fabd2b48d7a8caa5b2709b170ef3cb35b69cb01e90403cc931bdf3d6f13f246fcd49ec9f5710a8fc6c84776b961cc7026138cc9f16071d59;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5203749e66dd552c1bf4bea38e55ba2cd6a5767e03d1429078645fc7387ad68aa79d3b808bf1c14f024d0fb3682479f1be38957b002f178118cd1fda1;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6859ea47e24f86d6d37ccb9dac9779a2745867e4017b9c11671d12ae7e5e418bababcd998b5468176fbd4dc3929bee42d1993b6c81a4e414781750d5a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hffd607b7c0abae49f0d5c48efcec4ec4a027936754f8f6aa966b78fbc5b3c53aa5904d1acb2e56e310a562dec81a76a80e19db9f34077f78b55ee4e72;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hef049ee006b92905cf786b7179770c4f3f2cc1c31e62319beb47cc2c6e31e193ca132201479b014f00f4cb3e004f36c9462733ef9cc18fed7a388174d;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf529a203f080e30750d9bf63de83a157faec86db750f543f1a6c2a0b8c36ff941356900fe45ee9dddaf40a8c8188ba01b7599ccb6813a8adbfb31f697;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1dfb515af9ee05e8428ce1b51edb3089d121e73d57f0df62943eec6fac838efdd22b851a59c7e4f48515f338299c27c7af770b9d01d017345d6af59fc;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h59eff9f35004358e9729a998b17bb02d368d78b7f01f02793354a625efa27aeba6d87e6b1dcf50d69a72c78d71526932488f5432c4822184d751946c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4f4a1218743ee1397cfd7eb2a5479565a393c6dd9ca99dbf950d5da18f438644a21ee8fc3edc138746e8a1ffc794366b05502f022360599722abdb1c9;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h34d16862ab932d9d30dab777dbfad46ab9b4259f3bbf23bec11d95300b13df2747f2f4b1dbd96510002cbc3835e05e97f037364d8ff3b514909323975;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5691c40d19e4b10a1ae2ead846335e9d3ade9a619da8520558fdcd6e03e5fb52a17ae207330fd5d25579d565ac34ea5bb9df03c2e507e56f95b0c14d3;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc7e603831b17bfe1ea11316a29f9f2dd136526ddacfb638dd47821c1a91affaab30236c040551309670f6ff033cc5f0728c0944f03fca6ffe8ff536f3;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hcadb6785d9e32128c24c746e0d484a707e0ce39e7c835e6039022841ee96773461ccc310e739b9b5e1c880188e5add6460c9ea97ae3c0f2e0022c1ada;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9db99015459e3a4519ecfcd7f057ae77d6e3ffcc8eea435d399929600aa498161ed048e28fcf902972fb030202d76812e4e802b968fd549d19ebecfe3;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h53ab33f3c95b908fb73a0ac9ebf9daee7c5276541178ad9de50bf2c90872b3ae877d2683184c4f10bae03d3457748ca58abf8929b4cf4e3a6cc6e75f4;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hcc38ca0dbf0a0107f29b4eb2bd3285d2526502b0a824e434d2b0108b60900eb36ae123a33c8589baa261a564f93ad0e012ccc51ecd53832fa7fa22b05;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbcc45b03c6503e63a9f8fe20c72b032c486ae7357043bdd39210898b2e2aa58326f1fe089736cc7840187b4941a86a5da0b475cb4d852506430abe092;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h30bbc033c60696696fea8a2fa4a775cd633d90cf0edf0d84e80c96ce9ab4ea93f3860bb2fe0c784c8b37ff9de86c3287fcc2aa4091f745556f0d40870;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h46da9606638b58d6ff27dfcf289b91df0a6a2947a4e0ade7613c8e9ec61bd6dd1fdb06b9f7660442ab9f9f37d5a5dbbd2ed4efda926edca9d2a1befb4;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd18b0355b26ef1be2a85b6dd5834afaf54a8eb064224a174a0d529648388ec22ed4980179e4e83eecb6a4a627bec96898a900d75a86744827c976dcb4;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h84014f6338fcb23bec3fd6614430e17b6b2f7b0f38a8d574f337448316eaa3a63e7ef9749231bac80e22e5f76edbad88efc6d5ac6f0168a3c3ffd10d4;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9d08eca3f1b940e0d829b29a79ba5bce7052dac80019c27ebd5bbe4211f850b87ef93c0e3bb12c3c321a02dba52727a99779a8955a96c84d4a060aacd;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7adf648e2b9c44201d771dfea364373d9af141ecb421e5ca0f165ec28caf17cdb29f8c387730dcac76d3d28dc18b94b920e05ed65312effbb19f31140;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hef4f0745b0d2935faf545033f2e876155509b94a913069234001629e8b7d4c6c64a96286e8280f5ec01c3beadeecc0b91964f73db09e1781684f32404;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5d6b48ee962cf7ba1a5845de75c40290887070688036d48b6e0330b88d7d7b2f6c56ae0e655427a3acef3a09de0a3f84afecd56615e61c02c573b888a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf7f26983bf260fd62462d7a7994cd02b6963b23b03de2515edea1ee354a78d53dbfd2cc6d25fe356d8d87e7aad93a4badda87b7a3416e7240749aee6;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb9f6efdce30b1c713332e25269d0079344738a691db12aaf7efa4361b20d422438aa649adf3787ffa16d15df2d0d572b864eb219ae3d41d7cc9ab2aba;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3beb8efe491e6f730e1614159dfa12aedd08e3f023e6bc61c363bbf02dca2d710e156786afeeb008c999f3cca30a1219b921cb682a80b0ff70456ece0;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2e3fdba353244d1dcb6e84b9429708c5e51837a3c502054c6e213e3848d014f56bc5b05b209e83959e47e52ef1ef77a88af2e1bb879690433d176e04c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2e16cdc1a88b07eb0472c8402c24d391a20baf71e285368b70c623da2bed49e3a94c9eca3eb93fd484b2efa35c35c608b13d9ef1a52e51f36a74b3cdb;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4c845b585c1eaa57160c356e032afa51f7b540be45985dda744ce61afce8835dc1511277c5312451247839f213eb2f9a0c6fff1e063bc54abfa4ed93e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3b86bba955df53c7f03d448693ad385e1997203c3fc9df49c255e05b54efe24a8f257242dcf15e7ba299d430d03e0c701f25251bb3ad9b90bbc11a2af;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3c7e290da64da52ddd06f2c87a21a02e2ea9572ff335037b1c541e98437ad3b0b712bb32433041bab746784d2da8b1ff82c67a21513955027479fa929;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6440ae3b5c5b824b59ff1e9e1e26f7e7f81436d98b4573243651c156a988a28de13f7f0ea25a74db376d4b700f9e47bbeca294a1de3fcfacf11306a58;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdc903ca87e2d3f1aaac2ca064a802ea48a931da8a9c07211019e4cba10c36f0813cafbae830ba5980264b53cead217e67c2834beeae04ffb2b2448b97;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h813264165626f1b71cd920dbb99422352d5456866f04f1714b6037185311409a3e201c52d9be8177a28be169e0da502027d662c40e8d0b9080167d395;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc1e9ad658d473023decc401a326b5681ec4d56c9aaf705ece9791bac60bebcd09c8d04d01aad21d56f7e2a7289fadaca0e21741808983154e9890654f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h50eaf8cd702000c9e71f9d1065eeb5ee3b6189a11c65c832b6ef07994e2ba3512d920e1e94595c2a1c450377d961c90476b89c84b301d3ba8015b3c99;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h61110fdc8162f19f8e5d8491c6fa40cdc65c36d3c8411daa0d31fcbfde87d117923bd19434e2a8ddd60708ee2bf801dee443b88aa8208f49e9f96a702;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc5163dbb13fed0eb92a3874209eaf9d719e9573e8a1b091a7b6a9988013347301020a43e3b2df61ce657804ddb6b4547dd7ebb0e81a5457c2640c185a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3edbcf99707df33a7a1605065918525f2f654bceebfa280d1a2844159cc0723f54846850fed613f9da8ee88b60b2d4a49a44a1a6442daaa6b7f9d7dc3;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3903c5e60c5dfdd72bda4b902624162fd09c5960d5087a92f9ae4b99c652ddf3d824166bdeee8f205b2d1d9e36b66ed521f071578186528e6371ed1b2;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'haf6a0454bed7e2cf9a119b87e8ba12152be9acf11e0f7eb385c43aef639d0ad09f2f4a7162705675f5f624789b7c055326955f9d0e3ba4fa5ea4f9b6c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha6ae5097873339888495c470530ad5d83fdc5eb8e955c6ccf58f069e103d5b7ae41be3865b12f509081f078678f51c16f0ce077affc1b017ff080ae6a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h56a3e3ddf822480e1e98d6859aa162a32d4b78ae4c0f4de24a58a90d721968dc98d3e937b6df6bdc11e355ecba72420208c8430605fcf314c50d27e45;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9d358e9c348bf58ecce85463b7d94c512dafa4247151e49fe459873f310bd15a0f729205b2dc259b56f25368cf580622ff16207894207cb3b7c9e89f2;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h37f38707a27f9f590dcfcb1f2996c612171633b603143d32cd7b0baab1af0399dd8805eb103343f2d1f28a47beb43b0280d0ba4d897d6eee0c3f3ac06;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf80974d91fdeb135554eea4eb297d557897dd5a986d383eee86f2dd6b3dda479c8cb0bcfff5839ce14aafc52e791087723d2c2732a3c35a12dd45f9a9;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h518eb85c3791bf1adcb3e3d8888a9838092271995a6b78e74a9161aff9f40b2cb971a1cd472fd1f3f6461f0a76646932f3e2059511f84763446350d4c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8fce8aad9607c5f7170d974ad9c3a4e38d675ef0523d374e212543848eb0430cf0283864a3d6adc33f293fc8d7d2324b2ced18382d97610e3e4f16635;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7ccca63f9ba5bf88a10f0b27c857aa4dfa7292b38153da5b3dea692ce448902e1a0d213f16475ab2cf0b24d4cd546a0dbcc53167b2ac491f64bc6e4a6;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3eb454bb8ae059a81f0feb98f7ec48833485c6335a1821e06acf733a0231772480b3d6b90998c84be991637c7e6431becac538d0b36456c7d268ec0b6;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h27dd92230300ca0c659e315653db98f60b0da24b98733dc525cfee5c1a1aaba9da89dbeba24652f6edf7a4607630cd5d756f8e6441d3aaa42b824dbc4;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h43e046ef5dc773ce720347bbe64095140fbfe83917eec75d904aac8cf3f1fb2989ec9dd7e9b8502386fe2d792fe6fd9f8ab067c83ae62a5441d7dc26a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8ce78488333317e5d4e6b80b6309dc9954b874e36d9bde3bfbbda39f15f0d42a6555d6a87aa6562a66a0d6f09c52bc71ea75b9cba0175861acf0ef82f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha9c2ac09758038ba81d19df4cb791288ceaaa4c0a753565760a764e715df7af5f1a3d3b6e05e4a2d77976bb9424730add4d5d1dd34fca7e5e7a0656ad;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h68168d7f41b6aba78ac9e439009bda49856d98df4662275a5f62228df5a275a7e4adf5ed71605789f189ba732d1dce2f462b90f613f4c3110104726f1;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc5aaa4e5a0678e06e70ffc0ea8e4300a1fb24e16b7aca97734de093f3022d584ce4740e111aa84c0c42071aa3272310614e916b8ca77aadba92c8342b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfd8836e31698c0aad9aff6bd856ebf6643700cc45c2a5ece27054bde50354c39d41de0ec427025bc970533d9da703fdcf63f254d9517f4190d3f35c7e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf44e1b07a5d3571ff5426ab1d674f321e9bac694806b76782b1af40782a7bc0242fcbfd90ecaf70704614d66aa161b754472366ef2d1fb636d7ea1e8f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb626a78432471d2492c1980cc61d53e42c9913b9c002435726797190d01d9f9cf4ac0f5a288b0d052e25195ef2bcd9501424957ac9c4755a312373290;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h37d7306e00a6b4e88c7e5e714dff00b6f9c78a37b593fad256a903fb1f1c012c199a645f202b3103abab93882eaf94c65b2f328b4b73b3f266496b20b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd1d2a9d76cbbd8d572cdcc153f04cf16272429bca58ee26efa8591947eaf742e0ca5821d99ebf71ef0d3a8a350201235c4e57ff445369c0c3690e437b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h46d02eaf3f30e96a0984bed62ee9c2e52abaeb603928c305c2497217f01d23b8318a51f6ca976c2f0338822934afdbf4aab23fabcd3b2bb39a32720d2;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h74182d3b682c227e6e47f254cbaeb34caade08cdeb1c0d4d54970deab36fc2bc4dbbd87ae9dffdd18f75161655d8d8509c7dc66d420024e3cb589a9b4;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h53ac40d91b82349e209855494cda6c16c7c53388d8d5de9834d83cf2b300be14468fb4657b4cceecb2257489d12b9769f7576a9cb1fe7c19589b58353;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he0dc4f7a70ee231729b474c53faaea04ef6573e8977f0fd0ae6da48ade805a3f53387253b1af0f3e322fecc752ed9cfa9ec3fbcbf92d6c36746aad6f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd91ccf588d03044aaedea98a1a3e5f4efd2c4444927a72785a1f96fbf44f17ae73c6e89402dc651a1fb6e8ff7adb99c86e28ffe6dd8ad61e52484243a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf6194485741186c62ababa08d605d82b65c22582b8e532c15c5c9f5f113eee6107f0bc2e9f13834d32855289be21e0c4f4d0f4164bdc2ef67512d96a4;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1f3d0424bb16a1e1e667afff685c1096dbf426863ff4d66e17f4d0533eb125d1ccc351c2c96d5e2033eae4450ab455b36fdef14bc328d9fd2a6c3fbc;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h341dd1a644d32cc4cf260b43bd75796aab2b951de7656ec672bddda63e00109b1252213520136ccc0484e60a2be2aec6c79526c62b0659ce663be437;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd174307f0aa2862dfcbce320de94b5b65cacf634a6bfabb1515bba5bb7383161f14dc4aec4e8c4b9cb0118b74ac8a12e1ed16ec776399d6d8e5eddd67;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfb9a9f5c6dd8c029573924f9a2dcea20468a1fb8fccdb771e8296191f2585422b189abbd8c01ad01611516a5188d0d7de0cb3c65ec6f1e44d94d34e65;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9757349e0e82c4705ba9927586a47a9307863091a46fb864a48b276f6283967a47b9c5ce88e5c0388b9aa4a806ee2f345c64553489bc90ed407b41cbf;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb7f36864f2d01b7ff8920f30964abd30800705dd2ba3d20ab9ccdf8a59e9555b2472603e418efe50c999385d2760cee0285675d153374af2f16bd3842;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5e5b8d2aa377b48cd62958ba60bdf581aaebdc5741ff8df546a68397f37fb7788b3d0677e4054cc510cb93b74e33f37df5a48aa2f805b773e7329c216;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'haba5773f276d00148d327119fac9d02b3c9668eaa391934be438036a3f7298fb89cade307b9c6f5dece9e5cb745b263fc807875710be3de1317defd2d;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he61df26ba6b0d8fc95cc473d77c01b71bce63e126d7043d313feffcfb174e174e8ead7e574a88f45efbe2caa9b944757d2fb37fe9d1554786459c0a01;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3fd5b066b203f5be278219fb4c06afe1ad1a9f0a05190f63ccb6141b501f299a031b2d1336ffc3140d261761d8bdd725ad81bc3b14f15bc07c0c19277;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h38e95d7dff7aebaf0a47ee82fb80901fa7d57384d492be363259cb1df544835dbdcf0ec2ecb2cfbcdb6804b82233fef0afa78e6ddcd110eb4d7c9cb91;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h986228cdcce38e6be4c30f5ad87ea3f3f031351070a97c429b1f09c103093c0a23916e0b7ee948bdaedc296030a86ebe644c68448f978fcdf252df6f2;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3857c01e4e3e84d185712dc2a0e83a65da937791c6ab05ef5682be33c11bfe8357f9cf9bb7759a1cd2a0cff2e3085a9bce7422db4f161e2ec7a88b3d8;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h766fff424982d4fdc874042057f5e79f950f63190c96b56038dccd7fbb681dbf2510aa7f8632699673854d0f10867148c4e536032f3d32ba14088abd0;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha8df472c74e3c3d36dfce48533e2a0af71ec41e67096cae12085418c139aa5d3da76345171a40a8c9d2fb456926c8488d0341f326d89aec12141202e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h31111e5f1cfbc8475178bb00645157c4e568baea165721ff67b4eced82dabc5157493729fe59eba7af626a7234ef5931fa1f6d134804b7263f33d44d;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd79a00dd0005c0173156ab2cab6a188d0d8da808d1255f55e1a8692165bb5b97f9cf82ab34298f69cd56054e7d0ddf34dba6064b490bc4d110d62df5c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha2573c05981547846d4fec95bc49ef470821f3450daa0e9320fc22c6cee42a7f09abc04685c73a1966b77a8e36fedccf1e6675e34aab2f223e444bd78;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbe434fa14d0c7965d5a5d2692b3ef6a1e1ac86ca3166cdac68363cf1ad940694ed860d1738e79a65567a8d0693e1459bc226106527695de813c7b92f9;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb4f3d83ff7421bd95c634682221a4fcd9172b797fdac042bd90d6868d234d206e7c7e5dc2c9139d5807bc5b03e967c10682ba3ccab05cbb9ba09bb006;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha62127e09d25a35527c85d88fcf9f47b509f27e12793a3d779f06ec58837776eac9dddf92232c50d91f88b39ed96d919dda3d835f44f52b23dfe9e44c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb06006caf37cbf3e19ab1178ae20f54e10de3ab7119bf481a0b5bb63a7ff9855667fc6b0abc1d168666f7e2fc07e1dbb413ea33babe1efc1217e0cbc2;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h94dcbd6e4bde2b2d9feb627441ddef338d14813c61f740477f7370ea2a004d852bc8889be62f115873317f92fafb7bf7e0af492f6f4255a511d0e4e5c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc29627531b575ec1cf0d6eca002a3d9515a29b99785db462460b230f9783915bf49f7642bf20a5030e4fb1706a1bc19db0aaa986ff513160b6623b7a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h857ea438638c89e333b846349cdd668d634c56d6304bd9afbc511f89311cac611fee2c8de5ef5536f1203a8071f78c0bcdba8fa6e030dad42a3a74a7c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb81cccb868f8929ff45a79fc518e41907bacdf349d9f86fb715a15430ecad265472efef6b8762e52ad9303d0ad991fb02b14fa1ab2ef2b2dc95f3e0fc;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb7352f676605abaf037d19da8a1a869ec4bb02c2468515cab005d23e9d00c4abc670291b831e2bbb4dd4b9e0855793d03bce29a5f539613ad258c2f66;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9c32016d9ec5f305b7408f15ac47c17b6a0a99b689a44a4d52187b1ae0f145267f0344ee91c8c378f6c16748a8785c0c68b74a8202114647a6c21941d;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hef8aaa146bc34912fc61756b6024363711c3b0e76e1d4f3afac38a0162bccc7b23d1444eddcf8c31c01f7aed5b10e70689468a975ce221a0a28e933f2;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9e38b74b5f664d021774b093ab458c50c4be35034875d1ad032e604b8078c1d1867886dbc50c3bf745efdc10828b8ccc49bda674c9275dab6fe1a8fd9;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h68b0b0209a7354aa84e4838f0ce3f3bb1ba94f3fffd839da5a55c2e870b20c517a21b978da7ecf4a1f864e4477adb8c1fa36031b1e0ac6054c7e24d29;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc0c93415b76047f0da77feb1b11f6f66cc9988d977c275d1442c98e387d79ce0f0aae325efac09d20eaefbd64b0702ea3fba7a1bdec1a9ac448f57a89;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf6625a626f7e8340c81bb1e1615a0b13557a6112cea24ac87d4c65c627d235054afc431d5c3cd435701b7dd3d94685f71a95502762d2b3664a5383d71;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h813551094b54ea1cd6711a70778c1d24b1c7efab77ef76ae4c3e16c55664e2224911812adf3d410da8287ebab90769f6cf96bcc42e6cae824818286c5;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdf0931cb696faa820e5f8b039b2eb11979e2b0af4f6486938e4d0e4169a43b5029aa2338c43a5e09be0fe4d40ffe4bcfed75a759f687d76e6c858efb9;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h450d7ef98b9f5d9612bc50e3fc5170fcce2c0c9b170829cf9a5215da12a36c785b2cf330a1719d68f88db0afa9a9b33353fd2d840147328921aa11ba6;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'haf3eb23702e000acf8cb2950aee8d338fc2f58ec18871de2779b5a8adb6f018778cb92da0a0ba42c75cc98713929f288963be6156a89210d5652e4547;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hea27de41b3f1189dce3739d2efdba3fc2e10033d9d0e0b10838d09c95a256aa4013306edfdcf5ffb112505f35d11e83d1582d21370a7ed683c8fafe8d;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9a13bd49ad405ea75ea294b3d478850b27ff59f7a95336cda259649d4e5640d3d44212fd3f4399c27e0aaf32eaefb3fbfe1dd63020a465a052bb1fb98;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he25db748b2ed3ccc1a26b24325e128b212ee89cca1a061bac9dbcdb03a20d95dcfede6abbedf0fcdcd31a535c6cac3bca6c5e9170bb83a74813831869;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdc0e9cc217fd640500d2dd213e7a5afc468ea385a0e2d17a12e698c33db6702d8c29797817e7cd5935f6ec3853b7f96ee3d144ef8ed541580718a088;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd0ea2637eae6e290724dece34fc72471d4387d9c0d0694b6db0368ec216e1a4fae2690bbe65fef392e1c3ef36e6f552f2063dfdc7790e8dfafa769b3d;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'haf26ef129270d8f6334cfe215f26e3f6b9d715955c79292a13de755fa7ab1a8b31a79f481c42912c31915f1ed01d6fb3e669711907b7e8a6938c91da8;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h75017fba7c310bf068e727743aebd5dbbfb4e9317c375faaae1225b4a18cfaae5fb85799df6b4ba0691e12f2a464d9f829f3eff8b134e46ed9a8103ac;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he435a8ce78d78b18fbd80cabc4e1147d20d6abfecd3b3df0228b7817465acf682ffcdc4dec03e2075cce4932f50200aa3edff4a3d3e6942ef4645bf8e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc76a3fe7512620cc60c544da667cc2371d1551626d7b7183919c963ecf5e00db0c170422a5d5a0f05d17b345af06364f125e267d9da0ae9139daa58e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1d9a0e2c6738e185aa8a081def13cda3c0c4c7cffd282793174f7c6c444f1682bd370094b540c0938f02b28b59903aa48b8531da443a2cd19563f3e06;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h443615f50a87615a9c9d741fd14b8b4b851b772872681bc6904bbebebf74245b786727789fb384153e04582c6bba72c48bbed53ca58aaa1b68addb6aa;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h56b50b0295e8455724351468e2f3b3ffcfd06a43576ef99f07a231f64ed6a0c157ebe45bef0b876deb71b66603daf1af58479b3b9945f8a97b83f0b75;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hcacfa6bf7abfd5638bfeded7ce5f57e4f9bb7adb5e0ffeb5e6ff5ae05d6f312cb67050dfa9b9d5fb5bef7a71ea2b1ab1ee5bdd7f456695b25c6e58e73;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4110400a45c31016902674da38c1db1e8bcc80595316b6feb6340f4baee66cfae46184c41ae423c55941ffa025a27ca9fe7e3682c823ed9755d67dce2;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb19fbb8ce0a669a3e8e36a75b5d223827b92b7f2f708737d9004f295629581a7195f1f1e8391cb7c78bdde4c8ba5d734922292f0e7cf72949816e30b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hcdcedc727d4a76fec19092a0ccdf589abbb4c67330f31e085bf2c267bbb3a516ff8b43e7ce2810d0cf98758c8e2399aac5b4c89d847b2ac2c4c409a66;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h40e1c21136ae8d9ebd7624acd4dccb9d27909ece7878c8b735f43256e2eedac5633272eef53e3430eab140df61d3a1a75a932f8074d26bc07719f82b7;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3db08c5116c998c4dd905a1ce7b0f45c98210c5202257f743a6ba067d511d343a6919dd03cde02dadf6b3ad31773a6e5bc914dd90a10b80d7f2a75a0d;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h806aefd647be51f0904229b9110257f3a93336e7cc7e238a5abd98b6b55fb3b0b090c4fd8f4030903b1e1c908d19657742b13ccc15e3d35777bbe0d51;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf0a92baa27de4c984e7fc96fef35e29e8737b224cee4cfcbd4a4e72e382dc26648bb70c3141db97d08e9d2ac9602bc711666a0c4ff1114472364d8492;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h12f1f9deed5b9f35fd20c0bd4da9f13ee9dd1761269b2ae539d5a0110fca179c1d769cac62eb42e785d872d73b95c23a04cf4f069f10584250f2c7784;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h74246eaece61644ddf1b19ab50e0c654ea51c1df45413eb0487fe76f69070eaf18b93a5367bb3e40335efc996e83e23757fe372f41938db8d5bedad56;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf2eeafc04808506d9cefb2b2acb524537fe6c072b10daca660c7d4dbfb614d69a36b3991d8baa1bcf17319be96506f615386f0418984dfe91ba2f35f2;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6dcd173ac2d236a1a2a9b92e6bda97218c237770d492a9279cadec995968c5aa0038240d25e4850057fb510d0cf9744be6a1273c67d68276e44eee601;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h52a9bc42abc2bd2a522a83e05b12f3a0375a49e63c32706e9e966b9678ef005530ad9e2b2e6975c29bb820594bf7de02480bc2fd45aaaad6ce9401edb;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd3ea5636cec7622458d84a2f74b315e6e67f0c98c3dd2359b8b3bf5fe21b01ec13a38691e612df257c67f9083f142844ce1ee8e336d416ba4a19b1898;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6df66bd86cd58519c2c35db1f6db126fae356880784942a5c440f850a22195febc9f54b3538a17bf3e56fd969693652ea961037ae0620b81fc7d5e41c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1c274c5667dca13155691b4934572ab202be47a2a1de404c1a822215bc9f42b3eb1f9a798ec49b9133cb8cb05f00db1601e203875b9a7e5c1249ca5b4;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1b73936f9745b7da56a551a2baf01195ad0e48619da9f58151dbb62634e73228110b590cbc22fde01096b0d0e901b1c42e195e110096b19b78ca400b3;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h793183c018e43ecf3f5e3b039d807ccce902442b68c36bb1a0214cfc114979ecd1fbb5ea207a52e66fd8089faf956d722900a38bbe20516237d076bd7;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7d94108b339f79a863c5c24492c81597a3d043bbd297a07ef2fbfed201cfc229df095c7b5417ae0bb7a6197b6720d8fc9f7bfba3d0efaca87b339a966;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6612acedacdeab1176ea18ed73267c7d0b12c5e9790812ad461a8a635569e27fc9f86d70a344e2c8d3a4f0cf1800173ab7667d802e93d9ed10c3b32f3;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h258e310c9ff6ef4e3f619e39e9e96f402e20a17fe2cbb45e900a75095a64987814212cbd2a5bee3ab6e482964e94f4ae802d3b563e37edf06a9cde71b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd6846e88caff5de9e3a2cdae32f00d078146217186a77b2a6f1ac914b8cb58e00c9cd22841c7f3749de199821d849422f6f65b6ac10cfcfabaedb6f5e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbfd690b71e9ad5063917a4c996609498cc34dbd2c889bfde56a8ec47598d160d4b4c2042b020c931dc8dfe7259548c5a4457753664f4bf3bb9599ef50;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7a6183281688687dae73754881ec419bf90db4b17986391cbe3da120ff94b48007d3a2fde262a5c0b29f7a9c02d0913a561d73630f79da26eea9325fb;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hcd1e651db36298a184494efd2d32bd430d9476d94f79287be03e925cbf37fcd738e10c628cd636d883bc101370ebca8a9b1141bb49bed5f9b1fb61deb;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3b7eb9fa975b9c4ce0417f0e81804f263a21476000c5a081b4f62794c210a241e99f7e11a2872b8b59b8da8342440bb2e115e905c0ab5ddb7869cea88;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8552109a6e720b00349835d260cd8fc62712b9dc5b3066d5203d37c51d011ead6dc4359dfdb0fde2a5a7b031fc70b6e2c438dcf4c7ccb9a5053e85e4a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h98f233fec401502ffd2793d3268f35c54dc089e53254cc635471561e816847252e2e1a24d6db74452b486f4e8f2d2e8aa05e6a3561afa21cdcfd4a1e3;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h86e88d39a9c4baf2aa2bc29cbce12aa761e19a61daba3785b3046f3f95ddc9a43f8eda0e18f52da9e77f5887f3264f1e14175a3a61dd9136d2b9bbf92;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3167aaad42aac95b4ed234dbb0c3bbca7ba51bedb9e4ae807e2ad4d1cec397883b1a73e870cc787003df9e1720d81d0f64baaed4e85d7d389ce3f8346;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9dfe0720328abd4fa1af08f7d63fb8a4553fef106e7d1f92cc30b1ccca40197538481e0bf3ccea723a80e101fdf537fa0ddc0d55e3193e9adc4fdb1e4;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h650f8ccbe699aadd538a55eb562b1997ba44bd0cd32ca56b04d9ee193051bc2c0224b0e5c97b4466eb2aaee94e72f606bba473f94bbfa23596d563667;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h91299a8149a16166de02f409c025874ffcedf38b04603de73f14ef1e3b71dd6760abdc5dccf9ae45bc90d9979b826734d989467e395ed09458f443a05;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h67c961dc62a5ff80dda870596f887af304097ac34c6c849576aad54940f26fb9866360c9d7bdfe80dbb7e2065389e40ac52c74b5da0f12b652d72ddc;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8120ff09f9697fdc27834d179b9c494293014a587ba17151a5384bafc222d66c6cbe53e365443300a103af7135527a1ab0d5f5efd0e04ae2a1668ee94;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha3561f3aa104f3c6f6536222b603907d7bd0433d0e4087d840b88c2dcb5e6060866f9689f21325458e0e0d0d9573b6c3fe62f660d8ec91efdcae4c86d;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7cfff72494e3b22bb249e191db442bc4dd454cf7d662421d895502f1cb10c0d9614fee96bb39e150dfbdc301e30558ba3ad0ef1e379dc8cd943db71f7;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h91ab2dbdbecc73d5025625a7f30eae81fc0ef41592d9663dc4315c5db3bb9397f5e2d59c3d9208c0dbffc07e832fbc150079888f0cbf7a8af3f3c9736;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6803f579b53e37b837db091b58b51c69c53c80aa718c14c64c489660fd81c1ca38173cd6d0234cb916be61c824e164b64f3bc931b08c9c81d65fda9ab;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h680894e5dd8d706fc6fedde6d2b086b546a58f0baa8e6b5ced78fcf3bbac615832343245ddf0a5fcca449c527c433fa78dfaad5746e05d513055aec2b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc0bee02dbb31f7938e0b03d99f0989685b899091f60dcd2d5ad1fa4b645b0f34697a97235d32641b9fd887eca9250e9b15628e90b23608193ec54c3d1;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4a731607df8cff2e9b06a334634a13f0e3cec0f897c81db97efa116e673a546a9ab524d2589ce8604f6ee454098017ff6e7ded9aef29dce45432260f8;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc6ba5f305d5f02e2b2b4c510148c2998e4078d7d4050496b183436fa26fbab21883670f4b5377ec7387c8755fef64ab972e7bd33af853fc12dffb24b0;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hac083c30df34d1296e369495c8eb20069c1c0a8ff7bc91d811f4fed51917167749792a2a7d9590ca4260906dd51a6a1ed79dc04eb59b6c83fefce2f52;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hcfb50db496dbc0ba69eade6c5579ab9f00dad8cd080d1bd3a0c71e038aa17cf90054acebc3c032b8a9d309228865066195d222f06bbd73162d17ccf14;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hde4547ace6e6400a76e52e522312b27d93dc805be23b517fe97a3d8113aa1474d6d769d77f6d9b59f13f6e52c7e41684bef1f440ff0cb2d52debc8813;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h27c3a7abd75662710c9480efb36b83460af7cf3e8fba650e8a354381e944e61a052c6e8e26f6beaa60d29bcdb108ca1af7cd565afb88b330364c56680;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha29292f67934e4e1abf054b955a8f21ab4fc3827c2110338779fcc6ffc9d01df1f5f069ec1a8299dedda9390301b3bfe11e78dca5b7877db56ea7e09b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdb59a992563048e3c6d2584d33e09ba7d738072fc82bd8043a75d05c5e7a3bc6f2bc9a138d1285fb244aa0916b78fb62dcbacadb693e976f8a1f18322;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf04119ce2d1eb40889db022b47a5a43568516247c28f112303ac606e982b4c14e4d1cf50395b4a6018a21f5b7c3d37f19839cacc670a3581aa8a993d9;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h74a67cd71bfb9e90a7352eef581efbc58a6b0da7ca49b7aa6f7b9e116aea0011a445566c421d2b6468fa3ef22ee9112072e2e2846ba7bdf4e33e0d40c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbcafb73a7479fc0578e7768230f704bd08fa3a18a826ef6f6de5559bec97d2d7975ccc5590781d0dc7c58c301dc0758b32f10a29b56edeff589ef3199;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7d7fb7af10ec3566bea0857b2933ba6f06807878b84d5354d490eda3713bae3dcf377f91979d95980fe2745f17dcb61c96c54e9a3283f261caae747cf;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h819945c53c7b3bc36f93c38c67e4d877e81d3144aa39f767342bf134c41360b5591670dabee71f0f9438ea90f1435a379db56ea816f33fe5c77a667d2;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h276e1561f78a1849ec4eaed98e29a102a6ec3154fec38ef9da85b647b6a837cf5072d0f3d3eb1040955d2171e89bdb2625ab9f8abfee9b80435394a11;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h18f030d3865a409f2d170d7d5342bda2a007561e346f7762f751b4e7abe276ef2b1de910a61286a3dc66cd57ebff1c3867c20aa9a323a889987713755;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he522b34cdca1aa1c0b9e2c507966548961aa0d12a126dd4de57a13b208b1aac25416054d845c0b40f05223e45f909150f6281e6635813c4f2b8ed5378;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he0184d5167eb3174ca63001e710a545ea2e13d1c594b5d1fba3ce8205e6d6d66d7c65e77547f4a1bdbc6238ebd913b2e607d04cc5d01cecb12b541ef0;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h33fb55d9e9da02ff5d23abf8e1ceeee5b0a039da44cdbb70af93dfd485411007ffba20043761a23df592c0ccb6a73076d4ba0156c0829d154a296893a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8302d28d73ccd55fa39a3d892b08635db82febe50c6f2f2591378f3f31cf1823bafae51d890436b8d973b2cdd14c2e2776c57315d4f6af79c5d9ea390;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd14b8e896c9ea3b953ca15618a405704c9327af4288652732946401e7268ab2000d6acd4784d44790fc29b5611d275dcf766092030ed2b608b02cc017;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5ee1b1aac1ae7911ce83c2fd10cc406ee572810db78512d4a69ff69929246b558f1614e2d870cfd44145f6635b8411a47c53ed6f11d8212f95f8a84d6;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h860d8844196c5ceeefc90f2d755ae0b738175a16c58d23cbaf5e09355f08294092382132e41de83c05755edfcec897343523e0630ae8166f3fa722165;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha78d01b8d54f9206f85a8cb7553b5e01bc57b23b0d95c63c06e01c58fce0ed9026468d5846c13ffd47c62f307765ecb42895889b6ef6a53719f8a86f9;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbe58a1bdf00dd88ccda680a1a538b082f640faf7a2ea0d574b4b69154e1ec4d816250238e772e6fb026afeb6a6c514a4981168877e113829c724842f0;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3e4ca4818fcca007208a6e60a2b444e440ff512c6d1e2ebfc039ed5f74af47fc8a28f1da99164bd0119e0ec3b666649e772bb0e33744f17b2ba0261a6;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8fcf47dfaf38a865b97d64095aa33f22c3c0719f7ec29ae386cdcfb8f1fbff644bb5199808c17b497173059a987cf66908ad9b3959a59f1c0bad15b93;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h44d09adc156b1402b52c4fb1bd60f64c90d2e1d1baf54d3b3e367d45f20dc6a29c815fa8a995ec8faf1e05c6406a160bd9ae7497b6008d0166f809c2b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hafe7d9a8f03125e8d50d395b5226989a7731ff4a5e24c5f5537fcd92f3f9f7a2573af25ce0a7d7570362773782aee9c58ee08288ae860c6158a236062;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd0131d3fc3540fb598664a282663378fa8d3e1fb95d36c7fd2d23413845404cc71fe61ca13c36d62895c8f690d1ad82f537604e02d1b7650f08388596;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h853347dde1b40c6642b9af14a3999a00d92a3087de0c971a94df875eec8ddb68ff537cacb8a2df7485c45574373230f98f57821b45c756c6813253db2;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd496dc1beebae727103bb0a3835b462ddca57d14b257642a4750ef5601855d021591b08a7beb62edeb1ce73b0cb0f394817d4d1f0f890d574726193a8;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1be0a636c798ab2bfbfe54ab1aa4b4588da1a1b675b521f158e2bb78a96a61a47a5705f0080bc48800ef32bc94aca0d6404fa6eb0a10a544ade156309;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbf41f02eafc0cb23d8d7cfa6666fa4560e9acec9a2d5476d709924066be62469732cf9ed2a9fa8bd4362cab440f62dcfae1749eed7c54713388052529;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h99d7c7a6a1c7d6de566b0f9e965ee28cb7c327f1c1d9a11e19d41109f8e02e4f82471e2f12e7f661d7795fa8e8382d9ed98170b84707964316fd1a0ff;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1e827ffddf1f3e8b20cc067d3b79e63416cc46ba8de5c8365a4b923b10ce2630835c46bee467dc462336eccc4dc6b13a404b3f6c7ded06f143a720d05;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h66d6b65020dcd642f64930677bcd966d7dd31841bbdb556b89a602d2a76ede670e86e191327d4c9282581e8f4b90e9bb9940a90284b9c6880f2c2ac1d;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h79a138cf6c6601178baea28348eb4444384251246a46efe35c43bdba6ba67d3fc898b262094d67fbcc154db6480b187e032064f1fdd96c6d08f8c27db;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9b4503a476df76ac00b14ba1235d05efbf67af78a5109688535771b6b0ee57b0a18bcf8c569d43bd0261aecddad2eaa7f60cb610f5413c5ecc35a4f92;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5fe59796784d7d4c1cd376d573adf30910436bc851067c1c4f34e4d1ab62a3000d3f6e6c6ba47c5659c48e1d087755909a32f8696bc38d7a452c61ca2;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb3fb249803e287fc9ffc61755241ba47429a4bd2307413f6977f75dd9ec7036ccb9998d104a46c84687e99e8e90122231276ce6e007f8498f51846ad5;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hab511e35526e041e77f9ac948113da489668fd4fd176c51f87e571d53f94c4bcdad00c73b0a6075c3021eeb7ed5d86efa1a4e5c0772f4c16683826564;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf8d2bd0208f41e24dc114b150b5d2fa9c0d68bfeb4cd4cba2e2edbee47304aadc430278b0e92bb1b812102cc723a20dbc8a1f34f8c09057e4ef391db9;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h93127b4d3fea5d3836e289ad22fb0dcd9bdf65e20fed54ed8a91f4f5756b56dae211020e3d8db08f2e49fa7ff8d4281fc9086ff15770620ac9abccef4;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2ded807e60c4aded36b6f435dab81581d8543eefa4373a0976b83668bd69e6fe99c05d28f8bce35e36171d2b0e7b828b1c330cc2cc82970dfa27e144e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h95f590cfb4ea837cb22b785a6d3e7189d5d5485a622139c514aaa2b026478e4aa2ee6b8d003f74e5aef548cc768f69b5dad8b11795f99e46eaddaa546;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd3dbee643f72651cc4507441c8c4eaf60a30ef52bd6fd4c52061f2c9481847feaf902f367eb3be74bac1929b9f2344f14f4a35b47e5ec5dac64cb51f7;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3c2f5700506682481ab8873e75800de9b63ce2ad04a98b864873413bfc8b88c5233fb3d910b7a12f3122efebc69a1246f5e05d1166cf765c5e0a3bae6;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf5f4ca3692cf5b6bf8a60f722df48bdeaffa7ca1c0b1f6fd01997b901140eb8fdb2becb5c7ca2c0ddd6cc03d418f698ceafb81d99b95f7a8edf7b7669;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfdc1928ad1f660efa0ceaece8f5c9a23f6392c37bcdf096d3d0df76fb6a619bfe0ee098946083902131188a3a1119fdea5147742aaa0ff1cf6b4cef0a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h498c808308d29f990db9abc72cf2ce8c908454c83fd5c480da78f680f67f598e7f46e4d57dae2d31e415f5543f381006df6b2bd3f3f3bc5ed98156785;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4b2b3b20bdcb9f84dcae42045b99e48f402387d41fb02652dbd2af2d9929f9de58540507d46b1a632ddd0c5aac5dc52f6d7e7eb92835922d520e291d6;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h567769712ca88f0183bb6d762b5e40007b8c63c708a8fc7a943e5be535184b43b8a8c4d9f824e558277d7545c3233e35c43f0e5b6d089e7ce3ee0c7ca;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha3f12eeecac41022663d9c794207b67a8758eb6d0abda2a2192a126944e44b781317d88bf50a2e4c2d20c96a59d0f152087628fcb9f5b7f6dbb1f04a8;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9554641e6302821de58452ab40241050f3543402155cbbfe44b795653d193045357094db2b337113d5b4d80f58cd2ddc9d85d22463bbf64cd41ae9723;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd57ff9daf313d4b3045533d775a87d3a9680507df758f023d145ce9fcb005cbede6058e9a126069583eaa850bf9d2c3a68679efd65e06c1a81383990f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h91c93acb42f816886e8d00b97c0791b51cf4dfaf51233d777a686fcd70592286de24399df4f938925ee156c546846059a78dd4eceeac21a2c154a1dae;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7d0c517d4aec40cb1e4251465c6ab0be3d63f932b2e886d16ff0660d6a8cd01f827359975b34a7d5e288c3db2d5cae1dbffb1689d2b32098afc1742e6;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h309d07ae07841d5e459744a704af3f7aa66391948b67ed83b070b9ab859500816cf21c05840e2e49c86af66e080c2b9023f896660d301ae630245e074;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2df5592913a286699dc19943adfa6121c66f3234129f9f929fda6cc23431eb1f92366bc55f65d901f25899087d9100a59c3ea4ed4994b24f00a3fdc5f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4020225bfa885970a0808eae49e4b5809e1ffc4cc176ec9c6dfc227913bff897d177fb2fccff0a5f9b13e592780689da08b9b2ff75ea525955883e8ea;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1056c4a1b764b4e6828df57c966e2defcc96c7acb8cdb8409e7ee3e5ebf4f08d1f0e21bf46ad823d3b1d98aa0aa88fdb47ff3a91193e2e3833ff2491b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9310c7b36e6f5b1c3458d03f8ee33cb5c0c95e745e3f28e935d3726853aac855531565286f9335f2528a63646680ea029e89b900c704a58f3197dfa3d;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9406df896553dabcfb1745ade2f7ba6d91e54d687112bfb63e506750dc6f59ebb69fee19c65a9c4db74658a75024b4800d347ff48d70878fcbe4ece7c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf390f5eb5d6b6e4d18da373509f8d7f56ea400f73afd0421b9124a67be7f30b46c0925ae2250b02635d5b623c1c8671471e0866ee5018902b54964fd7;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf61d2af5e2e1fae5add68c6f4b67439b293de63e7749cb91c71808edc4a2d86d9db7e85597ca5d673e2eb098a54a3db1b6cdc0ce3badfb163868f3aa;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbfcffd80249f606b85e99ce7c006861e8514188cb969352aebf901e5bda5f0d992cfda63c9d9c19df7c22572b5f6d42462cacc05f08bf784fffc3e384;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h40cc2492c85f82540940aea10114a46f74e8d814d223de10ca08ca33a20dc371aec978f33097376cf1140d3f3a62964decf4ce05650cbd8b64fb2a8ae;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8287dfdb7f7a4fcf3d5d45d1097ba9cdf34305ce1d0906bfff7b9770508b40b0f7e4332f0900d7b4499f87cf9bbd39dcebd76a056a5bfdd062a62a883;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf67f2ea26824f0b97268edb49b2a1b9586fb0b2b935271ac63f3a27c9d890c5bcf13ba7c1f09e84fdf6a45754a1c758623e323e6380d279dd4bcfc04d;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd0eb2efec31bff03b2e2732a32aac17b94983006ec14291c36aac174b5086a6abc2533e9b76559c35f827032b1dfae6234a2c04e19a0c68d6ea627658;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4bd2233022afc141c5a6aa333a71187fd9c78dc1d5407d5884a674f8e7634d4d139c17a01bec8a7bed48822273c38e564e88483b4ce35dd132d2cb2ef;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he1ab1a1b79f19995589ed2977e4cb5cfd88b7389566eebe41b28a27d8161d413545de72591ef5c8c1aa0e873dcbeed5b412bffeec785cf12ea35b4183;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5e3ca9ddb2e11a3d15db05a920e1310463022c63a90729698c823b8e42c5020e28be511edb588732bc0e0cb9df2618293acc4dd7864d3017a86d28206;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9dca30b51ea698c84f12049c841f1e16f4754fa99b7df32c878e06dfa9b5862217c638e229f968885eb4daccb1794604e6277481a702789147b2dba38;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h74da40106b106e00a1b738ed0827c1777f579396cd589ca87c8f2102c6dd57503622b1708ac937f0361cd77d2796e197cf5197e2ebd7f170723cfc75d;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hcaffb78639fbfae409375d41d411ce8040e2a33ab942422920e3fa4f77d8d82b5a966adf503838bf3022d00ec6ab70dec37ffa111842bd42d86ccfe04;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb88300d7f10c7b228f59e80ff6d6c767eacbc668870c93a17b2668b3f48d164da23608b086ea85802af3bd661c161c69095636f9f498cda6828a90451;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h932068c13446d60e86b546b6112144d3dc7ec89f27eed46d8b643de3b80705c0a67bc85f557ccb011421cab73891841c8a244d36325aa9f8a0495a9;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc092ac34b2003eec70d4836ac5e9352425c46df5f654ea62f05652ba69df28ecac367efad6da6c02d88d517203c5f9892e4a3a9cb37b9763766a46bfd;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6015441d558fc4366a1a885c314640a824ef30abd7b51a5c0f7e35bcf61c0c6ecf3c9b1622ed21888d48a7f20d29a7cb26389a02daa7376df261eed5a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5ba13fdd19ef8894185e9e88acf3d0cda4bd5c35a41805d41b71a5dd062884ddafe53f4d2656cd6bd57dbd38d6f1fc8a1bf94065773d59114f2b95563;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h41e18467f3f45f90d475f6709bdf588d4f5da94bc548eb7065820efd89dae90905d3758fffbcb6221c7c2957a76f3683471367f1003d3aea2dacead17;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf3b16bfb4357d322e94577e9934f8ac3345e42d441fa558e5b5a0cc0e4b02a53f10df02158239819782469207cea30df1c50c324b59eecb04aa278bad;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7baf8d8a0d3d7df671e9b22d3067ea931553fbac8dc6d8ee4c1104059c6234ffa576651148d6acf20f9f46d65df5a0c7970c777255802372f2bd13559;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9e5ce8cb11d2d31fe68b65f2319bbe79367da3db97d3e95cabd80e96fb26a7cd2def925b3f5ea82ab943c50656212cef28acae5345a85a8070ed19fe0;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha8fedd51ecf530b080c6bf852e626ad841b670e2225c8d4c843ae58d653f5eb8f3fd6cf7f539befec98fda02212652647361fadf79fe1add260671fd8;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5c99cca591358525b20837b210a169997d1db614e75c5c58f7578f2b474c84a2e502b5529c66ad23fd9f905e4e100c5dc3d7510708f4709f6adaf919;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h173ac072c7652669c04b6849468ecb08bb6c2d62640d5b7b7e40873789410f0626ff8d3636df8924b10031b9278c01f793642c0650c1faf5355928a03;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8133c5d8a7ede65cad7098704839ef064ec992994eab526c2192fd42de28bfc92a711900eda00c4683610ea1b0af90a852ff0561997692f40d11836f5;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he651b3c023d7dfe87fb1715f16506823036d066b790cf56a5106429dea6d75660eebd97c0b5462fe100a05894eb4335154063418c959971051d90aea6;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h85741026402e4f0924c57d6c5c052a93b24d8f9870884ef2dd08b423c886dffae729d39517bce6f194d95a11525101c63cafd61c8f3d4b6e3be335577;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8d1183dd690956afe2350be72a4d7d6b2442ff95b76dfa196f2ee20ab9f5410578adab49053887fd70e33800a20e34bcdfe12fb8c8713d4d466aa16a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4a65dce6a4d6c7a08a1540a7045435090071f7c79562b78187f60276b0b4a225a27c7e85d25614fe836ea5c10daf05a300214b648e45711cc5543c91a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h31f49bdd8d7d48c1f0124042e651ca17c8ffbdeebf172558aa4c029cd3c2259a2f18079fd42f13734d04428a00f97124c7ce0ea85001e2949a31975bf;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd7cb2c132538c840c500a4ccce15148e2703a43f3e74a4b150d8d300462e13d790dc980ccc9eeca6620fc38f6d64bc8ab2121aff7b3a45277d79ba3ce;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h34cd3bf2a596d2b98ae4a7e398dd77eaab87a97e436fc614ee3a27a36be5bf8962a76ea052dbfc5cb679e895e60e315d208ef8473e25e333266eb4597;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h431e186e55e78faa1754b13eadd728e646bcc59c0efdeddef512788336e9c787eca60188f2cfffe6c9efcbc4bc12afc17d6003d0cbd849f4eec5654fc;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9a96803712fc38a597ad5b90dd18aba70764f05e4d72081799f90ad77dd5a230f358c1bf7369d3343a205bb660d282cf67909ec8683c4e9efb11cc5a5;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h278be48b811ae31e7d508652bccd127d3c252429f7874ba4ae2926553d381250153ab9f273762fca1107fd4807c856691ca00f4f13c34909728035cd9;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h61c90ed3890ec3607db4e1e2270ed64568a205d1644b5b2ffa6c6662a2484519f2eb370b6857a4179a215499dc492d5cc2adaeb2df75dedaabbaff421;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hec7286ba24d053579a46245c5c78ef2225c010feed41ed021a7348afbd8adcd718485e5f99bbe99d971fd5f0016f5f0c937b3afb43f7fa182ac7ce00f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8116af5e205b47525b65fb7a8f7a80c34e1a9e5bcca35802734ca2f7568ac88818aa64dcdd92b7e031224dceaf415b4a2841edc01ee84abbd07ed27a3;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6eac4290d7220cde11931fcd86d5a199f64de2843000eceb6ad3b047849f7ea1b1255a8bd5b9693bad5f5be2e953463c8c6c9fa9d21ee4e9f076afd34;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he2e7ff79df204bd0cd2bab8795fc2a9d889bf9f9192bb3be7e12f999801b7879bfae5a641ce930490849a7b8dd78ce721a80bc1bb5aa3727538148081;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7868d312217a1b0af7f5a06a1a977ad0cd37c6c922cf63191a375e190292ed88f5e56ee7c8778adf53e513d45005a3dcf56a64d376daede9d6541952f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h866cd1a20bd409c3f2c29301e58514b3d1d1ce234310aa203a44711b6136b1d42db3c02b1a55518e047eec3a63aa5fd67a9809f4e3c557855a31ca600;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4ed24cab0c184742811b4e0a152b8d6d7b91d76e172207acf293d40a88e687ac0d5b53b318664e8b6b98776e30855338d1ff095f07b7741aa1a82375;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he75abf90a03da4563d35755535adaa18f9d455b89e9235c4c8e94aab6b1634f0caad9eb129cd37995d55b68754541cebdd92afbb8d3f2452a83c4604e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7efed00b7905ff26210f49986f15c5ac6ff0a7f04bcda3cc8cad60bdcaec7d9fcf6ced76c561eb2122bff7e295b0036a6ca7c92040a4b9fa296b49d22;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hac0fbfbe49194da515904a3b2be931a7a36e806fe306a699318505bedc265cd6962dc4e59071799af7078f236c9923c4cfc43078b54ab2b4dbb617c6f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf7699e0a0795afb2ec62e95417c61f11b6cf524a760721b7f396010663c6f7da128d8a70f19ff4f61b5362430d80881b917b8c5d7a59844fe640d4bea;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'haf2e8dcb138460ad261ef2b4965e13905b504594c561e298a04e247ca7a9e82ac30b5ca87823712e9c78fba8a4d2286e81c810d27025590dd8416c508;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h51928a92ceda0b40412d4f36111bd25b6c9b72634df169815094b1b2263c13a59bcb03a0b67dff3f301d88834d189f99e5d429c93b2e8b9e30dd0811;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd2c1f89d5f70c66ac9359d90101a84e52b4faa30aa75cc3c8554a579344086c8262906615fcd7ac6d539350288ff83ca033657c777544e0f290b762c6;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h30d965ad35bf8e79d1e766ff34f5bd425f0868caa8c6078ab247f059b293609da98770956df3dcb1df517a6c66f2a739c0138e99c2c4062458f2323b5;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h99017f547b1f47241fe013268811099654bc07a9f8ff1d99d51d2594c70e0b1a489bd5beef54de026ddc84da9cb6cecc19200121ed1e3d675d25e3d90;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h55e75e1855c27273647b1708a546d77d17767b0781e2c518431431ad57427739a8ea350956a3f6d335ddc12fbc649d658cc54abb6a94f1411370f1438;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h45a764af6ab07822ad3e93ebfce5294eee76579fecc71444ad78cf90c5f65417fabb0abe919acc10c39365d9f4a4ea612e05f40b18aaace8665dfb877;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h99337ff09168d186af92c8c3704309ae016379159f54eb145f90d73a0b0c5b17a18b5413638efc834e9858949188d7b7feedb9b0e5f2f3f6ef18ae90e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb1a47e75fc599df59dc9968bf1538af883001d60eaca92c2061f96148d98c4c8199328aa103826327571077948f6abf80ffda417610b0f7a453a844cb;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h880249ee0feeaffe3c70f16e301e21a33b580a18a86a46049c7e9b542120414c53821bcbb52b0ff13f2531fb3189692306d8a27d6b4fad01e1edb227a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9d50831e49415856433736475147e7028f2ff1e25ff81fa9b13ee8f935c4acb4d4ff17dcfa2253958e1ed900a056c1d47e6b9f1f590ca32ec4c8b9f2;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h162b05f740f2c9dcbc691c498ab64e360fda87a07f2960a2bb07ab727553e28befaca865428f1a201545578bc6b5e226c8ce0b43c3e6e65a725168a45;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h141c886d66038d171648b8a90b0dce2f833b5a61333deef391630cd635a191c58e2413ae9da54702254eec95f99145b9efdf6b098b40b2268823601e0;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8a10060ef38a0b08e817a568e59815c6dac2e2ab95eb835d4f863069bbc65f8e24ddfccc4a8a477ba836e1a6d5ff746217101ddaf1e719d5136c39aa1;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h19059d78d3aa28a3c1a9faac6ba816e80c678bf481fc09bdb27d8a899f3451a6acd19739f4300b7c75c3f3f791cd08e36021f142e5c77b5a9e7909b36;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h61bb002929dd28211db5d39014141fdf607c8fd9c897090fd3b7077933eeb635b83e4dac76a64db0abbf0b35eb458385e52f8ce4091a40c6c49b0c723;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h948966e3f9bed4021096bf17913a35113c6dd162f1d32eadafab06711536717b7d82593ff08efb75def2161f8ad231d9c479098111d1cfcf01885a575;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h560347e3c9631a76af4d225991cfa20efd50daefa68af3b05ebbf643081b6b6aec2ba5ce719ea14fa70dafe8d2c24057c86cf5445103ddf99567a7f12;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3b443675233ff3dfae148cde6f5e092306650e20355ba0e013480638575f9571de88a0fcf69d8d67dcd329d342e69a06c65a2a550355dcb4bffaf2373;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb4752edf0249cecda6faa7384d0700a5087e401dcffea5b4531bc128316c551a5165db6abb55104f37c940ab7b5653b5650dde20a454422b4ccae58f0;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7390473a451763e699bd94e378393c5a258cd33c962c8a00c8573f911f7930bbbd97b8d156f27b48a5127d04e251e8ef32e2b6e8c28b9b84553169ff9;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8bcf83fdd5973a7084198cb5a600dc880c07936b0c30f46c3664782a7b3b9d791031f10113b0fa1fb7e6e9e5d81127a201901869bac9231741d6c7ebc;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h337a17265356ef17647cd796a3e417c0196fa18028cd7a60ef7cf3aca0f383cb37213455a45a916a3944146f45218805f7b9dcbeb4ab836126b607529;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hde31c30b0a6f14f7f92aec94c7250689e7489743c7aaee3d87da1cb17c53219778a5d504880ee9be230cc3d6d6e5be08a2b4c597e7a621a8f966a145c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5839f88054f553e568ddbaf5ed560ffeee9144da6cd7373e07b3fdb27efb131b2a15ad5ac99da2eaa00cd1659847d6e2887e7549e62e224861b09c665;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7c4980ccd0bc2593f6532192af89ea5b89c68148a23f66d73f74c628c307c01da36044c2834db528ca844b117a5ceef2c26ba5bafed74880a3530ec78;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h263cd57fa3060c11672b6d20d2748de14a7032f091ddff1f1425be8d225bc8fa9b57ee782b8dea15e67fab79ee3c97750038fcc82918c14cab92f2fd5;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h56b4a25307d9398adffac933414aaa0d96a7e850377fb34e68e1b4fbbe3cd482eafb674787d8405c50daa7919e0f064f32fa351d92802a900b2c83252;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdcb595579626a7e3f9423c0bda98cbce8ba03e6c98720b5d8a8a564c29cd7f816a928427ca11cfca396141407c911290bfc850c55308a67e4854e2bc1;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he86121b14b2aab31c3ebd653941c6d7580113a6b47577fba30bd316941029774c8c3e070a4473b2464dfbb9c5d7113fcd965867bad8bbdb87ea9c4ef7;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf263632cb946acea1c78556dba5dc4a96219e08c07317e0a519c3522766d8dc7dcaf55e506b6df9cc08ba2a2e4772de8ed387439d377fbc1545ab045c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h484d8ec322f5aa202f7c08ff234166e90ae90ac30ac960eec88cf9ffb29a4671c8203ef31944f66f8409cc955369877d33b4fac6e17efb3ab830d073c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5a3c42e4297c0db48b757497a0799c5847bd24d5027c2a2ecd91c570da67a7b57621d76cd57f924585dd63cad7e6b988efb2542c9af5bf2a65d813155;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2128cd67eeae3ba9b8ba32002f555764a46b92b696e2123aa8fabbd17ccced16e2a3ff870212e22e550f3467c30fde1c7c571dc97367edec00c5647ce;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h61e1fe0d946406fe8a4749bb83faca139e8e3fd1c4f242d5aed7b3e5c80020e73f8f5a8423b6cf29ab22e22c02ae93d730e191a3bd1cab40c358afade;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5933185547617d7339cc1f6ea23015981b69e7a8d2fea33c237fb37fe880565e75c6983e92458780ebf32b7461c8dbac1695f2323b490d0cf18f311c1;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h90e85d3d3252ea640137792683d2e6be8ccd2fccfa95ea617959d7b8aaeb0f83ce6ede299b0e513134f73865518a331b9d1275f7ea82febf954d0c9f3;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5b06c401610733b5f8aad1e6dc7becc56002dd0c3363752d21abcc4c7921eb33bcb7f53fa138ee4129d4f68744de9ca5a371496196df3379a0d309ade;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h73bb4663c64d2576e092ff67d0af3497b99de888c8dd1b81f0b41ee9cddc2c422c1aa3fdc92e78e309b87ce37bcb317ea459857c68d46bd9b8f7ab5bd;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h329eef5029dd464fdcf94e6617b02e3deeee519cfd99dc8080d76bfb4ff83dc4524ebf72465328356ede88f0fc7bd9e0d929014262eabaf8aaecf626f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4a99ddf81836f8d5cf4bd0ed06ee625839796649fc530748b9c277ef1336baa07ae796e7567512f4822750ee250053af48ca97d3d8602ed4be9f1b134;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4322a94b958f514fb31fc45500830972e31027fb875ebfd14175c777c7cb4d0b740455f84629e76dd43870995c886b279027f59173693a58b19a110b3;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9346cad7e428330bd382f35bbaed655bbec240d21fb8ccceb31709a380b1c7ba553f2cda38e937a6d7b6535ddf0951395920783d810db5f25fe09cc64;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hec004f992b6bec87f8de5da64e077ca91d55018260174cff84b719f21777cea958b276ceef01a817f15974ba0725058c4b5ba6facd7e83bf877c8a2ed;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha583b7f37bbe426894019473fbbe032b8a0838ddabfefd71798b3e202fa673262542b7a3b9777eccb28b48a6c9832d6c41620a0577be3f771d87b69c4;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h65e15bcf189295a78adba4cf28b16ebf63120a14140f36fe6c927ca2a458b5064e848fcc4bfb897f2ad48b7fd01c252a5b1a10de799442477638430b4;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha98444cc3c312fd0bcc262ae98d5cb750bd6cc30a5ba4ade9787e5e6dbdbf009681e98094594aa1fa8450f8d082d85d15e766e4e8e962ca7222ea02f2;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2ed4e5dabce5bce9f56be5246a0a477f7cbc85716ed9b8e4b63f6a552639bfc122e8e29c51046cf4dfc0171ba8d5757a5d34e6cda6a79c8f2fa7eae45;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h88f695d0e8b694c67cd13f743f5d724457d8bbb7d9763acf0d03294815df7521c3e2d7f622a707e0901a54e6fcafc73a57fd0659eaea894ffb0bf1f78;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3fbbaf59f4d3ed30c7774addc288ce676878083b1d86fccaa699d30adc24ce4c3791c900abe6cfbb38b5ff0e70a85234020daa0e850e755f51c5ac7e7;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4d39443ea88a74a560f1ca5c1c934273a17fc79de3ffcb0e90180a029c455f46e2852be5dd3ed2a07122c3769317c44ece5d34eae9f3dffe10cca38f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha5bf268e068f61a7aec5686ac726c2f1f20099e97f0358114b8f0d0c95a31902333e7ccc9a20fa7e60168757d1a3cebe5a170e8af62217cf45822d1d2;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1c28e16158ccbc25384169d1ee3bf04b560ae85bd0e5d0f86a9993bf3a3894ebd1ed01d2531b56356c45b29552476aea9535b70e4e6c6aaed5094a088;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha938479f754055ac6f7ff9c2759815a9161c48cdac9e7fae28d0b11019332216e26a2297c24d26ff2d8a3885e5ca9fd3c41d4cb0545a1cc316be285a4;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h177c7f7f8af3f71edbd15a5c846a8d076077645c7edb8ea85138b7e7bae1f671b0f908d6ddc3c858cb3cc9ea340c760a83045f479edde28b845c7a778;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbdb2afe6c89af3aef17df37588f1d8cd1b4f6e9c0c61fea8bb69aaa3272dd74624b8e0d3190e14c8bca4271d8ad2d3ecd6f63fe2f5c93e219cc8571df;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc63aefa799851679a5f4f2ed66cfb30f54e65975e0b9174cafa51cd8ca4c1562b15614fba0b8accf8e4643458b7e107db9f82bac37150a6e0104003d6;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hba821397a9822f3ab35b69c0c8282a0a680d9c8ac3b5816a9a983cd03518a68fc83e78c76cd1260664d67d99dce428ee4b775ace7cf7780196ecb0c46;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha527357379bf04a8753913c8c4cc883cebf247722bc508ff232d6928f2e26ae8166c938eb9c786cd07db8a00f993a3beef4f68dc3968890b94098a863;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2388338d198ee88dd50fa75a1820c8d624dbc434e2e047f66a5270477bc89dda4b2f1910636c3c5b5368dec8bdb38c3f1d8de6f8aa5e3871c2a19f69c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf97ee15bc24e8b39279d6038a71b8ae8b2854e55afc49c2d811dd86d7b65525d01c32f3ef1bbc60566fd258e4826fc34af666db1d910631589dc8d45c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he7f520cb5d0f5ffbcf307ac40757de17f0be830409a4372b0f70233ecd27a60c160f21789bdedc23f3f07ca5232ebc59919377a83e1750b592fad74b6;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h581885a9757de381e650609f3639edad663c3dc885a0cbee707006a024a82515a48f948b97ebc45b836925a36ff19cdd38c97721964fba0ddce19b663;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h111d02619ead2d2d18693b01e7cc747943e7109f1eb8c3d0db7a8b7803bd3d83dd68667424cd159d0073ebb9f79cc51ca196ed47c9c14e0226c3a706a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf33e9dab85abd17f40a2c6ece6874a1794e72465d6bf73f53c3d1f497aabae028117842ac21dbcb5b257e11bd612e1f21233a670f924bffbdedb9e2d1;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h66230785b5624f91758cefe319584679e08fb76d6c92528d142bc8611068e2b9c96f4ad36ed00b161e18418dc571d8853ecbc8d3a08ee06088cfcc473;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb53dc2fc61f9f242e26a653aa7cc8256ab89e73759a59a534660529dc8001ff70158c14d2ee15ad4cd358f4dffff47b48d2c69f51e87990723d158d78;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf94a2e516fb0b4b408877e1cd60a9f5fdd080ba55f30617f38f6ef59bc35109142cd32f61895e07ca3047acff5dc6085d02e106421c20f1c8fe0b723d;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he565b2ed507596ec83e7ab34a8173353ae1715a3ed7f557ce1a8ebbc619265c944011e37ac9ce11d546e12e856e82275e464092a9ea4f2839528457c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2a604a999b513e86f155b3b12338ed516eab17d85ec5f3c6fef8d83253ddad5f790bf5619286e4cb9c271f9d7177163939c0d2d9924997d4864fac3c6;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdafd19a68fe397b5560f3d0b4a5ce90df7b99fb7c8628a91c793551c8f84c0f0fae4fa0a1a9ba2ec04a7163f666960ddf47a249caf3644982ddff61fb;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h141084fbd4f8efeb8bac0cf3223590d13bed3621cfe195dc931499cb8fad336c0f506cf8f7083af3465169d7e65a5c959aba8338fd75b2fec486bec47;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h37a7f2d85606d91c7df7e6c47c4bba90dcea6b91a45d8d5ed3b372a4134c6c60728fe7a560b6f027368f79c7285f9e15b9432f4bb41f2a874086341f1;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h55073fc7b15b5fb01889d5e0ee4de9e4cce23d8a1fa335591fb02c605b8416c2625ba8169fe4638b5797c04e73bc45064623b6cb0212e79b29592aa4f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd9c304cfb66f086af8f79c68867564f74166d75603daf82a6905ada187f09a7d1d5491dcdde95cc267bd98c425236aca87dbe823e7d5445d95f5362b4;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h18f83634d09475ed928ad7578da35afdeefae5023660e0059ea5c9dd20a433b788b927b8bba109b1babe647c80d6ecccca87b220d2f99dcdf81b4e363;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4108c78ba4cf5f02e01957b1e92410161c8d49fed4ff6e3a4e2b5d1e118efbef742b4f50343dc01c3e31539a8b7e91c56f690cae52c251196ad9a4164;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3909c3eb0d5b4dc54837e833474d0801fd2b135f4690047ee9df73d38ac96d7392404bfc0d44a68efbe59ee88a6ef97a2e8f498668570bc9499316099;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3611ce5b54b27e9ef389daa932fcee82b97cff79230fd68f27f6e4882a51b608443de9677e474dd493d759147ef9a6cb1100d9ab7acfa1b10a9e81e18;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h57e82d253ba2cec31de23a29ff584bb2f066100ff72afdbce6c0ce8244dd8989c77313df34e60fc0ce0dcf475e738b5601e1704053d1dd3f96e97c7dc;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8f93c7737865b7a64b888ed1b2ab7c2eadb65b8c7d0d45c80af28dd38e85d7dd62bea8d01ea5fd4ab7394d5dfbbcd6ae3b4d91a8dd1914f52fc1089cd;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h851371760f99f27b1de2c7026cdec7ba0faa291552b3dcb1fbeb3338cc5a5d51fbd66522a3367dfdbb878bc73d25ae65d1f22310350a3d998a7dd03e2;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd0ac95138c293a8ce990fca8ad1dec45be00181590ab58f8c1f701310d71ed57f3778b0f38d80cadcd8999dc67c02862293eb2f7af3bc77d10cade36b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h18f8519754ef3428c21ff2a168a2475a8d92ac1bf38673abb344d3da9ccf069511ede2f913f896e85849f1fbc3bf9a73783c3c522483f513ffa5f859;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdc7f111321fb133decbff80c1214bfdfdfd01fc3a892911bdeefaff33703ed2ee67b1947357ba8830eb3bbc0efcbe1a4d1d56de4914789aec39afb4c4;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2aeaba27d690d83b076210633a0f24d298a4262e687871ff7da81a06f8044aab44ea755725ade17dd92e8efc62d78ee0205f17bdd3e0f070b9a1fd32e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h44f95caaf6f64ac5a34c8e5f53ba5c0d673ea7e5d9e9bb5c91c9bc46e2c0763870a1d8f423daa48528942e84787845e2edf87360cbef287e6cf4ce1e6;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6823330b3bfe960bbce431dd3d4e17bf33ba07789369ad5822142a38abdab2a3d9e05a4b48a0b4d87f2abc512c2df82c82deca9c01620e92d1307d122;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h881cf38f177fed5b0bd33784013c5ab6552ac2bdab51add9e31b33fe2d6595934790cf5167fad98fe4c0d33828c6e60568632ab2265fa1dfec8cb2df6;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd448d2234845733265d556028a0df251a064e057a17713bab2124ba801a46a737aae670b57ee3a06a6b1029ead92a292363ab5f3a4583480b42922cfb;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7d2e398d1b98f817a3b000fb0aa7cfb1f883f3005a4b0df833dab126e21844d95cb2320536e3c8178ffa84937dbc862b8499b20f3700e3a7bb9f0378b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbdc42938430fe8b04d4301ee115c266fe3960cb2f9cef5d695adf3765a7f4a81bbd2badcdaacb089b618c4c04132f319c0cc956b23e2f9c3411ef7641;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbac3c4292aa09b6c9ab7d95a4441fb16e7573dd9260254d5096185c0bd16b269534bcf5869c9c7e05c2a767a7c1cbbdb8e82b3ae8d9e2d2ce440028c8;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h44f094f6c1d8a2855f08ee7f3528c811743d5391f25b97370f6042485666a457e5d61b7c7cbaf9713f7f59c567da7acb364893913f5bb0c64d5c6ad2;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2fe5599c6614cd390e3cff713785cbc05a69a8ad24c03def3bff295d528819e241dd54e0419449034238078f0050ff42862bfd8654e597cd3b8ae27fb;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1b4e0507fe1a139d615550b150594dacde8048eb16a5e9dc7eb391887d8fd825f2a06947f7e06b7f3777f04b480137faa694ef93434d40efc82a5c02e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h70dfedda27dfee44beb7b58c701ec635eaad2640931fde75e38fc554fa9187356bd15202f4d6d6ca48bc221e61250795bba2a9ae78561928dfa4b1beb;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc34ea4db7d2dca2d01884adf4d7abcd0d1335d0062979a4ef375cf2afce1231e7136276283f38d01785b73ae28b29b29fc0b4fe20f94f5bec279e1433;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdb815c55b05ec345090633c61a87b03ae7906485d60c020f620941c9d48f0d2042187ab2449b74b02907ddda4358dc908a20dd65862bd911ba606aa72;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha82374d0ade1fab459e3595fcbb48ea0082eb315ade21e87c19b3049fd2daaf67c8a53b6b0cfb8ee5f61a1da90c4fad241b9c8a45f772d062b9bd619a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha88a16942e889f5eab344c2a2e64bf8ea5109a2aa097fc4687edfc217115f1ba1eaabc0a788915b91a69c7c613d3666fcf354e13e660b750e4124d90c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he55d5c3bb4c7bf1510fdb4332b08ff9b1239988b2e725b0e4e955b9b5c8c89c2921d3a0b037ab90e5386266c0bbb3d071a7422c3038a3c88dc475ee85;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h36035f8340748597acdd3daef9c149e17e689910d91935f898dbe8ca3104bd89f807d2cee4acc8db0bc7fb395f9871fba1cc156eb996575e056b5403f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2790a5f68922c1237207b3109e9fbea2dbde52da1f0be7448ce7fc7c9230e0261653404032ee58cc05cb447c7f779b0c3ea2e88bd70d7e90edaee450;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha95dc03da82488e36567638befb553b76456f45bee98ec3d713705944223630eea8b2eb116dcc51a97efe1d00133023288993795dcfbc2e6517eef5da;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h82363efb18998f096c666522641651dae77dbd12dd4f765a3803e7d3573b5ffcb3b49cf8abac5ebcf408428341a8809b9c4d67976624b47f68935b3f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9d587b3c1ade814fa6c9c36f89764a4071d9e139a9238dce2a0ddbac4b432aa0cdccc7a9a5327fbe6faeb1e0e31db04e2d10dd53243844c055b7a985;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5b256d3ca38d5eef4f763f157946ad931fde058308fb1bad67339e7cd582a25bd121b39be31b3217683bb309881addd659a5d0441767eac359f736362;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc94459744ba70a1a9d4698a31583122857b4eee7b747f69da08588fbad9268e9a8620af6fb79f5be910af5dfca9629badac01eba6248fb0c813cb605e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbcc83a727d246fab9149e15f2f0dd42b79ed667fbe7a59a306802a17e41d3bad979c6c16b45d1701b776ef5038186bccf4e74567d80c0bf736539556;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6babbc1263fe52294a30d51d9fe7888807b544135e5fa9bbb4a5ac169e7411661dfe95b8601325b9fabc044f96ec87b939abb1db10cceab56c06dcd19;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha32adb1887dcd1eccad0cf0f8500bc6c82b68ca325cd24ea445239826933a109b62286402d7f416cb88394d4f4641402eeb4db5453da334f5543ff95e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h21eeb26b5ec93ae8465a6b0eba7ae9b0d05acf7cdf444b6f1a839ac8dc1cf169be5ee94dcdb7d38863358a0156e455b299e8fa839e730f9ac605d90d3;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hcf8e9ca27828779e9922f6e11225537413049a74fa52dfce2561dc4c67bd860e833ec28c99a995a7f518267e84b9b2bfad9484cd9a02cbaec88e99d20;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4895d1d1dfd33dc734340baa13fad6086e99665bc5b463d3a4d240935eca06b64c2b09658e951b8e988d47d40608c35e64f322359fb3ff73c8ca91490;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb04f601b4b3764546c63b3a08751d70e92c432439f84a6f5b2a205cc53103867a3074c1c7ca861da6d21d9aa23c67555018ec420407ecb4d13a478e96;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h649b1f69d46710131c83757e2f7024a4b6c86e0a110116d55d180eeddd715870b1c1d032d1683ee37bc93d382643bbe366a6a06513b2f80744eca85d6;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h693f2905f13b59ee77826b2127b021987d5e16fe6e9fab1180cb48b9c2c0456378b176f2592b94af435715a335d8bf4918c129f617dc80f9e439c73ae;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc54b5a066923d1e51e5b838515cf88ca8c8c93d5886aaee616560279ffaf12bba6c5c99e77224db4de4b920c862d3de904d685b231885d61326fc24c8;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd346da235941eab5019f001cce19c6e65d9831d5188684c0dab4bcfc084e145874f1e8892fb91de139274e264ba0df6f12d0779c6453592e79cb91f87;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6233b0a74f817dca7eb0f9db2779aa4b9d2d2560809e58e0117e3b4341c0cf5fb40a2583e59ca988c1710ac74187406d2991096a9e935fff96910799d;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1cd6ec3d9c139ee946a0206840b621aeb23c947efa4e5b2a31c2fc789402aef50348a6aa833715f00f6d8d90524e50fd719e4104e725d9781006b96e3;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf05fc56d41b89bff5471af362645e0cc64e34bc92e4ef286c82a86f296539a8400cee27bb87fddab20399e76fc90b45e1fc1611f1a7f27203725b6324;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc3e44baacbc47cdf5b81fdb86be5e1ef5502344c68e334214dd8020e5128f3bc352394cf9b724e15adfe02e827b840569ba8520fd56c6629eeea84907;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc026e00afe24999053a19737c1078465ef6e656d1b74b4a030c1c46f2b0759e853b3cd176d3dfc3a5caed6d6e348a2b30618c65b0b73a39aecdd7269b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1eff148bd2678f5a9f0b7ec399e228ad74ecfa36e01ee83bf3da9fa0223e7691f80f8a1ca2d01e441aff9c118b495172d5679ddb65bd8d86760b6a0df;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h87b8f015c69b98fafdb5216a927c22a598c51617a888609bacef94c3eb278e474084ac5105771712ee8d7ee7d4491abbb349e0779bff60ad050dd6adf;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h92d4071a7ffd3357144fcc5a3acf8628675a37b7726ee572cb40a8fc242aee1cd306b5bacfea6e9be4c0a56ab10a6ccb473989e84e56f77d6cfc3c57f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h508db955d0ebeb42c69f2b57a050bcd6374e71d3634a877084116c21511fffb0867b88ff5e94489cc958f1eef55ccd1aa766363e170c71a68f322797d;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hcebdf9747f933bc83a1a3d5faa24b7a4be5ed739dd29f1d1f8f1b4690598344c14793f99e0dcdac44d998c84232b619a210c6c1ac3ce7ecb9d7e48ad4;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha8cf034c5cf348f6998abb821b759584fe1b79d09351e0564e2358a754148f3b7794e983bdc49b2b451d8d9de7697436a0c93e3ff7032f2a6d1ac4b24;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h98938b4abee15df04762eafe22391ced788f10750cbd9504dc16fd1574e5dc110a86b70943ae3de9a3353803fbc628fb92440741045e80de8a47ea801;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h49eae5a35be2c61d80ea276e11cba01db0d736cb96ad649cbfd77e1476eefdaaf3bc3189d44e5a1bb89f829edd799ce0f415eadf6ec6487516ba5ccb0;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc6ba5042f81edcf2c907f47fe66ebbaac0faa9dd384b298eb0cda98e3973d31bbf36eae0cbd026585de1d8e85760ffd2465c89b2d1cf33212a6791d60;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hcb10f3d8c3f8eda49def8269a9ab67469ccb63081b35d696cd992c7fd8ab017921a1f6780997d873fa80ea34eb7a8910f7704302e122fb7baf79ce5cc;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h21ec198d5a4f9742c274b0a6ac6c0a591b6b03ffcc58d6fc809c350f733d98b9d6cb58e81ee59ce2f65c5ba51462c69d8b4070cd1a7333d381b29800d;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h55cdfe331066617708b12fbe964096aab14de9b7c049e0119fcfd9ed451321d281503b20f045a369e40e7b7a2195cac0ecab410b998a6f0c4a563ec07;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8ee9ba0fcbb3ccfb64d8bd01ec89578775ba423e4d27132fa567a3adab6b5b51c93d6bf7f724d98c93a0814515a56349044b65b8f3ea09c25ac63b47a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4b0bd81bb79408e7df5b836dba7e2c134e931f0af3e737c8d0c66578e3bc5d29e691ce9700b5bc3cbfc00e61039538733ce246a7724a1176eba82ba01;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd5b121ad0da9713cc18c876d3e5f8b3c9355fff4eace32b16bb25330fc663457077ed0d31ade6df5b34987f1b2e40059105e841cf7d86b37b2561dcac;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc2e601c1d76a0f10e6acc08c7994aa52ac2eeaa6aba0d8adeb825a1468bd4d9813c80cd01df1c22121d537358a3c17e930e9faaeba1ec8a147a3a5b1d;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb7b7a5c559a702d33cb2f9f877f3cfa6d803f5edee8195c5532eb07082c07d6e682d195344b899af027c7e72a296751700e593d541f3f31df82425fd9;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h30f4cc6526835d15953572231038d0ad8de249e0b70aa5b6445ed01b1271b307a7b2683c6ea06cd145be16f2833f45a304fca5047712715153bf3ad8e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h294ba83d736d5e5881ef94c0cce929f73c12056767fc3541b49f3becd213b9e8c0d534eefee7f58ce4ff9d9521c5c0339c3f553030e82f2375fc0c207;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfdefe08a93d17ee509adb379e63cc3b30a089c1546b485730aa12822dafc69c5007a1ff0558fae919367fff1a6f5eda5aef3c334c088bb289a51a838c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc0427e4b7e1d44b90c34bf793c86b5f7150fd5dec794fd7b4f6031fb74306c85779ec38c86e082a3333d1e78b24fd29d71a864e9476dfbbf22fb898a5;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hefed2738df768f93cd2b43823745d244ed203b4834d6213274be6cd96677d78eb06a92c1103fdc143f89a06c587c776023cd752062fe9c28da61618d0;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfa3f9883bac20cdd74dc21fd69051ff4ecc081309a1c78360dd8edad7ec87355ce9c9001e07a5d73f800b595953f5e97a2ee86fa08348fe810bf1057d;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'habcfad1f555b5963cb0c2931d43e1b2a755a106381fb3ae293bef77caa2b18037c1a38b6a09797abce2e2f29a86b70d4bf44a3f1592d05e262c01ec67;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd9ea71441a3d00d0c9f0c2f0d292708c54fd7ebc61e2a929eb9bfe2967144c49728acc5d532c2a7e44d656532d80977baa6690f2dc67ddea3eeacdc0;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc0ed67e2a19722c164b1d52ab8247ff2a7ad88e372b0477bff868f8d95da31aef7a6eedd687ff979f4d0ac538fa2011d6cac35d682f2e369a541ec81d;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5134858a11c7b3408cd5c3f41f0de17b41e9eef29da48a8e60efa0cbce2b7fe5cf7da185e4383a36b0958df57e62796b88a2360cc566cac80e528c3a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha924facfea536adb9cc42151f762d209d4e7224179f91c59c319f0c0d093021dd0623fdd2f1c2a6e79f483a94e634ce85e763d34b9cc605afcc5aa074;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4817bb7c6739f6d8fb31ffd8cb5cfacbce7ed23e47eb53fe8ef45dcc4af38ebeb63bd957d1bb7935b355e72399f8cdd795fef3cf9e65b39f14957a2d7;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha6dd8bbd044bf2427b10721ef2deae2d4ad2dd40341733b0811926985c9fe037abe52ac93afa8c313ae7bf788c46c3a99b0e7491d5b51e374ea10c540;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h84d5388423a9963a08b55d1b98a32f08e521b838eaadd70585af8ee3b176425511a7276c71edea66e47dce44e8210828b8b58aa959fe0a84148da7407;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha9d2bfecbac5f94cac7cd4a80204253b99f57c67cf78fd8fe554d13e0aa04871ab61c7aa0dd62fd99155080c64d162da75c26f9c14ac64aaee0ab12b6;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h813e579245933d681851a4e29ad05dc370f3ff0bf53fbfb736b64e52a53a06dda79fd8729fd054ef26540024a385b643274516529e0d1cec4cadf6304;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2c39a67d3473ef8b9de6bf199e33413c7b913500da1f073318979303a1d47700207aa600a34f6392bd6127424589b0fc103fa50b32d67172cc13f0528;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc0766bb1aaceb77659d97303a92f3b066f4f5e08026257faa1254f91e1afb9661c6c6b659aaa120ad9f3f6f82d5fa5b3e5c31708ccafad314bdd4aa26;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc4401f46c8383e3d83925f91008af71e5d75538dbc9c8027fcafa9c5cb4036ee27191b1e117be2ae7215a55c836e388dc24c4ff93a4393b1d3b02eaa5;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h10c725281a5e1b58bb059ed4b218b885ffaa66dfc2d0e956cf083a60546fcb063a4f899c90c3b10b5abfebc8a5d45a44cd1e553dad65393adc42c2250;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd6683e59778fc7bdbe8c7fa303953040b557588b68a54da52dcff4be71dcfe08e822198567054b1438c21a2183da65290c8bdb3e2e5f99677b0c03806;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h131ca77c029c980f7caab25f071d25cfff50e8508ff9420646e217d3e1606783158d46da8688af0af375204610102d68a85c5374304e2372c6681c1ea;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf715ecccb2cb9ebf0833aa89febe2463e3f0314a8e5801fb5f30678b0a6b699c12c47f96077177f98384609256369fca468e1d59dac5dc5f1eabdd73e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3896633baa9c7d81d3a7856ceb4ff45cb166014ba55da4ec761e0b79dddfa4d037550dea47c3a9912f22faa191d768c8cb8e0ed97a5caf9ffe56ac1b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdef32907ce0b4af861969c5829951483fe493b2c792c65370aedd9c81d674144270b63ba6113ca91f41d2a5467accc6d6be362736c14e3813829682ac;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hed7afe4bacb91bea0c72d0e5b80cd44aad6b3b362c7769c89564937cff7334e74f664ac0951afa1ff241fbb88915caf1a955947b0a8bbf5cfda82eee0;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h52efae8c0fbd6b2b58ef3e6600ca2becab15bb02f739e99983357229119715317bf71b41212486c65a5a0028fd514f7e6624239088633d3f045879e6b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h437ef4f9ba1876e8f9572e3247a4d67290d58d60f3a8473eaaa44765bd25ae2d27a40a1b731e182c56d67c2492198b297f0106e802d6bccaaad243bec;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7601b36c7f31a71d24518b33698b1fa6fc11dd61db2d4856433962e465d6da0290f5602ee2f74a894f05da4e279660a642704a2a52c8ec22101f3bba6;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h65cd17024749a53ca61103b57221a035bc9280e68db131730bc06033d36e76defff9dc7423461a87d597b45cb7f5c4e5393281b298a4874cc05e9d56d;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdc09c6acd150036179419a9e04cfe658989789c705e016bbde9ebb51be841a5915ddda6810191f025d57b93335852a4a640cbb5c55dad9d50695fa41d;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb64f002d0b7d52e1dce4e661871d9debf819d6839bc13830b1f291e2d35b5c55db946c670f2c338e6503acdab23f34920f17f8f381cd7cb8385627de2;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9fba0c1e3d2b35c8d59fe53a9b142ab8c90aeae188882d1f6eb5923f664dafce8a265608e892a90925beed182f9480a481967f63c0163a442e5ed69bd;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2de56be6f3c71b90ab834104e4e3431246859baa3832fe35c0358914dec27c1e0bc77e5dff18813016663c9819c4c8e9e7a21159655152ac9f0119fc2;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h37a8cb74c6ac26f79dd2b62e99a4bc7f07b2a29f4455d9f082f102122d07fe9911609ded6feee096651af17abb6c50bf25d313b89c0d56722bb3ae86c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc42f90a88e49b6054cbea512bf7d66d006a3c340c3346e953705214fc591b12a2efb4df43d73e767649e520200db073a8e5394e857772d110b796c4e7;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hccc0514afe28451aa283aeeb7444738baaa8dad25819c7e0399fafc6a15082770907584ad7ec77d327f07026aa9be85bbbb3b76464f4116e0acb434be;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h58c26e438249a3a8ea0d541509059ad8a9e63f958c45917fdfd761888248d1ecb08152bd3cd57ce17b034b90284d519ed38a03a8d18e2346ee1cc062f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hca86d59408c09d08d7c242d92b56a891d68ec7b5714b81746b15c9a8ea303b0a8207db24bc930ac4f4de63d00b94b057ec596c5678d2daa1d7e60a6a5;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he12cd203a806dc365f7d0959fe5fcd45a5721674ff6f08160b12a56e428f3e213adf776962ac934119166aa517584baf46263cad318a4a550f68629bb;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h62a03a5c8793a106b1052337ab4399382647fbc389a39480a40f148cbbc1103b9e8c530ca3277229f4caf011568187068ebaa84df4912173b3f2846cc;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7fd5af88424beba0192ba6ef3e181cdabc3f918bced748cec4d91bf7014454d43176071438c6c7750409ce67f45349e75e44932cbb16ff771181a7b53;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5cd44c16b441e72ca5ec8e2967c71679c8196fe2b6220fcdbb3db69655375edb5da42076274b6af9e20e395d3a0a75af8531a70263de70804d6305bff;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2c8b928868368585c26464d692b24b49e06f1f0d36a68614578bf69706d516ded7764705b375f94ad94262666796af5bbff56faa39e93c7de99158283;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h16b692c7c59369dbc57b1ff1089decf371f70c98253736e028364f44cdc4e3f39d674486da91f912202f78a7fe9a2b7088d17e69a78ed4571001f65fe;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd61793ee5f360ce93962bff5e3e83642892be24c7b6f88cfdc3131065f691165b71a3ecf6b7cbc390d8506fda02ad393b80d37f34dfc8711ac03b3e1c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4e83f003de63208e5135618cb533db739983712fbeed0d0b24b0bd8680f3b05f6a99979bf5aab15b9668aa937f707e3884f6dd04b05e167c81831785d;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h14cc5636bdb210897a4f593b1042b719a192cc8e40c20c7574d6e162183ef44a4badf6de5e95385254f19e5a4bcb6bf79969fa4efd618ada989fa2094;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he718f0afa8aec7debcd22718b72068f7d0c32cdc6e9a1f3ca850ae8f341563ec9510d265f107b12d8aa99a2b2d0579e14dd992cc4a13d5efc2710f6a9;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h29845bb9c50a302e1d1be6870512b9348e12593e8a6d86f31cb877774e9fbb22d0ab73ed8fbad27d12b79af38dfe13e73639eb75dec14eec25fbfb0cb;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2079528712e2db605c96970db02bae26ef610375fcbe0235a0ccdd9717643ef60b6147a29da08337ee28bad15c35b88c3907c5ededcce89d1012a9123;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd090567a47b46bcd573fa1aa8c0ed8fe2b4ec5f0611b7100edecf3078e76f2e3e40bc21105fa2d6c4db9a98fdb883cadbf819430ca332d0d64f1562cf;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h462bf01caf7aa5e81a2b32374a43cb6a9c01179426985c5cd13d75435556a4b972e894c9e8c19b414a177705a2fa6dcbafded27fdc3f78a26e7535fc0;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h377554d5302699cca07518b68afbd43cffd0dd87fe0f175364ed42a36d00858e8c1667aeb787b9b4a2b1d57801a836aeeb22f3c6a55aebccc52a3d13a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4f601cbdf301bb7c108e5b91b54acae6012b076a341bc85e3653f843d5060dd6a7beaa993e83c6db331e2a72d25b3894d3430d98f90773fb432211300;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'habff3968bbaa8381e95e75336896709f9d214676141557456d13d052fae628f7fb334dcc25735638c6270b5484ee8c87e04d8e99dc9e9104b9a0ed697;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5e35962ff18693dbf9e360519da7773ec521393e069bda03c1b60cf6a0ed571974033c369860edb726fdd034e601ad6fdeac478c747ec2b7dc80e566f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he628027d407ad048bd8b94346bf10d3a269687f0b8bd1a597213c41285bc705697b8709c797840268c41f8270364c4ebc2e04eb4e33d4b0f5a9b770dc;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h98da0403020692c1c9438366a4605cdbf4f2eb2bc441799b12288ae43ac5e5026d8fc2fef4819757f5d23c55d2cb240fcc5bacba90a1ef7ed9fb86345;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h205557cbbb6eab42f7bfdf4ce1e3d410e1f0c248ec1a1e60367380bc21a512ae71d255f020850adb8d6f2c6cf4a6b797c1ace7653f498dd815e0157bf;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h23d95b9795a8a968ac83ca8d1743e7f8dce91992c5277e3bd84dad14fdd3ddcdd740bc54e3877f1a63144ba8211d684739ef22524abdbe72746ed31d3;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2010942482315c807c429980127b90c7229844638ef4e2da2c40be65baae51b27ffd84d05250a34d9f24056539ecca0bf069ed4b8e40d64dcbc46c45a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h97183f4ece670da90065c7fe8cf8980a327d7dafed8a77d2e2156ef47c6d6578b324d9de272e1407b9543b2551544dd6d0bc3a9e38ad25ab114c59094;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd0822da58234e34764338057360aa68322cc2f7db5abec7bdc4029bce604dc287380821d86ee91ab8e55da54f59eb4aee7c58c0f290ccd1df8a680d0d;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hcde8d084e780f8c51a1fc75d0cec4cb68934c872ca8e80e23f8746c09435b54d0d3688e67230ee872ccd0f198a22e56b185d211868bd4a1824bc725fb;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1a9b9f2cd6ade229e15373c60ae383a13d923a5cbe484a1bd0454e3eae2722bdc9a17dd2c98f451d05e819885e896dbb2991c9464fbedcbea71c05d5;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h184fd3a4c8d7dc6dfe697d0798beddd97d698dfa1572afa2226cc32350036f06d1cf3b69a502d6741cc5fae0ab2d57a9b0c4355893e7dcdf6c3e1dc2;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5bf91aa6c5c6ba3756c6d9594167d4b6a73ccfe61401bde31eb5cc5e9ee2cba78ba8bf6f16570833ee28d56c1aeef882def4ba2dc45df2092937bdcbb;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5f180a3928ab12867820f6abfd5e8b085884bfc14309e0f993a156eae20b5ee9cedff05763ab830d2097053f4e3224baf9385ae7a51d7c0fd53355dc4;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8a73e2f3b26cace045bfd26f5915511605a460df3ab703f39aea61babd00d5590b49fc944ea87beeac54df310239e2dce408ddb9e72ba0cebc8420504;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9ba0de9fb701846b31f0d9d852df46b31057995ec6c26bff120f64acc2750a04b6018f63121890a8db8b6220bd953d80239df1ee68ba85895d804fefd;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'heeb5a6d2731fb0bc7960091a314c421418a1300cbba3ca9b01379cc5368c90efd8ab338a063200205801ed59783326b04266979fa22eb8b9dc85d500a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfc9fe655a699393628223d31c1e7c59365f2741aa3d49cdc60f52026fb82394a9ea637fc37a89243f794375e1fdefcc15cc156f45ef4f8f4d41606ed2;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6e0ea1bff5ad3e05b4a5e76b427babb74ab8c05061de397112a6bb0923b96e83a69c375c3a9b352df811ebe0f62cfd363d6d28d058d427fd81eab2348;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h646774e6d255d9ff733e531dd676e6c02bab287c6443f4ce7c89a3a85ed1b959401803d0c522f010b83da4f3afbc33036454769191b3aaf40feb09808;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd817303141060ff97dc7572a65ec47b50914e0175ad98b8a196b78e025bc0117c4519c7e0c755d1311c548c6a1c6d0989e44c84dc2b37d82a2a6e14ba;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2f72bff0e6da1182902f07ef4bfba8fab13341fa8f0a894f55a11af1a146b544fd00c379921dddaf5f84217eb6569a0949a531e80e63651128ff0ce89;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5d8d0c56835c4941aeb2e73b1db35e1abfdf40dd39118bec6ea95e28571e82daf62b1eb201d3964d63887429280ebd2a4b1a16c1a279c7775c7e74979;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3f496dae6d159c5cd77b810bc14a156f8d203a8db11953975302d74b1a07bd9cdfc88027a17a47faa518cb247227b6e6cd0a8b4c2e39f4a5a99889373;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4bc9cfa7caac4b9c292a1423888eb069b75cc44de1e07f0ee643dd0f7ad88203716268f8022ea39f94f895ebfeac6b3fa87d72de8c957677a38e4c3e5;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2347af19a08fbf5d81b14c1f90334b533e45db13161af4f5cd0ba39cb9a7d078bc0e03e199d1a8bf639b335b6ad327067aa512255ae3a16647dd7eb2e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4df78192f5897923d8669665c90779ee2b2a4d6c69163a0a438e701822565dbcd1e99e5afecb00bedfc7334e82e1451666a16a7190728d1abc8bfd361;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h68ebf2ce8b21c2cf81d9b5eb3f7e4706d8173e009791bd78cb4b19b1a45a1208deacb35da326ee4050854bec045892e1af51ac4e3c61976f5e5397d1a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h71813a160763813817ffaf3144141bfa09fa33137bcaaf1f8326fee322426951f31e7542aae86d48e764011757837d992c2a35ff797604c5b6e82000e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd9cccfec1525c5e55db33d6ecc6e13b3a6eb4d13ca0505299124efd9ba4f58b5e08843c0fc458a17ced9844ebb5c281f79937e3181c3507adbf1da22a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf4e293795f3bc0a361a7b48f0f13af0f6e9b455cdd06d3bcb0a3dd4275be464c581865839c1f7ddac7124b2b6db0760b686b28a48be173c642ad8ba41;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h156744c0c2aa3bd880429f7dd63c1b56e62aeed32a5417c56ff5e4a98e3bc508a686abf075ae5e5f0722492297aed167edad5c805a3cba2ab8b11caa3;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1b0f38c3b1788b8212f7e2c4edc567bdd5688cebb25f7e58297826ac3bc11843b4069e6c6c15ea7bf4a3770360b1236a09a0cf1527ed9e6d7119dd25c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc5d20eb8d16eda527640c3aca0bb21d3cce3c2908024fc01a35def220d2379f9cb3e7d77c9897187f036a96327f4164402b2da8a87706657c64df471;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7e6c425438af639a357d61e624f60b049bd2a01aeaebc0ed4c7cd08b6f4064b9051a5c871e772ec87bcf647f8be13e9a29e987a757fd247a8551d92cf;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hcd7a75b183483b3422775ee0bd47136856808db6709deabf321276b8a611995efcb28f5f1d106b33e9b617ff2b9902ab0990c27d3d068dc7267b4c457;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he6c3e977f0019115ab0cba69533c64e8652d231fa4b70a5e4afb69dd7e0e82b4f2b66a4339b2684ed0004f7cca17918f19fbcd1f38013fb512eba6543;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he02c861d92e12d210bc4d35524e9050f2315d4b25f340b81455173bbed48aa90c26c1bb0b53a94c66577dd142dfe34b6e8e8bad0295dd1c064aed3637;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h15415031bcf24e79fe7a603e316b20907877708b8cd8911bc4485c402a71c0a718dae930707010e5aad8916cae705c2b1e7ab1c907ffa9bf79b90f6e1;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2fe277a554b95a19f6f9197a6f456b363112759ecc7fa38fe072886652cec07015cf008dc9c472b5a1a840c6d07523dae08e9ebd74e4c788a77f19f33;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6092d60ffde6937ca926b2796e03a8d2616097818a736f3e4fd9822a47b27c3e28754a67ab9214dda430b918607664573b5f61ef8a53d469b3ff23af8;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha29779499de201fdd3b02c8eb263ce7588b9aef9294812044aacf291cb7c69cecdd48129d44c4de1d1dea60af9cc4331668a50f288ac12a048cff94d1;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb970467cf7f36578a85cf351afa56c10f8148cef8cf894d70b03b24238a33a3e9acb0512433583f2f348dcdbe83ca2cf6d45c89c462c6ab71d5cfcb10;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7801a862584848adab99b9655bda39c88ddee2cf0615dc3702243085e2b45afc6f6a63baaef02b340998211a5c6e5e896fa3fe09ea37e800e4e3ab37;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3a44c914d3b9dab5d5affc4c8d2f665e386cca97fee57e1cb5843cb9e274fc836a89722eebb77679f776d88dd3e15d9af456fde853b5b8d81dc5bd6f9;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfd181138a07d96ca453508ef771fc774122e358076051ba76bb4c8fb10f924b9f6a3d06113ed926dbeecda4747f40576d94ee5dbefc033636a8b0c623;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9b851fe0bada37cbe4977bbd3e7e36525df8aee1c32b44b5a507baced31aa649ceb4adaeff9a552f7ff2fb10b09caadf68b76e948018fcafcc2c4b351;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfe37f2e7ddce43d7d20ee43a1ac8079637ff734ea685150955d5a170db8f18349bb73accc817e9ac0a26aa172fe7fb58878467046403bf31a6348619d;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9fc981fd0a9e6b5c3b6036c7112b596f311a0869baf81e1c28cc5a08bb36b2099422961c1b8cfdee5bf3a229130a53208bc24190fbafe4ea64f4e04d2;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h88d440e406c06ccaf71469722ba9f879621b4f661fabdecdce7c226a931ed8c4c89fe1ec6051412b15b5707949bd64d5757b6ad98ec1fb5b4d3ce56a7;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h51c3c85585e2c293e2828ff8ddae63c4ce4d0015916465010b8cbfffcb85b65ccd3e706b1d86ba7d96426f32b6e6e97643059127b6bc905ecf2554d5a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7fe392d13993cacf1d38e22864615218f6a24ede2dd930066ea3cb7ea504e59c212f99fc19b03c9c22b6c990e9e3070fb652f9276388dacf6d8e1744f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha2af87febac86477419cc8669b7e0c0d5b5aec9a04c96bc8cf05c741145d87c67b9b5be7ac819fc23a7d327d93efd4cfed1d91a1131a8f8abfbfd1d59;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h99908dfa8d21adeccc1ade5195da5745059549dec72674b8281e84f998eeca0a0a36d1fa62ead39102d362ab20b197cdf05203a443f6c0bc684f08a4e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h64d3c4799fde7074ed9a80798bb0561086aba34d3f5fe1f6db0bf3b08b5a3f9c85e9d52681966491277519d0683b8a3b12cbc78c769bfa4208851a38b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'haf5952b31fbfcae7030f86000ef0924aef385b1b9927d8cedb7c5d0ac42635c96370eea507b35f687230585d337d3dd39437d61bff75a11d4d773db00;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h455d535a4053a91f6b5dbe5fae04d5a566c94baa7208a1ae6acc92ae0b64ecf88c9c7dc37be770a16c8ce2995f3ba56963d10b25c926c455e65f4f8e7;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h48211edfc0824ca57d1cb58f89aae0c7e8faa085323a301b7a18bbb41b25fc804aec10c82c595bb7e0a0764f07d7f06c777c9b44d22148753dee24db8;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha414e8bbaa8f452387b715b3027f3a2febd875c981e2db19e3db018a8cfbb5e36fd6708d4f7755c1422c51f759f59006bbb8d01440a699e0a0008bb98;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc2f4a0dfa47e1df534f88f0b3efd23be0dd362036a64a7fb25ea46da2db89da9ff4b79a071ae61216e7d9c4ee9b10a10e08ee21e9cdd7cf2c6782bfbf;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdccba0bb1dc5f0562865882b069fa3767c198f4039082c77dc5e0600bb536de54eb70d69ca26188a7a9e87670a80320ea0e7561d1526e9189e0a2ee80;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha98517a96fdc70f0f246043a602dddb1f05448b1168351068c75066502900e817a0fe270196ad3e5f767f9590ed411a65023a268ed919102f32cff9c7;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc1935c8d71182a8debe1089e74cf733121ccd1e09f0d886517da0a22f6229485368c4cbaeb76a0369185f7f90bec13e517f0a883ce215d3b8e311467f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc323023aba239792ac4dc74c4d133652463023a0afd5cadcc44a50da097d29ea8ce796172e6df5ffee0dc18f677a67a5c095877a8cb3380ac3afbb46e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb72937852d243e7e0f12090d6fe539e7ebf32cdf434f461f1f1fdbdb776670c869572f1773e6281b169d59c3cab6f04e651af0105d7db4f69ae71ecb4;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h54765425e83bd83cae724ae302cf409071082bc809f78fb43ee085a897a130f3536826d4500cd1f923f020da97185c99dc67e00dd41f2ab9e8f4b37d8;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h915534c11636f6867b1452935e02ed77118b042bb88d786bf2b519917b8c9a3b19f3feb0cb31a53206364b9d91e4712e6cb39266123049683b280a408;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h66016d97dd0713f2280f33c80b9f40f2a882d089cc8b09f82a93f3b9d5689de8568406f33851c60b56003072304b19e22ea30d39e7bec54647903dfdb;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h392607a0321f4de9c80fc805033d8bd84bbcc8b313993c78e7b8a1482a21f2977434a7f9bc0faf6ada3de78e79ad3000b337a6c9fa016d0a6d0ead644;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h889edb1d3614e775cdf6cac91d310df4581053ea8ebc29745770459d7b8df948a3a23c882ec3adc1141e2d640e7eb66f571f2a777d00705581f7e97dc;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6919bfeefeb9ed198558fa047f8274db20d1f06d0ca7084043871add0b5666a71c696feef2f6a8617b75a4ebc7a48d49a29e9bae768941b7b9e4abc27;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd534dceb0ba47c194fdffa6c6b35a5051f89c3e554d7b50cd52f00cce4927f2316c94756bb3500474f8861f8edbf67b4d7542de80ee19d596aa0db3fb;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc5dcac150eceb1530c32ed3a43e9d8c015c9d41c13aa02538919c43aefb7c32217abc6b3694074461ac08ca35449a2bfbccd17a1302a4478c349b350e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc8317707416a11a89b32d2748d4cab80949e2bb1183f4eb571a68198b0eeaaf76fe0607a68f2f009542da0ae7dd78dbb47140fd9896a1ed2edb20f980;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'habc5e8c82ae12ade5e4bb14d57ec88355014db331d0ab47da4f96ee1c5ccaf6a8c99cd71cac2088330f5424a860ed1055a9114e2b24f4875d4de9f2a6;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hcdba336de71052469e09d83c04ec4aee55bc9a1729047855f1fa011ece96e42fb110bfe8cfee8f246b7608ea84ec2f7dba9e1742d47212b4496e51249;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hde83ce1b4297ee765c7583864ed87e79a9decf72241e5dabed9b3ffde5d82a1f30ff71ae0fcd5cc3c731a9e2774f8f849f6f3ace14acdfaa1b9822b4f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2754bf618a0c1773adcfacbbd811fceee25d407e4b10e43cea0b4c4c0d2892aa023e0a55789df470cc59fe5f4c4c706cef569393999d6eb383c3ee7c4;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h21bec287c69c54a9b06561aefe8458c2dee094c18c18423d7fdff727049e83bb64d2c6f0583c299a5059086d588f2f8f25c5502d2bdab552bf5f55e50;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha9b408df28a60844ef44586ea8907044e72d1682f71e31cbfd69cbd9fd122bc9ea79ee365c7945a4551e1aff5f7ba26d03d70cfefdc2d6ce0ee141ba5;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9011dc6b28aa54733c73cf57eab3afcdc5cf9df5995574fd97152087577970ac67a9b74648970a51f321d8de8fa23aa8ff63e1403feaec120b672c5c3;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h520d78169677b7003e1ed76a076dfdb12b2958446abdb720cd5ca0ed70770bf69b529025ffd52fa14f42cd1598f37aeb139bbb7d96f62e34df89ec437;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc4af8421a897877edc7152cca4529c182c807fa660c30d9203d9ddbb7e64ef7010c6ee0034e9e21513d739b258d94c2f4ee3d063d22177ddc5741feb8;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf4fdd0a8b2edad35b5e6237148017ad62e3b5aef1872544364cc5abe0203097f7951427405f9d0e440100297fe469f7d3657948d13faed98d84fe76ce;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hca495847a12301718d1f385647a5c699d6520160c34d7d435a95d68e42ab9a72cced86aed885b4b0d9a9ed52cc95eca7bc23c566f103a684e2edcb6f6;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2a367cbc5d79f452578a4653fc73176514388fe54bd0e76400ba2ff578a78ad407b8921b38d74b7482c394527f5e700db7f6e66f09df5bbb9084f2e19;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h11fe8417fe6224b9d897e8ed0c754754b4eb6bdb3c0bbe061d384925b91c3e3e85a10fa06d24da776150129ec2629077aa6417d37ddfacacedcdfdf52;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hcde97301b24bf855d48ab44939488ff1c4d872d37f7f5ff14c37e25b0ddc79b24d3783e167881178bd38fd78945192c75d19d80503db2526b4ef435b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h98f722c9f9f35a6c0b947238d1eac0250658d75301947cb1589010aeaa7b2a819a45f9ad9a327e8da16c997600ceafadec906ae0f2a4c305086dbacf1;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h67596530ae5327c5fe59545884c70b73aa1d7235781f2aa94faf0ea73e6e139d3ef1722ef9cf16ee09b1ce0ca166dfeab79699b7b58fd03d15e9b6c54;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hacc4d481f3e1f6634b4a4c4aba78620e50d9af48c59ac3ed4911eb89edec29154ebc37ee93ed7c5bccbc10f7d69a84860bba35d85a7d46adbb860b16b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he8bce9748479cbbc5aa9901972f7b173fdca0627c3525127d23a6fcc5a7228ec59b1c9758c4a8c42c4e4113722656ab446600a3b199b1459c3556171f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h64c1ff4b67db2483c7a9da7a7f6e41d0db36fc08d94aa164dbe9002a5310b10738a5f4104327bf32d9406a988e195d21d74e3997a497f4ec8747495c7;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha648948382e7c744113da3b15954f74befd8be2765e370696fa7cb6f798572d62b200f34eac9c022e481d8df70839e61e6c8229f7b25a861a6427363;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd79d1499860d1faa12d76d311fe03f58fb4e509e9a4907f181c2cf4ef8d0bf56936f8cee7168873712c5ff42097ba171f76d99b825d6e9396f54a2512;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbb9f40252b91211b2b673b70126bf538c1fb3ba4b13df4208ac5b722686ef72f42f3a833244e8ad308d1536fbc8b1fac0d36c9ea9b3cbc529f2ede68b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h57bfb0d6ec169705bf184c4a510bbefdc45585239bb0a4f5f6d7d4d8f6243ec48b99d24fe258bfbbb002c5690bfb2dd8e034d9f228e672e2daa18e37e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h594162892729e1ee37a6c0fc0d8d63a5e8412de6d48fc47a24e87670693134c68469f17bb98f931d5793f86c255afe246ef49dcc97767cc77b010a159;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h30fea38d5a55fe200ee63bac5c82d63945ac6141805c0871d6fbc187ffd4870d0022292dabad0f531bd5f6c42f8e0294926f6986e1233004d7d14d8c4;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h27beed97f0f5e8ab80ce4b0eff00e2402ca035787ebf0bff45fa3b1679097ff849accf6c32a941027fcf8c3e349fdf6883e7526223bd9cfa7e0aa3f76;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h211151370559d36f15874426d57c35d9068b73cdaf55f43e4d22a1ebc74b69fc97e5deaac78a75aba18fdc5d9f6909d9b9e3f0505735e1e26a49bb79e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4903cff448318776dca2b0fb9454ae06cb975fe259d87cd0a251dde53bec55b0d429b91d3155c3e727aa57ea99a55c14c655da0924135c2288901a96b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hce0314c7572fe6a77b26322b00ce5546e0cf58cd60a0043a48c7ebfc0325222300ebb4a4171414b7e674fef352c82868ece13088db47edef499a592c2;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h637ff7c0247c248bef0c48a933f8ee1f596ec5a8f2b0397bd48575b5953f3483fb6ba2bcd3a043be282265d89d98402b8589e1fcc5cf23329c761134f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3fdcb750bb7dca52eb7943a1dced5acc5e0a705282616eaed81994e39fceb32e917607d4bae33db018fc0b4c31f59c71068d29d2929b9427035e6ec7c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h21af2b85adb6b4a80f9db8eca865959cdb1afd9ef913f7969f16a39bf8df8662e64c2881a9fa42f323fc2b156dcf1d93ce9732c9832099cf9f38e04ed;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8105b2775a3008c884ae8b8b2558d9094d69ff6e7e6a8a4faee608caa43287feccf4d02cd70e0ac060c3cc86471031dd36f18be95a92ed8f5ca92eed7;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2366c3ad3801fb1d8f475ba357b36ff1b8cdca5276ad99c3c6aadc63d9b0239998b1e0490fee8564c688eeb550ac7b9cac3c04379a05aa659f0daf9d9;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h980391c2f5a192ad537b57baf768902f9cfe71a81d68c9509ae8184ea7c1537b9c5057c096bae7150a48637fd6d1d41b46d25538c642173a65d63c879;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha56873825c123fc4f0deac800e0deff267f10ba5a4251ebacb1223abd61c96ce9b9989f87d0eba4c092747c9ad07b55dab4e3ab3f1254e7e992adb392;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2a3b79e915d91c0fbcd60b24b1a27a0d8bd7ea75ddfed0d3247be8a943c7b78b5b4ef359ae5d0c71793a73272ff86ecf26a00496959b0a7983ca8cb99;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h733ef0056f59acdc621dadbeec2b9f03a8d58873bb748df7ed77ed2f1718fee8d8b5aa97eae917a4e0bd2647a708d2f0a5b0f41c1cec5b7f49387246b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h443c677fa3dbd94c677e5fbe4d15f649086842e9830c37703736986746de51e03b5886a27f2d1ab478b5a3782df874a71a74ae59ea9795924b15ef545;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6ba1c98f39e3b5f9b2d767ef451f3b5df1c197652ec9106e56ea35fd1613533806266c771d80f74e81a69c14e0cad7c296449b0656e469aa8a1e32131;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he251496a6b12352b192ac3e96603e619d812e0a414daae46449d60daad6d9fd734a8973e46ba1dce508e77482a8efc60e0daa4297480e14b35254dcc0;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hde99098eaee18ad8b6f75c1e7a893dfa001b2c8c71c263853b2b20fcf8e31b6594b26de36e3a928b029fb4f8b679a16ac58ca43a8816ced9e823aa8b8;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3c3f52b36a4fdf208763a2c23cc05276e5744bc1119df81e396c1b2415e5f5aa357832de87b31655bbedea91d5cce11731787aaacba8a1848b0f1d4d8;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5e865af26b15ac5a2d624cf39bc6975cf59e24e46dd2d57f483bc3b2f18d14bba429a9e6598873363613996fffe5866f51c8278084bc8dd9272b258f8;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hef1e2e66549c453d261ab588cdb99014edc92bb2bc1079d33e731c8d917d13786bea6ee0a095b4599a88b1c23e4fd9bbf12a94b18f056adcb87f3b510;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5d0fdd21209223283052d6e35329773640479c911fc762049b98a23afb6bd02236f2999a9e2bf4ab325c31e6a9bfd71e965f5e74eccb75afb53eadc5c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hce52a2a705b8120e2b952d8d08d3d4a69cdc1d908a5f0b9a2c642950984ccdd80f4e2e979baca411c7cddfd160fde2fe452d87e319f8fb00646f03911;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5a640b4c2937769a221581ceb6a039b66ab4fa8f26c421e8d0e8a9778387b6724da5b752bf4b863cc0702db231257bf4a27868628c135bc72e6627686;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfac5e0267fe309c7109ee79c1f92435fbb44dbe2ee5825f5d3ed277b588ba1a51138671a3e7ccb91dabd76122ab41c449c173b4a368b2a2d52f361d43;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3899025cd703f57953d9b3a76ae68566e45595cf343fab8b45518b1e86c200b4dcd7225e22f5e506580d2f79f7d7dd0590d19ef783b80deb001569fb4;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd716c45bdf90ecaa76af31140f717eb898ebcab8427b36be54dd5ca16cd8e8d9907818476981df676b1091c7d4801e213276ad6c551066e9d4d8d6232;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hded41d944a846f100d21a8f26e714716d2870dcb23c6f81b020bf89d005c60e2673472e1c538efe63d597e156cbfe459990aff88123779abe47a1b827;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc14d3a89f58a5850fa28e1a317903fdc8bd354727a26eeb880fad4aa5cb8c3db7cddb0078761f9e9ccfa420fec66001d0e3dcaf304d77a4dd819d38e2;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5a58b1df27d66df2176c12b508b058c8e037b544b71da02e8eafcbe412aa770e09f60c2355b29159ec501cbc9ee89a7cfe8f32a9cbf56c5a158086b09;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'haa5b2d87c7a783e4eded643205042b579f4fdc1deefcb29bbf9ff6bc0d82c0c68100d22c49cb2f1625a1d69f5a32498816cbec825256af13378c9f9e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5cf0f87844804673910698fd9e7d0331449f7f1025710ed5660069edcc9c6f51f6dd032683bb8aa0c39a97dc1930eaebf9ce65a25ef7b26f7bc5f9ed0;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h841e976131e537a3aa6d28a3e698cfbfbe2108d21fafd2ea1c273e28acfbec9dae671db3d77bf41f32b5ffbf6fb332b5e487e4c8670b58643ed36024f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h76f2fa961632d552eab06036164d4b2895995f34f6c506aebe66837bc30deed6577dd98b414df5dd4b92c476f074c59ab82a90aea0e92dbbf0d6d954e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h25e5fadf138672bbb56c648b7b1c9000509b2d29743ed82563ec0ffebf19474c582a268656f48dc308667f283de7c13f640cb590aba78629f4ad7c237;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2678230e9d8685d948d86a78fbbee4622cab71f42d33a80591dc4130e34493a37cb1fb804c420e291c125750688ac90adaaf8553c59fc429a8fe80a72;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h663845bb370add141def72bb44e9269d48e3b7237f6fa4b40a38955ac3a1ef1513b551971ec98af457a8208f6d9054f838ca8d4c8f17d303290f2d7a7;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9e042cab49c5113f8927603b8d38f4f5b58bbec5fc9d3ad3911339bcc6a899b3ae5e16c7e9d0d72fb0c9398a968f2a46d7b3b7dd08061ec509759aab4;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbe4755a482da03241c069c02daf50927fc8a8cfad53182d54bd04d1096158e91237637162d99567c100b1a10b65e5b2fae3eda2164e55aa4cf9b8dc70;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7fa6b997b3149fceadd75bcc2405b9842cbece094c0a73bb4e81a1bf5396d7c3f61037f4b78af1ad2afac3a9b9e70c7ce88c42d8995c111e86c222268;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h559b07e4a1d7260094d00cd53b78b2d27c593040043ce34662115378861a5ab18a0c714b954d3744fdfdfc12cc4dfa722b6652a817e31dc980230f68a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc29efb71c6e8c644b4eb3c722609c5107f88fa6c0ce2bff57df1c123ff47fcf189d737182c9afb040b80a5f3be8579ee4b7029e63315c691e5e739481;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd585f74fcfa5aa5f9da1465654e893d71e910e457d13593125c5f94500b2d7f4fdceaff78a187478627a6d1f885f107a29a1c3f69e9e54091fb769490;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h69152de17fcaa33336cd41bdde044e543be594d3cd9437f1d1528d73b7335b244a4f295ac4b02ec8d1c36618d51be0c5dc355978921ee544a297e62c7;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb0e6ae537f2f84ac825c7a6acf58a2814c508507e1601f9d9b52074a85f3213fada4e848f6f6335a21b4dd2d69cbf4233b3b8ce5cac41b7445981d364;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he0a2011d9606505b0bd6feb2e4af35a12d7ea38bfb17c228db7d0fd8ba3ead0abcc8cbb9fe1d2da6129eb342988d2351a082979ce9b3704e84914a1bb;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9939d318a4ecd72570ca2e9efb4a979babcf7035c2d49a0af57f336aa2350362275b98845f6755b8cf47323f183ffa2847b6f2fd8c302d93b4187b5c2;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'heca7086521d8809b1bfed312b6706f68bfdef5f590971f48450bcdffcfa3733c8854a398798ea09609ee83175fb7cacee0a5e7c95a49a1a6f0a465fcf;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6ffccf34bc89c302eb7f750b4d103600e5a1ec00ba3e965164701b6967bb91c804b128c99125f6393bb9c83b4273f09e06d3bd31a6a967e73295c667b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc4bf264d0c4f97ded938c7ad746652415f87fab1793b5f0d4c0178c8e5742bded045eda9fd49f03b0812d9c5d332b30ad399711b1ded63d448dc423dd;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb461bb4694533f99e5e82460c5e435bc5927c64dbfeb4de3b6f15688b6a7f489ff91fb06c0812d368c8e6c0b398dffbd0b234037e07f369c9fe0c5bc1;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9f23e05efb56b50883f819d3333f9fbbcd6260c96821e38bd064af5465813b1fdda527a4298d152ed557bd3d2ce6009d00fa265dc13368549b028b886;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hed3e6f441ab0bdd518f92ec0bf519b55c676f9d23a2c2aaa309594fdac7ae511c255901c545dfdf9888047f3737d619cbecb4010028b36d117a5710a2;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hcd19b5bfed57c17f781890e9c36c3f0b420523a366fbdc3f13f1ecd244fe01e2bb439c9b5993fdabefa5d9794ecf043341ee509abe354c9200e6e58c0;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h610233604903418b583fd205711a8f39da6ca2d521cf1c2deb86a8c50d93074a5716a1e7f17b35ebe0f5c5098b9710256952275f3697847bb0c88bfc0;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h113b3f51777c78a158b4d1d819a019e77c2281c262bdb05e0b56826d2a26ef1ae2fae95122dc51518a291dd9d86c11a285bb97e6c0d5f66909b875e6e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfe1ac6142079ea87bbb52a6dbf9c9c2d1bc1ce5279d47b7b75b11ce02e43c9543ddd85ae6ac56829edbd4d90ec7c6edfe6ed3d52422311da9a385a2d3;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h489b4bec65bf3bb0b2c8f5f1c18b7e3e51110dccb2dc6ef2ea3d11babf49cdadf2f5ab8433f2c5b48f24b921a822ff838cdb82c5d4ae62ecb97e0c3d9;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc879595a4c1a2416355af737d77f82669bd85d68ad6650cef97176225b6e3a5f0178a4167398793849e91998d9c2cc11376c781bb8e04189e00df8984;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h698473d8a7e27bdceb48566c0f44cc175a54112a697275663f17c7a0eefa777bd5b9ef56b8b876fd01885f654cccdab32500b1305f651fcb50ea3830e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb2ac35155ea3f026d00ccf8b155d0b213ec71c9091b8743d2fba99aeaa7a82e217907fe2a408c2a54d97ab712026447dabc11ca74ce1c418898eecc10;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9e2d676a070bd87dac43800e1fa8487466a60e3d6a67bb4b404f350d1ceb1e6c8c9ec86c6b81c04d2f5594778313892c54deee59040265bf21d4df759;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc9332bf6a7a39601f246261c0289deba68c3ac2b0684f6581b6a78e36be2a7158a7206fb3417199be463f1fc7c52b64f52b58e8a1f48685dfbd88a87a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hab39a6fb301a2ea86a36cc515edf9d1d7ddc2d66e60bfb1aa6465762d3dfbb457c0b57a8debcbdd923b2d02c5d49563917148e6ca8000bf7408713dcc;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h94adf34d44e529ade28fa9cce62297eeaf76b2f95e25309a127fba9364d4cc762d051ba25222562f899152ba5770949803b72df032dc86d33383ebac0;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he4bb78f04e386c928132a9f4e4e2a85c55b917ccf1748e784c42e4ada0d0ba1b236f24935b1f458d18c3971c2dabdbe159561933b2fca1ee41d93e3d2;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7881af7bb0e714abeec5de1cef696e621ba01fdf1b001cba9162a39c3d639b161b21953ef175e3e6f4737244e54945eb1feb87186059ccf3e4a56d7b2;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8f56b3419b3859c207278afddc103e28e719e1610a7262e2e61079572195e1e0506f5e5f52d7ee38d8be1d26fb410f467963e9a7e54763f2cb54b104a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3890fc53065af91c7171697232046d1bf5a42e37c42e416f72656e46a58b38919c73957cb9918901b5ab7ee6157ba95bb94623529be8b91fd309a9893;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2d661488e9b39d9c1f475020a654d496fe6dae176db2254bc94b10a3b8ea947fb84b86be76bdb3d272d3a0685b0fd56dc0dff9394194c9f18527a4460;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb0541930bfead5472831b649191c85fc76a49a573ad29548cd353ac90e21754d0a51df320aa17bdecf4c1909dfb6a1cb44fe334ec67eccb721e979084;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h20721486f7e03e3d369a470018daeb9e8d00fee906c73e24e2b7bf6c6a6c658ee2f9ce40b101d9689ad60992f107f0b553cfde18d65f04e1b04391877;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9559fd91dc624136850575de445968802b7039afd8652e84007539b9af3e9e24f48784473913e682ceed1596e8052b10a86135c69341afd1686f9a1cc;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h53113829a1fd89dd74ae6475926c9221f26c446fe091efae1738ab66a4c2d21136809a3366226e39f125d8af16040739255939b37e4bc657cfe7e2fb5;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfcc3210f2ba622e25d687eb5c00919692a2eb13d784679aa8cd603426156849685c0a0ebf2bf8ba4bb30ad5ea379da9c8f6c8f7fe2991a476888d3ad0;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8471af3b1760e8ff2700229bbe4c91c5531df321edd28e9729d4655f2baab4ad193b0c4bbba1ab9259ce62168daa453d6bd03fd720177f17d05fe3fef;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h59a7ac388af6acdaaebc34d9d9ad9b83db1046ccd3177506f8d097382cba0ef49d15b1826d831ae6ab9cdf2c652732368281eb974fa516d7f2ec6dbbc;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h506dfe11b0fc5cc1b0c8b068288635da2dcff4c2bfe9f413120c3e7714b19d0aa7279d585a5355d8ac50c51c73aeabc8514ad8dd8cc115467cdfbbcf2;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb4bcc5b73743a887e731b66b46b7113f29c263d88ab838062ea5eecd110bf17b2c6d9931b1012574b1c77c78b2393bf1db9b19ab39d9a673d358def0d;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc2e2e1672b1f1c18a9d75cd6e61873749cbb5209a4181a59dc4684fb38f9288d6f1deb039caaf2e23a21261d201121433bc793b665c73e5d5a736c234;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5e824090287452fb3925ab7cc5253211502857f3bd2c9ca597c4613d58aea071ca4ad063cbcb90f5e4e7daf5885e6d4e6ed664b7b3f2bca17e2dc16b7;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'haf3eddb74d9f3f5732ba64ac40e07662879032d82e8e26aec91f448a639fdabd9b98e70ca0b0faef78dbfd969170157b9883174664b1ceaba7a4b7ff6;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2465926e517bf79ac082260fc848e912ed5f097050cf832e12da3dc6f1dd4e96c59ac64043803c392e96b5f432276bbaeaa8f248db5d907f0fe21af5d;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha9d04da4964bd466832221c5f1ecb3dd6744f6fffe53e3842556b6f9d6492edafee199250e0e67a7e396400029bf1eb1dae3e4a3bc9bb9b83c2f6b732;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1e44a7938c1b599534135c072bd3ec04eebebe754c14d5a929ceb543eb566037db893174b267bcf984d311fddb337d11e33ce197639ce9512339c9486;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3f11d7ef19eca9dba620271037618de1c3927b357313d8f66135d418ae7518279b1b694bb8a21d347fb64077e5d86e4bf9445b8cfa79b8b9d6bd9cdbe;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb22a8517f5eb819a952809bcec8294661c3d47620f37271c09ad9ae58135f1a4cc6cd0c8045c61ca2845446c5d639474e1fb794f8d86b5a8d51c71ae2;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha9d6b54a67dbe22700be94469836e0fb1cd7f2c009b6ac4c6a70ac119d7f8db0c95ce493d96b75686051ce589e9f602122422943b4fee4399040af836;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h77c43b1a03840639bf1577d6d6032e17b093dd4370921058e9b18f4854ae679fae88a1e58e8fc4a58f42a6e7685b39b239ea08840ec29cc13c087663;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha5b04db54ee793926eab56c223ddfe55409aecf9e2e6dd57f7401e4dc2f102bd9b464877a89f377160fb9b7c852599e8a95d4df1a201698d67658d0e3;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf229aa700fb6cf612191dc8d4690e599a35d1d88529feddffb60bad8cecb83363bece2eeb7ec8a9b560caf2aeecabd922f20eea69bb7c350477e71dbf;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h38a8d18c5dcaffd3381f88433e02c75be683ea708b6360fe8bb546385d6ca1a3d50a02e6bc865ad66a3525b36f364c322bf3539c2f4f2a7213eef81b4;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3ce3d09e65fb16fe4ea96be7a1025aa211a849f85c81f7d3151ad60956ee93cef7f9919414ba0a27bbc2a7e2d1eb86b4c24e7e51de7abca723a0403b5;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd0cc666142b34f5d08019db27d6dc4cc272d044bc3fa5123eebcf86fe0c8f0926fa1acf8040a9b5bfd1cbd429bd105d0eff4f96b9c17d839c6da5a8be;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h730761b99a3806d3860b9e09426d50fbc4bf76aca4e073b3a2f302ebe030d834ca2b3153da6dd1f461827c437a543aae1815e728f439f51e14b99343e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h164718d4d96483131ac52bfccf863f85def501dddb0847ec8bc53e0b584edc7b46eec6991b61182ef35fd360f616011266c7e5b8596ae38b3e1be15c0;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h61ddbd1c5691f62d69c2653b726eec07688f200a78d1547c5aafa63b6707670ec624aa0f0785d83c50a0262ddae965e9107b1abe44df0b7eae5eed75a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1e4224f8b6e127384d994f61405076a5b589841ff98755c23cfd8eaec4f4dc009e1cb700a335e9c2cd5cb6369546a7c591b3c81341c91d9c13b2e3c17;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2c758521aecade9753fb8cbb99681b754d93eed7f3a1409d7b4bc9fa6cb028116b364c2acd3a7e1e39f05d8935033b1d5be799172e212108d1a45546f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hebd7bf1d5ebf3030dc94b19b51c0b8006f43176b4809eb0da1fcaa36408adf6e6cfada61a84646acfc7188fc22c589eeac670164c78b67c8b6a882c20;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1fd6df492b63c8d5822fa54450d4bca5edd795e97597424ad27808dee8d421f897cdda7dbb4b27b1a039358ede3ac242012cfca066b4b62c04c39cdf1;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hcf920c1d8422829174d098909c1da13767b297ce8e30547dac65749f58b490cf4ab3e23d20ddd781f67b7cf265783d1ce8de93389055babdc46a22f11;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf11c3edd09db93e1bab934758cb84cd67c085dfcdadf073ecb8c83e771e07b95102925d83923200e8463b257647f1afd124aa44703674e78aa2519bc6;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1d6687fb11bd9f934dd2741c093730d3ee6dbb0e476ab4189f5188c09a429dc2071f3539d665a1ce9f77ad29c5fd0954e8f98573f709439be8fdc1e7e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5bd1d00cec48aeb96da47fc85cfbe1255d75c72808974d8e05774b36361625906c11666f0ef3443559d640961667e09a0ad5fadbd4a143e7d8fcd0a58;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha911cce667b4bb386f42b64a97eebe330f97b18805aec4cd5e2f1c528e6fa91ef39c3113b8feb29dc356317725bfb3989dc003c4b064cccbe10c53be;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9a3ade318ceb58b650e7a5f9ee8a962dfb39573a7b56ff4d97d362804a23256bbd7b3ec6799f8480d3516d2780d2222cca1716634d66792f305872bd6;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he1b463b5cf5ba5c6cab13aaa97a08e8561c16cb33cf33473674a4829d04a39da5b4265b56b67df01b3dc0b1d42f024403741b2d3f9b0a6eba75dd855f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfefc01ab34790baf560e080ebde59df042c88e4b70013e74c8464d87ed6f0626c7ce344fd62a89924689345aeb55785204ecf4cbc26aa0626fe61e945;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2dc12e2339842a4b26ddb412012d01775abd54927fc879f12119eadf03eae27170b9833a9f275eb9ac45bb0380f940408bdaec85e39c016d584b47199;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc038c9b554439b7d2360509d5694810f23f346edeccc915093742d7ffca7b51b191ae7ef504d536618c5f8d81b8f2862b9111c76ccc82dab0608c5d0c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h63e82700d039831f60c99b9933704954d3e7eac0d90a52d34d86bdc095ac2b1dade9c4899789d279e4ec24ba49105b8483a37051e6a20dbe70468de36;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6b8ee39dbffc246f46bd8946f253b9930f9590aa49f751299ce4340c84580fedfda3113d5742b1a05a9017c7b5db8bbc232706d2ed05ac9b72c6d386b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdc2d5c919621234c241fe5c61013ca70a9b9c47fdadcdf00e4343dc28d1df5788bf5d50c634df62aa65045b498f17c86cf42d520388b416437601bba4;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h567e89645e412b0ccfe29f1d00e9309de90ae8df884c37ec1baf2a9f5abf0015ec70d1c7025d40d4a17914c8fad1b921dde3b802509c93c21a2db2eee;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd726027f234784523ff2817fd61879514a7c89344d68d02f753d24df0ebc0ebc464bfec113c03bc9b85fe6b7786dafde389e9aecc2de2bdaa3f900e03;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbfbc4411d4b069d0ac3d92a4a9ac74e41a1b774f6eb2013aca469ecc7d4c7bb98aaa8729f8dc6ae854feaf7457c98f35b73344901d56d302310959eac;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h20104c30a9eec353a5019b9f78349b529db626dcf1a33e42c3cf42cc6671ac6126332dab1b512aadd21b110b49accb6acae3124b0a9e99135a5d5192b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5aba5c99fcf100748ac66dee68c99f0a54cf8bf86ecf508823c929cf66da5b98eb80f698cc7d141ebb993c0f687d2dad5e69ead52f7fc51569c022003;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8ea867c48547501e46f21465dad10af97f2c0d51898e9ff98d4ba1bc76fba8fb40771b5399706e47053140603a9c2fde4c4abad4c0d38205faa7946b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h281879d86b5cacf0accd4840f5d645a1762c3a776576188996fb9e7b95eccf2c9f854b21d8871afe84c78339646c6a35426d544d13ef232f4c101c20e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h839162c66f3b46ea6df460f2409a64194dd3f8386fa282323fd41badfe265631be301c5ef4556e6aa502a5a969d65f53d5d1cf1f0fbc7081df3a370;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4633f00d8b3886cfbdd0f5c8ccb7311c418e461158d1cc76cf7d50966b891be69870d5297b2af4913236ba11a82e235453d4615fa0ce2cb6cb7803423;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h61fd6092f2b26466f224b4956d47cdb259d839257541a0fc697237d1f74643c6a72e3630f4e8ebd1f8ad5ef6749978004a8dbaa06e34ccf1df073d74b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd0da2b1945cda2c4092c5f7d905c27a226fefc1afe6f61c03c0ab1417797fd6bd8990ed93affbd860157b4a1fb37ed3c407ad4b93ec0f7e21bc40cb1f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h554b9c58b6a83640a260453ef01a82b13347223121a8184468af97b31730c3613073ac3b13c9c27fc2da7ed8371514709e9b8323e5ae11e60072f1658;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6de485ed771bdbc73c23373ddf2a2070ea9f9af07c5d7186c3babc3761f07a138721dad2275d27ae65ce5b1c8ba03cc42fa43bbeb0eb395327b13d956;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hcddc4a4b78b8885ef5c8f75eb631034bfb05066082114a3cd17c6863ee6202f733820f259c16c472bc49e6c8887ed92b216df9ae6c4c75d10ab654cd6;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb87a45b88c142d6be1842b3dcea7bbfb91d29966f86faeed61dac4a20c17779a2e5c486ae9c4a384056e4e616c0a91a814d194e7dc5fa9b399ba892a2;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha7f24b1bc2abd9491813b0c5ba09e7e9cd94ce73bc7900bdf66710553d8db91bcbf5c8e70028df87dbf914562b36d4842f55fe6ffe7407003fc459f2e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha2d771de5e8e350657aea8025dabb53d2df3f7c0d6221e491975c42d8e97c3499ab4c9643bf8cb2de656fc627a5aba7f8e7e20cf7ac436814aa8ee205;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd1b8663a83d2cdb46d274089bf0803e9ae79f789e7a55a207a1b4d68d6039d50f75e6ed42be41de0ecc99787c2114087ebc3f66496c66fd831e6725f7;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1a0f56300bc32d722a716f0c43ae8a82c9bcaff37a2925a397583f2849f01b0e57bf440698344b5fc5b034e2687d817993c4684bb84aae39a10fa2c7a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h584a78bd8b8986a16bcdb38aff66a511a9e0b41ba6e7f377914a24bd8d335d2c0189e0c7c3203edabe78c59e2215d02fc2eba631f5cd892b1654420d4;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf108ee94335f682150bc09527429bdeeabb7de9a5f024a549d57e28f15f66cb64f0545252ee53970421c5c19d0cbc7791f207a2230c56a3ba3ca6575d;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7983de9868d3e4618596872d7dbb2fe4a479d2454abb7596c1649d563de828fc18fbd632d140bbbb6c8ea4add35bbc2710675d5e134ffff613218be6f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4158dff4b35e58d176a01562c4449a7bde25459a81a6aa618fcfbb6a96bb530c1974d494f162a68f3040376bcd76576100d45bd66c6267851eab17971;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5ef4bb732d1b396526b8aa3f5fb21965f26a3fea04c96e28f22a9d2513e16d997201ef90494779d6adfcbf1448d233ea074a3be8815eb1779a46c27bb;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he6e202ded5dbf0a86965b8b421416b5104d76c70c4915d1d37e4286a49b8ae6709fd20b716eed1926ada7ee555814862d70d3306352066e1f233ca5ec;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1e306938ea92876e7371cb0f14f637a3c50bca56fbd0398a30fdeb90898cda53febf686c83979ed21f344079f13aab0b19e28eb758a373e8adefef185;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8fa340821f25e50362f4bc2e733216e28520346c2b0060ae80e43924e966b6002d293b4d698cf0631d0c3d345836949eb7d1d23db91cb7942e52bf13b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h65d01a9527d81c3084edcbcbd39a2f22d2b16d0320b79ac2ea6f2bcb6b35f4150d1c47c9ce64e55bd1cf36ad00b882c63cc081b0906f016fdc48d00bc;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h69c27e9372400eaac345adab4eeadbca99acbabffe38b216df5f0118b8561564f53ffaff271294ca3e35c7f1df6e84f80ee27136025ea26a0dcb4e261;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hcaa1789a8e6a55ccf12b787002587f4a878b5b7962292dc0b7563609af8f0911742f6892da7dbead3be36c95cbc9480afe68a9346e71b89a543de48c0;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd47be0accf8f96e6c40a0301eff1864c7fa0fd4732904a0f3d4fffbfa8243f6d9ba12bbb7fcc77a787b80d7037072c49a5d6075f6e965c95d406668d5;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9df6c9ce89339915ae04798e9edcb5a7c2857e1da66f446b9ccac2d1becfb5337537e28170197fa8d20df352bc4c00334bc127e60f712407b8195a311;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h328b8efe90ef8a1504fa5a03af5e11f14a3e04e7aad91277e657bbc05d3f13af2bd21131f4a0ecfaeab03eb3d4e1f4da6b15f2be3e40207295989808;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3da003536fe72f7745c10ee47ae1ac8e80d2de35d0883b8664d91d4027300ab2825b9e05fb96e9c9c90612367567fe5fe232f7d00b8370d91bcc48ea2;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd47f3543c8f786d8809aff61e121ccf85d84c250ce8358554144a5d6d16af940b30fb17348474209c530e25cf470562b3ff32a375705bc129e72025f8;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd2dec22a7c000d8d3e1f6bd47d94b03ee0f19ceee71c12139058a4f6b96181524a7354b5f6e2c19de6ea9c71106a4daf7ee52a4a150d38a8f7838232e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd6e61d856d9172ca513ab836a468122d456c29a33a42b9bb2baca51db378c0d5931def88d1e307bb80387b2743c39fe26dae6adefc75aafae517e9ffa;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h87b5235cf1f99a72fa8c364b7e2e98fb3e590a9d8f1a94f9790fc75df822685349d0eb4baa7ed40573b5fd2bcd84152a7a081cf139f4911f05a4e6d2e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3b5d8cb4d219d5ca636505d46f98235379bd88d53073e5efaf5e7c2c306628686803db56a6f01804b5f05b5ac2caa7bad62cf4d57c3a05932a30dd4b6;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h176b56bcb004307b4c097879b5b928d9726b69708b697f54a7f1d9bdd2e56bdd8c6f0791e62128dfdc0edee92fb12c43db646c504ed4a67a2eecb4c9c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h59cf5ae914415e6bbe8a44b354ff21709b2f387bcc7efb22f88cca26163203eaccfec06f0398b6eeb6f6c2b7893c4628c7e65d3cfe1cace000e4b858a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h96c6f530fe8b2fd1a3b5dedc7fe65734b280ec73b40874671ed5368706f09f4321dc0ad2858f4fd504503ae34e9c91ab059b785b666e79b20ed2c49e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc9bb39a95a0e48b8fec3180625831394071a380c4f81951377721fdaa1c28902cd12bdd35edfee6857d09b85e38acdc491ea9b5698ae4b0adb899176a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd268b30a61613e18c2a4268bb0508657069725e14b15e875e97971c8d963b09a8513964ea9fbfc305ebd47507c882a31d3d4da193e797c53ac6107a98;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hff5443cf1a7c98aa027e2e6239582e97d68c99db8de26910221a4891286f047e30be2d6c08c037b359d06c0637dce22584295a7b8c8864944e9dc0f03;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc1c7f7c1ea64a767e3f9a9bb9107eb0f18d8ee483ec210e509d9d811617a3ce949a424f537b26ee1b1f9c49eff00019677c02c436126e8dd2004c612;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h377369356c589be823f0876b2d26ef5cc9fe5228c1f70dc4d348826a07e337d5785025d0ff5e020679b68278797f41d31af8fcd582b072657247367ff;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h673804ee348a71be8da8d4d421cee282665966ec8f2aab50c89630c87a294a52462f7c8a0171f2806cad493ed1a3fc6f3d5bb5bc4aca520c9513b74c7;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h273dc00629eaf08e01f4f458ed5d3e7657a3bafa57f3f9ccfbc8b4dccc9520a2636573ef32d45450126553907454fb676ab27675fe0112d3c9123808;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hee03873af2b2d049885e73b7df9c5b63365b5190fdf6606dc0c6eaad2d76ca2c693512016a82091fefaf131da40da193f29e2d9f7e8818307eb78934c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdce0a3cfbc7538e175012e7b3baf8c8b020593360687c79060316087bee8fdbd72be06e688b5db52a93a2238fc60a5b90946da67f569e89fe522fb2b9;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb0ef64f7a589434f0f1bb1d74d72befde1900f1372dfbb223dcf51c9dcce60affd7995794dd69c8c2e8e75d78a08edc3f4dff44d83ffbe69763d39444;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd0bf9639cde49b6e4973d87bb35913571b6ab3cd6f3404517d6ff2464bdd1a2e703759721a777b5b6c423d30b70e1ed51d6ed40736185dcea2efac286;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd4bd9db8653f5027b5f0d423382845cb27b38bc55c6d4e7e4a0a51fa707127ad66abc876b9e120018f810c43ddfec2bbba158e2fd29f86a8207902007;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdec66ede20ee069aab222de04845a38e5bea769be329200104802eaf905576c9d5780b87b4bd7441b342b73cc68f4c4e12b3cb92cb90f8a7f6918f885;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5f1d55ad89e44188692abffaecac515914d7e164504bc2c7690ab5bcdf6bd244e549f72c2c2330f280032d1f5a608c5ce83060f6fd2780efca76c61df;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h19caa2e9af9bde72c40d48e8ff8a749fcfc02404ebd6cb66d17a6ae5fbf0296dd2bd0fd568e4f7c0398df8d2a276298057ba40fdb70faeef0b58eb8ae;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'heb14fc1f40a0159de86ab25cd47cee565d058e4c003b7c106d86520690617c365069225c5971a1ff29e92379efe023a005a8143ee91a46011a709b6f5;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h310291561966f309094dca031b41957d87a6a34b37fd39ad01a6322d8050f8eb3ccf3c5335385ca39ce5d1dca70720622e1d5da84f9e2618b4d1fb03c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdc996c499197e6ce16cba10ea6dd167e68356dbae49016ee367f6f257d602625430174fd4e8e7d8aa5c4c07c04e22c50bdb77a8abb2e2c8e58382630d;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'haba7f838f0c567c4f9da9e80bdfa6875b77e3f7a908946e3f74a27eb3cf2e98e91e997f0b2b1a0d9ca5ed30a4aac9b0b377e0bd5cbbc64a8af753fdfd;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha30d4699d318fd070b159ae90a4ad6a1edc13c9ee0f3fd4f1df3e9c8e600a811f5806c6c3175e265fe153396fb035deb62b5ac4b9daced14e19cdb167;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8fc4316b4e4ae0e4252fd1206557e6e5c6026a0e528691f39a0500509c69e1ea69e006a5dbd67cd63c2ef54cf5179f60420d23651625c91c104da838d;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6743708e00a86e3eb9de8e2e1fd64fbf516d6ad183f35c01893747cc4988afce3738530828c509eba596b9ff94db142686a92c52584ee20a20128889d;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdf1c5e4a774df9e0fe0b8603c8bdc750dfbf0e8def447392b1a779dc881186a957034049bb58612a5e9acd2caee2513426e8137fc0622cf2f6a75c82b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h72f123b0b87b6e9cba70df8f870359c6b95deaeccdd4d00df734cf7e7cefd47cde1d312c5d53c88f3fe3a3aed71800fab64396608a17441d677ce22da;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8528c5ed4158080768f5c7bc899eab92048982cf5fd652fa04b6c649f712734ad14c71ab06486c1068df28776805a3838908b582ff7f7dd16ecaf3e1d;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hac5c6b80e4ff7ceb91e2576f126b3f4cc443357f29e386d75219824b3a1eb0e22deb3a58a7c0b0cd034262d76309aa35964e35b3c4d60fa392f7996a3;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h323cf918e30261f2912b174e824456b92d45c48cb6ed0f8217285839ba85baa3a6b14adc6da2f3a7a6564c66962c74260d7735d65cfd213c23600a917;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h15c25e14bc073ca3472523f0a425299b386a1a186299d55efd0babe659fcd8634ee65bd45c61f521b37d06a02d4bb995dacedc8c145a7647186a21f6b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h88076723dfc2f1c262b8e60d5f3ebf794498b8b5d8dc085fb7bfdd9f1cb6a92128e2efbf4ba55dde6ff904eec5ca0e57ace1a6ddc19534132b822ecda;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfdcb80808b5737b57f9d9b2ee52c7d461a8c1ec7e2282ac4fca5febab3afe92ee37642c39b92b4116b8e9d05027e8694b3ff1d7e3f58449b7aa0aaa43;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7b56081238c85cdcac71f1fc47b63f500b94ae1feb3c64fc6894a4d7b93ca33dedbfce78d20c49520deea374cedd556024c632e1ed68b39ef7140a2d3;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h73a30320813f5d163ae18e12216c424031e96f958fd1f12e700257a26eb9c7727616fac081c4fa589950cf2dc3522ecb39af50596082874edb922b229;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha6649ca4940a25a885e870e42feb6123fd66b0d2307afe5cf6ccfc236ffd9e1449e4a761f07070d9a8afe1c508aa559b0aafbd1588f0160f0561a84c9;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h67de220c0c074e69fbf2dcf34e530fb94360d77c8530629d284fc00158b2d6fb3341a2354f15acdb9f60601164d612e8cf284e431005b03911d8103c4;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hac035d3114b8605598b5e3eff8c3c0b2d5596edd1217d8d61923530efa8799fbd911df3a38265bfde13adbfe9ea0d87ba7987bb7a0f626c827779eefd;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h91f85ded7cfb443c51248992eb995ca92ed6cc0fb56a09d64bc5fa52660942ef871e3d901ef32c0e093463095fe6c31476afa549ff5b522a970194d12;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h82013dd5db47459b00cfedff08b80e3f7456f71985b25db465152ff145bc70ae6f09ea050b8a4ac9d09db4dcd274bd3af2129386275e0779ba9a0442c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdb325da6db6655e757cb19ae59981565e7c568bdedd3b1001f7c536d8e5973d6895dc6b534fc3527813d234ad70dbb7aac8ba5d036aa83001f7dbace6;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdf1913c90a397d08a5fa4ecdda241412130352719bb5e72105fa485e5662893eb89918ab33dac3581857da864553fdfffea0ae21f084a9445f48bf323;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hcc9503c7bb822567fa265a7ed4db5887db6c14fc03dee4cd0ad73c1dd73f72bd8135e038d65f4b70ecb855dfcda54ccf47509a58fb066b57d2e414abc;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'had38ff613e802ebdc0c987741fcd4b2cc91d8e91806e2a4a293ada722283671f4cec60e7c60e1f33c7db1aa0a3cb61601632b51ecd25e912cd907661f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5df007180416b2e1a3480b1660780a457038714267f9e5e1fe908dbdb586fc1ba7c1b32dc65ef97ba6389195b388d30f5e24239a3bcae7472e77aa836;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4a95bdd75d3d517fda35f800303a9bdb463895d65bbd137f471b594c9bfe90811aee88ed12ed9c736328488b27f86b342c386f1956dff4a1d52a1be31;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6abb7badd476a7148752a179a824ac6693091b41e91e6cb023af4c9f976c25aa716f6ce45124a3a4094e68aeb3703e454ba24cdb6e07f08f8e7c36515;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hcb0c8c0111ef4eec90076bfabc3f8b43569d628aaad4874b8dbccdf436c196a895e017de79a9dab3bfbb9a9f7c9ce3eb85de0d1cd522dfea97755b49b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5f2a5fd3c09720cd854a7d0e1f8c8eb594feb3ca31d3351e63320f7637b9aba918a579f70f6b75443fd91975f5c7be0b373c613107765f08a800f9de4;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfcb3cf69613056403981863ec93a3d55ccb4f10c6f18e9459daa0b307c1c3b323380d4bb3aaae1a699032097006065d5b6acfa347db0eea4480c319a3;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h50e934d07eb15b0385b68bc0ff8016f86b9d656cedcc1e6b2170df9782edf8a97c8d6277a124928806afe51abf3f1681bb2bab0ea5f1c760e9a6d2754;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd20ffd2cd70e2410a8451edf0bb74880e91e16f04e115886863c9485112d4ff7f81b08ced564243b47295700c06926e872c7f8cb1a06745af70e92855;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7461dfacdad27a49a82b23477bea1d0117a65272782f421e43a8a35634d160db2385fefcdfe2fe56d913e371581fb06cddae0eb6bedd4486cb5fc64ad;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h94870c6bfa73f8cc5a111800e3e9b8d17e99b33d6ad5586847a870eb7d1ead997ec83349c6328ed231e0310d69f9b710f7211efa2666e3c031b2dce80;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h91aa4bb0eb3e1a6e87967d1ee7f02f6a70f9e6fa48785a0a82c2d868b7f453e4678f2f8ab9d5682a67134328939c56677b1fce69722a52379ae433645;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hec37ccd70fa567c77cfb4681631eca44a014ca2573ac5e22fa21753fb95ac0db6b0dbb99ffc174edc376285966de71febacad6afefd59cf10fa299655;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha2296b27df20fb1bd78f24bd65d40406dde8b8ceabb5078cb7f042e1551afd526228c7f839bbbd45ec89c196a0407d4874038f234581c6eb320346073;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8456654cad6991f4afc90371dd23a2e1a907798f597bb9e58f1e81c178064b2672308e3dda6478bfa5d4e41713aa4e096b6a3ce71562de49bfd2da64;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5ce6c496b0c5b6f96ddb581583827ce836120327a9e60c0de460ca5e5f74d0a017daa74b4b8dbb595f3e6ed91781a6b10b6faeb28c35e959162d64c0;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7ba0be7e7c0000cf24a51c4dc892be022bcabe8954b49cdd11226d74f5113e61104f3cfd2863b3320c5103bd64c18a41c2afeef3b43350b7cac04d3e7;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h30ad0b847ed5f494c7a60f99ee12e7c2dc424fffc778789d38c798bb61c2531f3465049a52e58a5be9e0ced8983ef82344f61e9097f63553e5d6867d9;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf91659a3d1d27c944d5a6ade329fff237c5a9f1ad02dcdc5a3c8c863a065bbc92dca19f688c88f108b7076395feac7667383d062078e73b248c6df492;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc3d2e6a922a29a49b2d9bf06cb70dad1fc8a2baffad94c44209ff4b0237765532e9c8a3e02afeac7f6ab23a0e86fce36c6649da27b62392446a5e2f6a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h52e0ae44b5e88f5bb476a79f40b76ba10b4eeb608a31bf2c66a9acce5593c45a5f800a89d3e00f86a957e7e4c36b409793f0d041d6e342e5a511a97f4;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb77a26e33ea99cfa749a056ddcdf05cf8f32821c44d5faf699c25fcae054bf543258bf3dd8342e54b7a37ea3404d77db742d21ef65dc0d97434667f46;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfc5101d8c1f9342758cf03c70ee827bbe0bf4d8cc1d974fc0518c50896bd93c14299040863c2d210c6ba92c7b376b58a6ba4a4bdfb10c6dbc075822c8;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7d89ef3b4f0cdca29dbbd8d79d3265976d1a919c37a7cf6b04f23dc8664d6450ed3db279bc56c978d17525b50f40601a00c91a0adf88655d76c8bf9b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc2bbb2b0ce295161d0674b191c52806d3be3a8ffe8e82a4501146c62db936a7440da3dcf0f13fb9d278e94c84fb0e134a6d2dcedb5ef186409347866c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8c69f74c53f6723e823ceb77507ddd43e22bd8e1a7e58d9aa89e17ca152d874ee47e59a3f6543d084e1294bd97f57a336509f0f004b2dc461088e29d4;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4868b93ca9add6a78d2c5cf5feadc42a21f18e5dd45718d1af97446a96466de509b50a24cae232488866760f5b86cedc6cdacdc444a8565d3d06eaeec;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h935926f2e9f773776c85ec1ad3ee13ee98d17f743769952dd6c596ec0f801a882adc9d6a1074686fc9665b380b56dd46c09479cb1fd54e1df65da9fbf;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h62b1dbfb198581ce0b85c9cb08ab273e1d504b276971c688a18d93fef3b830e3f4f1c281b6f97941706c355a7730493eaa658400cc23325aeb466a4bd;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h80db77065479b34612fa14a58d2875c3317b00aef059a4e29737b07024a82c02be0c173985b5064028f8b7d9c7f72684206a94d4fd9cbcfc2272f9c6e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdefb343b8dbeaafc61cc06a786c975ff2e7de755ae08ae7c809e8463b190cb59fba4e4c0fe3a77a67014f5de29e3b2826c75d7f4037fe8b600dd848f5;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h179d843e75f152b7a98fb1fd11d517789ce65cd21803ca4dfc30b06710f057ad6ea500dbc44ea2eb81822756cbfb656121ab18d2bc112ae354c010e1a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h55c3e760dc2e75aa0ce3a3c01e7fa42ece1291de099c8d90efb035fa7edf0c82190f2e9f2451e946cac0375b7b3d983271be220e0c0916d22d44f82c0;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h76b76a3d71241d39003aadb980c57d89d283a7b1b9e40b944c644d4f2a45c3bdc8988140673323cb055a18f7da19f2663a1b9fc8ed05234a4ed17c8de;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb2f56be248592f5112ddf59c51459bfc8e59937715fbfc51426832d7c9e5524f74da2a3060aef66d18cf47155946342f176611d8f3df4bfb57b2d0e10;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3c2de3ae6323a67740499b63a4e9c3c24c6a997029c84a057c6a05b79345e8a707668b8368edc7fb77a99cfdfd012871c7a3ae7690c6542764feca3be;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he978ceb24608792be3d37b9a9274228e8cf33be4a52d7263d67ef1931e6ae6748e8f20e9cedeef7ed128fcb4c60b76b4ce56844e2e477c46cb6735ef;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdd4b13fe25b170faa63e27629abfda5a21193547b60345e8b5d2bfe8107e50f044c2ff28fe9b5339076a2ca8bdfbf9c7b2ad0a29744cedf8b25854bcb;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc57eb5a92eb2f63f8a1959646724c751374cf4b8aa932aad6fb2740442b87ed66bba1d49d843b599331586fe7bc5e12911082de87272541fc212908ae;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h11a008af20c43bc1178570708a8d5fbcce64b7b367ac286ebbcc5d62aac93715d994f2d1804005f96ce1cf2e22ee2a66e1128c360591d873b852ff1cd;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h203a340bcf08b350d2796377311ffa89c4070943e5e084fa9bae888257aa5c18299716ef5efbacd39e924f8d81eae5f4c3b51ba29c17bfc8b44098cd5;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc58526db71611123dc26a5d06d6e4b8965d5025b84c81a1a65b9328cb8446b7b323df3344489c3bc702bd637f3c2911098282502f89e646e8630d5dbb;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h50ec5cbdcd1baaba89e172aa7df48a63c831db8b2851969f7f20cbc2f8de7a00bd84ebfba9bf90a81140f7ae0131f5797460a9807498f5b06d436ad26;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd16eb08f0cf959d6630dd46fc05af13a43e7adc8561ec718420fcc29a116c08d85d23c233574ca7aede14a12cad593c64acd647eb0084ba93dd652835;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb5aa008b5e760e31624b9528a0cf4884b6259358c9415d63718b727aa4cef61656be13fc45b8308e887abb10a9ce267039d54e679ab22ba276b320cd1;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc54393ef746c47bff75a92d296d0ba354eb9f5f9e6ce0ba4333eac03b719495fe12f027f6344cc4cff4ec68ebcd2a303fb9f92e1a3e7d126f5de91a82;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4888b8299068d770161f229822359872970b4d54f2b93d3c187679ffa1108f4e0cb301c3e6bf3664e64f8372e14648d40c2759a14c08f38bd64b80fd7;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6ad695d0f152a1d519ada138ac03b6246f4b93abee202a1464541a843270e7d24ffba3e8d3f1d9c0e427d11b03e6dfbf5c162ea5047261689a96a10b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdcd5e3c61135657185c62c46b812a5e19dc6f922db6d34ad205fc50de62dc1d853b728ab700d3ffd0ee433849e8029308d4e5f1b10389ce9685965cc9;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8bfac2d9d51e39cd5729f08c761958fa34541892f2da53fb87072bfaa82701091b33bb1633b3da8a32f2f42b36e8f987e38e56d3ff5ab77945a779423;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h355543655db5e4b59e942284f92d515a45b04bcd0fa0b8df7147ea1252b7a34e26ba04498c3e35cc81e256203430648b4acce0b8181e5804a295c6b3;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h547cdb766d2ba9e8fa3d12e743547a90c08a8fcdbde89e98cab0e632dede163341eced2278ded8ab92437229b2c9e92f136435be3033e88814a4c7e01;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'haa4d470c769213ec2f5987bc8c5b0ece61810745b3c7383de8f38856124429c6e70f6091fcc420f410eb1153c41286d642841bafe62c5a304b271e9e4;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3b831ba79e677d799b503a2d75f1b710e40c8525ac3cb70dadf419fa2f05eb8abf4c052348d7adf5f17669dac387c8fbf756eadf603ada835d1fd8362;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6bf6a73fafe84c7d97a4a4b0b8f3db3106e5b89d178888128bf22e04ad5f0c154d03be7a61633fe02b892b14cb1ffdc038bf1deb1a879e4904b57be03;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5e38ae950bf149724f5ea535f7711bb3f494308ec4a80e4c1c3e54ded1440f0e207287b91fd52544ca9307a6ae8a4d616e0294bdca9b45687a1adfed;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9b5ee4bd586d69f35745bef5c58267ec4f10409eae6611a62ab11223c9b13a4fdd3ee670f9ce1eee55f6267dbdc6a98b9c2c34311dbfdc4f3b9907fbe;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3b5fd8b93f396bc77b189e29ec8ac415cf6b2294f39064e923b7e3b8d3f60848fc420bd28c5fdf452122b475fcf1fcd419472f54b64043df2e5d66fe1;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hed1593b98486f5ad65eaa5be75ba14935b3b72ded1668d03b14449cfcf9246fd4be0f9c9d1921b8953a3599d181effc082f723a6d051c47ee65f8308;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1920cd9fd87af9c37829aa0d703f15f5fc9cd374624841470f0a871afdbd1c5ce046632ba3b997e31b598e9ff4df20cb0e4f3ce63e8c3d0968b629b64;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hcbcdca9e8976862f6e45e608043f9bda4468187dbc3f99d83d9c02effc664fcc5dc032bd5af3431c1b69722c5709e64de0bd053392aadf7cc8b6021cb;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha2d338e560140801fe34a5320973aa8896d6f6ae98c9f753dadfb5fe71f79eaf8bb13720ec85cda211838799f16fdedb40a3bbbe5db58788103a60bbb;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4a8edc8df1aa345a31bb83f04cbd941ef8450eff8565ce5aba6a8f84acfde77b22c0dcdca03ea9ec27ff52ab361b054a78d674e5eac5907936736ddcf;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h115d3ec805c4308f5750db7175a66dab365068343da8cb75aa99756a12ed8aab6025fd6d2f0a1455eca299acb1a427273cfe542260c3c46cb83a13ad1;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6c79fecb951200875211ad7e0415b6ad0337e74d342b1da7d1a52beafc514e4afa75bcf9a04b56f8c8830685a1db32bd58f872e4e0464a5c492dc443a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he687ff78482b9c808c2380fba0cc72d5570d850f2978329f1572dd9a26abcba0a479e536dfa61f7f13f7df87b12fa3a25e6fc4ebe8923305d2d4d1f17;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5aa7ceb477c82f1ae7faf0c3ae79d064292ec855a97ea3b6c8723e9985e0943da74b126c7e774c640690c4b7b9910ba386f8d43dd7bacc2c77cb533d2;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h14c0911130e2d085dc7d233047164b41f5f2ae8eee37c26152c2614c92dc9ed971c97bf655c118f5f959812c32958f103db99689003e8dd2f1bfd1123;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he759f84d4696757dcd337d4ab7aaf8dc7027a7ca7767402fe51305201c62a9e943dbde36a8952699163084009802fc2385e35be528435fdd21d8d88ed;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1d5a47ce9413225c21636c12a83d7c4bc9c0c899a1690e853ce4dd1a7502c328eb4bde16a4cc67f4606a4d45da6baca9eee5e443680a2282b07268eb6;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h28f437721b77d74fa5bc108983a33b8f26803be4117a6ff8891c0e73c6765c88a047389f43ad42841c377647ebc232aed97662fa966e9054e958b1c0c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hcdf37a0d2dfc46dce3d39339d0d83ec1993aea72c70b0161dda5f256b32fe8e50e3097b25dcfc4c12b5e402adfd47fbefba608684fcc1b84964c8bd0f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h73c15e4f5164c35d8f799e27eeaa19aca39bb57e9cf0cde501f178599da4531d1e533aba1fd8ff0260706ad5350c1ef1f42df03eb6cb18ef6e8833c8e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf20e0589605ef8c56cc381832c8420b16c996a5027d54e3615fa067f0d438a9fde578d90473b24ff2942355ca19ab06b5193a0122cd1c878b4ba87e2c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb2183fc3797340972a313bdad4ef34bc16e817401d00d8cd30d9aff259aeba3725d7ac0c3f3837943b46df31452b6cdd7d45f8825dc50432b253c70e8;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf86f94008e5a17040a9b58d584a5e9a02c3346b8c8ab6727789eaf9a50b51b1117cc78a2075b147706bbfc86bf62842fbe43b51e20937cf8af982c8e7;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5f242a4386b1fa086725f75e5abdd2f18a435c0307b6b54cb603a60c0e34cc11ab25ab717e5e6b8beab493f37a6f67a7fdc717ee21fbf2f20f41e29ff;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdc83c2d2dc46457f74112a52e507a6ebf15155a34fd5f81471f1ea17feab6da1a7685c7878a67dfbc745a70677cfc8870d11f6766a0d74ab4e2a478ef;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd4c961bec4aafe7c095407c3593500e115418f12da1cdcfd87755712a4ed67b260d09796730c33faabd126f86428e1e57b97e830bd06f2e198a47be0e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h35c6c4868bc5856174cdd8f4e191b4ba1fc0f32c574140997570f8dfb41bb4ced4d5f555ff82abba51518b339ebc2cfe9d626fd5cf1c0c9ed75dfa7a9;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h37e2be708d4e190c5665ee373aab11de87520faaffbbfee9b917fa2bdc683a887628d90c03012c07767bf7d876a2b68b1fcafc7dee1f131ae3ec1f2b2;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h99ae3d3c1cf9e7ed829f36e129c395e69dd886ac6b17212bce389163ba1b82b82d8f9b85ea527efa80214878ec1ddd2e3dbe6ebfba60b854f96fd25cd;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd6dc44df8a0642e2e88b93adc4ca272c644126a0dc7982b619cb68a55f41fba8d3979eebcb38451f5899c03a38ee05ebbc8a5b2c973abc11f0aa6ebee;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'habe97d844eee3b3b0b955fd8a1fdb942e01d145d14cd9ecdd32694cc653963a97793eb323c0ebb90f74d7d0db73acea72241972b749022f743f943841;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'habf025f622a1a8de125cff0097479bd470cd2e93c19dc4bda4fa203c67f7ccc8d041e6d2273edaa93f4ec567f46a3e4bbeb97a65f63837d87397521a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd1d2c0b19464382a348b056fa3644b23b81b94e67de7b29b0ec35c1462c741c20da465a827c2584c1dc64b9c28aa6ca405f5156ea716cea06ce3b8833;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h98639bd5994e426fb3edd67155f28a41100778e3f78735cf25925f7d0a632cb9f2f2f594ddd99be25954773a24082b4064a90f7741f52a71abcbf13c5;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf470625bb30139b6894e157c4ef475ae0508c43ede31b62750f1f8908fa03b669a0cf96e0d74bb6ee7a6d541ee4651f0f55a3373383b9fed20d1ab0cb;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he060afff93241092a1f1304e3ad3df44286a8e10ce53afd7779a458d9f4c160918ed101730f6ac834d6fbc6af36a308829abecfc1645dba552a7ad660;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5758a50f5af465ac30278fa6466d3c5d92366961dd3ad4df85db9c4a845c01ec38f085fdf92772a81d27ad48e66da2d95f648411a02ed81149becd99b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf0b7d0cc27dd53fc057da539f549d801cf978643071c63aeafd2b9dbf147b86b010b05967cc1bf330cf2404ec929d4eccf29119451284da7e9cb90182;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h527b58a56e4ef45f3b24dc78d3ff71ae02241ea57fd4fef74ac622f29174562e1fc65ebbfaa7b98587a39c07343de7c288f45e111a7808550e79d3b77;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h60ed5e45dd5e02f337b0026c1d347a69fb4f5502d38f7a5402b863375876a413cfc6fa13526776412b74cf044f7976e86602d7e567c0288b1a873b3c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb795f1c1c5167d5451e8eb9899863db9f466197d50c5661dfa37ebde528017b144ae5478e56b36d1fa701170ba87c903c447e240fb5113d062048c3c0;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9d251cf9aacc073c0d9995eae5c238d3292fb30f1da15fa177a087b781ac05980de8006c2724929b66ee86bc764298a01f26e1459e1a32518bbff16e7;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha07739a9776d444bd63e7b3bef88e29ae90099d9a88069f79fbc98aab68e5c19e2e46cde5ea4cbfa85e5a2d121d964db044453086bbcf4f69fa5c955f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd9da8e21e74149382e4d40403d5e1a93b40445d8d581bc083c35dbeece158ee935210c011d6f14c9b8a266c1fda76c822f2f5df0ba4e9ae1567225a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9878cbceb91d2e0d2663d9ce761f0dfa51ec6e94916f69ec84e11b67d48c30ae019389ca4fb3e4a70f82452d3997ca27d20cb55f7e31e9c0afe498407;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbdec99abada11f072e2d30b5690ecaf85576be6e3272e6cede76a430b8d27d0b885f98221d466690805dbdb01fe1fd8128e4fee8a9a0afa1eeaee9681;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha91a91d1454922303f0e1ab22e7bb4d7d55f5304b0e05e94940983e1929a4dfbdb93f904d4c0d3f9d55d105ed138aec40b58858a8ce88664ced685548;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h121d747358f2ee5991253ab8eac4593d0424220e5a88e8ddd0636eb629169a59a133f677ecfa023978b1588d0657188bd63c74c359b48a695cb02046;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hee297117f85451601796391f2fc8f42206b1165aea1d8e49fd41719b797f716d16cc88db578d926a650b4c0056152d57d6db705f2482d5843fffd5ab5;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8d951fd09c8cae5e9d3362bed9ba0558307c7397af1832b8f9e4d7e12a4a6fdc8c878e896154c6b7e70987df386567ac91ce4bfec5ccf01e16623bcdd;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h99c1affe10246daaefb95be5902e0a54061708833e6fbb2c8c41485e0e36e30e82857052c7ba9051d34b07a484cdf62e2b986f600f28ced8abcaec55a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he1f35ad3b4ed6eb5ee4673fec74c82b96cb9cbcfde363e2b9d7b2f2ffa044bd01c9df45fdad81f67cd83089e8e6e4e279c83a17ba4ecda715225249ad;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7131d6e34008b10971799b048173b10ceb7eca91581bbe7403706a0b42d46b87e2f34f9e32c379e39fc54351bf72932f46f09940e2c02870a56793a33;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7f62ace2361d81b9d783ba1038e15d7c963646de495762c471c9cfcaa78dd8327ff4288d7194ddc5211bc9fca261c8098603ff09c72b8f44c03207176;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he8fa9de1a819114804583203b75ed74a5ddb928844891bdbd102be23056e8946334694b527c1a7d621403b629174c48dcb80b06e2e677713f2269be91;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6cca776f406b236a84c2810d901fada674669f473452145bf445dcff9a1b0d639ebdb2d6ad66f33683251481ef049a170372fde4361c589479611cadd;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9681d3d6ec43fa7dd13531d14194936c9b941fabb92efa4acb1454376566b6310d5c34dd8eb2f29039413adfad7a37b9bd691aeb18ac39949e7bed963;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha4989347fff8801e1fa9b15e9ba4348c0690a67729384f70c5dca395b7cf07bc31f4b8423a5ca6d87ba0102665d818f39deb6086ce5e7e7d2b40148dd;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbed8fa9632810f3c34e9fdff5c594ab3c9d8030c7c4c40b960d72b7ea01b0ff466e999bd6c4448bc5173d008b7fbe7a3074ff9ed8f573331e1d0f3672;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h15bfb0f0e4eda7f756c51bd3ae37e50a9d22d45b9f0f054954ef121a663d1ea01fff83d90f16ed03d908ad2175448665431717b1cf7644cfcb38efa01;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9fd59f3b2ee3903d6638b6bc3fc576cb225119e6b6860c6b97a111bd1e03acac0256a998315b13b96107932b6b94cce2b4373810c07d123d08f049771;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hde1b821fb851be59e21e771a462a661f8cb3f10dc014b4533cb86e9054e785b6fca014615a208074ae888b710bc5d04451b0cd4199ef82589f978f676;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h16a1a2e419520c02d13be3958303e4ba1f3625200428cb22a8d716d80cbdd267f80488680860c54496ec594cc1bae3ea6fece64ce07b83bd623291da;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h541466a3b413249a2f2f0ad7a6abb4024b3d8c677bb7782a6b923ea7292a6fb179a3fd875b82fbdb21c7790f0a060c23fdb8f31134af31ee420513b01;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h18411005ebb13bbe45103091994b5e85d8b2b24a798507abad86bc950f3215b1113be8ef739225f1eac848604c31524c7b49d8ad7bbf9721014b23726;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8375b295d0d539f66664369e21ab354ae58b0d398092932322286bf559cae3bc1fa4efbbd4126e9c0ae138abd1fab5668c8dffd6715fea1de37738866;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb38ec72497497b6dbf95aa0975bc03461be30eb18a5def2c602d3b666d3588e45ee01a0008310f20294b1b68b0dbc15c7bfe1b41ac9ed72164565dd6f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc5d8306f92825fcb25cab0ab32e9102b50c5fdd04d9a7008acb2743de7ac84ebd17eaf7d8003e58672f2cd842a50f270b4d9a265db8627dd0dc838946;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h25be35345b49421f7079f56183d521dc2b3ba587e7adc9e52b95920b67ba32b9f4dcb56a6bd9326a97ff0b529cbda741c17cc7300eb8f01d1f81ea156;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd4df021cb89ff2a9c4f6bb0d2f1e1e230cb9de3e1d459b317195f790c7abaaaa5738d6b41e5a7b8e64ff34b22b57fa7c09834a8afc105adf41acf4c2f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h903ca065602423b8f295b9cf7f59a3d70237f08b2bd445ba01fdc54997920a5dec1abb3e5956872f2f09676a84aafb4cd853c48932fc55b4ea0885313;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd2941009096f61935b6c5084d1107d1a5e987e9c6fb92e1d95380ac6a9c123e2b9d18d0496bf8c081aab4d801f9f3b844c72cea02db7ce98c719e5f77;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf4e3da4501d8122a9349a1525bac1b787cd4dbbd974a146addb9ed77657511b90103da4fd1687dc0ff8f13dc30a86cef6e1af26d4d2a5a28199baed33;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h274687ed8672d15e2e4344482518100fa4f39bdd72cce0d13e5add1c3f496639b34befa806974cf2c540411f08f9fd1e42e033d0fb0df3340b3d74f5e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf656d02d51f47b213f934c6ad2162043419ecc3e525ab8ea476126b51706672c0d4f23f384fd4970411ac488e9fd740da8c26156672209304e52b7f06;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he741ced5967cd7513cb6a2b9bb03743c66d9ba96fd4a750b9929b8c04b93a430e66a8fdf232a6b9cbb1efc643e47f877979f055f2b173e6c8dce30f0a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h12c82a8ec42859d4471cfae1777252e82c09b3d4361f0e5e3297419ac74fcfb32c87288efc3d7b8647ea6618da39b192511355e628d43afe43f10b95b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6456f5aa4ad4f78ad3a37feb764d55f4a4bbcb2c2a323a81f817ee7151c12a047c998791cf38fd42cab919f6307e92ffb04ed28e7d25cdd5a2bd25fbe;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdefe984f6a9494d1d14ca07fe656e0dbb7e57884f3a84458141b77c407507cd687793702730a97d18dd3535d43ae37d59a4275dac6c1bde17d9dd60bd;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8fcf690390650c09dd291d99a587660d318b0702d6323112068443cf896219043feae4f8a679661e8dd1878f34ba0ec1cbc025d1249b5bc0361ada2c8;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbc6c8acd37a2a5f00396dadb49eb8e1df78a569016e94f944f88ef31e749d69030cbb2d2558c7d4b6ce0f1888392516b672b40e9dc46076a2b58d864a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h87c54d739b1e5a7d1d85916977673faea43f667f8a4fc2a894b3efbaa54a7591c16fdc6cff229c7fb0c9373e0d9a8d6d24c474bd20a0a8bb40f3277d7;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h35a6897767042aba8e7fc1d38351e6451f24c33d21a44e877fdf7016b80cd0cb7043b261f521764ff8fca0e176660c52db2eba961394dd179c45b7064;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'haf4efa24dccaf3e88317831f7f102af6a635ba7ab961d22a6e4429e9079b592afd3d1d870d91936ffa91636572c37cc4283560526fca545afadd1df50;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdcdaa49da092f15d0b87a23a5eb0a975d742ea3ceee52cf3becd7a8dc4fdc96eb0e417fdb152e9bd632d1eecd3b383f878655aa5d38baa729c1bac68e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'haeac2d5c25a6c0d03aee9cfa75bd584c412877cebd36e483df7d61a4607e927792d1f44eca9a0997d5809ae5a8957fac1537414f9a35f1f6bf3c72276;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4133ea42543c09eab5571115bec72f8d4a178c913c21ba5d05b16792061e47b538ea5e6b5640f95f564ebf29ca8ca357c1389ad9c6d837a2e16b8c47c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd6044780179f4ac51de02bcf82c5bd7139edafd8c483d0d11814a8ac191d7c4e555040c190aece4ec69f9c93b1ddc82064c508b3bf824fbb4944100e1;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd084997fd405481c6641c520e11857570ab004e6b5f2cd8b3171a845ab131586b4bce1b06a09046148c702630724eb21c9d9ef21b39e8f9e83bff446d;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9fd04d00744e59ea830b51192978ce3162b652f57e3d65597696be8d5ed158f7b98523dbe335fac87c5be19859a88aaedbe282fdfebe6180197d3cba8;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha8e9f19e48180a5ca562120408f70726323e1a8f1fe37180813e98838861f57ac89acd716191ef45e2458737f952e91455d2afe22c5e4ed1bc41df083;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2a42a80fe29a75d40e6afa154efeb74fbf5184e89c3a58034192436d99d1eca43723198fa33d85995b9ab89c3efd9db95f8acf269f5bcc8199928a3b2;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h967bec89514e1797b5160b3df6f775c5941f54978ec77ea2b38e7179770e39528208bb071813943f5862b4d0574dbceeade8f181e82e5974394204b1c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbc1149954f8147f5f3dde14d5ad590e7455785d78e670b4d6d18c4da69a2fda5ab7f398cad858afe12ac4441bbcb02758aff6a1d396a8302fe8390b5;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha14738e3efea66a0f9be94b84c230a935a54a635544721b9311b9cd78e151c2cce171de14fad59664e28124ca1d4a258d2fd0ecb764d572a43944bfd3;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h267c3cebc264f85339a75634f9a3820eb1efcfd91513e3c4ea3cd8928b8d87c0a468fb2cda33cd46fce52da8a42b0cb06e8ccb2e31b15cc02ea4e7e19;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h84547d525b23e9101d7dc014d9f7d57ddbe2e00dd9f6f786915a73d93a19bc358641ce3d2ad4c78f101b82e715129c67a83d7e30d7b800406919920ce;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4f828656bc4918c7026af0d310d67f142a26ccbdba04fb18282452b72d2562335ba7481c26870084ebf79ad7c8871ba8fd60e6253637fe76a44456d09;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbed0ffc09b0d7f845e2060621ed66007c418ee88b5c537dc52b778714dbe2f09b483e57603c5bf83808f91278fffea0ad80d2bd1de51aa5c0b0a53d81;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5ce6bf0e6ec4e5c386ea25ea3f69e206c96c0c5445ddbd2040a62128db3f2df7c1d03dfe5b8d1dc5c0961a956c370e8c9686787425a4dfa514d1a7ccb;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc3736aef775d57c4b74e5ab338fe03da01f871821457f8efb3b1e74acce19a5bcae494f85a23af59162a79abbe9f9969958c349035a9160b3c75b32d8;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h57a62ada0391700894063660ebda877665fac5c74b116641d99fb7c4f9ecc3e7aa6aba9885c10dfb1df632e8c8b988f7fc2c5d86444cbee8833fe84f2;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2283f4cc0fd2c78d9d037baa89924245177615e00f1129ecce8d459be3bf55c18e6854e575dab3834f3cd0dcf5b671b4926289fabc17a127ea34e4bf3;
        #1
        $finish();
    end
endmodule
