module shift_register(
        input wire clk,
        input wire src0_,
        input wire src1_,
        input wire src2_,
        input wire src3_,
        input wire src4_,
        input wire src5_,
        input wire src6_,
        input wire src7_,
        input wire src8_,
        input wire src9_,
        input wire src10_,
        input wire src11_,
        output wire [0:0] dst0,
        output wire [0:0] dst1,
        output wire [0:0] dst2,
        output wire [0:0] dst3,
        output wire [0:0] dst4,
        output wire [0:0] dst5,
        output wire [0:0] dst6,
        output wire [0:0] dst7,
        output wire [0:0] dst8,
        output wire [0:0] dst9,
        output wire [0:0] dst10,
        output wire [0:0] dst11,
        output wire [0:0] dst12,
        output wire [0:0] dst13,
        output wire [0:0] dst14,
        output wire [0:0] dst15,
        output wire [0:0] dst16,
        output wire [0:0] dst17);
    reg [63:0] src0;
    reg [63:0] src1;
    reg [63:0] src2;
    reg [63:0] src3;
    reg [63:0] src4;
    reg [63:0] src5;
    reg [63:0] src6;
    reg [63:0] src7;
    reg [63:0] src8;
    reg [63:0] src9;
    reg [63:0] src10;
    reg [63:0] src11;
    compressor2_1_64_12 compressor2_1_64_12(
            .src0(src0),
            .src1(src1),
            .src2(src2),
            .src3(src3),
            .src4(src4),
            .src5(src5),
            .src6(src6),
            .src7(src7),
            .src8(src8),
            .src9(src9),
            .src10(src10),
            .src11(src11),
            .dst0(dst0),
            .dst1(dst1),
            .dst2(dst2),
            .dst3(dst3),
            .dst4(dst4),
            .dst5(dst5),
            .dst6(dst6),
            .dst7(dst7),
            .dst8(dst8),
            .dst9(dst9),
            .dst10(dst10),
            .dst11(dst11),
            .dst12(dst12),
            .dst13(dst13),
            .dst14(dst14),
            .dst15(dst15),
            .dst16(dst16),
            .dst17(dst17));
    initial begin
        src0 <= 64'h0;
        src1 <= 64'h0;
        src2 <= 64'h0;
        src3 <= 64'h0;
        src4 <= 64'h0;
        src5 <= 64'h0;
        src6 <= 64'h0;
        src7 <= 64'h0;
        src8 <= 64'h0;
        src9 <= 64'h0;
        src10 <= 64'h0;
        src11 <= 64'h0;
    end
    always @(posedge clk) begin
        src0 <= {src0, src0_};
        src1 <= {src1, src1_};
        src2 <= {src2, src2_};
        src3 <= {src3, src3_};
        src4 <= {src4, src4_};
        src5 <= {src5, src5_};
        src6 <= {src6, src6_};
        src7 <= {src7, src7_};
        src8 <= {src8, src8_};
        src9 <= {src9, src9_};
        src10 <= {src10, src10_};
        src11 <= {src11, src11_};
    end
endmodule
module compressor2_1_64_12(
    input [63:0]src0,
    input [63:0]src1,
    input [63:0]src2,
    input [63:0]src3,
    input [63:0]src4,
    input [63:0]src5,
    input [63:0]src6,
    input [63:0]src7,
    input [63:0]src8,
    input [63:0]src9,
    input [63:0]src10,
    input [63:0]src11,
    output dst0,
    output dst1,
    output dst2,
    output dst3,
    output dst4,
    output dst5,
    output dst6,
    output dst7,
    output dst8,
    output dst9,
    output dst10,
    output dst11,
    output dst12,
    output dst13,
    output dst14,
    output dst15,
    output dst16,
    output dst17);

    wire [1:0] comp_out0;
    wire [1:0] comp_out1;
    wire [1:0] comp_out2;
    wire [1:0] comp_out3;
    wire [1:0] comp_out4;
    wire [1:0] comp_out5;
    wire [1:0] comp_out6;
    wire [1:0] comp_out7;
    wire [1:0] comp_out8;
    wire [1:0] comp_out9;
    wire [1:0] comp_out10;
    wire [1:0] comp_out11;
    wire [1:0] comp_out12;
    wire [1:0] comp_out13;
    wire [1:0] comp_out14;
    wire [1:0] comp_out15;
    wire [1:0] comp_out16;
    wire [0:0] comp_out17;
    compressor compressor_inst(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .dst0(comp_out0),
        .dst1(comp_out1),
        .dst2(comp_out2),
        .dst3(comp_out3),
        .dst4(comp_out4),
        .dst5(comp_out5),
        .dst6(comp_out6),
        .dst7(comp_out7),
        .dst8(comp_out8),
        .dst9(comp_out9),
        .dst10(comp_out10),
        .dst11(comp_out11),
        .dst12(comp_out12),
        .dst13(comp_out13),
        .dst14(comp_out14),
        .dst15(comp_out15),
        .dst16(comp_out16),
        .dst17(comp_out17)
    );
    rowadder2_1_18 rowadder2_1inst(
        .src0({comp_out17[0], comp_out16[0], comp_out15[0], comp_out14[0], comp_out13[0], comp_out12[0], comp_out11[0], comp_out10[0], comp_out9[0], comp_out8[0], comp_out7[0], comp_out6[0], comp_out5[0], comp_out4[0], comp_out3[0], comp_out2[0], comp_out1[0], comp_out0[0]}),
        .src1({1'h0, comp_out16[1], comp_out15[1], comp_out14[1], comp_out13[1], comp_out12[1], comp_out11[1], comp_out10[1], comp_out9[1], comp_out8[1], comp_out7[1], comp_out6[1], comp_out5[1], comp_out4[1], comp_out3[1], comp_out2[1], comp_out1[1], comp_out0[1]}),
        .dst0({dst17, dst16, dst15, dst14, dst13, dst12, dst11, dst10, dst9, dst8, dst7, dst6, dst5, dst4, dst3, dst2, dst1, dst0})
    );
endmodule
module compressor (
      input wire [63:0] src0,
      input wire [63:0] src1,
      input wire [63:0] src2,
      input wire [63:0] src3,
      input wire [63:0] src4,
      input wire [63:0] src5,
      input wire [63:0] src6,
      input wire [63:0] src7,
      input wire [63:0] src8,
      input wire [63:0] src9,
      input wire [63:0] src10,
      input wire [63:0] src11,
      output wire [1:0] dst0,
      output wire [1:0] dst1,
      output wire [1:0] dst2,
      output wire [1:0] dst3,
      output wire [1:0] dst4,
      output wire [1:0] dst5,
      output wire [1:0] dst6,
      output wire [1:0] dst7,
      output wire [1:0] dst8,
      output wire [1:0] dst9,
      output wire [1:0] dst10,
      output wire [1:0] dst11,
      output wire [1:0] dst12,
      output wire [1:0] dst13,
      output wire [1:0] dst14,
      output wire [1:0] dst15,
      output wire [1:0] dst16,
      output wire [0:0] dst17);

   wire [63:0] stage0_0;
   wire [63:0] stage0_1;
   wire [63:0] stage0_2;
   wire [63:0] stage0_3;
   wire [63:0] stage0_4;
   wire [63:0] stage0_5;
   wire [63:0] stage0_6;
   wire [63:0] stage0_7;
   wire [63:0] stage0_8;
   wire [63:0] stage0_9;
   wire [63:0] stage0_10;
   wire [63:0] stage0_11;
   wire [11:0] stage1_0;
   wire [19:0] stage1_1;
   wire [23:0] stage1_2;
   wire [24:0] stage1_3;
   wire [27:0] stage1_4;
   wire [30:0] stage1_5;
   wire [23:0] stage1_6;
   wire [21:0] stage1_7;
   wire [28:0] stage1_8;
   wire [30:0] stage1_9;
   wire [25:0] stage1_10;
   wire [21:0] stage1_11;
   wire [18:0] stage1_12;
   wire [11:0] stage1_13;
   wire [3:0] stage2_0;
   wire [4:0] stage2_1;
   wire [7:0] stage2_2;
   wire [9:0] stage2_3;
   wire [11:0] stage2_4;
   wire [11:0] stage2_5;
   wire [12:0] stage2_6;
   wire [9:0] stage2_7;
   wire [7:0] stage2_8;
   wire [11:0] stage2_9;
   wire [12:0] stage2_10;
   wire [10:0] stage2_11;
   wire [9:0] stage2_12;
   wire [5:0] stage2_13;
   wire [5:0] stage2_14;
   wire [1:0] stage2_15;
   wire [3:0] stage3_0;
   wire [4:0] stage3_1;
   wire [7:0] stage3_2;
   wire [1:0] stage3_3;
   wire [3:0] stage3_4;
   wire [3:0] stage3_5;
   wire [3:0] stage3_6;
   wire [5:0] stage3_7;
   wire [4:0] stage3_8;
   wire [2:0] stage3_9;
   wire [3:0] stage3_10;
   wire [5:0] stage3_11;
   wire [5:0] stage3_12;
   wire [2:0] stage3_13;
   wire [2:0] stage3_14;
   wire [3:0] stage3_15;
   wire [0:0] stage3_16;
   wire [1:0] stage4_0;
   wire [1:0] stage4_1;
   wire [1:0] stage4_2;
   wire [1:0] stage4_3;
   wire [1:0] stage4_4;
   wire [1:0] stage4_5;
   wire [1:0] stage4_6;
   wire [1:0] stage4_7;
   wire [1:0] stage4_8;
   wire [1:0] stage4_9;
   wire [1:0] stage4_10;
   wire [1:0] stage4_11;
   wire [1:0] stage4_12;
   wire [1:0] stage4_13;
   wire [1:0] stage4_14;
   wire [1:0] stage4_15;
   wire [1:0] stage4_16;
   wire [0:0] stage4_17;

   assign stage0_0 = src0;
   assign stage0_1 = src1;
   assign stage0_2 = src2;
   assign stage0_3 = src3;
   assign stage0_4 = src4;
   assign stage0_5 = src5;
   assign stage0_6 = src6;
   assign stage0_7 = src7;
   assign stage0_8 = src8;
   assign stage0_9 = src9;
   assign stage0_10 = src10;
   assign stage0_11 = src11;
   assign dst0 = stage4_0;
   assign dst1 = stage4_1;
   assign dst2 = stage4_2;
   assign dst3 = stage4_3;
   assign dst4 = stage4_4;
   assign dst5 = stage4_5;
   assign dst6 = stage4_6;
   assign dst7 = stage4_7;
   assign dst8 = stage4_8;
   assign dst9 = stage4_9;
   assign dst10 = stage4_10;
   assign dst11 = stage4_11;
   assign dst12 = stage4_12;
   assign dst13 = stage4_13;
   assign dst14 = stage4_14;
   assign dst15 = stage4_15;
   assign dst16 = stage4_16;
   assign dst17 = stage4_17;

   gpc135_4 gpc0 (
      {stage0_0[0], stage0_0[1], stage0_0[2], stage0_0[3], stage0_0[4]},
      {stage0_1[0], stage0_1[1], stage0_1[2]},
      {stage0_2[0]},
      {stage1_3[0],stage1_2[0],stage1_1[0],stage1_0[0]}
   );
   gpc117_4 gpc1 (
      {stage0_0[5], stage0_0[6], stage0_0[7], stage0_0[8], stage0_0[9], stage0_0[10], stage0_0[11]},
      {stage0_1[3]},
      {stage0_2[1]},
      {stage1_3[1],stage1_2[1],stage1_1[1],stage1_0[1]}
   );
   gpc117_4 gpc2 (
      {stage0_0[12], stage0_0[13], stage0_0[14], stage0_0[15], stage0_0[16], stage0_0[17], stage0_0[18]},
      {stage0_1[4]},
      {stage0_2[2]},
      {stage1_3[2],stage1_2[2],stage1_1[2],stage1_0[2]}
   );
   gpc117_4 gpc3 (
      {stage0_0[19], stage0_0[20], stage0_0[21], stage0_0[22], stage0_0[23], stage0_0[24], stage0_0[25]},
      {stage0_1[5]},
      {stage0_2[3]},
      {stage1_3[3],stage1_2[3],stage1_1[3],stage1_0[3]}
   );
   gpc117_4 gpc4 (
      {stage0_0[26], stage0_0[27], stage0_0[28], stage0_0[29], stage0_0[30], stage0_0[31], stage0_0[32]},
      {stage0_1[6]},
      {stage0_2[4]},
      {stage1_3[4],stage1_2[4],stage1_1[4],stage1_0[4]}
   );
   gpc615_5 gpc5 (
      {stage0_0[33], stage0_0[34], stage0_0[35], stage0_0[36], stage0_0[37]},
      {stage0_1[7]},
      {stage0_2[5], stage0_2[6], stage0_2[7], stage0_2[8], stage0_2[9], stage0_2[10]},
      {stage1_4[0],stage1_3[5],stage1_2[5],stage1_1[5],stage1_0[5]}
   );
   gpc615_5 gpc6 (
      {stage0_0[38], stage0_0[39], stage0_0[40], stage0_0[41], stage0_0[42]},
      {stage0_1[8]},
      {stage0_2[11], stage0_2[12], stage0_2[13], stage0_2[14], stage0_2[15], stage0_2[16]},
      {stage1_4[1],stage1_3[6],stage1_2[6],stage1_1[6],stage1_0[6]}
   );
   gpc615_5 gpc7 (
      {stage0_0[43], stage0_0[44], stage0_0[45], stage0_0[46], stage0_0[47]},
      {stage0_1[9]},
      {stage0_2[17], stage0_2[18], stage0_2[19], stage0_2[20], stage0_2[21], stage0_2[22]},
      {stage1_4[2],stage1_3[7],stage1_2[7],stage1_1[7],stage1_0[7]}
   );
   gpc615_5 gpc8 (
      {stage0_0[48], stage0_0[49], stage0_0[50], stage0_0[51], stage0_0[52]},
      {stage0_1[10]},
      {stage0_2[23], stage0_2[24], stage0_2[25], stage0_2[26], stage0_2[27], stage0_2[28]},
      {stage1_4[3],stage1_3[8],stage1_2[8],stage1_1[8],stage1_0[8]}
   );
   gpc615_5 gpc9 (
      {stage0_0[53], stage0_0[54], stage0_0[55], stage0_0[56], stage0_0[57]},
      {stage0_1[11]},
      {stage0_2[29], stage0_2[30], stage0_2[31], stage0_2[32], stage0_2[33], stage0_2[34]},
      {stage1_4[4],stage1_3[9],stage1_2[9],stage1_1[9],stage1_0[9]}
   );
   gpc615_5 gpc10 (
      {stage0_0[58], stage0_0[59], stage0_0[60], stage0_0[61], stage0_0[62]},
      {stage0_1[12]},
      {stage0_2[35], stage0_2[36], stage0_2[37], stage0_2[38], stage0_2[39], stage0_2[40]},
      {stage1_4[5],stage1_3[10],stage1_2[10],stage1_1[10],stage1_0[10]}
   );
   gpc606_5 gpc11 (
      {stage0_1[13], stage0_1[14], stage0_1[15], stage0_1[16], stage0_1[17], stage0_1[18]},
      {stage0_3[0], stage0_3[1], stage0_3[2], stage0_3[3], stage0_3[4], stage0_3[5]},
      {stage1_5[0],stage1_4[6],stage1_3[11],stage1_2[11],stage1_1[11]}
   );
   gpc606_5 gpc12 (
      {stage0_1[19], stage0_1[20], stage0_1[21], stage0_1[22], stage0_1[23], stage0_1[24]},
      {stage0_3[6], stage0_3[7], stage0_3[8], stage0_3[9], stage0_3[10], stage0_3[11]},
      {stage1_5[1],stage1_4[7],stage1_3[12],stage1_2[12],stage1_1[12]}
   );
   gpc606_5 gpc13 (
      {stage0_1[25], stage0_1[26], stage0_1[27], stage0_1[28], stage0_1[29], stage0_1[30]},
      {stage0_3[12], stage0_3[13], stage0_3[14], stage0_3[15], stage0_3[16], stage0_3[17]},
      {stage1_5[2],stage1_4[8],stage1_3[13],stage1_2[13],stage1_1[13]}
   );
   gpc606_5 gpc14 (
      {stage0_1[31], stage0_1[32], stage0_1[33], stage0_1[34], stage0_1[35], stage0_1[36]},
      {stage0_3[18], stage0_3[19], stage0_3[20], stage0_3[21], stage0_3[22], stage0_3[23]},
      {stage1_5[3],stage1_4[9],stage1_3[14],stage1_2[14],stage1_1[14]}
   );
   gpc606_5 gpc15 (
      {stage0_1[37], stage0_1[38], stage0_1[39], stage0_1[40], stage0_1[41], stage0_1[42]},
      {stage0_3[24], stage0_3[25], stage0_3[26], stage0_3[27], stage0_3[28], stage0_3[29]},
      {stage1_5[4],stage1_4[10],stage1_3[15],stage1_2[15],stage1_1[15]}
   );
   gpc606_5 gpc16 (
      {stage0_1[43], stage0_1[44], stage0_1[45], stage0_1[46], stage0_1[47], stage0_1[48]},
      {stage0_3[30], stage0_3[31], stage0_3[32], stage0_3[33], stage0_3[34], stage0_3[35]},
      {stage1_5[5],stage1_4[11],stage1_3[16],stage1_2[16],stage1_1[16]}
   );
   gpc615_5 gpc17 (
      {stage0_1[49], stage0_1[50], stage0_1[51], stage0_1[52], stage0_1[53]},
      {stage0_2[41]},
      {stage0_3[36], stage0_3[37], stage0_3[38], stage0_3[39], stage0_3[40], stage0_3[41]},
      {stage1_5[6],stage1_4[12],stage1_3[17],stage1_2[17],stage1_1[17]}
   );
   gpc615_5 gpc18 (
      {stage0_1[54], stage0_1[55], stage0_1[56], stage0_1[57], stage0_1[58]},
      {stage0_2[42]},
      {stage0_3[42], stage0_3[43], stage0_3[44], stage0_3[45], stage0_3[46], stage0_3[47]},
      {stage1_5[7],stage1_4[13],stage1_3[18],stage1_2[18],stage1_1[18]}
   );
   gpc615_5 gpc19 (
      {stage0_1[59], stage0_1[60], stage0_1[61], stage0_1[62], stage0_1[63]},
      {stage0_2[43]},
      {stage0_3[48], stage0_3[49], stage0_3[50], stage0_3[51], stage0_3[52], stage0_3[53]},
      {stage1_5[8],stage1_4[14],stage1_3[19],stage1_2[19],stage1_1[19]}
   );
   gpc615_5 gpc20 (
      {stage0_2[44], stage0_2[45], stage0_2[46], stage0_2[47], stage0_2[48]},
      {stage0_3[54]},
      {stage0_4[0], stage0_4[1], stage0_4[2], stage0_4[3], stage0_4[4], stage0_4[5]},
      {stage1_6[0],stage1_5[9],stage1_4[15],stage1_3[20],stage1_2[20]}
   );
   gpc615_5 gpc21 (
      {stage0_2[49], stage0_2[50], stage0_2[51], stage0_2[52], stage0_2[53]},
      {stage0_3[55]},
      {stage0_4[6], stage0_4[7], stage0_4[8], stage0_4[9], stage0_4[10], stage0_4[11]},
      {stage1_6[1],stage1_5[10],stage1_4[16],stage1_3[21],stage1_2[21]}
   );
   gpc615_5 gpc22 (
      {stage0_2[54], stage0_2[55], stage0_2[56], stage0_2[57], stage0_2[58]},
      {stage0_3[56]},
      {stage0_4[12], stage0_4[13], stage0_4[14], stage0_4[15], stage0_4[16], stage0_4[17]},
      {stage1_6[2],stage1_5[11],stage1_4[17],stage1_3[22],stage1_2[22]}
   );
   gpc615_5 gpc23 (
      {stage0_2[59], stage0_2[60], stage0_2[61], stage0_2[62], stage0_2[63]},
      {stage0_3[57]},
      {stage0_4[18], stage0_4[19], stage0_4[20], stage0_4[21], stage0_4[22], stage0_4[23]},
      {stage1_6[3],stage1_5[12],stage1_4[18],stage1_3[23],stage1_2[23]}
   );
   gpc606_5 gpc24 (
      {stage0_3[58], stage0_3[59], stage0_3[60], stage0_3[61], stage0_3[62], stage0_3[63]},
      {stage0_5[0], stage0_5[1], stage0_5[2], stage0_5[3], stage0_5[4], stage0_5[5]},
      {stage1_7[0],stage1_6[4],stage1_5[13],stage1_4[19],stage1_3[24]}
   );
   gpc615_5 gpc25 (
      {stage0_4[24], stage0_4[25], stage0_4[26], stage0_4[27], stage0_4[28]},
      {stage0_5[6]},
      {stage0_6[0], stage0_6[1], stage0_6[2], stage0_6[3], stage0_6[4], stage0_6[5]},
      {stage1_8[0],stage1_7[1],stage1_6[5],stage1_5[14],stage1_4[20]}
   );
   gpc615_5 gpc26 (
      {stage0_4[29], stage0_4[30], stage0_4[31], stage0_4[32], stage0_4[33]},
      {stage0_5[7]},
      {stage0_6[6], stage0_6[7], stage0_6[8], stage0_6[9], stage0_6[10], stage0_6[11]},
      {stage1_8[1],stage1_7[2],stage1_6[6],stage1_5[15],stage1_4[21]}
   );
   gpc615_5 gpc27 (
      {stage0_4[34], stage0_4[35], stage0_4[36], stage0_4[37], stage0_4[38]},
      {stage0_5[8]},
      {stage0_6[12], stage0_6[13], stage0_6[14], stage0_6[15], stage0_6[16], stage0_6[17]},
      {stage1_8[2],stage1_7[3],stage1_6[7],stage1_5[16],stage1_4[22]}
   );
   gpc615_5 gpc28 (
      {stage0_4[39], stage0_4[40], stage0_4[41], stage0_4[42], stage0_4[43]},
      {stage0_5[9]},
      {stage0_6[18], stage0_6[19], stage0_6[20], stage0_6[21], stage0_6[22], stage0_6[23]},
      {stage1_8[3],stage1_7[4],stage1_6[8],stage1_5[17],stage1_4[23]}
   );
   gpc615_5 gpc29 (
      {stage0_4[44], stage0_4[45], stage0_4[46], stage0_4[47], stage0_4[48]},
      {stage0_5[10]},
      {stage0_6[24], stage0_6[25], stage0_6[26], stage0_6[27], stage0_6[28], stage0_6[29]},
      {stage1_8[4],stage1_7[5],stage1_6[9],stage1_5[18],stage1_4[24]}
   );
   gpc615_5 gpc30 (
      {stage0_4[49], stage0_4[50], stage0_4[51], stage0_4[52], stage0_4[53]},
      {stage0_5[11]},
      {stage0_6[30], stage0_6[31], stage0_6[32], stage0_6[33], stage0_6[34], stage0_6[35]},
      {stage1_8[5],stage1_7[6],stage1_6[10],stage1_5[19],stage1_4[25]}
   );
   gpc615_5 gpc31 (
      {stage0_4[54], stage0_4[55], stage0_4[56], stage0_4[57], stage0_4[58]},
      {stage0_5[12]},
      {stage0_6[36], stage0_6[37], stage0_6[38], stage0_6[39], stage0_6[40], stage0_6[41]},
      {stage1_8[6],stage1_7[7],stage1_6[11],stage1_5[20],stage1_4[26]}
   );
   gpc615_5 gpc32 (
      {stage0_4[59], stage0_4[60], stage0_4[61], stage0_4[62], stage0_4[63]},
      {stage0_5[13]},
      {stage0_6[42], stage0_6[43], stage0_6[44], stage0_6[45], stage0_6[46], stage0_6[47]},
      {stage1_8[7],stage1_7[8],stage1_6[12],stage1_5[21],stage1_4[27]}
   );
   gpc606_5 gpc33 (
      {stage0_5[14], stage0_5[15], stage0_5[16], stage0_5[17], stage0_5[18], stage0_5[19]},
      {stage0_7[0], stage0_7[1], stage0_7[2], stage0_7[3], stage0_7[4], stage0_7[5]},
      {stage1_9[0],stage1_8[8],stage1_7[9],stage1_6[13],stage1_5[22]}
   );
   gpc606_5 gpc34 (
      {stage0_5[20], stage0_5[21], stage0_5[22], stage0_5[23], stage0_5[24], stage0_5[25]},
      {stage0_7[6], stage0_7[7], stage0_7[8], stage0_7[9], stage0_7[10], stage0_7[11]},
      {stage1_9[1],stage1_8[9],stage1_7[10],stage1_6[14],stage1_5[23]}
   );
   gpc606_5 gpc35 (
      {stage0_5[26], stage0_5[27], stage0_5[28], stage0_5[29], stage0_5[30], stage0_5[31]},
      {stage0_7[12], stage0_7[13], stage0_7[14], stage0_7[15], stage0_7[16], stage0_7[17]},
      {stage1_9[2],stage1_8[10],stage1_7[11],stage1_6[15],stage1_5[24]}
   );
   gpc606_5 gpc36 (
      {stage0_5[32], stage0_5[33], stage0_5[34], stage0_5[35], stage0_5[36], stage0_5[37]},
      {stage0_7[18], stage0_7[19], stage0_7[20], stage0_7[21], stage0_7[22], stage0_7[23]},
      {stage1_9[3],stage1_8[11],stage1_7[12],stage1_6[16],stage1_5[25]}
   );
   gpc606_5 gpc37 (
      {stage0_5[38], stage0_5[39], stage0_5[40], stage0_5[41], stage0_5[42], stage0_5[43]},
      {stage0_7[24], stage0_7[25], stage0_7[26], stage0_7[27], stage0_7[28], stage0_7[29]},
      {stage1_9[4],stage1_8[12],stage1_7[13],stage1_6[17],stage1_5[26]}
   );
   gpc615_5 gpc38 (
      {stage0_5[44], stage0_5[45], stage0_5[46], stage0_5[47], stage0_5[48]},
      {stage0_6[48]},
      {stage0_7[30], stage0_7[31], stage0_7[32], stage0_7[33], stage0_7[34], stage0_7[35]},
      {stage1_9[5],stage1_8[13],stage1_7[14],stage1_6[18],stage1_5[27]}
   );
   gpc615_5 gpc39 (
      {stage0_5[49], stage0_5[50], stage0_5[51], stage0_5[52], stage0_5[53]},
      {stage0_6[49]},
      {stage0_7[36], stage0_7[37], stage0_7[38], stage0_7[39], stage0_7[40], stage0_7[41]},
      {stage1_9[6],stage1_8[14],stage1_7[15],stage1_6[19],stage1_5[28]}
   );
   gpc615_5 gpc40 (
      {stage0_5[54], stage0_5[55], stage0_5[56], stage0_5[57], stage0_5[58]},
      {stage0_6[50]},
      {stage0_7[42], stage0_7[43], stage0_7[44], stage0_7[45], stage0_7[46], stage0_7[47]},
      {stage1_9[7],stage1_8[15],stage1_7[16],stage1_6[20],stage1_5[29]}
   );
   gpc615_5 gpc41 (
      {stage0_5[59], stage0_5[60], stage0_5[61], stage0_5[62], stage0_5[63]},
      {stage0_6[51]},
      {stage0_7[48], stage0_7[49], stage0_7[50], stage0_7[51], stage0_7[52], stage0_7[53]},
      {stage1_9[8],stage1_8[16],stage1_7[17],stage1_6[21],stage1_5[30]}
   );
   gpc606_5 gpc42 (
      {stage0_6[52], stage0_6[53], stage0_6[54], stage0_6[55], stage0_6[56], stage0_6[57]},
      {stage0_8[0], stage0_8[1], stage0_8[2], stage0_8[3], stage0_8[4], stage0_8[5]},
      {stage1_10[0],stage1_9[9],stage1_8[17],stage1_7[18],stage1_6[22]}
   );
   gpc606_5 gpc43 (
      {stage0_6[58], stage0_6[59], stage0_6[60], stage0_6[61], stage0_6[62], stage0_6[63]},
      {stage0_8[6], stage0_8[7], stage0_8[8], stage0_8[9], stage0_8[10], stage0_8[11]},
      {stage1_10[1],stage1_9[10],stage1_8[18],stage1_7[19],stage1_6[23]}
   );
   gpc2135_5 gpc44 (
      {stage0_7[54], stage0_7[55], stage0_7[56], stage0_7[57], stage0_7[58]},
      {stage0_8[12], stage0_8[13], stage0_8[14]},
      {stage0_9[0]},
      {stage0_10[0], stage0_10[1]},
      {stage1_11[0],stage1_10[2],stage1_9[11],stage1_8[19],stage1_7[20]}
   );
   gpc615_5 gpc45 (
      {stage0_7[59], stage0_7[60], stage0_7[61], stage0_7[62], stage0_7[63]},
      {stage0_8[15]},
      {stage0_9[1], stage0_9[2], stage0_9[3], stage0_9[4], stage0_9[5], stage0_9[6]},
      {stage1_11[1],stage1_10[3],stage1_9[12],stage1_8[20],stage1_7[21]}
   );
   gpc207_4 gpc46 (
      {stage0_8[16], stage0_8[17], stage0_8[18], stage0_8[19], stage0_8[20], stage0_8[21], stage0_8[22]},
      {stage0_10[2], stage0_10[3]},
      {stage1_11[2],stage1_10[4],stage1_9[13],stage1_8[21]}
   );
   gpc606_5 gpc47 (
      {stage0_8[23], stage0_8[24], stage0_8[25], stage0_8[26], stage0_8[27], stage0_8[28]},
      {stage0_10[4], stage0_10[5], stage0_10[6], stage0_10[7], stage0_10[8], stage0_10[9]},
      {stage1_12[0],stage1_11[3],stage1_10[5],stage1_9[14],stage1_8[22]}
   );
   gpc606_5 gpc48 (
      {stage0_8[29], stage0_8[30], stage0_8[31], stage0_8[32], stage0_8[33], stage0_8[34]},
      {stage0_10[10], stage0_10[11], stage0_10[12], stage0_10[13], stage0_10[14], stage0_10[15]},
      {stage1_12[1],stage1_11[4],stage1_10[6],stage1_9[15],stage1_8[23]}
   );
   gpc606_5 gpc49 (
      {stage0_8[35], stage0_8[36], stage0_8[37], stage0_8[38], stage0_8[39], stage0_8[40]},
      {stage0_10[16], stage0_10[17], stage0_10[18], stage0_10[19], stage0_10[20], stage0_10[21]},
      {stage1_12[2],stage1_11[5],stage1_10[7],stage1_9[16],stage1_8[24]}
   );
   gpc606_5 gpc50 (
      {stage0_8[41], stage0_8[42], stage0_8[43], stage0_8[44], stage0_8[45], stage0_8[46]},
      {stage0_10[22], stage0_10[23], stage0_10[24], stage0_10[25], stage0_10[26], stage0_10[27]},
      {stage1_12[3],stage1_11[6],stage1_10[8],stage1_9[17],stage1_8[25]}
   );
   gpc606_5 gpc51 (
      {stage0_8[47], stage0_8[48], stage0_8[49], stage0_8[50], stage0_8[51], stage0_8[52]},
      {stage0_10[28], stage0_10[29], stage0_10[30], stage0_10[31], stage0_10[32], stage0_10[33]},
      {stage1_12[4],stage1_11[7],stage1_10[9],stage1_9[18],stage1_8[26]}
   );
   gpc606_5 gpc52 (
      {stage0_8[53], stage0_8[54], stage0_8[55], stage0_8[56], stage0_8[57], stage0_8[58]},
      {stage0_10[34], stage0_10[35], stage0_10[36], stage0_10[37], stage0_10[38], stage0_10[39]},
      {stage1_12[5],stage1_11[8],stage1_10[10],stage1_9[19],stage1_8[27]}
   );
   gpc615_5 gpc53 (
      {stage0_8[59], stage0_8[60], stage0_8[61], stage0_8[62], stage0_8[63]},
      {stage0_9[7]},
      {stage0_10[40], stage0_10[41], stage0_10[42], stage0_10[43], stage0_10[44], stage0_10[45]},
      {stage1_12[6],stage1_11[9],stage1_10[11],stage1_9[20],stage1_8[28]}
   );
   gpc606_5 gpc54 (
      {stage0_9[8], stage0_9[9], stage0_9[10], stage0_9[11], stage0_9[12], stage0_9[13]},
      {stage0_11[0], stage0_11[1], stage0_11[2], stage0_11[3], stage0_11[4], stage0_11[5]},
      {stage1_13[0],stage1_12[7],stage1_11[10],stage1_10[12],stage1_9[21]}
   );
   gpc606_5 gpc55 (
      {stage0_9[14], stage0_9[15], stage0_9[16], stage0_9[17], stage0_9[18], stage0_9[19]},
      {stage0_11[6], stage0_11[7], stage0_11[8], stage0_11[9], stage0_11[10], stage0_11[11]},
      {stage1_13[1],stage1_12[8],stage1_11[11],stage1_10[13],stage1_9[22]}
   );
   gpc606_5 gpc56 (
      {stage0_9[20], stage0_9[21], stage0_9[22], stage0_9[23], stage0_9[24], stage0_9[25]},
      {stage0_11[12], stage0_11[13], stage0_11[14], stage0_11[15], stage0_11[16], stage0_11[17]},
      {stage1_13[2],stage1_12[9],stage1_11[12],stage1_10[14],stage1_9[23]}
   );
   gpc606_5 gpc57 (
      {stage0_9[26], stage0_9[27], stage0_9[28], stage0_9[29], stage0_9[30], stage0_9[31]},
      {stage0_11[18], stage0_11[19], stage0_11[20], stage0_11[21], stage0_11[22], stage0_11[23]},
      {stage1_13[3],stage1_12[10],stage1_11[13],stage1_10[15],stage1_9[24]}
   );
   gpc606_5 gpc58 (
      {stage0_9[32], stage0_9[33], stage0_9[34], stage0_9[35], stage0_9[36], stage0_9[37]},
      {stage0_11[24], stage0_11[25], stage0_11[26], stage0_11[27], stage0_11[28], stage0_11[29]},
      {stage1_13[4],stage1_12[11],stage1_11[14],stage1_10[16],stage1_9[25]}
   );
   gpc606_5 gpc59 (
      {stage0_9[38], stage0_9[39], stage0_9[40], stage0_9[41], stage0_9[42], stage0_9[43]},
      {stage0_11[30], stage0_11[31], stage0_11[32], stage0_11[33], stage0_11[34], stage0_11[35]},
      {stage1_13[5],stage1_12[12],stage1_11[15],stage1_10[17],stage1_9[26]}
   );
   gpc615_5 gpc60 (
      {stage0_9[44], stage0_9[45], stage0_9[46], stage0_9[47], stage0_9[48]},
      {stage0_10[46]},
      {stage0_11[36], stage0_11[37], stage0_11[38], stage0_11[39], stage0_11[40], stage0_11[41]},
      {stage1_13[6],stage1_12[13],stage1_11[16],stage1_10[18],stage1_9[27]}
   );
   gpc615_5 gpc61 (
      {stage0_9[49], stage0_9[50], stage0_9[51], stage0_9[52], stage0_9[53]},
      {stage0_10[47]},
      {stage0_11[42], stage0_11[43], stage0_11[44], stage0_11[45], stage0_11[46], stage0_11[47]},
      {stage1_13[7],stage1_12[14],stage1_11[17],stage1_10[19],stage1_9[28]}
   );
   gpc615_5 gpc62 (
      {stage0_9[54], stage0_9[55], stage0_9[56], stage0_9[57], stage0_9[58]},
      {stage0_10[48]},
      {stage0_11[48], stage0_11[49], stage0_11[50], stage0_11[51], stage0_11[52], stage0_11[53]},
      {stage1_13[8],stage1_12[15],stage1_11[18],stage1_10[20],stage1_9[29]}
   );
   gpc615_5 gpc63 (
      {stage0_9[59], stage0_9[60], stage0_9[61], stage0_9[62], stage0_9[63]},
      {stage0_10[49]},
      {stage0_11[54], stage0_11[55], stage0_11[56], stage0_11[57], stage0_11[58], stage0_11[59]},
      {stage1_13[9],stage1_12[16],stage1_11[19],stage1_10[21],stage1_9[30]}
   );
   gpc135_4 gpc64 (
      {stage0_10[50], stage0_10[51], stage0_10[52], stage0_10[53], stage0_10[54]},
      {stage0_11[60], stage0_11[61], stage0_11[62]},
      {1'b0},
      {stage1_13[10],stage1_12[17],stage1_11[20],stage1_10[22]}
   );
   gpc117_4 gpc65 (
      {stage0_10[55], stage0_10[56], stage0_10[57], stage0_10[58], stage0_10[59], stage0_10[60], stage0_10[61]},
      {stage0_11[63]},
      {1'b0},
      {stage1_13[11],stage1_12[18],stage1_11[21],stage1_10[23]}
   );
   gpc1_1 gpc66 (
      {stage0_0[63]},
      {stage1_0[11]}
   );
   gpc1_1 gpc67 (
      {stage0_10[62]},
      {stage1_10[24]}
   );
   gpc1_1 gpc68 (
      {stage0_10[63]},
      {stage1_10[25]}
   );
   gpc2135_5 gpc69 (
      {stage1_0[0], stage1_0[1], stage1_0[2], stage1_0[3], stage1_0[4]},
      {stage1_1[0], stage1_1[1], stage1_1[2]},
      {stage1_2[0]},
      {stage1_3[0], stage1_3[1]},
      {stage2_4[0],stage2_3[0],stage2_2[0],stage2_1[0],stage2_0[0]}
   );
   gpc615_5 gpc70 (
      {stage1_0[5], stage1_0[6], stage1_0[7], stage1_0[8], stage1_0[9]},
      {stage1_1[3]},
      {stage1_2[1], stage1_2[2], stage1_2[3], stage1_2[4], stage1_2[5], stage1_2[6]},
      {stage2_4[1],stage2_3[1],stage2_2[1],stage2_1[1],stage2_0[1]}
   );
   gpc2135_5 gpc71 (
      {stage1_1[4], stage1_1[5], stage1_1[6], stage1_1[7], stage1_1[8]},
      {stage1_2[7], stage1_2[8], stage1_2[9]},
      {stage1_3[2]},
      {stage1_4[0], stage1_4[1]},
      {stage2_5[0],stage2_4[2],stage2_3[2],stage2_2[2],stage2_1[2]}
   );
   gpc2135_5 gpc72 (
      {stage1_1[9], stage1_1[10], stage1_1[11], stage1_1[12], stage1_1[13]},
      {stage1_2[10], stage1_2[11], stage1_2[12]},
      {stage1_3[3]},
      {stage1_4[2], stage1_4[3]},
      {stage2_5[1],stage2_4[3],stage2_3[3],stage2_2[3],stage2_1[3]}
   );
   gpc1406_5 gpc73 (
      {stage1_1[14], stage1_1[15], stage1_1[16], stage1_1[17], stage1_1[18], stage1_1[19]},
      {stage1_3[4], stage1_3[5], stage1_3[6], stage1_3[7]},
      {stage1_4[4]},
      {stage2_5[2],stage2_4[4],stage2_3[4],stage2_2[4],stage2_1[4]}
   );
   gpc615_5 gpc74 (
      {stage1_2[13], stage1_2[14], stage1_2[15], stage1_2[16], stage1_2[17]},
      {stage1_3[8]},
      {stage1_4[5], stage1_4[6], stage1_4[7], stage1_4[8], stage1_4[9], stage1_4[10]},
      {stage2_6[0],stage2_5[3],stage2_4[5],stage2_3[5],stage2_2[5]}
   );
   gpc615_5 gpc75 (
      {stage1_2[18], stage1_2[19], stage1_2[20], stage1_2[21], stage1_2[22]},
      {stage1_3[9]},
      {stage1_4[11], stage1_4[12], stage1_4[13], stage1_4[14], stage1_4[15], stage1_4[16]},
      {stage2_6[1],stage2_5[4],stage2_4[6],stage2_3[6],stage2_2[6]}
   );
   gpc615_5 gpc76 (
      {stage1_3[10], stage1_3[11], stage1_3[12], stage1_3[13], stage1_3[14]},
      {stage1_4[17]},
      {stage1_5[0], stage1_5[1], stage1_5[2], stage1_5[3], stage1_5[4], stage1_5[5]},
      {stage2_7[0],stage2_6[2],stage2_5[5],stage2_4[7],stage2_3[7]}
   );
   gpc615_5 gpc77 (
      {stage1_3[15], stage1_3[16], stage1_3[17], stage1_3[18], stage1_3[19]},
      {stage1_4[18]},
      {stage1_5[6], stage1_5[7], stage1_5[8], stage1_5[9], stage1_5[10], stage1_5[11]},
      {stage2_7[1],stage2_6[3],stage2_5[6],stage2_4[8],stage2_3[8]}
   );
   gpc615_5 gpc78 (
      {stage1_3[20], stage1_3[21], stage1_3[22], stage1_3[23], stage1_3[24]},
      {stage1_4[19]},
      {stage1_5[12], stage1_5[13], stage1_5[14], stage1_5[15], stage1_5[16], stage1_5[17]},
      {stage2_7[2],stage2_6[4],stage2_5[7],stage2_4[9],stage2_3[9]}
   );
   gpc7_3 gpc79 (
      {stage1_4[20], stage1_4[21], stage1_4[22], stage1_4[23], stage1_4[24], stage1_4[25], stage1_4[26]},
      {stage2_6[5],stage2_5[8],stage2_4[10]}
   );
   gpc615_5 gpc80 (
      {stage1_5[18], stage1_5[19], stage1_5[20], stage1_5[21], stage1_5[22]},
      {stage1_6[0]},
      {stage1_7[0], stage1_7[1], stage1_7[2], stage1_7[3], stage1_7[4], stage1_7[5]},
      {stage2_9[0],stage2_8[0],stage2_7[3],stage2_6[6],stage2_5[9]}
   );
   gpc615_5 gpc81 (
      {stage1_5[23], stage1_5[24], stage1_5[25], stage1_5[26], stage1_5[27]},
      {stage1_6[1]},
      {stage1_7[6], stage1_7[7], stage1_7[8], stage1_7[9], stage1_7[10], stage1_7[11]},
      {stage2_9[1],stage2_8[1],stage2_7[4],stage2_6[7],stage2_5[10]}
   );
   gpc623_5 gpc82 (
      {stage1_5[28], stage1_5[29], stage1_5[30]},
      {stage1_6[2], stage1_6[3]},
      {stage1_7[12], stage1_7[13], stage1_7[14], stage1_7[15], stage1_7[16], stage1_7[17]},
      {stage2_9[2],stage2_8[2],stage2_7[5],stage2_6[8],stage2_5[11]}
   );
   gpc615_5 gpc83 (
      {stage1_6[4], stage1_6[5], stage1_6[6], stage1_6[7], stage1_6[8]},
      {stage1_7[18]},
      {stage1_8[0], stage1_8[1], stage1_8[2], stage1_8[3], stage1_8[4], stage1_8[5]},
      {stage2_10[0],stage2_9[3],stage2_8[3],stage2_7[6],stage2_6[9]}
   );
   gpc615_5 gpc84 (
      {stage1_6[9], stage1_6[10], stage1_6[11], stage1_6[12], stage1_6[13]},
      {stage1_7[19]},
      {stage1_8[6], stage1_8[7], stage1_8[8], stage1_8[9], stage1_8[10], stage1_8[11]},
      {stage2_10[1],stage2_9[4],stage2_8[4],stage2_7[7],stage2_6[10]}
   );
   gpc615_5 gpc85 (
      {stage1_6[14], stage1_6[15], stage1_6[16], stage1_6[17], stage1_6[18]},
      {stage1_7[20]},
      {stage1_8[12], stage1_8[13], stage1_8[14], stage1_8[15], stage1_8[16], stage1_8[17]},
      {stage2_10[2],stage2_9[5],stage2_8[5],stage2_7[8],stage2_6[11]}
   );
   gpc615_5 gpc86 (
      {stage1_6[19], stage1_6[20], stage1_6[21], stage1_6[22], stage1_6[23]},
      {stage1_7[21]},
      {stage1_8[18], stage1_8[19], stage1_8[20], stage1_8[21], stage1_8[22], stage1_8[23]},
      {stage2_10[3],stage2_9[6],stage2_8[6],stage2_7[9],stage2_6[12]}
   );
   gpc135_4 gpc87 (
      {stage1_8[24], stage1_8[25], stage1_8[26], stage1_8[27], stage1_8[28]},
      {stage1_9[0], stage1_9[1], stage1_9[2]},
      {stage1_10[0]},
      {stage2_11[0],stage2_10[4],stage2_9[7],stage2_8[7]}
   );
   gpc117_4 gpc88 (
      {stage1_9[3], stage1_9[4], stage1_9[5], stage1_9[6], stage1_9[7], stage1_9[8], stage1_9[9]},
      {stage1_10[1]},
      {stage1_11[0]},
      {stage2_12[0],stage2_11[1],stage2_10[5],stage2_9[8]}
   );
   gpc117_4 gpc89 (
      {stage1_9[10], stage1_9[11], stage1_9[12], stage1_9[13], stage1_9[14], stage1_9[15], stage1_9[16]},
      {stage1_10[2]},
      {stage1_11[1]},
      {stage2_12[1],stage2_11[2],stage2_10[6],stage2_9[9]}
   );
   gpc117_4 gpc90 (
      {stage1_9[17], stage1_9[18], stage1_9[19], stage1_9[20], stage1_9[21], stage1_9[22], stage1_9[23]},
      {stage1_10[3]},
      {stage1_11[2]},
      {stage2_12[2],stage2_11[3],stage2_10[7],stage2_9[10]}
   );
   gpc117_4 gpc91 (
      {stage1_9[24], stage1_9[25], stage1_9[26], stage1_9[27], stage1_9[28], stage1_9[29], stage1_9[30]},
      {stage1_10[4]},
      {stage1_11[3]},
      {stage2_12[3],stage2_11[4],stage2_10[8],stage2_9[11]}
   );
   gpc1163_5 gpc92 (
      {stage1_10[5], stage1_10[6], stage1_10[7]},
      {stage1_11[4], stage1_11[5], stage1_11[6], stage1_11[7], stage1_11[8], stage1_11[9]},
      {stage1_12[0]},
      {stage1_13[0]},
      {stage2_14[0],stage2_13[0],stage2_12[4],stage2_11[5],stage2_10[9]}
   );
   gpc606_5 gpc93 (
      {stage1_10[8], stage1_10[9], stage1_10[10], stage1_10[11], stage1_10[12], stage1_10[13]},
      {stage1_12[1], stage1_12[2], stage1_12[3], stage1_12[4], stage1_12[5], stage1_12[6]},
      {stage2_14[1],stage2_13[1],stage2_12[5],stage2_11[6],stage2_10[10]}
   );
   gpc606_5 gpc94 (
      {stage1_10[14], stage1_10[15], stage1_10[16], stage1_10[17], stage1_10[18], stage1_10[19]},
      {stage1_12[7], stage1_12[8], stage1_12[9], stage1_12[10], stage1_12[11], stage1_12[12]},
      {stage2_14[2],stage2_13[2],stage2_12[6],stage2_11[7],stage2_10[11]}
   );
   gpc606_5 gpc95 (
      {stage1_10[20], stage1_10[21], stage1_10[22], stage1_10[23], stage1_10[24], stage1_10[25]},
      {stage1_12[13], stage1_12[14], stage1_12[15], stage1_12[16], stage1_12[17], stage1_12[18]},
      {stage2_14[3],stage2_13[3],stage2_12[7],stage2_11[8],stage2_10[12]}
   );
   gpc606_5 gpc96 (
      {stage1_11[10], stage1_11[11], stage1_11[12], stage1_11[13], stage1_11[14], stage1_11[15]},
      {stage1_13[1], stage1_13[2], stage1_13[3], stage1_13[4], stage1_13[5], stage1_13[6]},
      {stage2_15[0],stage2_14[4],stage2_13[4],stage2_12[8],stage2_11[9]}
   );
   gpc606_5 gpc97 (
      {stage1_11[16], stage1_11[17], stage1_11[18], stage1_11[19], stage1_11[20], stage1_11[21]},
      {stage1_13[7], stage1_13[8], stage1_13[9], stage1_13[10], stage1_13[11], 1'b0},
      {stage2_15[1],stage2_14[5],stage2_13[5],stage2_12[9],stage2_11[10]}
   );
   gpc1_1 gpc98 (
      {stage1_0[10]},
      {stage2_0[2]}
   );
   gpc1_1 gpc99 (
      {stage1_0[11]},
      {stage2_0[3]}
   );
   gpc1_1 gpc100 (
      {stage1_2[23]},
      {stage2_2[7]}
   );
   gpc1_1 gpc101 (
      {stage1_4[27]},
      {stage2_4[11]}
   );
   gpc1415_5 gpc102 (
      {stage2_3[0], stage2_3[1], stage2_3[2], stage2_3[3], stage2_3[4]},
      {stage2_4[0]},
      {stage2_5[0], stage2_5[1], stage2_5[2], stage2_5[3]},
      {stage2_6[0]},
      {stage3_7[0],stage3_6[0],stage3_5[0],stage3_4[0],stage3_3[0]}
   );
   gpc615_5 gpc103 (
      {stage2_3[5], stage2_3[6], stage2_3[7], stage2_3[8], stage2_3[9]},
      {stage2_4[1]},
      {stage2_5[4], stage2_5[5], stage2_5[6], stage2_5[7], stage2_5[8], stage2_5[9]},
      {stage3_7[1],stage3_6[1],stage3_5[1],stage3_4[1],stage3_3[1]}
   );
   gpc615_5 gpc104 (
      {stage2_4[2], stage2_4[3], stage2_4[4], stage2_4[5], stage2_4[6]},
      {stage2_5[10]},
      {stage2_6[1], stage2_6[2], stage2_6[3], stage2_6[4], stage2_6[5], stage2_6[6]},
      {stage3_8[0],stage3_7[2],stage3_6[2],stage3_5[2],stage3_4[2]}
   );
   gpc615_5 gpc105 (
      {stage2_4[7], stage2_4[8], stage2_4[9], stage2_4[10], stage2_4[11]},
      {stage2_5[11]},
      {stage2_6[7], stage2_6[8], stage2_6[9], stage2_6[10], stage2_6[11], stage2_6[12]},
      {stage3_8[1],stage3_7[3],stage3_6[3],stage3_5[3],stage3_4[3]}
   );
   gpc615_5 gpc106 (
      {stage2_7[0], stage2_7[1], stage2_7[2], stage2_7[3], stage2_7[4]},
      {stage2_8[0]},
      {stage2_9[0], stage2_9[1], stage2_9[2], stage2_9[3], stage2_9[4], stage2_9[5]},
      {stage3_11[0],stage3_10[0],stage3_9[0],stage3_8[2],stage3_7[4]}
   );
   gpc615_5 gpc107 (
      {stage2_7[5], stage2_7[6], stage2_7[7], stage2_7[8], stage2_7[9]},
      {stage2_8[1]},
      {stage2_9[6], stage2_9[7], stage2_9[8], stage2_9[9], stage2_9[10], stage2_9[11]},
      {stage3_11[1],stage3_10[1],stage3_9[1],stage3_8[3],stage3_7[5]}
   );
   gpc606_5 gpc108 (
      {stage2_8[2], stage2_8[3], stage2_8[4], stage2_8[5], stage2_8[6], stage2_8[7]},
      {stage2_10[0], stage2_10[1], stage2_10[2], stage2_10[3], stage2_10[4], stage2_10[5]},
      {stage3_12[0],stage3_11[2],stage3_10[2],stage3_9[2],stage3_8[4]}
   );
   gpc7_3 gpc109 (
      {stage2_10[6], stage2_10[7], stage2_10[8], stage2_10[9], stage2_10[10], stage2_10[11], stage2_10[12]},
      {stage3_12[1],stage3_11[3],stage3_10[3]}
   );
   gpc135_4 gpc110 (
      {stage2_11[0], stage2_11[1], stage2_11[2], stage2_11[3], stage2_11[4]},
      {stage2_12[0], stage2_12[1], stage2_12[2]},
      {stage2_13[0]},
      {stage3_14[0],stage3_13[0],stage3_12[2],stage3_11[4]}
   );
   gpc606_5 gpc111 (
      {stage2_11[5], stage2_11[6], stage2_11[7], stage2_11[8], stage2_11[9], stage2_11[10]},
      {stage2_13[1], stage2_13[2], stage2_13[3], stage2_13[4], stage2_13[5], 1'b0},
      {stage3_15[0],stage3_14[1],stage3_13[1],stage3_12[3],stage3_11[5]}
   );
   gpc606_5 gpc112 (
      {stage2_12[3], stage2_12[4], stage2_12[5], stage2_12[6], stage2_12[7], stage2_12[8]},
      {stage2_14[0], stage2_14[1], stage2_14[2], stage2_14[3], stage2_14[4], stage2_14[5]},
      {stage3_16[0],stage3_15[1],stage3_14[2],stage3_13[2],stage3_12[4]}
   );
   gpc1_1 gpc113 (
      {stage2_0[0]},
      {stage3_0[0]}
   );
   gpc1_1 gpc114 (
      {stage2_0[1]},
      {stage3_0[1]}
   );
   gpc1_1 gpc115 (
      {stage2_0[2]},
      {stage3_0[2]}
   );
   gpc1_1 gpc116 (
      {stage2_0[3]},
      {stage3_0[3]}
   );
   gpc1_1 gpc117 (
      {stage2_1[0]},
      {stage3_1[0]}
   );
   gpc1_1 gpc118 (
      {stage2_1[1]},
      {stage3_1[1]}
   );
   gpc1_1 gpc119 (
      {stage2_1[2]},
      {stage3_1[2]}
   );
   gpc1_1 gpc120 (
      {stage2_1[3]},
      {stage3_1[3]}
   );
   gpc1_1 gpc121 (
      {stage2_1[4]},
      {stage3_1[4]}
   );
   gpc1_1 gpc122 (
      {stage2_2[0]},
      {stage3_2[0]}
   );
   gpc1_1 gpc123 (
      {stage2_2[1]},
      {stage3_2[1]}
   );
   gpc1_1 gpc124 (
      {stage2_2[2]},
      {stage3_2[2]}
   );
   gpc1_1 gpc125 (
      {stage2_2[3]},
      {stage3_2[3]}
   );
   gpc1_1 gpc126 (
      {stage2_2[4]},
      {stage3_2[4]}
   );
   gpc1_1 gpc127 (
      {stage2_2[5]},
      {stage3_2[5]}
   );
   gpc1_1 gpc128 (
      {stage2_2[6]},
      {stage3_2[6]}
   );
   gpc1_1 gpc129 (
      {stage2_2[7]},
      {stage3_2[7]}
   );
   gpc1_1 gpc130 (
      {stage2_12[9]},
      {stage3_12[5]}
   );
   gpc1_1 gpc131 (
      {stage2_15[0]},
      {stage3_15[2]}
   );
   gpc1_1 gpc132 (
      {stage2_15[1]},
      {stage3_15[3]}
   );
   gpc1343_5 gpc133 (
      {stage3_0[0], stage3_0[1], stage3_0[2]},
      {stage3_1[0], stage3_1[1], stage3_1[2], stage3_1[3]},
      {stage3_2[0], stage3_2[1], stage3_2[2]},
      {stage3_3[0]},
      {stage4_4[0],stage4_3[0],stage4_2[0],stage4_1[0],stage4_0[0]}
   );
   gpc1415_5 gpc134 (
      {stage3_2[3], stage3_2[4], stage3_2[5], stage3_2[6], stage3_2[7]},
      {stage3_3[1]},
      {stage3_4[0], stage3_4[1], stage3_4[2], stage3_4[3]},
      {stage3_5[0]},
      {stage4_6[0],stage4_5[0],stage4_4[1],stage4_3[1],stage4_2[1]}
   );
   gpc1343_5 gpc135 (
      {stage3_5[1], stage3_5[2], stage3_5[3]},
      {stage3_6[0], stage3_6[1], stage3_6[2], stage3_6[3]},
      {stage3_7[0], stage3_7[1], stage3_7[2]},
      {stage3_8[0]},
      {stage4_9[0],stage4_8[0],stage4_7[0],stage4_6[1],stage4_5[1]}
   );
   gpc1343_5 gpc136 (
      {stage3_7[3], stage3_7[4], stage3_7[5]},
      {stage3_8[1], stage3_8[2], stage3_8[3], stage3_8[4]},
      {stage3_9[0], stage3_9[1], stage3_9[2]},
      {stage3_10[0]},
      {stage4_11[0],stage4_10[0],stage4_9[1],stage4_8[1],stage4_7[1]}
   );
   gpc1163_5 gpc137 (
      {stage3_10[1], stage3_10[2], stage3_10[3]},
      {stage3_11[0], stage3_11[1], stage3_11[2], stage3_11[3], stage3_11[4], stage3_11[5]},
      {stage3_12[0]},
      {stage3_13[0]},
      {stage4_14[0],stage4_13[0],stage4_12[0],stage4_11[1],stage4_10[1]}
   );
   gpc1325_5 gpc138 (
      {stage3_12[1], stage3_12[2], stage3_12[3], stage3_12[4], stage3_12[5]},
      {stage3_13[1], stage3_13[2]},
      {stage3_14[0], stage3_14[1], stage3_14[2]},
      {stage3_15[0]},
      {stage4_16[0],stage4_15[0],stage4_14[1],stage4_13[1],stage4_12[1]}
   );
   gpc117_4 gpc139 (
      {stage3_15[1], stage3_15[2], stage3_15[3], 1'b0, 1'b0, 1'b0, 1'b0},
      {stage3_16[0]},
      {1'b0},
      {stage4_17[0],stage4_16[1],stage4_15[1]}
   );
   gpc1_1 gpc140 (
      {stage3_0[3]},
      {stage4_0[1]}
   );
   gpc1_1 gpc141 (
      {stage3_1[4]},
      {stage4_1[1]}
   );
endmodule
module rowadder2_1_18(input [17:0] src0, input [17:0] src1, output [18:0] dst0);
    wire [17:0] gene;
    wire [17:0] prop;
    wire [19:0] out;
    wire [19:0] carryout;
    LUT2 #(
        .INIT(4'h8)
    ) lut_0_gene (
        .I0(src0[0]),
        .I1(src1[0]),
        .O(gene[0])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_0_prop (
        .I0(src0[0]),
        .I1(src1[0]),
        .O(prop[0])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_1_gene (
        .I0(src0[1]),
        .I1(src1[1]),
        .O(gene[1])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_1_prop (
        .I0(src0[1]),
        .I1(src1[1]),
        .O(prop[1])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_2_gene (
        .I0(src0[2]),
        .I1(src1[2]),
        .O(gene[2])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_2_prop (
        .I0(src0[2]),
        .I1(src1[2]),
        .O(prop[2])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_3_gene (
        .I0(src0[3]),
        .I1(src1[3]),
        .O(gene[3])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_3_prop (
        .I0(src0[3]),
        .I1(src1[3]),
        .O(prop[3])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_4_gene (
        .I0(src0[4]),
        .I1(src1[4]),
        .O(gene[4])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_4_prop (
        .I0(src0[4]),
        .I1(src1[4]),
        .O(prop[4])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_5_gene (
        .I0(src0[5]),
        .I1(src1[5]),
        .O(gene[5])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_5_prop (
        .I0(src0[5]),
        .I1(src1[5]),
        .O(prop[5])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_6_gene (
        .I0(src0[6]),
        .I1(src1[6]),
        .O(gene[6])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_6_prop (
        .I0(src0[6]),
        .I1(src1[6]),
        .O(prop[6])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_7_gene (
        .I0(src0[7]),
        .I1(src1[7]),
        .O(gene[7])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_7_prop (
        .I0(src0[7]),
        .I1(src1[7]),
        .O(prop[7])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_8_gene (
        .I0(src0[8]),
        .I1(src1[8]),
        .O(gene[8])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_8_prop (
        .I0(src0[8]),
        .I1(src1[8]),
        .O(prop[8])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_9_gene (
        .I0(src0[9]),
        .I1(src1[9]),
        .O(gene[9])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_9_prop (
        .I0(src0[9]),
        .I1(src1[9]),
        .O(prop[9])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_10_gene (
        .I0(src0[10]),
        .I1(src1[10]),
        .O(gene[10])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_10_prop (
        .I0(src0[10]),
        .I1(src1[10]),
        .O(prop[10])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_11_gene (
        .I0(src0[11]),
        .I1(src1[11]),
        .O(gene[11])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_11_prop (
        .I0(src0[11]),
        .I1(src1[11]),
        .O(prop[11])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_12_gene (
        .I0(src0[12]),
        .I1(src1[12]),
        .O(gene[12])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_12_prop (
        .I0(src0[12]),
        .I1(src1[12]),
        .O(prop[12])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_13_gene (
        .I0(src0[13]),
        .I1(src1[13]),
        .O(gene[13])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_13_prop (
        .I0(src0[13]),
        .I1(src1[13]),
        .O(prop[13])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_14_gene (
        .I0(src0[14]),
        .I1(src1[14]),
        .O(gene[14])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_14_prop (
        .I0(src0[14]),
        .I1(src1[14]),
        .O(prop[14])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_15_gene (
        .I0(src0[15]),
        .I1(src1[15]),
        .O(gene[15])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_15_prop (
        .I0(src0[15]),
        .I1(src1[15]),
        .O(prop[15])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_16_gene (
        .I0(src0[16]),
        .I1(src1[16]),
        .O(gene[16])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_16_prop (
        .I0(src0[16]),
        .I1(src1[16]),
        .O(prop[16])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_17_gene (
        .I0(src0[17]),
        .I1(src1[17]),
        .O(gene[17])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_17_prop (
        .I0(src0[17]),
        .I1(src1[17]),
        .O(prop[17])
    );
    CARRY4 carry4_3_0 (
        .CO(carryout[3:0]),
        .O(out[3:0]),
        .CI(1'h0),
        .CYINIT(1'h0),
        .DI(gene[3:0]),
        .S(prop[3:0])
    );
    CARRY4 carry4_7_4 (
        .CO(carryout[7:4]),
        .O(out[7:4]),
        .CI(carryout[3]),
        .CYINIT(1'h0),
        .DI(gene[7:4]),
        .S(prop[7:4])
    );
    CARRY4 carry4_11_8 (
        .CO(carryout[11:8]),
        .O(out[11:8]),
        .CI(carryout[7]),
        .CYINIT(1'h0),
        .DI(gene[11:8]),
        .S(prop[11:8])
    );
    CARRY4 carry4_15_12 (
        .CO(carryout[15:12]),
        .O(out[15:12]),
        .CI(carryout[11]),
        .CYINIT(1'h0),
        .DI(gene[15:12]),
        .S(prop[15:12])
    );
    CARRY4 carry4_19_16 (
        .CO(carryout[19:16]),
        .O(out[19:16]),
        .CI(carryout[15]),
        .CYINIT(1'h0),
        .DI({2'h0, gene[17:16]}),
        .S({2'h0, prop[17:16]})
    );
    assign dst0 = {carryout[17], out[17:0]};
endmodule


module testbench();
    reg [63:0] src0;
    reg [63:0] src1;
    reg [63:0] src2;
    reg [63:0] src3;
    reg [63:0] src4;
    reg [63:0] src5;
    reg [63:0] src6;
    reg [63:0] src7;
    reg [63:0] src8;
    reg [63:0] src9;
    reg [63:0] src10;
    reg [63:0] src11;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [17:0] srcsum;
    wire [17:0] dstsum;
    wire test;
    compressor2_1_64_12 compressor2_1_64_12(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13] + src0[14] + src0[15] + src0[16] + src0[17] + src0[18] + src0[19] + src0[20] + src0[21] + src0[22] + src0[23] + src0[24] + src0[25] + src0[26] + src0[27] + src0[28] + src0[29] + src0[30] + src0[31] + src0[32] + src0[33] + src0[34] + src0[35] + src0[36] + src0[37] + src0[38] + src0[39] + src0[40] + src0[41] + src0[42] + src0[43] + src0[44] + src0[45] + src0[46] + src0[47] + src0[48] + src0[49] + src0[50] + src0[51] + src0[52] + src0[53] + src0[54] + src0[55] + src0[56] + src0[57] + src0[58] + src0[59] + src0[60] + src0[61] + src0[62] + src0[63])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13] + src1[14] + src1[15] + src1[16] + src1[17] + src1[18] + src1[19] + src1[20] + src1[21] + src1[22] + src1[23] + src1[24] + src1[25] + src1[26] + src1[27] + src1[28] + src1[29] + src1[30] + src1[31] + src1[32] + src1[33] + src1[34] + src1[35] + src1[36] + src1[37] + src1[38] + src1[39] + src1[40] + src1[41] + src1[42] + src1[43] + src1[44] + src1[45] + src1[46] + src1[47] + src1[48] + src1[49] + src1[50] + src1[51] + src1[52] + src1[53] + src1[54] + src1[55] + src1[56] + src1[57] + src1[58] + src1[59] + src1[60] + src1[61] + src1[62] + src1[63])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13] + src2[14] + src2[15] + src2[16] + src2[17] + src2[18] + src2[19] + src2[20] + src2[21] + src2[22] + src2[23] + src2[24] + src2[25] + src2[26] + src2[27] + src2[28] + src2[29] + src2[30] + src2[31] + src2[32] + src2[33] + src2[34] + src2[35] + src2[36] + src2[37] + src2[38] + src2[39] + src2[40] + src2[41] + src2[42] + src2[43] + src2[44] + src2[45] + src2[46] + src2[47] + src2[48] + src2[49] + src2[50] + src2[51] + src2[52] + src2[53] + src2[54] + src2[55] + src2[56] + src2[57] + src2[58] + src2[59] + src2[60] + src2[61] + src2[62] + src2[63])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13] + src3[14] + src3[15] + src3[16] + src3[17] + src3[18] + src3[19] + src3[20] + src3[21] + src3[22] + src3[23] + src3[24] + src3[25] + src3[26] + src3[27] + src3[28] + src3[29] + src3[30] + src3[31] + src3[32] + src3[33] + src3[34] + src3[35] + src3[36] + src3[37] + src3[38] + src3[39] + src3[40] + src3[41] + src3[42] + src3[43] + src3[44] + src3[45] + src3[46] + src3[47] + src3[48] + src3[49] + src3[50] + src3[51] + src3[52] + src3[53] + src3[54] + src3[55] + src3[56] + src3[57] + src3[58] + src3[59] + src3[60] + src3[61] + src3[62] + src3[63])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13] + src4[14] + src4[15] + src4[16] + src4[17] + src4[18] + src4[19] + src4[20] + src4[21] + src4[22] + src4[23] + src4[24] + src4[25] + src4[26] + src4[27] + src4[28] + src4[29] + src4[30] + src4[31] + src4[32] + src4[33] + src4[34] + src4[35] + src4[36] + src4[37] + src4[38] + src4[39] + src4[40] + src4[41] + src4[42] + src4[43] + src4[44] + src4[45] + src4[46] + src4[47] + src4[48] + src4[49] + src4[50] + src4[51] + src4[52] + src4[53] + src4[54] + src4[55] + src4[56] + src4[57] + src4[58] + src4[59] + src4[60] + src4[61] + src4[62] + src4[63])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13] + src5[14] + src5[15] + src5[16] + src5[17] + src5[18] + src5[19] + src5[20] + src5[21] + src5[22] + src5[23] + src5[24] + src5[25] + src5[26] + src5[27] + src5[28] + src5[29] + src5[30] + src5[31] + src5[32] + src5[33] + src5[34] + src5[35] + src5[36] + src5[37] + src5[38] + src5[39] + src5[40] + src5[41] + src5[42] + src5[43] + src5[44] + src5[45] + src5[46] + src5[47] + src5[48] + src5[49] + src5[50] + src5[51] + src5[52] + src5[53] + src5[54] + src5[55] + src5[56] + src5[57] + src5[58] + src5[59] + src5[60] + src5[61] + src5[62] + src5[63])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13] + src6[14] + src6[15] + src6[16] + src6[17] + src6[18] + src6[19] + src6[20] + src6[21] + src6[22] + src6[23] + src6[24] + src6[25] + src6[26] + src6[27] + src6[28] + src6[29] + src6[30] + src6[31] + src6[32] + src6[33] + src6[34] + src6[35] + src6[36] + src6[37] + src6[38] + src6[39] + src6[40] + src6[41] + src6[42] + src6[43] + src6[44] + src6[45] + src6[46] + src6[47] + src6[48] + src6[49] + src6[50] + src6[51] + src6[52] + src6[53] + src6[54] + src6[55] + src6[56] + src6[57] + src6[58] + src6[59] + src6[60] + src6[61] + src6[62] + src6[63])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13] + src7[14] + src7[15] + src7[16] + src7[17] + src7[18] + src7[19] + src7[20] + src7[21] + src7[22] + src7[23] + src7[24] + src7[25] + src7[26] + src7[27] + src7[28] + src7[29] + src7[30] + src7[31] + src7[32] + src7[33] + src7[34] + src7[35] + src7[36] + src7[37] + src7[38] + src7[39] + src7[40] + src7[41] + src7[42] + src7[43] + src7[44] + src7[45] + src7[46] + src7[47] + src7[48] + src7[49] + src7[50] + src7[51] + src7[52] + src7[53] + src7[54] + src7[55] + src7[56] + src7[57] + src7[58] + src7[59] + src7[60] + src7[61] + src7[62] + src7[63])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13] + src8[14] + src8[15] + src8[16] + src8[17] + src8[18] + src8[19] + src8[20] + src8[21] + src8[22] + src8[23] + src8[24] + src8[25] + src8[26] + src8[27] + src8[28] + src8[29] + src8[30] + src8[31] + src8[32] + src8[33] + src8[34] + src8[35] + src8[36] + src8[37] + src8[38] + src8[39] + src8[40] + src8[41] + src8[42] + src8[43] + src8[44] + src8[45] + src8[46] + src8[47] + src8[48] + src8[49] + src8[50] + src8[51] + src8[52] + src8[53] + src8[54] + src8[55] + src8[56] + src8[57] + src8[58] + src8[59] + src8[60] + src8[61] + src8[62] + src8[63])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13] + src9[14] + src9[15] + src9[16] + src9[17] + src9[18] + src9[19] + src9[20] + src9[21] + src9[22] + src9[23] + src9[24] + src9[25] + src9[26] + src9[27] + src9[28] + src9[29] + src9[30] + src9[31] + src9[32] + src9[33] + src9[34] + src9[35] + src9[36] + src9[37] + src9[38] + src9[39] + src9[40] + src9[41] + src9[42] + src9[43] + src9[44] + src9[45] + src9[46] + src9[47] + src9[48] + src9[49] + src9[50] + src9[51] + src9[52] + src9[53] + src9[54] + src9[55] + src9[56] + src9[57] + src9[58] + src9[59] + src9[60] + src9[61] + src9[62] + src9[63])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13] + src10[14] + src10[15] + src10[16] + src10[17] + src10[18] + src10[19] + src10[20] + src10[21] + src10[22] + src10[23] + src10[24] + src10[25] + src10[26] + src10[27] + src10[28] + src10[29] + src10[30] + src10[31] + src10[32] + src10[33] + src10[34] + src10[35] + src10[36] + src10[37] + src10[38] + src10[39] + src10[40] + src10[41] + src10[42] + src10[43] + src10[44] + src10[45] + src10[46] + src10[47] + src10[48] + src10[49] + src10[50] + src10[51] + src10[52] + src10[53] + src10[54] + src10[55] + src10[56] + src10[57] + src10[58] + src10[59] + src10[60] + src10[61] + src10[62] + src10[63])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13] + src11[14] + src11[15] + src11[16] + src11[17] + src11[18] + src11[19] + src11[20] + src11[21] + src11[22] + src11[23] + src11[24] + src11[25] + src11[26] + src11[27] + src11[28] + src11[29] + src11[30] + src11[31] + src11[32] + src11[33] + src11[34] + src11[35] + src11[36] + src11[37] + src11[38] + src11[39] + src11[40] + src11[41] + src11[42] + src11[43] + src11[44] + src11[45] + src11[46] + src11[47] + src11[48] + src11[49] + src11[50] + src11[51] + src11[52] + src11[53] + src11[54] + src11[55] + src11[56] + src11[57] + src11[58] + src11[59] + src11[60] + src11[61] + src11[62] + src11[63])<<11);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'h0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'h25592f9183768c042e3d7cae7eaa3b70afbaff1d01c3c62f760b27a609f0c00c89d13ac765889dfe352c86a4f3df759c882804e8492b3993ad518bca7327c1b4e04f651b42f1726689a69ff3e440adcf81369c54f34c09234b2199a169595337;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'had9dfc361f366b6e103cf1b6fa69b5d4889fabe7a3c2fb0db2e2f5ec9cb7a581bc96a07e64bfc7bffe5421175c7ae9e227acf29dfa39e93467dfb59bc90ffefee61a0043f8928e17b523e7aa7ed0842e62aeaa0c397878c7e19abe3944144dcd;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'h75aefc0ee602c9e00a2f3c4a8e37167266dda4d444c942271d0bec16a720f34ab837ffd28d125d2f1e843a076ebd3d1e943038cf73324a71a61242c5f198842183b6e52644b1932ebe2a18055b5f7b7c7bb03326573155279b0b78acbe882d99;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'h16bd12cbbd586d2df74014665fd987560faef45d6ccf375c9fd680cc4651d40781937cd23e5f80a84966c07e76fc4aa6356c4a8528c30e46d8786590e46f6a60ddd7ede0bf0dd7ac0634db8e2022f0421113c302123551827afb30f8c0d347ab;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'h2160c9c468ac586a86a9672a52028fb5421584fa941968ba33581fe664b46b9f770e8382d7752007d4700d2ca10efa813867ebc1f243f44c5c2eda860e2d3642ec7597da881f202bb8f9005e01a98ccb45e2ea312e6912c7582d75a439034fcd;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'hd8602f4c2c318de51a1456607cb35c9d70edce902c4d0268d2488aedc81a7141788da7da3436fbaa8b23d3339f0d46c0c7da4a7136b10f745d05197f2ce1a48b7ad8d81b374a3b48880df2f4973c0fd0a74579e6f50f36041cea05541be5017d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'h2f61e67813c20c485d9bed3ff56249816ce430e8f0fc11583f8005add76d3b6522c0f660315ed2537dfa2c4cdbfcb519af0b9cbcaa6021aa07b6fc31bebb4f7a673462a0848e393c8328445e78b9fb972afcff4c62e94528439c6ec1221c7b04;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'h101921e43edef797aa1d03ee22ae854d2b8193a0f99063f4256374e57a6cdf69dfac427dbbfb6d2ec101121efe9ec8fb567e15e08cb66c654a8e391106df853e772e0774fdcd70c4d9138006aa8b867d9debb1884cab68f85c9f876c0ecc0852;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'hb71363eccdfd2ef1e28de4832a7741b492aa7efb932ee80a84fae96193816ccf5f1ffd1833c6fe30df3bec157752af44aff45e8ce8c4e5f3b94978bd631a69a3255bf38734ca0a3480ffa5e76821b18ab3dcf6e371215448b820f9267202455;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'he1063fce22b25e83eff320e501205049c6bf3789d8c18b1e7eb8509f73505156518f34837d6f51a8e0336627ae83c7a42364bc41ec18f9358c58d9fc969cb4ea015fee2032d5b70be473a25c0d4009b5e5724af13c84d9a7154a3ab4c399fc54;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'h31851996850baff03ec86a1c110b26baed2b059012929ac93829d2aa4d7092ced846bf17dd9416210d3bfe5c873481941dac750172402ee9c3c04ea8b54e58c412760f48c2d7d52a58a2f984f48bd26c7afeb5b77313fae542eb753cadaeb362;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'h2f37e9d66643b993228a5a7e893bad751684c81d02255609facfdb30a903dc5ec6523b7ce73b48e22ac9a6ddb346ad419564c07a4b921bdcce61f11e5fa9c7ee29270953c774cdf1dfcf39a3a612a5a1c7b49fa2bb2ec02ae78a1c54d2ec4118;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'h47afdb2382becb3a2f11cca168b5fef6f2ba3c7c1c608a8be5d78a6d321cf9dda36b095e8aee3fb3603be89b41e1eec3c354fd3cc27b135fbfb307397cfae21ee748da99c7ed38e4eead04452463b242816b15af39835e1a902a0e80c4aab19a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'hc04a42aad31cbe2d2991aa224facdff3a0c916589097ff912820d6d089e5d838df256b5ec0827cf6ab35bb9d353c07dfc13d0ba11332efc573f048cb6aad4f3234fd614f2635de5b6e73ca6ea7ecd658d00e8af81ff0f3404cf81ba7b9944f12;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'h7515f2b3e1c9d3cad0c7b4de70612cb94ee233266368d09c26cea71d7a0e6f9893afba5a7e5bd8bd7526058feaaa6929d6ebfcf0233bf91ef10a714c84c4097c24e2698533b438f5abff74deeaa5c101fe5d12fbf21325591acb28b7b402f79d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'hb6255b7c1a1c4c74fe56c1e7af974c97abf09ccc4926b08379bd1ca18e9422814513ca69667f13232ed682270a4ac4fab83c8dc4dd3dc8c2284d8c65583a974817ed8bee0998c7c24c051be922e526757b53733bb827ba365c3ee3436725c23d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'h18179fa00452de292020a22015881338422b3b438672230636cf264918a9e7f5f00f672c2bfd78dc6348f002b53bc36c8b6faeaa88d3216f4e0e2baf825c966b897dc99819f7028b8faf1fadbbb82a967c6b4f1e52153e30d3f1aa8b4ab6db4;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'h82c1181a448d505a0eef31aa093657f1f7603d1293ffcc9522dd0d65ec3cf3398c6f5843105fade30ab89f3fd0b064359a729a64272d42916ebae649d6c563f63774ebf934ea299638a26b526be9aeacc90823793ebba55e9fdf01052afbf6ab;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'hc3d21553ef57a83d1507005d8da16ad21a34e39cb8a2fba8f68b3e90e2cdee65770c7d87c2400ebb3061be91c1b5edc18e8d1b6e1b2a774289f747dadadc3b8fd9b6fb4c135d7529b71adf90390dd62f5d54b2efabe3b1118b14834f3c3aab8a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'h71ee075fd78ad10f533564abbaf5c01b28c1af4b8a4482a8094e5e3503372f912a773c1d7f0bc26b06b7550dccc4461795db8dd435b07be9b418b16b3da53c3bceaa4f3f84a01ddf10b2a25fadfbfac72620be0365e1cf3652f6e61453f32a57;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'he72a99af527bd56a5e5c6ffab59b4cb37e8fa14f1c705b92cbd4a893aa78737f8a08b086b61086fb263f312d524bc633c2b1d069f4befb74ef1134f2697ae7f1f5ce7d30c7acbc04bb27bc2f6735b5e3f9f6ecf2262b935ce56d5b59d64f612b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'h2865f2d19cae4810f2a89e9141147cc3848b3891ff89670d127b6c54fbd0132f6781923a72cbb1238d04a2e66d37ebc8c2c45ec87afa6a6479ce263cb6834af2f69c98a3649c217a02bc544b5333fc04ee7fdc033e9109a43073902c4db246b6;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'hdf7c6115422bb1aec0e4ec67d66b8e4f55cf9f32182302903013a852e47bfbe4b8f97a277b092ea569755f8f60200413a3bdcb64600b058a4353b4e59f5e42abc7054afa958d7dc988f19479fcfc14cf6ca23dd790efb08406b565fd09710b5c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'hc4d83b82860adb6931671c0f877435e0ac616cf1968e731c5cc0a717767e10417e69de003f74fd24fcb71ea5c0366354966d9669c5496a76f36e085aea7d486254e0202f833d97e358f004155911ef364fb373f63cced469d9b18426a0aad458;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'h378fb3d498740f6910e09e57d0a156e6d483abbaf7b4bdb2a9de0f13f3c5c4a6c03b4b9a02891eccf7603c953e5d00dd6dd4bd4618f2560f97c7ca80421edb310990c873c4073a3d380679d0d0c2affaf007d306a41460c81f48a72118116122;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'hd36bc20804ec28516a7b685f6e91e41bb4a50b86ec4f6d5f68c0990df0dca3b495b0c0480f3d9d1021450278e14af4e7089472b7a8c4b22c329992a3bd3ccd48342a25568be4f07dcdf0699e76f6883447f28e32144cd9246f564566dfb947f8;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'h28fa8a923172ccbc0be0a72da563221fa393722643aa812fbe7912600fb334fab7efc7f55c634fff5db5ebfc7aa650a1880c6459810f266d91b93adf44e8099b47cc35bc7e3c12445d8c7b401bfe332e0055c823112c912efb89135658a0e70f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'h582df674d6637562bdd90d0290a8cdfeff4bdb265f11a29e024f13f9f5173272cd5c9ea42feb13f483542dc1e6ec88881e0786fb17f42577f7647e4a5154e5ca3badb9b5849f36437784bbbb94bce562edfbfbbea68f8dd20c68c7cde0a90008;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'hb4adb9473be7d767f82578de53f85e983b2d147e4f58d2732b28c049fbbf4b9c99895fb07c27680d14876a02805dcb35d549516cd7671d9e9b8f4c1e105eae714fa3be312226c47d1c56e905068504c200296b528faa7a667224bdf1b623890b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'h5460c1d2486d8771c32077fb0e9a5c5f742b237fa87d270b2770dc1d073073a65d57eb15bfb45f8aa935b3733cebeb94be5c6e537eff24bd05129e2d9bbbd00e23e1a060d2dd3bdd29ee3aeec788d68306db3138c2bf5a5bef166aef3f4c589c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'hb7c1d1edc22af77b2d7d50d807450f69f9388a6439d06f5fde468477fd771c586034c413ee606dacfd0eec5d5031f8a246d9630c3f77110d653487a7a8503d2728a7f799d075d0513b31846949530abe5c1e357dec4a4192be0cd743ae1048e2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'he616a1f17cc83a207438d102e8e525df88f86db13de3573a41d545cb83d497f5053215126d86b421b57123486ddd23794a5995618912f2d989ab89d0ff80c0e53db2f631ad65b40b79a20d7a179379f299c46bd4af2d4508f79d9f47e2c21c33;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'h922c3578bc789ca4e43617fa3bb7ee97390c35dc9f38737fd1bd27a416fb7feed3c48d4ad721a97cba364df16ec31781311512c6faf164e19be750191bbf60d2d28833da79f70686dc39d1dafca03f35827d46a8413e23b24c40b2c1c838d570;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'h37189d4e41f1c4c058353bd27012c8638abaab33288374bbc3fa77665b6f7aaba3203f6f7389034c9d04f637876226427e3c614f7d74bed7786fc4cccd1bab5f2a792109c1368ecd336a3fd17f61a72e8c80cfef871a6db661e8fddb9274c71b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'h9d16a368c6672ef707029cf9d42b286e7b2c78cf414505f5c6bd4826bc5f74da1752ad38f3cec749015d62d2870fb16e1c06f9b86ebaa516d894c94ff69e9e7e6968f6f44f02797649e810c25edff817392add1bf540fbf4b0c3199cdbc045a9;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'h25aa4bef60272c5f0073f549c2b3ffc7e382e8c15d502fad6779366bc6a03e0a253085c5c83e4ac817360b966453ece18df560077026d1a5c08a9f165f25244cfddc2a145530cfad4c247c42337f931bdbcd4bc146ea317dbc8d6812e23c4ad;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'h98fcf904b4d547d369eab29d8e06a67bd9a35da85c7b1a8b55db2f39ae38b32690621d16a538506906c0827ec183b3e9262fab4d17caa606ee25743be0a61d2700eed41cce3014cf10e47faeba0a91a08f986fcf445934cab7e862090ef3caf;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'h52ee934f7b70c042ff266ba3f457fcc52cd825274f662c730bf0368b88bcfe6a6b9dd3588024c5fad1293df10850a63346756c4e4fc6c639c63479d5a9da5be080bfcd65c036f6ec01009cb8e681d3b6a1dc60b5401d8835ac0f070dc1ecdeb0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'h8ff365452635b01a917650d3d7c3fb973813017e8ec0689eb0bf15753833373d2b15aa602f35aa71b444d79c4e4d026c001bff5ceb132a788413afea44814b3279eae238a4fde0bedeada42f28add4cd5c88d3d7731d8a31557402e727bd2131;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'h9cfbb4fd43cb0fedf6aedd76b824fe0baa26e1c5230c6d4dd3f2907765bb22c14ec270cc2c5b827c3ab973bb1f0161e6556d684a4be8d7337a3b427228ce48cf33b128fb81cfaebcc6f239e08f2c66edf7a4674b327956e9d5ed2f4c9cb003ee;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'h7a3c720adf05fe0c8ef490be6d3971e17a0d01aa18c3065c6275c9eaf1cbad462dc1a2d7354004531cd858e9c5ef70022dfe7b8eb6ecb244c5fb3422934b1d3fd6426c92ec8f709b031c334ed77c2e148eb04b6fc1f7cb817f8b44aae39a620d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'h678086ac23e7bd9dec3f1d3976f708c34dc3de8fa0f9ebf7868fa0bdac2d59c020ed0f0ba1c809164998b70a77e092da9cb0bb6f77d080f0fc761c8c2f024dda9a7ff5fa333260bfc8de35d76b09751305850937a54bf3b594948e13455b8c30;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'hf4903851029f89a050aeeef6c1fb54cc50f3dfcc63d7d40f9d79815b9e57b5797ecb96df3624a9f920ac42ee8aa2acb0fc7a1ceba456e772506b615c91cb18c0575b9788b3966c8db02359850f6fa4575dad6cc694fbb4321ae437340a28f38c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'h7f12bc968e417f1724b1322019c9537a9b4fb3dcdf2808748b5ffa54699b15f2173a506a80f15d39b32dea64f5325ef37ef727adf23141d44963b2bdae78ff43f5987d4a5ddc95531bdebac8b0269aa0dd2463731976902fcdb11b325201e766;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'h4541abeaca09f5cffa5926ec31af35e3e09d2a07451c165bf9e40856c17145ed52e8d9676d8d6e753ecfbacbca6a0dd14eb290014092efc9ecd775f48038de6bb61558aed3e83d6fd8643b5e2fed0af695704c630a3d09757f85ad9ad62d1f67;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'he018aede62d979f6f81dbe70fb2332184d2b33050dc63967bba4e0a89e58cc42fb01ba8cc38c6e6acd361b8332ccf82b750e71c3bd2d553568b2d7785fe2be8f378a15a2775fe5a03fb40a23596bd9878f1000dfb70d28fbbbb2e8793b0b157b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'h95806142cfdfdf955955a01de52482a1182bc8517e10c11c1bf4bf046335d00aa768d5dea73ed84a0ddbf78beae4e90d28399adc5cec7bdd2c8667e1c9543662dd1cd09a45611ff2841bd77e058018d8a1bf21418e886ce12dca3c84d1472a3c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'hd8440064da3e9faafdb9a6a89399d2729ae47855a50ab7347d9b9510aa602de45d2e6b023b0b28c81a1c8ad98b575c8b55f05a53776a24d1aa08a32ffcd21e60508590b1c2c4147747cd4619525e5ecd0412b91106896cc33b91ca73a9f890b6;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'hb5ebfb9ba5f77206a9ea016a85d0c8fd2e68f1c5169208cbf1b55bcbc16aae8dc3d6df97d2aeabb2095a8279088fbb6f286bcfb47f760a160a92e4ddf61fccff3871405fbfed9cfe0b4cdc77b318a26faa792f9c3f73b6a331125158d831792b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'hc9352dc8107f849d70136154f0d3b1ff02ed911a5fd9ace15c9afaa51d757b2efce5f9da91567812828fdac66ef29a51bfe67a26b538df37bb973dd854beab2c33e33b0217e9e2965c8f563d805e7a9e502302a6e33ef2131f9343210220058c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'he0f14eb7d0dbba07e0b77e53b1f7dbba716c92e66a3313349a1b1d3114a787d7b93113709e776cfce1fc4a1b0a591234cb0597b71e529028941b85f271242dcaa0ff3a602954f855ad8147377b2470d49c15179b192ae2547fa65477c7f6e6c0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'h13ce4b24e6ec2bf25ec9e7136d785a40f8b7b561e29a6489968d3fa6d7e866639e7ef499b291a072c437dd89b9a26cb7cce342ac93055b258a502f609c0a334cc68822bf6f885f116c8d6161e1030c33b754685f47ef2a54775739a9571d74dc;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'hbb1016ed0aad39b95496668a408f1417e75dd005b8f76a7fb8952b5888277390624a148e38475d729ed6d2c7fed9d2054beb550f9fbabd74d8874c437d8ba45c60b3b19070c40d44b82bcb03f9b425c08b55c41c0e74a8f7fa4991aadc2eddde;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'hc7b6654ce63d72bc1449cf2415e25d6ce7d47f984e99d2a83aa50dd404b0491b58856aa39866fef1ef17a2aaa0961b4dad5eda6f50a064731aa7f5ebf3f7032afd246a1867738b5047863788e8345b39772faa6c5f19b10835c528f6c2082545;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'hb41735d5a5201c57600b128452ecb7a9ddb9830b6c5cdda3fa7d499f6c5fcbe50b7251122291772e298344feeb69d8c434099b81f4e2e1c83dd40fa7b83e99439fa0c604526e4514ca1097eab97f71925533088372509d638d89edb6e35e605d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'hbf33821c9e56ca254f57603fe7dfe20fe098ece4190513ece2f9198938291e3298d849289c25f637064dc95f64555a648f8c4af198cd44cc0a3fc404e1d8cd2539604da16b5885e958d06c9b32df0fb7e23d25cec0fc681ecdaed56c14e8098d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'h12014f89e411e5718470ca4a71371609c716ee2d6441009a1d52aacf8ed96f761fa010ab59cd7c9482f90f81ff6481581baf207b1c47ceb143ae53532cb4f01dfb2fe861f383290c1c2dee41c4a1e2494df6ccffb7df262c2f5d3b79e108b786;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'h9dda580b4b33bca3121041d6b4f6727e23c9addeab86aa69270f8fc00f842c6d4656e6fe583faf0896e89a1d40201b4f95fe8e3d39be30fd21dd64c9e597c4e78681cd36bf71664c7a83beccd175daba36793df02ddbeaaa9ecea94c5606978d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'hfba7469cafbe0ddedede6c58f3d2644f9f4c3c2342cb5c95c63c3490d1d6754c5c1a3cdc55acbbbfedb41763a6c84c6ed28086f672267dc62e6dc133c91247c812ae37bec8138259668159d5ea721018e865ae1f3f65fd3184829972c2f52d97;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'h989744f8a763cf28cf35b64f38974e2386fd52c9ea1df552ed456a019502670ba0a502acb0db6a2067b0b3722b5aa61d27c9a92ff391918059cea96b3046dafd041706b9d428e9608d4819b56c3cf7b537c62c887ae06c2db9a98c9573353908;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'hf810eb3770d1ce2f0a20ec04e3f7c723813d89e8ac95b06118e1abaf70307b69bab6f2b5ebc669a83615c9ef7c18748352ac84da4309dc3cfeacafcaa0d20a922e2d8bee71ee1042dde78133124e2c2265e21a8c8b8d9ce196b5fb44f8b4cc;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'h6a0949f96b675ad95b86e398c35cc7ec5d47a4a7c9515b600b53c67a26c3281b680d3580383a9065852878d8a641d9b22a417b5f6ec3e45a0bf0fdf67709d2944ac4fd9bf156c0ef076df8f7a9825b273ce4d8ab95feca67ab7b6c988335da7c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'h4b26fd654a3f42cb734f8c694886870368c876f2db81d950f69016da324da191ae8374de053678cbd959e94499233e539634b359c52d661a0aae8eb4b12cdade585bd965de03254dd87d66f6e9286b3eacd656895078587cba79b804aff35b5b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'hc13a110dabfc048475266dddf5daf8f10c99bb897f8c11199b8d751e9b04197b68ac3adb25a5c9152b4df464f4085b941e3a810e868cc1842c3a88c2d371319a12f6994d545ab603cafa036db4d727ad123098f9b331900533edf3a463554772;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'h1602017c2e6b9d4a2adb620b21f227681e4d692285a9f504bc4c504f5ed73ca198b86ff85931ed373c748138cb6655178a2a59e056290f99998e8bb92107441e888129504e9980ddc9cbf4762eb206c6a73b6e3ee6a0316916c0189547b739f6;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'h89603ac62a656cc3bbc792950a0a0e5416f4c040f0609ff0af452f99109db28ba71438d789643c073a1e23584b86a2ab0a6509b5da6cd470f3d6be75494466fe4dd66789c1e9b275e854e84a6745ceb769885ee17d46da331d97967858b0668b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'h8b9962fc5eef953b6c57dac8263f59df00b0e1db0bb5930083624eb41bbc9f538a75d74dc41e79e03e108301a8d42634a56801126425e2f0501026e418f73c7515ed52e46e46717182224e9da846fbb033f032520bff8bfe438cd96dc8ecf6f9;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'h859bf9132d68cd3c351a02722755211a2e224fcbde08866d2422ee7df9b6d935642b969b4b54534e3a81e7f61000825c26a58d5146b34b2940c443717e0d084a75b66efa25758e34cb86d6b5b188ea398aea45b7532100ee94a128bb9a5978d8;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'hfb0c302b51bf0b4b8ea36d785ed9315f7bc3dd153d238b40136841d21503ddc11689f3074e3c024f74141510ee03edec90d61d5d45efa65a18d728935d80dc09a2ded17fb03cb75091dfd26ae0509c30e5bd51c862fc1582c52de121504ea6f8;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'hf84b7cf9682cff5ff954df9369d2030b8cd538e8f5371f92abae03adb511c73ec32122dd29264849f15186600209d76aa833267d0e114afdd240b984ac0a03b7ac1ce813a1e11c6e2d076b822656f0929f5b47f59d646ca4386b4a0a0f395e36;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'hc3df1955980067119b7abbf6ec72641e2e0fb8eaf1ccfa6b43c9d72f659c22f81b94cfba5083fc60204d20a108199f3ff76796e291f2c87f6dcb0e63095a615413e3afe8163c658bf1b807a49c53863d5ee19c4853f485f61421640b6ac0f381;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'h6544470eb590297cf24af0cbc89b29d9ab0794e8ae29442b9e23e1f66192208933557fabd276d74fee1932e3aa46959d3f3ca23a7e298e2dc98e9c532e1de10a0a0c2702bc322c0f3c20e00d9de4d8aee2db1104d7c70923b1ca4781e32cf1bf;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'h5065e87b674c9c29abfe2ac6dd4f47c14e0237e39a1ad1416d151da323a92fb81e79384ce95fc934d172915822f146e4b66a800c78f43592672a0f3783d7fb6351b05ea6f1b60fda2c48590d87a1c235de6cd7eab8571a0bbb448ac8240bdcd3;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'h99d3acbaeb01c2fc9d6bf7bf99a7ac53255799fe3e62867ff011484db8a1913865baa561ff9c7ed4f24d690d0910ff74b6febd974b8695d058cfdc1736c92c92d9d92e8c718780d7681ec7b9f06c9e264160c81fe33a8e45db9d73a5ee00a6f0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'h129dd0284c8649ab6d35e6bf36e5c9ff81f778fc35611ae9c0e6c038e4ed5a8aafe830882fd3d036a005a98997f484847b0aa9fc4c9e68a6638ceb07b5a621d06390896a268ba9f81449976fbde7c6737025f6fc6c44a74edd6654db2b5a1325;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'hda9bbe638e3252029bba06bbd08492730bca1d74b878f701b6f9e58a4fac838a814a5a012375404eafb2a70f355c56c5ca405709ef7a9743070b8a188a400eceeada34a5a11302bcc6955b498e44d4ba3005f2802939b41bfb932f34cc74362d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'h5b52a585d4b10b15292eb670ad06cc29d3c33944ed715964473e1bc988dbdfbbc819d10477d4864555369a4096a2ca7c0da27deb8133dd50413b11cde7a46d6d96e459ec14445f0daef79582e75971abd81994d6c625b613af075f2dd871e316;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'hc359d8de317602879fc951b8b0ef2913dbfa79de4aa919b1b91a6a85a1f90de88619d81cdc95cc3ad37eea6477adc84c2b26ca1b0b5c6406d00343a9e790f441cfcbe93fcc63415773d1a48f53fea3ebc34e38720f9a06af9873de9b1f4dd4ae;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'ha8ec31da1569bda0cbd4eb859378ed8b8cce83de48085c83dd9c16f543c8adec4f8f650185bd39912d8fce677f422d8c3b2486869ea9916c175f80a846ce625fbafcac909be42c69eeb4832d5a8662f8c9bf60a762bb611c57156f415fe82e49;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'h38f550fe727223713718a768044f26b87f581fe13907686aa7da537b47cd629d8e415bcd03a8282553b58845259558c68afa5bff42b6ff7189c09a6a05a3a70a11868b22e522c809297f136f3fa1857702958815af365af8c52bb3bda390e706;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'hf8c2989b670cb1b25d5343b47c8bf53475c9a2ff58f5adb4f710c07e2cf98059748ab9b9ae74fcfe5cd2293ebadbe12087dcea2833e92eb1f93d21095e5eecfe80ecf101f1996f77cf0d85760462f72ab2196b3081dd04a1ad58a8bcac9cd04;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'h89575f111f1ee713458a6cef0ba457ea0f34d433e15416629bb6cab423164cdb33bf6926c038206ab68d116f108fb90e51643f62ee12276dc8e4eab2ae9f4fd19d2bbca17e5a6c678a9d7ce99afdf4ad1ee4e167609538f1a01b0b5c210aeb4f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'h24f72d9639b6f137e71beb73b7fc6188b831db1492552946ff0ab1718f5daea78c20fb3b7b7d4e160b63af88876a320c566926b01a94d8f39bf8cf86c3d55e436bc94d54697fd52bca1be9ac3dc41f0c9c16b8fd366fc25d6603c1a4a47d2c90;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'h698bf89eb6a0b7ea467275cd179fca69a9f6995867421b8ab74eb0cfec1fc53a5342b321e4a720a574cccf8ccd15c523c8cd6acee3de30b9f12ac44c3cc7d440b3693da4359b8b0242a584dea503431bb7e6ed3ac13a0a51886cc567841be959;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'hd0ebe5875215a86eb0d68ed5751ceb7eb46e3454b724e27e5860ececd8aaed1987a359ef98932f9b3ed0d266c05ab35bff5c87b335df641d10d49d32a09d3a9e7881378334ac9e009d760aae581af5495273f5c73f5048b604c24dace37f4e59;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'h7913dd6125b0fb65ce4e2bcb7898361d90aa4f56c52b7022ab86b87c04813b9da469eb69ce725ece940c3f4eb4e534b996f300c580175af5ca2d7793370fff211a6bd6853c77fc4064c2ad6e24c39dec872014505bafdfcd9084ce011a06534b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'hffe5070e3bda758d029cd4114375395911b9aea6f8ffaf9ba0d4e5dacb8f7f195afce4c2cc836e37e84776fc28814d6610bb221982fca9d8dc89f5d913973100e6c70e89643f04ab0613fbc8d87b1a03b3c3f78b067e784eeeb22c8e0f0c4461;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'h2fd3f4743c04f90960e94098c2e33f27679a0683c08be8f5c5033ab1e2ac33f69b1fac383ec8d1056677105971625c3e6faf96608301d74da3012fa101f12ed1eafd7b7350e9a1344be82e37d79bcb545b7505df371a719c94c51fef60683c4c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'h41f0e2b3dbf9fc5891bc3f92f653e10ffd6a295f3172b51d15a4786d8c7899fde03c79573180a71822c7cc9a93edefe9ed4d5623b1d7059f4600e55701a6577a2e53c6781e58df688f11eb04681c895fd532c611fb48272f40ffdd853e28071c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'h585267d175046d16a59e54ede9b084187edea021c666ad66e61f3e11d4689248282b5c5d13d33bff6a43122567cd2c387208575bd947403d3c6d323596c78b9fa2c001a431eb631649d3c1be28632065e9bdf0d3dbdc0001389959b1fe4b1252;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'h975d13c928cfd8a5e97b0ef9576a69314109986bbc99dfa1316a4ace1da06682611b145e78a422e2a520202d56b488569bfc993ecc4b2341cb3df1a4721de16b0f0bee30127639d92799369ef06d5377b6d946bc244b33a3383204c8fa182bbd;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'hdee519e87b5c0dd8725fb891457efbadf47ead2cb3ab7b8ce31efb9e03b299b1a10bd15a49929608b4b6adc5c5a2516fafeeb0e9e740a4800abb662d45fb90cfece8148e32ba9ac0142398871ceaacdbde13ddff23335342e89eb0f1f4bc537e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'h862cc78b6b7231a97db2c27b5f79dc596c2eb8ad983344a423971d844ceb365e0016325aafc5f209769c3bcab6239bea98634a425ff1350907d9bc382dd2a888614e7190c398abcb735642f77cc33b7cc928eb2a5a788fdc497fdebfccb3a4f8;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'h1e63404b2909bb425dce5da670f6f15e0ad739fc7ca0d0d627661f59636134268f528b10eae961d37117c7765ca851584677b57e514ae398fe1c0bac717396f87aba9d1c0255bed1127a7f4b064989c9798558ff6330e7bfccbff14abc85de9f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'hf308602d7f48af567f6ab67e6ce0e4cf5273154f1828b2b5c9c55ef2c954d7b1ad99d34b6ccde55f50fd25685cffee3b3ac81c31761caa85b03b784b1884dc31939fb4aa682d42e2b503e97cc5e6f52da4ce2411c9202f1898167dbe79526147;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'h12216c9f9fd24d37cf742afcf50aeb5b41f508d77599c3ccb2acd2e500e76b468e9cc028a697e31ebf5a1254a757d58ef53c22be1acc44a1a0043d569542a6a54303c73dff826b0223a840781983018eca7fba5b7bdec769f4c8ecbf45b2108a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'h63bb3a07179483835b65ec6acbf93beb9f53d5597e4a965f42933726f1502b6548f3c2e369781acee8d8ac8e8bac461d1cf3fd92bb3d397313332ec550af8f3fec201998222c79de40f8694b74182d6f80c491a24d5295c8cd2e791fbd698595;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'h8378d90320680d5466becd872b7a36e5a8a426a9f32d767fa5ecf2201579fa8f1dda1628b644b8a0824d5ddc06d6885fab623209ae043366cd3cb743e6b5f366c8b1c55871e0ce373ad12392798ff59a8a1c3ecd4cd013539a355401165dd55;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'h173c36a8fb06904d73d2c3780c8191ae306f6405e386c2350700c5b1cd02a3c502451b52dcd2bd711ff81c4ce60e3823eedbb95a6ba1086c36168fa401814fd9997592c202493b09491c0343cd0468e7e09b24591abda0f6d8af0a9466ace7db;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'hd78082c9d6c959aef142796182fe72188e0dc5e132f55f1f4ec14dc83d9a3d697a1c6f0bc5af8867ad64e951da2316b3271920f7579daf9bb9ee177a3927dbd376aab3b4ff532c8200a7452205485422eddb701d9a4ed81b40fe0ec0139ec4b8;
        #1
        $finish();
    end
endmodule
