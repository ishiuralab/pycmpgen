module compressor2_1_64_16_shiftregister(input clk, input in_data0, input in_data1, input in_data2, input in_data3, input in_data4, input in_data5, input in_data6, input in_data7, input in_data8, input in_data9, input in_data10, input in_data11, input in_data12, input in_data13, input in_data14, input in_data15, input in_data16, input in_data17, input in_data18, input in_data19, input in_data20, input in_data21, input in_data22, input in_data23, input in_data24, input in_data25, input in_data26, input in_data27, input in_data28, input in_data29, input in_data30, input in_data31, input in_data32, input in_data33, input in_data34, input in_data35, input in_data36, input in_data37, input in_data38, input in_data39, input in_data40, input in_data41, input in_data42, input in_data43, input in_data44, input in_data45, input in_data46, input in_data47, input in_data48, input in_data49, input in_data50, input in_data51, input in_data52, input in_data53, input in_data54, input in_data55, input in_data56, input in_data57, input in_data58, input in_data59, input in_data60, input in_data61, input in_data62, input in_data63, output [21:0]dst);
    reg [15:0] src0;
    reg [15:0] src1;
    reg [15:0] src2;
    reg [15:0] src3;
    reg [15:0] src4;
    reg [15:0] src5;
    reg [15:0] src6;
    reg [15:0] src7;
    reg [15:0] src8;
    reg [15:0] src9;
    reg [15:0] src10;
    reg [15:0] src11;
    reg [15:0] src12;
    reg [15:0] src13;
    reg [15:0] src14;
    reg [15:0] src15;
    reg [15:0] src16;
    reg [15:0] src17;
    reg [15:0] src18;
    reg [15:0] src19;
    reg [15:0] src20;
    reg [15:0] src21;
    reg [15:0] src22;
    reg [15:0] src23;
    reg [15:0] src24;
    reg [15:0] src25;
    reg [15:0] src26;
    reg [15:0] src27;
    reg [15:0] src28;
    reg [15:0] src29;
    reg [15:0] src30;
    reg [15:0] src31;
    reg [15:0] src32;
    reg [15:0] src33;
    reg [15:0] src34;
    reg [15:0] src35;
    reg [15:0] src36;
    reg [15:0] src37;
    reg [15:0] src38;
    reg [15:0] src39;
    reg [15:0] src40;
    reg [15:0] src41;
    reg [15:0] src42;
    reg [15:0] src43;
    reg [15:0] src44;
    reg [15:0] src45;
    reg [15:0] src46;
    reg [15:0] src47;
    reg [15:0] src48;
    reg [15:0] src49;
    reg [15:0] src50;
    reg [15:0] src51;
    reg [15:0] src52;
    reg [15:0] src53;
    reg [15:0] src54;
    reg [15:0] src55;
    reg [15:0] src56;
    reg [15:0] src57;
    reg [15:0] src58;
    reg [15:0] src59;
    reg [15:0] src60;
    reg [15:0] src61;
    reg [15:0] src62;
    reg [15:0] src63;
    compressor2_1_64_16 compressor2_1_64_16(.src0(src0), .src1(src1), .src2(src2), .src3(src3), .src4(src4), .src5(src5), .src6(src6), .src7(src7), .src8(src8), .src9(src9), .src10(src10), .src11(src11), .src12(src12), .src13(src13), .src14(src14), .src15(src15), .src16(src16), .src17(src17), .src18(src18), .src19(src19), .src20(src20), .src21(src21), .src22(src22), .src23(src23), .src24(src24), .src25(src25), .src26(src26), .src27(src27), .src28(src28), .src29(src29), .src30(src30), .src31(src31), .src32(src32), .src33(src33), .src34(src34), .src35(src35), .src36(src36), .src37(src37), .src38(src38), .src39(src39), .src40(src40), .src41(src41), .src42(src42), .src43(src43), .src44(src44), .src45(src45), .src46(src46), .src47(src47), .src48(src48), .src49(src49), .src50(src50), .src51(src51), .src52(src52), .src53(src53), .src54(src54), .src55(src55), .src56(src56), .src57(src57), .src58(src58), .src59(src59), .src60(src60), .src61(src61), .src62(src62), .src63(src63), .dst(dst));
    initial begin
        src0 <= 0;
        src1 <= 0;
        src2 <= 0;
        src3 <= 0;
        src4 <= 0;
        src5 <= 0;
        src6 <= 0;
        src7 <= 0;
        src8 <= 0;
        src9 <= 0;
        src10 <= 0;
        src11 <= 0;
        src12 <= 0;
        src13 <= 0;
        src14 <= 0;
        src15 <= 0;
        src16 <= 0;
        src17 <= 0;
        src18 <= 0;
        src19 <= 0;
        src20 <= 0;
        src21 <= 0;
        src22 <= 0;
        src23 <= 0;
        src24 <= 0;
        src25 <= 0;
        src26 <= 0;
        src27 <= 0;
        src28 <= 0;
        src29 <= 0;
        src30 <= 0;
        src31 <= 0;
        src32 <= 0;
        src33 <= 0;
        src34 <= 0;
        src35 <= 0;
        src36 <= 0;
        src37 <= 0;
        src38 <= 0;
        src39 <= 0;
        src40 <= 0;
        src41 <= 0;
        src42 <= 0;
        src43 <= 0;
        src44 <= 0;
        src45 <= 0;
        src46 <= 0;
        src47 <= 0;
        src48 <= 0;
        src49 <= 0;
        src50 <= 0;
        src51 <= 0;
        src52 <= 0;
        src53 <= 0;
        src54 <= 0;
        src55 <= 0;
        src56 <= 0;
        src57 <= 0;
        src58 <= 0;
        src59 <= 0;
        src60 <= 0;
        src61 <= 0;
        src62 <= 0;
        src63 <= 0;
    end
    always @(posedge clk) begin
        src0 <= {src0[14:0], in_data0};
        src1 <= {src1[14:0], in_data1};
        src2 <= {src2[14:0], in_data2};
        src3 <= {src3[14:0], in_data3};
        src4 <= {src4[14:0], in_data4};
        src5 <= {src5[14:0], in_data5};
        src6 <= {src6[14:0], in_data6};
        src7 <= {src7[14:0], in_data7};
        src8 <= {src8[14:0], in_data8};
        src9 <= {src9[14:0], in_data9};
        src10 <= {src10[14:0], in_data10};
        src11 <= {src11[14:0], in_data11};
        src12 <= {src12[14:0], in_data12};
        src13 <= {src13[14:0], in_data13};
        src14 <= {src14[14:0], in_data14};
        src15 <= {src15[14:0], in_data15};
        src16 <= {src16[14:0], in_data16};
        src17 <= {src17[14:0], in_data17};
        src18 <= {src18[14:0], in_data18};
        src19 <= {src19[14:0], in_data19};
        src20 <= {src20[14:0], in_data20};
        src21 <= {src21[14:0], in_data21};
        src22 <= {src22[14:0], in_data22};
        src23 <= {src23[14:0], in_data23};
        src24 <= {src24[14:0], in_data24};
        src25 <= {src25[14:0], in_data25};
        src26 <= {src26[14:0], in_data26};
        src27 <= {src27[14:0], in_data27};
        src28 <= {src28[14:0], in_data28};
        src29 <= {src29[14:0], in_data29};
        src30 <= {src30[14:0], in_data30};
        src31 <= {src31[14:0], in_data31};
        src32 <= {src32[14:0], in_data32};
        src33 <= {src33[14:0], in_data33};
        src34 <= {src34[14:0], in_data34};
        src35 <= {src35[14:0], in_data35};
        src36 <= {src36[14:0], in_data36};
        src37 <= {src37[14:0], in_data37};
        src38 <= {src38[14:0], in_data38};
        src39 <= {src39[14:0], in_data39};
        src40 <= {src40[14:0], in_data40};
        src41 <= {src41[14:0], in_data41};
        src42 <= {src42[14:0], in_data42};
        src43 <= {src43[14:0], in_data43};
        src44 <= {src44[14:0], in_data44};
        src45 <= {src45[14:0], in_data45};
        src46 <= {src46[14:0], in_data46};
        src47 <= {src47[14:0], in_data47};
        src48 <= {src48[14:0], in_data48};
        src49 <= {src49[14:0], in_data49};
        src50 <= {src50[14:0], in_data50};
        src51 <= {src51[14:0], in_data51};
        src52 <= {src52[14:0], in_data52};
        src53 <= {src53[14:0], in_data53};
        src54 <= {src54[14:0], in_data54};
        src55 <= {src55[14:0], in_data55};
        src56 <= {src56[14:0], in_data56};
        src57 <= {src57[14:0], in_data57};
        src58 <= {src58[14:0], in_data58};
        src59 <= {src59[14:0], in_data59};
        src60 <= {src60[14:0], in_data60};
        src61 <= {src61[14:0], in_data61};
        src62 <= {src62[14:0], in_data62};
        src63 <= {src63[14:0], in_data63};
    end
endmodule

module compressor2_1_64_16(
    input [15:0]src0,
    input [15:0]src1,
    input [15:0]src2,
    input [15:0]src3,
    input [15:0]src4,
    input [15:0]src5,
    input [15:0]src6,
    input [15:0]src7,
    input [15:0]src8,
    input [15:0]src9,
    input [15:0]src10,
    input [15:0]src11,
    input [15:0]src12,
    input [15:0]src13,
    input [15:0]src14,
    input [15:0]src15,
    input [15:0]src16,
    input [15:0]src17,
    input [15:0]src18,
    input [15:0]src19,
    input [15:0]src20,
    input [15:0]src21,
    input [15:0]src22,
    input [15:0]src23,
    input [15:0]src24,
    input [15:0]src25,
    input [15:0]src26,
    input [15:0]src27,
    input [15:0]src28,
    input [15:0]src29,
    input [15:0]src30,
    input [15:0]src31,
    input [15:0]src32,
    input [15:0]src33,
    input [15:0]src34,
    input [15:0]src35,
    input [15:0]src36,
    input [15:0]src37,
    input [15:0]src38,
    input [15:0]src39,
    input [15:0]src40,
    input [15:0]src41,
    input [15:0]src42,
    input [15:0]src43,
    input [15:0]src44,
    input [15:0]src45,
    input [15:0]src46,
    input [15:0]src47,
    input [15:0]src48,
    input [15:0]src49,
    input [15:0]src50,
    input [15:0]src51,
    input [15:0]src52,
    input [15:0]src53,
    input [15:0]src54,
    input [15:0]src55,
    input [15:0]src56,
    input [15:0]src57,
    input [15:0]src58,
    input [15:0]src59,
    input [15:0]src60,
    input [15:0]src61,
    input [15:0]src62,
    input [15:0]src63,
    output [21:0]dst);

    wire [1:0] comp_out0;
    wire [1:0] comp_out1;
    wire [1:0] comp_out2;
    wire [1:0] comp_out3;
    wire [1:0] comp_out4;
    wire [1:0] comp_out5;
    wire [1:0] comp_out6;
    wire [1:0] comp_out7;
    wire [1:0] comp_out8;
    wire [1:0] comp_out9;
    wire [1:0] comp_out10;
    wire [1:0] comp_out11;
    wire [1:0] comp_out12;
    wire [1:0] comp_out13;
    wire [1:0] comp_out14;
    wire [1:0] comp_out15;
    wire [1:0] comp_out16;
    wire [1:0] comp_out17;
    wire [1:0] comp_out18;
    wire [0:0] comp_out19;
    wire [1:0] comp_out20;
    wire [0:0] comp_out21;
    wire [22:0] out;
    compressor compressor_inst(
        .src0({src63[0], src62[0], src61[0], src60[0], src59[0], src58[0], src57[0], src56[0], src55[0], src54[0], src53[0], src52[0], src51[0], src50[0], src49[0], src48[0], src47[0], src46[0], src45[0], src44[0], src43[0], src42[0], src41[0], src40[0], src39[0], src38[0], src37[0], src36[0], src35[0], src34[0], src33[0], src32[0], src31[0], src30[0], src29[0], src28[0], src27[0], src26[0], src25[0], src24[0], src23[0], src22[0], src21[0], src20[0], src19[0], src18[0], src17[0], src16[0], src15[0], src14[0], src13[0], src12[0], src11[0], src10[0], src9[0], src8[0], src7[0], src6[0], src5[0], src4[0], src3[0], src2[0], src1[0], src0[0]}),
        .src1({src63[1], src62[1], src61[1], src60[1], src59[1], src58[1], src57[1], src56[1], src55[1], src54[1], src53[1], src52[1], src51[1], src50[1], src49[1], src48[1], src47[1], src46[1], src45[1], src44[1], src43[1], src42[1], src41[1], src40[1], src39[1], src38[1], src37[1], src36[1], src35[1], src34[1], src33[1], src32[1], src31[1], src30[1], src29[1], src28[1], src27[1], src26[1], src25[1], src24[1], src23[1], src22[1], src21[1], src20[1], src19[1], src18[1], src17[1], src16[1], src15[1], src14[1], src13[1], src12[1], src11[1], src10[1], src9[1], src8[1], src7[1], src6[1], src5[1], src4[1], src3[1], src2[1], src1[1], src0[1]}),
        .src2({src63[2], src62[2], src61[2], src60[2], src59[2], src58[2], src57[2], src56[2], src55[2], src54[2], src53[2], src52[2], src51[2], src50[2], src49[2], src48[2], src47[2], src46[2], src45[2], src44[2], src43[2], src42[2], src41[2], src40[2], src39[2], src38[2], src37[2], src36[2], src35[2], src34[2], src33[2], src32[2], src31[2], src30[2], src29[2], src28[2], src27[2], src26[2], src25[2], src24[2], src23[2], src22[2], src21[2], src20[2], src19[2], src18[2], src17[2], src16[2], src15[2], src14[2], src13[2], src12[2], src11[2], src10[2], src9[2], src8[2], src7[2], src6[2], src5[2], src4[2], src3[2], src2[2], src1[2], src0[2]}),
        .src3({src63[3], src62[3], src61[3], src60[3], src59[3], src58[3], src57[3], src56[3], src55[3], src54[3], src53[3], src52[3], src51[3], src50[3], src49[3], src48[3], src47[3], src46[3], src45[3], src44[3], src43[3], src42[3], src41[3], src40[3], src39[3], src38[3], src37[3], src36[3], src35[3], src34[3], src33[3], src32[3], src31[3], src30[3], src29[3], src28[3], src27[3], src26[3], src25[3], src24[3], src23[3], src22[3], src21[3], src20[3], src19[3], src18[3], src17[3], src16[3], src15[3], src14[3], src13[3], src12[3], src11[3], src10[3], src9[3], src8[3], src7[3], src6[3], src5[3], src4[3], src3[3], src2[3], src1[3], src0[3]}),
        .src4({src63[4], src62[4], src61[4], src60[4], src59[4], src58[4], src57[4], src56[4], src55[4], src54[4], src53[4], src52[4], src51[4], src50[4], src49[4], src48[4], src47[4], src46[4], src45[4], src44[4], src43[4], src42[4], src41[4], src40[4], src39[4], src38[4], src37[4], src36[4], src35[4], src34[4], src33[4], src32[4], src31[4], src30[4], src29[4], src28[4], src27[4], src26[4], src25[4], src24[4], src23[4], src22[4], src21[4], src20[4], src19[4], src18[4], src17[4], src16[4], src15[4], src14[4], src13[4], src12[4], src11[4], src10[4], src9[4], src8[4], src7[4], src6[4], src5[4], src4[4], src3[4], src2[4], src1[4], src0[4]}),
        .src5({src63[5], src62[5], src61[5], src60[5], src59[5], src58[5], src57[5], src56[5], src55[5], src54[5], src53[5], src52[5], src51[5], src50[5], src49[5], src48[5], src47[5], src46[5], src45[5], src44[5], src43[5], src42[5], src41[5], src40[5], src39[5], src38[5], src37[5], src36[5], src35[5], src34[5], src33[5], src32[5], src31[5], src30[5], src29[5], src28[5], src27[5], src26[5], src25[5], src24[5], src23[5], src22[5], src21[5], src20[5], src19[5], src18[5], src17[5], src16[5], src15[5], src14[5], src13[5], src12[5], src11[5], src10[5], src9[5], src8[5], src7[5], src6[5], src5[5], src4[5], src3[5], src2[5], src1[5], src0[5]}),
        .src6({src63[6], src62[6], src61[6], src60[6], src59[6], src58[6], src57[6], src56[6], src55[6], src54[6], src53[6], src52[6], src51[6], src50[6], src49[6], src48[6], src47[6], src46[6], src45[6], src44[6], src43[6], src42[6], src41[6], src40[6], src39[6], src38[6], src37[6], src36[6], src35[6], src34[6], src33[6], src32[6], src31[6], src30[6], src29[6], src28[6], src27[6], src26[6], src25[6], src24[6], src23[6], src22[6], src21[6], src20[6], src19[6], src18[6], src17[6], src16[6], src15[6], src14[6], src13[6], src12[6], src11[6], src10[6], src9[6], src8[6], src7[6], src6[6], src5[6], src4[6], src3[6], src2[6], src1[6], src0[6]}),
        .src7({src63[7], src62[7], src61[7], src60[7], src59[7], src58[7], src57[7], src56[7], src55[7], src54[7], src53[7], src52[7], src51[7], src50[7], src49[7], src48[7], src47[7], src46[7], src45[7], src44[7], src43[7], src42[7], src41[7], src40[7], src39[7], src38[7], src37[7], src36[7], src35[7], src34[7], src33[7], src32[7], src31[7], src30[7], src29[7], src28[7], src27[7], src26[7], src25[7], src24[7], src23[7], src22[7], src21[7], src20[7], src19[7], src18[7], src17[7], src16[7], src15[7], src14[7], src13[7], src12[7], src11[7], src10[7], src9[7], src8[7], src7[7], src6[7], src5[7], src4[7], src3[7], src2[7], src1[7], src0[7]}),
        .src8({src63[8], src62[8], src61[8], src60[8], src59[8], src58[8], src57[8], src56[8], src55[8], src54[8], src53[8], src52[8], src51[8], src50[8], src49[8], src48[8], src47[8], src46[8], src45[8], src44[8], src43[8], src42[8], src41[8], src40[8], src39[8], src38[8], src37[8], src36[8], src35[8], src34[8], src33[8], src32[8], src31[8], src30[8], src29[8], src28[8], src27[8], src26[8], src25[8], src24[8], src23[8], src22[8], src21[8], src20[8], src19[8], src18[8], src17[8], src16[8], src15[8], src14[8], src13[8], src12[8], src11[8], src10[8], src9[8], src8[8], src7[8], src6[8], src5[8], src4[8], src3[8], src2[8], src1[8], src0[8]}),
        .src9({src63[9], src62[9], src61[9], src60[9], src59[9], src58[9], src57[9], src56[9], src55[9], src54[9], src53[9], src52[9], src51[9], src50[9], src49[9], src48[9], src47[9], src46[9], src45[9], src44[9], src43[9], src42[9], src41[9], src40[9], src39[9], src38[9], src37[9], src36[9], src35[9], src34[9], src33[9], src32[9], src31[9], src30[9], src29[9], src28[9], src27[9], src26[9], src25[9], src24[9], src23[9], src22[9], src21[9], src20[9], src19[9], src18[9], src17[9], src16[9], src15[9], src14[9], src13[9], src12[9], src11[9], src10[9], src9[9], src8[9], src7[9], src6[9], src5[9], src4[9], src3[9], src2[9], src1[9], src0[9]}),
        .src10({src63[10], src62[10], src61[10], src60[10], src59[10], src58[10], src57[10], src56[10], src55[10], src54[10], src53[10], src52[10], src51[10], src50[10], src49[10], src48[10], src47[10], src46[10], src45[10], src44[10], src43[10], src42[10], src41[10], src40[10], src39[10], src38[10], src37[10], src36[10], src35[10], src34[10], src33[10], src32[10], src31[10], src30[10], src29[10], src28[10], src27[10], src26[10], src25[10], src24[10], src23[10], src22[10], src21[10], src20[10], src19[10], src18[10], src17[10], src16[10], src15[10], src14[10], src13[10], src12[10], src11[10], src10[10], src9[10], src8[10], src7[10], src6[10], src5[10], src4[10], src3[10], src2[10], src1[10], src0[10]}),
        .src11({src63[11], src62[11], src61[11], src60[11], src59[11], src58[11], src57[11], src56[11], src55[11], src54[11], src53[11], src52[11], src51[11], src50[11], src49[11], src48[11], src47[11], src46[11], src45[11], src44[11], src43[11], src42[11], src41[11], src40[11], src39[11], src38[11], src37[11], src36[11], src35[11], src34[11], src33[11], src32[11], src31[11], src30[11], src29[11], src28[11], src27[11], src26[11], src25[11], src24[11], src23[11], src22[11], src21[11], src20[11], src19[11], src18[11], src17[11], src16[11], src15[11], src14[11], src13[11], src12[11], src11[11], src10[11], src9[11], src8[11], src7[11], src6[11], src5[11], src4[11], src3[11], src2[11], src1[11], src0[11]}),
        .src12({src63[12], src62[12], src61[12], src60[12], src59[12], src58[12], src57[12], src56[12], src55[12], src54[12], src53[12], src52[12], src51[12], src50[12], src49[12], src48[12], src47[12], src46[12], src45[12], src44[12], src43[12], src42[12], src41[12], src40[12], src39[12], src38[12], src37[12], src36[12], src35[12], src34[12], src33[12], src32[12], src31[12], src30[12], src29[12], src28[12], src27[12], src26[12], src25[12], src24[12], src23[12], src22[12], src21[12], src20[12], src19[12], src18[12], src17[12], src16[12], src15[12], src14[12], src13[12], src12[12], src11[12], src10[12], src9[12], src8[12], src7[12], src6[12], src5[12], src4[12], src3[12], src2[12], src1[12], src0[12]}),
        .src13({src63[13], src62[13], src61[13], src60[13], src59[13], src58[13], src57[13], src56[13], src55[13], src54[13], src53[13], src52[13], src51[13], src50[13], src49[13], src48[13], src47[13], src46[13], src45[13], src44[13], src43[13], src42[13], src41[13], src40[13], src39[13], src38[13], src37[13], src36[13], src35[13], src34[13], src33[13], src32[13], src31[13], src30[13], src29[13], src28[13], src27[13], src26[13], src25[13], src24[13], src23[13], src22[13], src21[13], src20[13], src19[13], src18[13], src17[13], src16[13], src15[13], src14[13], src13[13], src12[13], src11[13], src10[13], src9[13], src8[13], src7[13], src6[13], src5[13], src4[13], src3[13], src2[13], src1[13], src0[13]}),
        .src14({src63[14], src62[14], src61[14], src60[14], src59[14], src58[14], src57[14], src56[14], src55[14], src54[14], src53[14], src52[14], src51[14], src50[14], src49[14], src48[14], src47[14], src46[14], src45[14], src44[14], src43[14], src42[14], src41[14], src40[14], src39[14], src38[14], src37[14], src36[14], src35[14], src34[14], src33[14], src32[14], src31[14], src30[14], src29[14], src28[14], src27[14], src26[14], src25[14], src24[14], src23[14], src22[14], src21[14], src20[14], src19[14], src18[14], src17[14], src16[14], src15[14], src14[14], src13[14], src12[14], src11[14], src10[14], src9[14], src8[14], src7[14], src6[14], src5[14], src4[14], src3[14], src2[14], src1[14], src0[14]}),
        .src15({src63[15], src62[15], src61[15], src60[15], src59[15], src58[15], src57[15], src56[15], src55[15], src54[15], src53[15], src52[15], src51[15], src50[15], src49[15], src48[15], src47[15], src46[15], src45[15], src44[15], src43[15], src42[15], src41[15], src40[15], src39[15], src38[15], src37[15], src36[15], src35[15], src34[15], src33[15], src32[15], src31[15], src30[15], src29[15], src28[15], src27[15], src26[15], src25[15], src24[15], src23[15], src22[15], src21[15], src20[15], src19[15], src18[15], src17[15], src16[15], src15[15], src14[15], src13[15], src12[15], src11[15], src10[15], src9[15], src8[15], src7[15], src6[15], src5[15], src4[15], src3[15], src2[15], src1[15], src0[15]}),
        .dst0(comp_out0),
        .dst1(comp_out1),
        .dst2(comp_out2),
        .dst3(comp_out3),
        .dst4(comp_out4),
        .dst5(comp_out5),
        .dst6(comp_out6),
        .dst7(comp_out7),
        .dst8(comp_out8),
        .dst9(comp_out9),
        .dst10(comp_out10),
        .dst11(comp_out11),
        .dst12(comp_out12),
        .dst13(comp_out13),
        .dst14(comp_out14),
        .dst15(comp_out15),
        .dst16(comp_out16),
        .dst17(comp_out17),
        .dst18(comp_out18),
        .dst19(comp_out19),
        .dst20(comp_out20),
        .dst21(comp_out21)
    );
    rowadder2_1_22 rowadder2_1inst(
        .src0({comp_out21[0], comp_out20[0], comp_out19[0], comp_out18[0], comp_out17[0], comp_out16[0], comp_out15[0], comp_out14[0], comp_out13[0], comp_out12[0], comp_out11[0], comp_out10[0], comp_out9[0], comp_out8[0], comp_out7[0], comp_out6[0], comp_out5[0], comp_out4[0], comp_out3[0], comp_out2[0], comp_out1[0], comp_out0[0]}),
        .src1({1'h0, comp_out20[1], 1'h0, comp_out18[1], comp_out17[1], comp_out16[1], comp_out15[1], comp_out14[1], comp_out13[1], comp_out12[1], comp_out11[1], comp_out10[1], comp_out9[1], comp_out8[1], comp_out7[1], comp_out6[1], comp_out5[1], comp_out4[1], comp_out3[1], comp_out2[1], comp_out1[1], comp_out0[1]}),
        .dst0(out)
    );
    assign dst = out[21:0];
endmodule
module compressor (
      input wire [63:0] src0,
      input wire [63:0] src1,
      input wire [63:0] src2,
      input wire [63:0] src3,
      input wire [63:0] src4,
      input wire [63:0] src5,
      input wire [63:0] src6,
      input wire [63:0] src7,
      input wire [63:0] src8,
      input wire [63:0] src9,
      input wire [63:0] src10,
      input wire [63:0] src11,
      input wire [63:0] src12,
      input wire [63:0] src13,
      input wire [63:0] src14,
      input wire [63:0] src15,
      output wire [1:0] dst0,
      output wire [1:0] dst1,
      output wire [1:0] dst2,
      output wire [1:0] dst3,
      output wire [1:0] dst4,
      output wire [1:0] dst5,
      output wire [1:0] dst6,
      output wire [1:0] dst7,
      output wire [1:0] dst8,
      output wire [1:0] dst9,
      output wire [1:0] dst10,
      output wire [1:0] dst11,
      output wire [1:0] dst12,
      output wire [1:0] dst13,
      output wire [1:0] dst14,
      output wire [1:0] dst15,
      output wire [1:0] dst16,
      output wire [1:0] dst17,
      output wire [1:0] dst18,
      output wire [0:0] dst19,
      output wire [1:0] dst20,
      output wire [0:0] dst21);

   wire [63:0] stage0_0;
   wire [63:0] stage0_1;
   wire [63:0] stage0_2;
   wire [63:0] stage0_3;
   wire [63:0] stage0_4;
   wire [63:0] stage0_5;
   wire [63:0] stage0_6;
   wire [63:0] stage0_7;
   wire [63:0] stage0_8;
   wire [63:0] stage0_9;
   wire [63:0] stage0_10;
   wire [63:0] stage0_11;
   wire [63:0] stage0_12;
   wire [63:0] stage0_13;
   wire [63:0] stage0_14;
   wire [63:0] stage0_15;
   wire [19:0] stage1_0;
   wire [29:0] stage1_1;
   wire [23:0] stage1_2;
   wire [26:0] stage1_3;
   wire [39:0] stage1_4;
   wire [28:0] stage1_5;
   wire [26:0] stage1_6;
   wire [22:0] stage1_7;
   wire [28:0] stage1_8;
   wire [29:0] stage1_9;
   wire [28:0] stage1_10;
   wire [23:0] stage1_11;
   wire [28:0] stage1_12;
   wire [32:0] stage1_13;
   wire [24:0] stage1_14;
   wire [23:0] stage1_15;
   wire [18:0] stage1_16;
   wire [9:0] stage1_17;
   wire [3:0] stage2_0;
   wire [21:0] stage2_1;
   wire [7:0] stage2_2;
   wire [10:0] stage2_3;
   wire [15:0] stage2_4;
   wire [17:0] stage2_5;
   wire [11:0] stage2_6;
   wire [11:0] stage2_7;
   wire [15:0] stage2_8;
   wire [7:0] stage2_9;
   wire [12:0] stage2_10;
   wire [17:0] stage2_11;
   wire [7:0] stage2_12;
   wire [18:0] stage2_13;
   wire [23:0] stage2_14;
   wire [7:0] stage2_15;
   wire [12:0] stage2_16;
   wire [5:0] stage2_17;
   wire [3:0] stage2_18;
   wire [1:0] stage2_19;
   wire [1:0] stage3_0;
   wire [6:0] stage3_1;
   wire [4:0] stage3_2;
   wire [5:0] stage3_3;
   wire [5:0] stage3_4;
   wire [9:0] stage3_5;
   wire [4:0] stage3_6;
   wire [3:0] stage3_7;
   wire [7:0] stage3_8;
   wire [6:0] stage3_9;
   wire [2:0] stage3_10;
   wire [6:0] stage3_11;
   wire [6:0] stage3_12;
   wire [4:0] stage3_13;
   wire [12:0] stage3_14;
   wire [7:0] stage3_15;
   wire [4:0] stage3_16;
   wire [2:0] stage3_17;
   wire [6:0] stage3_18;
   wire [2:0] stage3_19;
   wire [1:0] stage4_0;
   wire [1:0] stage4_1;
   wire [1:0] stage4_2;
   wire [1:0] stage4_3;
   wire [1:0] stage4_4;
   wire [5:0] stage4_5;
   wire [2:0] stage4_6;
   wire [3:0] stage4_7;
   wire [3:0] stage4_8;
   wire [3:0] stage4_9;
   wire [3:0] stage4_10;
   wire [1:0] stage4_11;
   wire [2:0] stage4_12;
   wire [2:0] stage4_13;
   wire [7:0] stage4_14;
   wire [3:0] stage4_15;
   wire [2:0] stage4_16;
   wire [3:0] stage4_17;
   wire [1:0] stage4_18;
   wire [3:0] stage4_19;
   wire [0:0] stage4_20;
   wire [1:0] stage5_0;
   wire [1:0] stage5_1;
   wire [1:0] stage5_2;
   wire [1:0] stage5_3;
   wire [1:0] stage5_4;
   wire [1:0] stage5_5;
   wire [1:0] stage5_6;
   wire [1:0] stage5_7;
   wire [1:0] stage5_8;
   wire [1:0] stage5_9;
   wire [1:0] stage5_10;
   wire [1:0] stage5_11;
   wire [1:0] stage5_12;
   wire [1:0] stage5_13;
   wire [1:0] stage5_14;
   wire [1:0] stage5_15;
   wire [1:0] stage5_16;
   wire [1:0] stage5_17;
   wire [1:0] stage5_18;
   wire [0:0] stage5_19;
   wire [1:0] stage5_20;
   wire [0:0] stage5_21;

   assign stage0_0 = src0;
   assign stage0_1 = src1;
   assign stage0_2 = src2;
   assign stage0_3 = src3;
   assign stage0_4 = src4;
   assign stage0_5 = src5;
   assign stage0_6 = src6;
   assign stage0_7 = src7;
   assign stage0_8 = src8;
   assign stage0_9 = src9;
   assign stage0_10 = src10;
   assign stage0_11 = src11;
   assign stage0_12 = src12;
   assign stage0_13 = src13;
   assign stage0_14 = src14;
   assign stage0_15 = src15;
   assign dst0 = stage5_0;
   assign dst1 = stage5_1;
   assign dst2 = stage5_2;
   assign dst3 = stage5_3;
   assign dst4 = stage5_4;
   assign dst5 = stage5_5;
   assign dst6 = stage5_6;
   assign dst7 = stage5_7;
   assign dst8 = stage5_8;
   assign dst9 = stage5_9;
   assign dst10 = stage5_10;
   assign dst11 = stage5_11;
   assign dst12 = stage5_12;
   assign dst13 = stage5_13;
   assign dst14 = stage5_14;
   assign dst15 = stage5_15;
   assign dst16 = stage5_16;
   assign dst17 = stage5_17;
   assign dst18 = stage5_18;
   assign dst19 = stage5_19;
   assign dst20 = stage5_20;
   assign dst21 = stage5_21;

   gpc2135_5 gpc0 (
      {stage0_0[0], stage0_0[1], stage0_0[2], stage0_0[3], stage0_0[4]},
      {stage0_1[0], stage0_1[1], stage0_1[2]},
      {stage0_2[0]},
      {stage0_3[0], stage0_3[1]},
      {stage1_4[0],stage1_3[0],stage1_2[0],stage1_1[0],stage1_0[0]}
   );
   gpc606_5 gpc1 (
      {stage0_0[5], stage0_0[6], stage0_0[7], stage0_0[8], stage0_0[9], stage0_0[10]},
      {stage0_2[1], stage0_2[2], stage0_2[3], stage0_2[4], stage0_2[5], stage0_2[6]},
      {stage1_4[1],stage1_3[1],stage1_2[1],stage1_1[1],stage1_0[1]}
   );
   gpc606_5 gpc2 (
      {stage0_0[11], stage0_0[12], stage0_0[13], stage0_0[14], stage0_0[15], stage0_0[16]},
      {stage0_2[7], stage0_2[8], stage0_2[9], stage0_2[10], stage0_2[11], stage0_2[12]},
      {stage1_4[2],stage1_3[2],stage1_2[2],stage1_1[2],stage1_0[2]}
   );
   gpc606_5 gpc3 (
      {stage0_0[17], stage0_0[18], stage0_0[19], stage0_0[20], stage0_0[21], stage0_0[22]},
      {stage0_2[13], stage0_2[14], stage0_2[15], stage0_2[16], stage0_2[17], stage0_2[18]},
      {stage1_4[3],stage1_3[3],stage1_2[3],stage1_1[3],stage1_0[3]}
   );
   gpc606_5 gpc4 (
      {stage0_0[23], stage0_0[24], stage0_0[25], stage0_0[26], stage0_0[27], stage0_0[28]},
      {stage0_2[19], stage0_2[20], stage0_2[21], stage0_2[22], stage0_2[23], stage0_2[24]},
      {stage1_4[4],stage1_3[4],stage1_2[4],stage1_1[4],stage1_0[4]}
   );
   gpc606_5 gpc5 (
      {stage0_0[29], stage0_0[30], stage0_0[31], stage0_0[32], stage0_0[33], stage0_0[34]},
      {stage0_2[25], stage0_2[26], stage0_2[27], stage0_2[28], stage0_2[29], stage0_2[30]},
      {stage1_4[5],stage1_3[5],stage1_2[5],stage1_1[5],stage1_0[5]}
   );
   gpc606_5 gpc6 (
      {stage0_0[35], stage0_0[36], stage0_0[37], stage0_0[38], stage0_0[39], stage0_0[40]},
      {stage0_2[31], stage0_2[32], stage0_2[33], stage0_2[34], stage0_2[35], stage0_2[36]},
      {stage1_4[6],stage1_3[6],stage1_2[6],stage1_1[6],stage1_0[6]}
   );
   gpc606_5 gpc7 (
      {stage0_0[41], stage0_0[42], stage0_0[43], stage0_0[44], stage0_0[45], stage0_0[46]},
      {stage0_2[37], stage0_2[38], stage0_2[39], stage0_2[40], stage0_2[41], stage0_2[42]},
      {stage1_4[7],stage1_3[7],stage1_2[7],stage1_1[7],stage1_0[7]}
   );
   gpc606_5 gpc8 (
      {stage0_0[47], stage0_0[48], stage0_0[49], stage0_0[50], stage0_0[51], stage0_0[52]},
      {stage0_2[43], stage0_2[44], stage0_2[45], stage0_2[46], stage0_2[47], stage0_2[48]},
      {stage1_4[8],stage1_3[8],stage1_2[8],stage1_1[8],stage1_0[8]}
   );
   gpc606_5 gpc9 (
      {stage0_1[3], stage0_1[4], stage0_1[5], stage0_1[6], stage0_1[7], stage0_1[8]},
      {stage0_3[2], stage0_3[3], stage0_3[4], stage0_3[5], stage0_3[6], stage0_3[7]},
      {stage1_5[0],stage1_4[9],stage1_3[9],stage1_2[9],stage1_1[9]}
   );
   gpc606_5 gpc10 (
      {stage0_1[9], stage0_1[10], stage0_1[11], stage0_1[12], stage0_1[13], stage0_1[14]},
      {stage0_3[8], stage0_3[9], stage0_3[10], stage0_3[11], stage0_3[12], stage0_3[13]},
      {stage1_5[1],stage1_4[10],stage1_3[10],stage1_2[10],stage1_1[10]}
   );
   gpc606_5 gpc11 (
      {stage0_1[15], stage0_1[16], stage0_1[17], stage0_1[18], stage0_1[19], stage0_1[20]},
      {stage0_3[14], stage0_3[15], stage0_3[16], stage0_3[17], stage0_3[18], stage0_3[19]},
      {stage1_5[2],stage1_4[11],stage1_3[11],stage1_2[11],stage1_1[11]}
   );
   gpc606_5 gpc12 (
      {stage0_1[21], stage0_1[22], stage0_1[23], stage0_1[24], stage0_1[25], stage0_1[26]},
      {stage0_3[20], stage0_3[21], stage0_3[22], stage0_3[23], stage0_3[24], stage0_3[25]},
      {stage1_5[3],stage1_4[12],stage1_3[12],stage1_2[12],stage1_1[12]}
   );
   gpc606_5 gpc13 (
      {stage0_1[27], stage0_1[28], stage0_1[29], stage0_1[30], stage0_1[31], stage0_1[32]},
      {stage0_3[26], stage0_3[27], stage0_3[28], stage0_3[29], stage0_3[30], stage0_3[31]},
      {stage1_5[4],stage1_4[13],stage1_3[13],stage1_2[13],stage1_1[13]}
   );
   gpc606_5 gpc14 (
      {stage0_1[33], stage0_1[34], stage0_1[35], stage0_1[36], stage0_1[37], stage0_1[38]},
      {stage0_3[32], stage0_3[33], stage0_3[34], stage0_3[35], stage0_3[36], stage0_3[37]},
      {stage1_5[5],stage1_4[14],stage1_3[14],stage1_2[14],stage1_1[14]}
   );
   gpc606_5 gpc15 (
      {stage0_1[39], stage0_1[40], stage0_1[41], stage0_1[42], stage0_1[43], stage0_1[44]},
      {stage0_3[38], stage0_3[39], stage0_3[40], stage0_3[41], stage0_3[42], stage0_3[43]},
      {stage1_5[6],stage1_4[15],stage1_3[15],stage1_2[15],stage1_1[15]}
   );
   gpc606_5 gpc16 (
      {stage0_1[45], stage0_1[46], stage0_1[47], stage0_1[48], stage0_1[49], stage0_1[50]},
      {stage0_3[44], stage0_3[45], stage0_3[46], stage0_3[47], stage0_3[48], stage0_3[49]},
      {stage1_5[7],stage1_4[16],stage1_3[16],stage1_2[16],stage1_1[16]}
   );
   gpc615_5 gpc17 (
      {stage0_2[49], stage0_2[50], stage0_2[51], stage0_2[52], stage0_2[53]},
      {stage0_3[50]},
      {stage0_4[0], stage0_4[1], stage0_4[2], stage0_4[3], stage0_4[4], stage0_4[5]},
      {stage1_6[0],stage1_5[8],stage1_4[17],stage1_3[17],stage1_2[17]}
   );
   gpc615_5 gpc18 (
      {stage0_2[54], stage0_2[55], stage0_2[56], stage0_2[57], stage0_2[58]},
      {stage0_3[51]},
      {stage0_4[6], stage0_4[7], stage0_4[8], stage0_4[9], stage0_4[10], stage0_4[11]},
      {stage1_6[1],stage1_5[9],stage1_4[18],stage1_3[18],stage1_2[18]}
   );
   gpc615_5 gpc19 (
      {stage0_3[52], stage0_3[53], stage0_3[54], stage0_3[55], stage0_3[56]},
      {stage0_4[12]},
      {stage0_5[0], stage0_5[1], stage0_5[2], stage0_5[3], stage0_5[4], stage0_5[5]},
      {stage1_7[0],stage1_6[2],stage1_5[10],stage1_4[19],stage1_3[19]}
   );
   gpc606_5 gpc20 (
      {stage0_4[13], stage0_4[14], stage0_4[15], stage0_4[16], stage0_4[17], stage0_4[18]},
      {stage0_6[0], stage0_6[1], stage0_6[2], stage0_6[3], stage0_6[4], stage0_6[5]},
      {stage1_8[0],stage1_7[1],stage1_6[3],stage1_5[11],stage1_4[20]}
   );
   gpc606_5 gpc21 (
      {stage0_4[19], stage0_4[20], stage0_4[21], stage0_4[22], stage0_4[23], stage0_4[24]},
      {stage0_6[6], stage0_6[7], stage0_6[8], stage0_6[9], stage0_6[10], stage0_6[11]},
      {stage1_8[1],stage1_7[2],stage1_6[4],stage1_5[12],stage1_4[21]}
   );
   gpc606_5 gpc22 (
      {stage0_4[25], stage0_4[26], stage0_4[27], stage0_4[28], stage0_4[29], stage0_4[30]},
      {stage0_6[12], stage0_6[13], stage0_6[14], stage0_6[15], stage0_6[16], stage0_6[17]},
      {stage1_8[2],stage1_7[3],stage1_6[5],stage1_5[13],stage1_4[22]}
   );
   gpc615_5 gpc23 (
      {stage0_4[31], stage0_4[32], stage0_4[33], stage0_4[34], stage0_4[35]},
      {stage0_5[6]},
      {stage0_6[18], stage0_6[19], stage0_6[20], stage0_6[21], stage0_6[22], stage0_6[23]},
      {stage1_8[3],stage1_7[4],stage1_6[6],stage1_5[14],stage1_4[23]}
   );
   gpc615_5 gpc24 (
      {stage0_4[36], stage0_4[37], stage0_4[38], stage0_4[39], stage0_4[40]},
      {stage0_5[7]},
      {stage0_6[24], stage0_6[25], stage0_6[26], stage0_6[27], stage0_6[28], stage0_6[29]},
      {stage1_8[4],stage1_7[5],stage1_6[7],stage1_5[15],stage1_4[24]}
   );
   gpc615_5 gpc25 (
      {stage0_4[41], stage0_4[42], stage0_4[43], stage0_4[44], stage0_4[45]},
      {stage0_5[8]},
      {stage0_6[30], stage0_6[31], stage0_6[32], stage0_6[33], stage0_6[34], stage0_6[35]},
      {stage1_8[5],stage1_7[6],stage1_6[8],stage1_5[16],stage1_4[25]}
   );
   gpc615_5 gpc26 (
      {stage0_4[46], stage0_4[47], stage0_4[48], stage0_4[49], stage0_4[50]},
      {stage0_5[9]},
      {stage0_6[36], stage0_6[37], stage0_6[38], stage0_6[39], stage0_6[40], stage0_6[41]},
      {stage1_8[6],stage1_7[7],stage1_6[9],stage1_5[17],stage1_4[26]}
   );
   gpc606_5 gpc27 (
      {stage0_5[10], stage0_5[11], stage0_5[12], stage0_5[13], stage0_5[14], stage0_5[15]},
      {stage0_7[0], stage0_7[1], stage0_7[2], stage0_7[3], stage0_7[4], stage0_7[5]},
      {stage1_9[0],stage1_8[7],stage1_7[8],stage1_6[10],stage1_5[18]}
   );
   gpc606_5 gpc28 (
      {stage0_5[16], stage0_5[17], stage0_5[18], stage0_5[19], stage0_5[20], stage0_5[21]},
      {stage0_7[6], stage0_7[7], stage0_7[8], stage0_7[9], stage0_7[10], stage0_7[11]},
      {stage1_9[1],stage1_8[8],stage1_7[9],stage1_6[11],stage1_5[19]}
   );
   gpc606_5 gpc29 (
      {stage0_5[22], stage0_5[23], stage0_5[24], stage0_5[25], stage0_5[26], stage0_5[27]},
      {stage0_7[12], stage0_7[13], stage0_7[14], stage0_7[15], stage0_7[16], stage0_7[17]},
      {stage1_9[2],stage1_8[9],stage1_7[10],stage1_6[12],stage1_5[20]}
   );
   gpc606_5 gpc30 (
      {stage0_5[28], stage0_5[29], stage0_5[30], stage0_5[31], stage0_5[32], stage0_5[33]},
      {stage0_7[18], stage0_7[19], stage0_7[20], stage0_7[21], stage0_7[22], stage0_7[23]},
      {stage1_9[3],stage1_8[10],stage1_7[11],stage1_6[13],stage1_5[21]}
   );
   gpc606_5 gpc31 (
      {stage0_5[34], stage0_5[35], stage0_5[36], stage0_5[37], stage0_5[38], stage0_5[39]},
      {stage0_7[24], stage0_7[25], stage0_7[26], stage0_7[27], stage0_7[28], stage0_7[29]},
      {stage1_9[4],stage1_8[11],stage1_7[12],stage1_6[14],stage1_5[22]}
   );
   gpc606_5 gpc32 (
      {stage0_5[40], stage0_5[41], stage0_5[42], stage0_5[43], stage0_5[44], stage0_5[45]},
      {stage0_7[30], stage0_7[31], stage0_7[32], stage0_7[33], stage0_7[34], stage0_7[35]},
      {stage1_9[5],stage1_8[12],stage1_7[13],stage1_6[15],stage1_5[23]}
   );
   gpc606_5 gpc33 (
      {stage0_5[46], stage0_5[47], stage0_5[48], stage0_5[49], stage0_5[50], stage0_5[51]},
      {stage0_7[36], stage0_7[37], stage0_7[38], stage0_7[39], stage0_7[40], stage0_7[41]},
      {stage1_9[6],stage1_8[13],stage1_7[14],stage1_6[16],stage1_5[24]}
   );
   gpc615_5 gpc34 (
      {stage0_5[52], stage0_5[53], stage0_5[54], stage0_5[55], stage0_5[56]},
      {stage0_6[42]},
      {stage0_7[42], stage0_7[43], stage0_7[44], stage0_7[45], stage0_7[46], stage0_7[47]},
      {stage1_9[7],stage1_8[14],stage1_7[15],stage1_6[17],stage1_5[25]}
   );
   gpc615_5 gpc35 (
      {stage0_5[57], stage0_5[58], stage0_5[59], stage0_5[60], stage0_5[61]},
      {stage0_6[43]},
      {stage0_7[48], stage0_7[49], stage0_7[50], stage0_7[51], stage0_7[52], stage0_7[53]},
      {stage1_9[8],stage1_8[15],stage1_7[16],stage1_6[18],stage1_5[26]}
   );
   gpc615_5 gpc36 (
      {stage0_6[44], stage0_6[45], stage0_6[46], stage0_6[47], stage0_6[48]},
      {stage0_7[54]},
      {stage0_8[0], stage0_8[1], stage0_8[2], stage0_8[3], stage0_8[4], stage0_8[5]},
      {stage1_10[0],stage1_9[9],stage1_8[16],stage1_7[17],stage1_6[19]}
   );
   gpc615_5 gpc37 (
      {stage0_6[49], stage0_6[50], stage0_6[51], stage0_6[52], stage0_6[53]},
      {stage0_7[55]},
      {stage0_8[6], stage0_8[7], stage0_8[8], stage0_8[9], stage0_8[10], stage0_8[11]},
      {stage1_10[1],stage1_9[10],stage1_8[17],stage1_7[18],stage1_6[20]}
   );
   gpc615_5 gpc38 (
      {stage0_6[54], stage0_6[55], stage0_6[56], stage0_6[57], stage0_6[58]},
      {stage0_7[56]},
      {stage0_8[12], stage0_8[13], stage0_8[14], stage0_8[15], stage0_8[16], stage0_8[17]},
      {stage1_10[2],stage1_9[11],stage1_8[18],stage1_7[19],stage1_6[21]}
   );
   gpc615_5 gpc39 (
      {stage0_7[57], stage0_7[58], stage0_7[59], stage0_7[60], stage0_7[61]},
      {stage0_8[18]},
      {stage0_9[0], stage0_9[1], stage0_9[2], stage0_9[3], stage0_9[4], stage0_9[5]},
      {stage1_11[0],stage1_10[3],stage1_9[12],stage1_8[19],stage1_7[20]}
   );
   gpc606_5 gpc40 (
      {stage0_8[19], stage0_8[20], stage0_8[21], stage0_8[22], stage0_8[23], stage0_8[24]},
      {stage0_10[0], stage0_10[1], stage0_10[2], stage0_10[3], stage0_10[4], stage0_10[5]},
      {stage1_12[0],stage1_11[1],stage1_10[4],stage1_9[13],stage1_8[20]}
   );
   gpc606_5 gpc41 (
      {stage0_8[25], stage0_8[26], stage0_8[27], stage0_8[28], stage0_8[29], stage0_8[30]},
      {stage0_10[6], stage0_10[7], stage0_10[8], stage0_10[9], stage0_10[10], stage0_10[11]},
      {stage1_12[1],stage1_11[2],stage1_10[5],stage1_9[14],stage1_8[21]}
   );
   gpc606_5 gpc42 (
      {stage0_8[31], stage0_8[32], stage0_8[33], stage0_8[34], stage0_8[35], stage0_8[36]},
      {stage0_10[12], stage0_10[13], stage0_10[14], stage0_10[15], stage0_10[16], stage0_10[17]},
      {stage1_12[2],stage1_11[3],stage1_10[6],stage1_9[15],stage1_8[22]}
   );
   gpc606_5 gpc43 (
      {stage0_8[37], stage0_8[38], stage0_8[39], stage0_8[40], stage0_8[41], stage0_8[42]},
      {stage0_10[18], stage0_10[19], stage0_10[20], stage0_10[21], stage0_10[22], stage0_10[23]},
      {stage1_12[3],stage1_11[4],stage1_10[7],stage1_9[16],stage1_8[23]}
   );
   gpc615_5 gpc44 (
      {stage0_8[43], stage0_8[44], stage0_8[45], stage0_8[46], stage0_8[47]},
      {stage0_9[6]},
      {stage0_10[24], stage0_10[25], stage0_10[26], stage0_10[27], stage0_10[28], stage0_10[29]},
      {stage1_12[4],stage1_11[5],stage1_10[8],stage1_9[17],stage1_8[24]}
   );
   gpc615_5 gpc45 (
      {stage0_8[48], stage0_8[49], stage0_8[50], stage0_8[51], stage0_8[52]},
      {stage0_9[7]},
      {stage0_10[30], stage0_10[31], stage0_10[32], stage0_10[33], stage0_10[34], stage0_10[35]},
      {stage1_12[5],stage1_11[6],stage1_10[9],stage1_9[18],stage1_8[25]}
   );
   gpc615_5 gpc46 (
      {stage0_8[53], stage0_8[54], stage0_8[55], stage0_8[56], stage0_8[57]},
      {stage0_9[8]},
      {stage0_10[36], stage0_10[37], stage0_10[38], stage0_10[39], stage0_10[40], stage0_10[41]},
      {stage1_12[6],stage1_11[7],stage1_10[10],stage1_9[19],stage1_8[26]}
   );
   gpc615_5 gpc47 (
      {stage0_8[58], stage0_8[59], stage0_8[60], stage0_8[61], stage0_8[62]},
      {stage0_9[9]},
      {stage0_10[42], stage0_10[43], stage0_10[44], stage0_10[45], stage0_10[46], stage0_10[47]},
      {stage1_12[7],stage1_11[8],stage1_10[11],stage1_9[20],stage1_8[27]}
   );
   gpc606_5 gpc48 (
      {stage0_9[10], stage0_9[11], stage0_9[12], stage0_9[13], stage0_9[14], stage0_9[15]},
      {stage0_11[0], stage0_11[1], stage0_11[2], stage0_11[3], stage0_11[4], stage0_11[5]},
      {stage1_13[0],stage1_12[8],stage1_11[9],stage1_10[12],stage1_9[21]}
   );
   gpc606_5 gpc49 (
      {stage0_9[16], stage0_9[17], stage0_9[18], stage0_9[19], stage0_9[20], stage0_9[21]},
      {stage0_11[6], stage0_11[7], stage0_11[8], stage0_11[9], stage0_11[10], stage0_11[11]},
      {stage1_13[1],stage1_12[9],stage1_11[10],stage1_10[13],stage1_9[22]}
   );
   gpc606_5 gpc50 (
      {stage0_9[22], stage0_9[23], stage0_9[24], stage0_9[25], stage0_9[26], stage0_9[27]},
      {stage0_11[12], stage0_11[13], stage0_11[14], stage0_11[15], stage0_11[16], stage0_11[17]},
      {stage1_13[2],stage1_12[10],stage1_11[11],stage1_10[14],stage1_9[23]}
   );
   gpc606_5 gpc51 (
      {stage0_9[28], stage0_9[29], stage0_9[30], stage0_9[31], stage0_9[32], stage0_9[33]},
      {stage0_11[18], stage0_11[19], stage0_11[20], stage0_11[21], stage0_11[22], stage0_11[23]},
      {stage1_13[3],stage1_12[11],stage1_11[12],stage1_10[15],stage1_9[24]}
   );
   gpc606_5 gpc52 (
      {stage0_9[34], stage0_9[35], stage0_9[36], stage0_9[37], stage0_9[38], stage0_9[39]},
      {stage0_11[24], stage0_11[25], stage0_11[26], stage0_11[27], stage0_11[28], stage0_11[29]},
      {stage1_13[4],stage1_12[12],stage1_11[13],stage1_10[16],stage1_9[25]}
   );
   gpc606_5 gpc53 (
      {stage0_9[40], stage0_9[41], stage0_9[42], stage0_9[43], stage0_9[44], stage0_9[45]},
      {stage0_11[30], stage0_11[31], stage0_11[32], stage0_11[33], stage0_11[34], stage0_11[35]},
      {stage1_13[5],stage1_12[13],stage1_11[14],stage1_10[17],stage1_9[26]}
   );
   gpc606_5 gpc54 (
      {stage0_9[46], stage0_9[47], stage0_9[48], stage0_9[49], stage0_9[50], stage0_9[51]},
      {stage0_11[36], stage0_11[37], stage0_11[38], stage0_11[39], stage0_11[40], stage0_11[41]},
      {stage1_13[6],stage1_12[14],stage1_11[15],stage1_10[18],stage1_9[27]}
   );
   gpc606_5 gpc55 (
      {stage0_9[52], stage0_9[53], stage0_9[54], stage0_9[55], stage0_9[56], stage0_9[57]},
      {stage0_11[42], stage0_11[43], stage0_11[44], stage0_11[45], stage0_11[46], stage0_11[47]},
      {stage1_13[7],stage1_12[15],stage1_11[16],stage1_10[19],stage1_9[28]}
   );
   gpc606_5 gpc56 (
      {stage0_9[58], stage0_9[59], stage0_9[60], stage0_9[61], stage0_9[62], stage0_9[63]},
      {stage0_11[48], stage0_11[49], stage0_11[50], stage0_11[51], stage0_11[52], stage0_11[53]},
      {stage1_13[8],stage1_12[16],stage1_11[17],stage1_10[20],stage1_9[29]}
   );
   gpc615_5 gpc57 (
      {stage0_10[48], stage0_10[49], stage0_10[50], stage0_10[51], stage0_10[52]},
      {stage0_11[54]},
      {stage0_12[0], stage0_12[1], stage0_12[2], stage0_12[3], stage0_12[4], stage0_12[5]},
      {stage1_14[0],stage1_13[9],stage1_12[17],stage1_11[18],stage1_10[21]}
   );
   gpc615_5 gpc58 (
      {stage0_10[53], stage0_10[54], stage0_10[55], stage0_10[56], stage0_10[57]},
      {stage0_11[55]},
      {stage0_12[6], stage0_12[7], stage0_12[8], stage0_12[9], stage0_12[10], stage0_12[11]},
      {stage1_14[1],stage1_13[10],stage1_12[18],stage1_11[19],stage1_10[22]}
   );
   gpc615_5 gpc59 (
      {stage0_11[56], stage0_11[57], stage0_11[58], stage0_11[59], stage0_11[60]},
      {stage0_12[12]},
      {stage0_13[0], stage0_13[1], stage0_13[2], stage0_13[3], stage0_13[4], stage0_13[5]},
      {stage1_15[0],stage1_14[2],stage1_13[11],stage1_12[19],stage1_11[20]}
   );
   gpc606_5 gpc60 (
      {stage0_12[13], stage0_12[14], stage0_12[15], stage0_12[16], stage0_12[17], stage0_12[18]},
      {stage0_14[0], stage0_14[1], stage0_14[2], stage0_14[3], stage0_14[4], stage0_14[5]},
      {stage1_16[0],stage1_15[1],stage1_14[3],stage1_13[12],stage1_12[20]}
   );
   gpc606_5 gpc61 (
      {stage0_12[19], stage0_12[20], stage0_12[21], stage0_12[22], stage0_12[23], stage0_12[24]},
      {stage0_14[6], stage0_14[7], stage0_14[8], stage0_14[9], stage0_14[10], stage0_14[11]},
      {stage1_16[1],stage1_15[2],stage1_14[4],stage1_13[13],stage1_12[21]}
   );
   gpc606_5 gpc62 (
      {stage0_12[25], stage0_12[26], stage0_12[27], stage0_12[28], stage0_12[29], stage0_12[30]},
      {stage0_14[12], stage0_14[13], stage0_14[14], stage0_14[15], stage0_14[16], stage0_14[17]},
      {stage1_16[2],stage1_15[3],stage1_14[5],stage1_13[14],stage1_12[22]}
   );
   gpc606_5 gpc63 (
      {stage0_12[31], stage0_12[32], stage0_12[33], stage0_12[34], stage0_12[35], stage0_12[36]},
      {stage0_14[18], stage0_14[19], stage0_14[20], stage0_14[21], stage0_14[22], stage0_14[23]},
      {stage1_16[3],stage1_15[4],stage1_14[6],stage1_13[15],stage1_12[23]}
   );
   gpc606_5 gpc64 (
      {stage0_12[37], stage0_12[38], stage0_12[39], stage0_12[40], stage0_12[41], stage0_12[42]},
      {stage0_14[24], stage0_14[25], stage0_14[26], stage0_14[27], stage0_14[28], stage0_14[29]},
      {stage1_16[4],stage1_15[5],stage1_14[7],stage1_13[16],stage1_12[24]}
   );
   gpc606_5 gpc65 (
      {stage0_12[43], stage0_12[44], stage0_12[45], stage0_12[46], stage0_12[47], stage0_12[48]},
      {stage0_14[30], stage0_14[31], stage0_14[32], stage0_14[33], stage0_14[34], stage0_14[35]},
      {stage1_16[5],stage1_15[6],stage1_14[8],stage1_13[17],stage1_12[25]}
   );
   gpc615_5 gpc66 (
      {stage0_12[49], stage0_12[50], stage0_12[51], stage0_12[52], stage0_12[53]},
      {stage0_13[6]},
      {stage0_14[36], stage0_14[37], stage0_14[38], stage0_14[39], stage0_14[40], stage0_14[41]},
      {stage1_16[6],stage1_15[7],stage1_14[9],stage1_13[18],stage1_12[26]}
   );
   gpc615_5 gpc67 (
      {stage0_12[54], stage0_12[55], stage0_12[56], stage0_12[57], stage0_12[58]},
      {stage0_13[7]},
      {stage0_14[42], stage0_14[43], stage0_14[44], stage0_14[45], stage0_14[46], stage0_14[47]},
      {stage1_16[7],stage1_15[8],stage1_14[10],stage1_13[19],stage1_12[27]}
   );
   gpc615_5 gpc68 (
      {stage0_12[59], stage0_12[60], stage0_12[61], stage0_12[62], stage0_12[63]},
      {stage0_13[8]},
      {stage0_14[48], stage0_14[49], stage0_14[50], stage0_14[51], stage0_14[52], stage0_14[53]},
      {stage1_16[8],stage1_15[9],stage1_14[11],stage1_13[20],stage1_12[28]}
   );
   gpc606_5 gpc69 (
      {stage0_13[9], stage0_13[10], stage0_13[11], stage0_13[12], stage0_13[13], stage0_13[14]},
      {stage0_15[0], stage0_15[1], stage0_15[2], stage0_15[3], stage0_15[4], stage0_15[5]},
      {stage1_17[0],stage1_16[9],stage1_15[10],stage1_14[12],stage1_13[21]}
   );
   gpc606_5 gpc70 (
      {stage0_13[15], stage0_13[16], stage0_13[17], stage0_13[18], stage0_13[19], stage0_13[20]},
      {stage0_15[6], stage0_15[7], stage0_15[8], stage0_15[9], stage0_15[10], stage0_15[11]},
      {stage1_17[1],stage1_16[10],stage1_15[11],stage1_14[13],stage1_13[22]}
   );
   gpc606_5 gpc71 (
      {stage0_13[21], stage0_13[22], stage0_13[23], stage0_13[24], stage0_13[25], stage0_13[26]},
      {stage0_15[12], stage0_15[13], stage0_15[14], stage0_15[15], stage0_15[16], stage0_15[17]},
      {stage1_17[2],stage1_16[11],stage1_15[12],stage1_14[14],stage1_13[23]}
   );
   gpc615_5 gpc72 (
      {stage0_13[27], stage0_13[28], stage0_13[29], stage0_13[30], stage0_13[31]},
      {stage0_14[54]},
      {stage0_15[18], stage0_15[19], stage0_15[20], stage0_15[21], stage0_15[22], stage0_15[23]},
      {stage1_17[3],stage1_16[12],stage1_15[13],stage1_14[15],stage1_13[24]}
   );
   gpc615_5 gpc73 (
      {stage0_13[32], stage0_13[33], stage0_13[34], stage0_13[35], stage0_13[36]},
      {stage0_14[55]},
      {stage0_15[24], stage0_15[25], stage0_15[26], stage0_15[27], stage0_15[28], stage0_15[29]},
      {stage1_17[4],stage1_16[13],stage1_15[14],stage1_14[16],stage1_13[25]}
   );
   gpc615_5 gpc74 (
      {stage0_13[37], stage0_13[38], stage0_13[39], stage0_13[40], stage0_13[41]},
      {stage0_14[56]},
      {stage0_15[30], stage0_15[31], stage0_15[32], stage0_15[33], stage0_15[34], stage0_15[35]},
      {stage1_17[5],stage1_16[14],stage1_15[15],stage1_14[17],stage1_13[26]}
   );
   gpc615_5 gpc75 (
      {stage0_13[42], stage0_13[43], stage0_13[44], stage0_13[45], stage0_13[46]},
      {stage0_14[57]},
      {stage0_15[36], stage0_15[37], stage0_15[38], stage0_15[39], stage0_15[40], stage0_15[41]},
      {stage1_17[6],stage1_16[15],stage1_15[16],stage1_14[18],stage1_13[27]}
   );
   gpc615_5 gpc76 (
      {stage0_13[47], stage0_13[48], stage0_13[49], stage0_13[50], stage0_13[51]},
      {stage0_14[58]},
      {stage0_15[42], stage0_15[43], stage0_15[44], stage0_15[45], stage0_15[46], stage0_15[47]},
      {stage1_17[7],stage1_16[16],stage1_15[17],stage1_14[19],stage1_13[28]}
   );
   gpc615_5 gpc77 (
      {stage0_13[52], stage0_13[53], stage0_13[54], stage0_13[55], stage0_13[56]},
      {stage0_14[59]},
      {stage0_15[48], stage0_15[49], stage0_15[50], stage0_15[51], stage0_15[52], stage0_15[53]},
      {stage1_17[8],stage1_16[17],stage1_15[18],stage1_14[20],stage1_13[29]}
   );
   gpc615_5 gpc78 (
      {stage0_13[57], stage0_13[58], stage0_13[59], stage0_13[60], stage0_13[61]},
      {stage0_14[60]},
      {stage0_15[54], stage0_15[55], stage0_15[56], stage0_15[57], stage0_15[58], stage0_15[59]},
      {stage1_17[9],stage1_16[18],stage1_15[19],stage1_14[21],stage1_13[30]}
   );
   gpc1_1 gpc79 (
      {stage0_0[53]},
      {stage1_0[9]}
   );
   gpc1_1 gpc80 (
      {stage0_0[54]},
      {stage1_0[10]}
   );
   gpc1_1 gpc81 (
      {stage0_0[55]},
      {stage1_0[11]}
   );
   gpc1_1 gpc82 (
      {stage0_0[56]},
      {stage1_0[12]}
   );
   gpc1_1 gpc83 (
      {stage0_0[57]},
      {stage1_0[13]}
   );
   gpc1_1 gpc84 (
      {stage0_0[58]},
      {stage1_0[14]}
   );
   gpc1_1 gpc85 (
      {stage0_0[59]},
      {stage1_0[15]}
   );
   gpc1_1 gpc86 (
      {stage0_0[60]},
      {stage1_0[16]}
   );
   gpc1_1 gpc87 (
      {stage0_0[61]},
      {stage1_0[17]}
   );
   gpc1_1 gpc88 (
      {stage0_0[62]},
      {stage1_0[18]}
   );
   gpc1_1 gpc89 (
      {stage0_0[63]},
      {stage1_0[19]}
   );
   gpc1_1 gpc90 (
      {stage0_1[51]},
      {stage1_1[17]}
   );
   gpc1_1 gpc91 (
      {stage0_1[52]},
      {stage1_1[18]}
   );
   gpc1_1 gpc92 (
      {stage0_1[53]},
      {stage1_1[19]}
   );
   gpc1_1 gpc93 (
      {stage0_1[54]},
      {stage1_1[20]}
   );
   gpc1_1 gpc94 (
      {stage0_1[55]},
      {stage1_1[21]}
   );
   gpc1_1 gpc95 (
      {stage0_1[56]},
      {stage1_1[22]}
   );
   gpc1_1 gpc96 (
      {stage0_1[57]},
      {stage1_1[23]}
   );
   gpc1_1 gpc97 (
      {stage0_1[58]},
      {stage1_1[24]}
   );
   gpc1_1 gpc98 (
      {stage0_1[59]},
      {stage1_1[25]}
   );
   gpc1_1 gpc99 (
      {stage0_1[60]},
      {stage1_1[26]}
   );
   gpc1_1 gpc100 (
      {stage0_1[61]},
      {stage1_1[27]}
   );
   gpc1_1 gpc101 (
      {stage0_1[62]},
      {stage1_1[28]}
   );
   gpc1_1 gpc102 (
      {stage0_1[63]},
      {stage1_1[29]}
   );
   gpc1_1 gpc103 (
      {stage0_2[59]},
      {stage1_2[19]}
   );
   gpc1_1 gpc104 (
      {stage0_2[60]},
      {stage1_2[20]}
   );
   gpc1_1 gpc105 (
      {stage0_2[61]},
      {stage1_2[21]}
   );
   gpc1_1 gpc106 (
      {stage0_2[62]},
      {stage1_2[22]}
   );
   gpc1_1 gpc107 (
      {stage0_2[63]},
      {stage1_2[23]}
   );
   gpc1_1 gpc108 (
      {stage0_3[57]},
      {stage1_3[20]}
   );
   gpc1_1 gpc109 (
      {stage0_3[58]},
      {stage1_3[21]}
   );
   gpc1_1 gpc110 (
      {stage0_3[59]},
      {stage1_3[22]}
   );
   gpc1_1 gpc111 (
      {stage0_3[60]},
      {stage1_3[23]}
   );
   gpc1_1 gpc112 (
      {stage0_3[61]},
      {stage1_3[24]}
   );
   gpc1_1 gpc113 (
      {stage0_3[62]},
      {stage1_3[25]}
   );
   gpc1_1 gpc114 (
      {stage0_3[63]},
      {stage1_3[26]}
   );
   gpc1_1 gpc115 (
      {stage0_4[51]},
      {stage1_4[27]}
   );
   gpc1_1 gpc116 (
      {stage0_4[52]},
      {stage1_4[28]}
   );
   gpc1_1 gpc117 (
      {stage0_4[53]},
      {stage1_4[29]}
   );
   gpc1_1 gpc118 (
      {stage0_4[54]},
      {stage1_4[30]}
   );
   gpc1_1 gpc119 (
      {stage0_4[55]},
      {stage1_4[31]}
   );
   gpc1_1 gpc120 (
      {stage0_4[56]},
      {stage1_4[32]}
   );
   gpc1_1 gpc121 (
      {stage0_4[57]},
      {stage1_4[33]}
   );
   gpc1_1 gpc122 (
      {stage0_4[58]},
      {stage1_4[34]}
   );
   gpc1_1 gpc123 (
      {stage0_4[59]},
      {stage1_4[35]}
   );
   gpc1_1 gpc124 (
      {stage0_4[60]},
      {stage1_4[36]}
   );
   gpc1_1 gpc125 (
      {stage0_4[61]},
      {stage1_4[37]}
   );
   gpc1_1 gpc126 (
      {stage0_4[62]},
      {stage1_4[38]}
   );
   gpc1_1 gpc127 (
      {stage0_4[63]},
      {stage1_4[39]}
   );
   gpc1_1 gpc128 (
      {stage0_5[62]},
      {stage1_5[27]}
   );
   gpc1_1 gpc129 (
      {stage0_5[63]},
      {stage1_5[28]}
   );
   gpc1_1 gpc130 (
      {stage0_6[59]},
      {stage1_6[22]}
   );
   gpc1_1 gpc131 (
      {stage0_6[60]},
      {stage1_6[23]}
   );
   gpc1_1 gpc132 (
      {stage0_6[61]},
      {stage1_6[24]}
   );
   gpc1_1 gpc133 (
      {stage0_6[62]},
      {stage1_6[25]}
   );
   gpc1_1 gpc134 (
      {stage0_6[63]},
      {stage1_6[26]}
   );
   gpc1_1 gpc135 (
      {stage0_7[62]},
      {stage1_7[21]}
   );
   gpc1_1 gpc136 (
      {stage0_7[63]},
      {stage1_7[22]}
   );
   gpc1_1 gpc137 (
      {stage0_8[63]},
      {stage1_8[28]}
   );
   gpc1_1 gpc138 (
      {stage0_10[58]},
      {stage1_10[23]}
   );
   gpc1_1 gpc139 (
      {stage0_10[59]},
      {stage1_10[24]}
   );
   gpc1_1 gpc140 (
      {stage0_10[60]},
      {stage1_10[25]}
   );
   gpc1_1 gpc141 (
      {stage0_10[61]},
      {stage1_10[26]}
   );
   gpc1_1 gpc142 (
      {stage0_10[62]},
      {stage1_10[27]}
   );
   gpc1_1 gpc143 (
      {stage0_10[63]},
      {stage1_10[28]}
   );
   gpc1_1 gpc144 (
      {stage0_11[61]},
      {stage1_11[21]}
   );
   gpc1_1 gpc145 (
      {stage0_11[62]},
      {stage1_11[22]}
   );
   gpc1_1 gpc146 (
      {stage0_11[63]},
      {stage1_11[23]}
   );
   gpc1_1 gpc147 (
      {stage0_13[62]},
      {stage1_13[31]}
   );
   gpc1_1 gpc148 (
      {stage0_13[63]},
      {stage1_13[32]}
   );
   gpc1_1 gpc149 (
      {stage0_14[61]},
      {stage1_14[22]}
   );
   gpc1_1 gpc150 (
      {stage0_14[62]},
      {stage1_14[23]}
   );
   gpc1_1 gpc151 (
      {stage0_14[63]},
      {stage1_14[24]}
   );
   gpc1_1 gpc152 (
      {stage0_15[60]},
      {stage1_15[20]}
   );
   gpc1_1 gpc153 (
      {stage0_15[61]},
      {stage1_15[21]}
   );
   gpc1_1 gpc154 (
      {stage0_15[62]},
      {stage1_15[22]}
   );
   gpc1_1 gpc155 (
      {stage0_15[63]},
      {stage1_15[23]}
   );
   gpc2135_5 gpc156 (
      {stage1_0[0], stage1_0[1], stage1_0[2], stage1_0[3], stage1_0[4]},
      {stage1_1[0], stage1_1[1], stage1_1[2]},
      {stage1_2[0]},
      {stage1_3[0], stage1_3[1]},
      {stage2_4[0],stage2_3[0],stage2_2[0],stage2_1[0],stage2_0[0]}
   );
   gpc2135_5 gpc157 (
      {stage1_0[5], stage1_0[6], stage1_0[7], stage1_0[8], stage1_0[9]},
      {stage1_1[3], stage1_1[4], stage1_1[5]},
      {stage1_2[1]},
      {stage1_3[2], stage1_3[3]},
      {stage2_4[1],stage2_3[1],stage2_2[1],stage2_1[1],stage2_0[1]}
   );
   gpc2135_5 gpc158 (
      {stage1_0[10], stage1_0[11], stage1_0[12], stage1_0[13], stage1_0[14]},
      {stage1_1[6], stage1_1[7], stage1_1[8]},
      {stage1_2[2]},
      {stage1_3[4], stage1_3[5]},
      {stage2_4[2],stage2_3[2],stage2_2[2],stage2_1[2],stage2_0[2]}
   );
   gpc2135_5 gpc159 (
      {stage1_0[15], stage1_0[16], stage1_0[17], stage1_0[18], stage1_0[19]},
      {stage1_1[9], stage1_1[10], stage1_1[11]},
      {stage1_2[3]},
      {stage1_3[6], stage1_3[7]},
      {stage2_4[3],stage2_3[3],stage2_2[3],stage2_1[3],stage2_0[3]}
   );
   gpc615_5 gpc160 (
      {stage1_2[4], stage1_2[5], stage1_2[6], stage1_2[7], stage1_2[8]},
      {stage1_3[8]},
      {stage1_4[0], stage1_4[1], stage1_4[2], stage1_4[3], stage1_4[4], stage1_4[5]},
      {stage2_6[0],stage2_5[0],stage2_4[4],stage2_3[4],stage2_2[4]}
   );
   gpc615_5 gpc161 (
      {stage1_2[9], stage1_2[10], stage1_2[11], stage1_2[12], stage1_2[13]},
      {stage1_3[9]},
      {stage1_4[6], stage1_4[7], stage1_4[8], stage1_4[9], stage1_4[10], stage1_4[11]},
      {stage2_6[1],stage2_5[1],stage2_4[5],stage2_3[5],stage2_2[5]}
   );
   gpc615_5 gpc162 (
      {stage1_2[14], stage1_2[15], stage1_2[16], stage1_2[17], stage1_2[18]},
      {stage1_3[10]},
      {stage1_4[12], stage1_4[13], stage1_4[14], stage1_4[15], stage1_4[16], stage1_4[17]},
      {stage2_6[2],stage2_5[2],stage2_4[6],stage2_3[6],stage2_2[6]}
   );
   gpc615_5 gpc163 (
      {stage1_2[19], stage1_2[20], stage1_2[21], stage1_2[22], stage1_2[23]},
      {stage1_3[11]},
      {stage1_4[18], stage1_4[19], stage1_4[20], stage1_4[21], stage1_4[22], stage1_4[23]},
      {stage2_6[3],stage2_5[3],stage2_4[7],stage2_3[7],stage2_2[7]}
   );
   gpc615_5 gpc164 (
      {stage1_3[12], stage1_3[13], stage1_3[14], stage1_3[15], stage1_3[16]},
      {stage1_4[24]},
      {stage1_5[0], stage1_5[1], stage1_5[2], stage1_5[3], stage1_5[4], stage1_5[5]},
      {stage2_7[0],stage2_6[4],stage2_5[4],stage2_4[8],stage2_3[8]}
   );
   gpc615_5 gpc165 (
      {stage1_3[17], stage1_3[18], stage1_3[19], stage1_3[20], stage1_3[21]},
      {stage1_4[25]},
      {stage1_5[6], stage1_5[7], stage1_5[8], stage1_5[9], stage1_5[10], stage1_5[11]},
      {stage2_7[1],stage2_6[5],stage2_5[5],stage2_4[9],stage2_3[9]}
   );
   gpc615_5 gpc166 (
      {stage1_3[22], stage1_3[23], stage1_3[24], stage1_3[25], stage1_3[26]},
      {stage1_4[26]},
      {stage1_5[12], stage1_5[13], stage1_5[14], stage1_5[15], stage1_5[16], stage1_5[17]},
      {stage2_7[2],stage2_6[6],stage2_5[6],stage2_4[10],stage2_3[10]}
   );
   gpc615_5 gpc167 (
      {stage1_4[27], stage1_4[28], stage1_4[29], stage1_4[30], stage1_4[31]},
      {stage1_5[18]},
      {stage1_6[0], stage1_6[1], stage1_6[2], stage1_6[3], stage1_6[4], stage1_6[5]},
      {stage2_8[0],stage2_7[3],stage2_6[7],stage2_5[7],stage2_4[11]}
   );
   gpc615_5 gpc168 (
      {stage1_4[32], stage1_4[33], stage1_4[34], stage1_4[35], stage1_4[36]},
      {stage1_5[19]},
      {stage1_6[6], stage1_6[7], stage1_6[8], stage1_6[9], stage1_6[10], stage1_6[11]},
      {stage2_8[1],stage2_7[4],stage2_6[8],stage2_5[8],stage2_4[12]}
   );
   gpc615_5 gpc169 (
      {stage1_6[12], stage1_6[13], stage1_6[14], stage1_6[15], stage1_6[16]},
      {stage1_7[0]},
      {stage1_8[0], stage1_8[1], stage1_8[2], stage1_8[3], stage1_8[4], stage1_8[5]},
      {stage2_10[0],stage2_9[0],stage2_8[2],stage2_7[5],stage2_6[9]}
   );
   gpc615_5 gpc170 (
      {stage1_6[17], stage1_6[18], stage1_6[19], stage1_6[20], stage1_6[21]},
      {stage1_7[1]},
      {stage1_8[6], stage1_8[7], stage1_8[8], stage1_8[9], stage1_8[10], stage1_8[11]},
      {stage2_10[1],stage2_9[1],stage2_8[3],stage2_7[6],stage2_6[10]}
   );
   gpc615_5 gpc171 (
      {stage1_6[22], stage1_6[23], stage1_6[24], stage1_6[25], stage1_6[26]},
      {stage1_7[2]},
      {stage1_8[12], stage1_8[13], stage1_8[14], stage1_8[15], stage1_8[16], stage1_8[17]},
      {stage2_10[2],stage2_9[2],stage2_8[4],stage2_7[7],stage2_6[11]}
   );
   gpc615_5 gpc172 (
      {stage1_7[3], stage1_7[4], stage1_7[5], stage1_7[6], stage1_7[7]},
      {stage1_8[18]},
      {stage1_9[0], stage1_9[1], stage1_9[2], stage1_9[3], stage1_9[4], stage1_9[5]},
      {stage2_11[0],stage2_10[3],stage2_9[3],stage2_8[5],stage2_7[8]}
   );
   gpc615_5 gpc173 (
      {stage1_7[8], stage1_7[9], stage1_7[10], stage1_7[11], stage1_7[12]},
      {stage1_8[19]},
      {stage1_9[6], stage1_9[7], stage1_9[8], stage1_9[9], stage1_9[10], stage1_9[11]},
      {stage2_11[1],stage2_10[4],stage2_9[4],stage2_8[6],stage2_7[9]}
   );
   gpc615_5 gpc174 (
      {stage1_7[13], stage1_7[14], stage1_7[15], stage1_7[16], stage1_7[17]},
      {stage1_8[20]},
      {stage1_9[12], stage1_9[13], stage1_9[14], stage1_9[15], stage1_9[16], stage1_9[17]},
      {stage2_11[2],stage2_10[5],stage2_9[5],stage2_8[7],stage2_7[10]}
   );
   gpc615_5 gpc175 (
      {stage1_7[18], stage1_7[19], stage1_7[20], stage1_7[21], stage1_7[22]},
      {stage1_8[21]},
      {stage1_9[18], stage1_9[19], stage1_9[20], stage1_9[21], stage1_9[22], stage1_9[23]},
      {stage2_11[3],stage2_10[6],stage2_9[6],stage2_8[8],stage2_7[11]}
   );
   gpc606_5 gpc176 (
      {stage1_9[24], stage1_9[25], stage1_9[26], stage1_9[27], stage1_9[28], stage1_9[29]},
      {stage1_11[0], stage1_11[1], stage1_11[2], stage1_11[3], stage1_11[4], stage1_11[5]},
      {stage2_13[0],stage2_12[0],stage2_11[4],stage2_10[7],stage2_9[7]}
   );
   gpc606_5 gpc177 (
      {stage1_10[0], stage1_10[1], stage1_10[2], stage1_10[3], stage1_10[4], stage1_10[5]},
      {stage1_12[0], stage1_12[1], stage1_12[2], stage1_12[3], stage1_12[4], stage1_12[5]},
      {stage2_14[0],stage2_13[1],stage2_12[1],stage2_11[5],stage2_10[8]}
   );
   gpc606_5 gpc178 (
      {stage1_10[6], stage1_10[7], stage1_10[8], stage1_10[9], stage1_10[10], stage1_10[11]},
      {stage1_12[6], stage1_12[7], stage1_12[8], stage1_12[9], stage1_12[10], stage1_12[11]},
      {stage2_14[1],stage2_13[2],stage2_12[2],stage2_11[6],stage2_10[9]}
   );
   gpc606_5 gpc179 (
      {stage1_10[12], stage1_10[13], stage1_10[14], stage1_10[15], stage1_10[16], stage1_10[17]},
      {stage1_12[12], stage1_12[13], stage1_12[14], stage1_12[15], stage1_12[16], stage1_12[17]},
      {stage2_14[2],stage2_13[3],stage2_12[3],stage2_11[7],stage2_10[10]}
   );
   gpc606_5 gpc180 (
      {stage1_10[18], stage1_10[19], stage1_10[20], stage1_10[21], stage1_10[22], stage1_10[23]},
      {stage1_12[18], stage1_12[19], stage1_12[20], stage1_12[21], stage1_12[22], stage1_12[23]},
      {stage2_14[3],stage2_13[4],stage2_12[4],stage2_11[8],stage2_10[11]}
   );
   gpc606_5 gpc181 (
      {stage1_10[24], stage1_10[25], stage1_10[26], stage1_10[27], stage1_10[28], 1'b0},
      {stage1_12[24], stage1_12[25], stage1_12[26], stage1_12[27], stage1_12[28], 1'b0},
      {stage2_14[4],stage2_13[5],stage2_12[5],stage2_11[9],stage2_10[12]}
   );
   gpc606_5 gpc182 (
      {stage1_11[6], stage1_11[7], stage1_11[8], stage1_11[9], stage1_11[10], stage1_11[11]},
      {stage1_13[0], stage1_13[1], stage1_13[2], stage1_13[3], stage1_13[4], stage1_13[5]},
      {stage2_15[0],stage2_14[5],stage2_13[6],stage2_12[6],stage2_11[10]}
   );
   gpc606_5 gpc183 (
      {stage1_11[12], stage1_11[13], stage1_11[14], stage1_11[15], stage1_11[16], stage1_11[17]},
      {stage1_13[6], stage1_13[7], stage1_13[8], stage1_13[9], stage1_13[10], stage1_13[11]},
      {stage2_15[1],stage2_14[6],stage2_13[7],stage2_12[7],stage2_11[11]}
   );
   gpc606_5 gpc184 (
      {stage1_13[12], stage1_13[13], stage1_13[14], stage1_13[15], stage1_13[16], stage1_13[17]},
      {stage1_15[0], stage1_15[1], stage1_15[2], stage1_15[3], stage1_15[4], stage1_15[5]},
      {stage2_17[0],stage2_16[0],stage2_15[2],stage2_14[7],stage2_13[8]}
   );
   gpc606_5 gpc185 (
      {stage1_13[18], stage1_13[19], stage1_13[20], stage1_13[21], stage1_13[22], stage1_13[23]},
      {stage1_15[6], stage1_15[7], stage1_15[8], stage1_15[9], stage1_15[10], stage1_15[11]},
      {stage2_17[1],stage2_16[1],stage2_15[3],stage2_14[8],stage2_13[9]}
   );
   gpc606_5 gpc186 (
      {stage1_14[0], stage1_14[1], stage1_14[2], stage1_14[3], stage1_14[4], stage1_14[5]},
      {stage1_16[0], stage1_16[1], stage1_16[2], stage1_16[3], stage1_16[4], stage1_16[5]},
      {stage2_18[0],stage2_17[2],stage2_16[2],stage2_15[4],stage2_14[9]}
   );
   gpc606_5 gpc187 (
      {stage1_14[6], stage1_14[7], stage1_14[8], stage1_14[9], stage1_14[10], stage1_14[11]},
      {stage1_16[6], stage1_16[7], stage1_16[8], stage1_16[9], stage1_16[10], stage1_16[11]},
      {stage2_18[1],stage2_17[3],stage2_16[3],stage2_15[5],stage2_14[10]}
   );
   gpc606_5 gpc188 (
      {stage1_15[12], stage1_15[13], stage1_15[14], stage1_15[15], stage1_15[16], stage1_15[17]},
      {stage1_17[0], stage1_17[1], stage1_17[2], stage1_17[3], stage1_17[4], stage1_17[5]},
      {stage2_19[0],stage2_18[2],stage2_17[4],stage2_16[4],stage2_15[6]}
   );
   gpc606_5 gpc189 (
      {stage1_15[18], stage1_15[19], stage1_15[20], stage1_15[21], stage1_15[22], stage1_15[23]},
      {stage1_17[6], stage1_17[7], stage1_17[8], stage1_17[9], 1'b0, 1'b0},
      {stage2_19[1],stage2_18[3],stage2_17[5],stage2_16[5],stage2_15[7]}
   );
   gpc1_1 gpc190 (
      {stage1_1[12]},
      {stage2_1[4]}
   );
   gpc1_1 gpc191 (
      {stage1_1[13]},
      {stage2_1[5]}
   );
   gpc1_1 gpc192 (
      {stage1_1[14]},
      {stage2_1[6]}
   );
   gpc1_1 gpc193 (
      {stage1_1[15]},
      {stage2_1[7]}
   );
   gpc1_1 gpc194 (
      {stage1_1[16]},
      {stage2_1[8]}
   );
   gpc1_1 gpc195 (
      {stage1_1[17]},
      {stage2_1[9]}
   );
   gpc1_1 gpc196 (
      {stage1_1[18]},
      {stage2_1[10]}
   );
   gpc1_1 gpc197 (
      {stage1_1[19]},
      {stage2_1[11]}
   );
   gpc1_1 gpc198 (
      {stage1_1[20]},
      {stage2_1[12]}
   );
   gpc1_1 gpc199 (
      {stage1_1[21]},
      {stage2_1[13]}
   );
   gpc1_1 gpc200 (
      {stage1_1[22]},
      {stage2_1[14]}
   );
   gpc1_1 gpc201 (
      {stage1_1[23]},
      {stage2_1[15]}
   );
   gpc1_1 gpc202 (
      {stage1_1[24]},
      {stage2_1[16]}
   );
   gpc1_1 gpc203 (
      {stage1_1[25]},
      {stage2_1[17]}
   );
   gpc1_1 gpc204 (
      {stage1_1[26]},
      {stage2_1[18]}
   );
   gpc1_1 gpc205 (
      {stage1_1[27]},
      {stage2_1[19]}
   );
   gpc1_1 gpc206 (
      {stage1_1[28]},
      {stage2_1[20]}
   );
   gpc1_1 gpc207 (
      {stage1_1[29]},
      {stage2_1[21]}
   );
   gpc1_1 gpc208 (
      {stage1_4[37]},
      {stage2_4[13]}
   );
   gpc1_1 gpc209 (
      {stage1_4[38]},
      {stage2_4[14]}
   );
   gpc1_1 gpc210 (
      {stage1_4[39]},
      {stage2_4[15]}
   );
   gpc1_1 gpc211 (
      {stage1_5[20]},
      {stage2_5[9]}
   );
   gpc1_1 gpc212 (
      {stage1_5[21]},
      {stage2_5[10]}
   );
   gpc1_1 gpc213 (
      {stage1_5[22]},
      {stage2_5[11]}
   );
   gpc1_1 gpc214 (
      {stage1_5[23]},
      {stage2_5[12]}
   );
   gpc1_1 gpc215 (
      {stage1_5[24]},
      {stage2_5[13]}
   );
   gpc1_1 gpc216 (
      {stage1_5[25]},
      {stage2_5[14]}
   );
   gpc1_1 gpc217 (
      {stage1_5[26]},
      {stage2_5[15]}
   );
   gpc1_1 gpc218 (
      {stage1_5[27]},
      {stage2_5[16]}
   );
   gpc1_1 gpc219 (
      {stage1_5[28]},
      {stage2_5[17]}
   );
   gpc1_1 gpc220 (
      {stage1_8[22]},
      {stage2_8[9]}
   );
   gpc1_1 gpc221 (
      {stage1_8[23]},
      {stage2_8[10]}
   );
   gpc1_1 gpc222 (
      {stage1_8[24]},
      {stage2_8[11]}
   );
   gpc1_1 gpc223 (
      {stage1_8[25]},
      {stage2_8[12]}
   );
   gpc1_1 gpc224 (
      {stage1_8[26]},
      {stage2_8[13]}
   );
   gpc1_1 gpc225 (
      {stage1_8[27]},
      {stage2_8[14]}
   );
   gpc1_1 gpc226 (
      {stage1_8[28]},
      {stage2_8[15]}
   );
   gpc1_1 gpc227 (
      {stage1_11[18]},
      {stage2_11[12]}
   );
   gpc1_1 gpc228 (
      {stage1_11[19]},
      {stage2_11[13]}
   );
   gpc1_1 gpc229 (
      {stage1_11[20]},
      {stage2_11[14]}
   );
   gpc1_1 gpc230 (
      {stage1_11[21]},
      {stage2_11[15]}
   );
   gpc1_1 gpc231 (
      {stage1_11[22]},
      {stage2_11[16]}
   );
   gpc1_1 gpc232 (
      {stage1_11[23]},
      {stage2_11[17]}
   );
   gpc1_1 gpc233 (
      {stage1_13[24]},
      {stage2_13[10]}
   );
   gpc1_1 gpc234 (
      {stage1_13[25]},
      {stage2_13[11]}
   );
   gpc1_1 gpc235 (
      {stage1_13[26]},
      {stage2_13[12]}
   );
   gpc1_1 gpc236 (
      {stage1_13[27]},
      {stage2_13[13]}
   );
   gpc1_1 gpc237 (
      {stage1_13[28]},
      {stage2_13[14]}
   );
   gpc1_1 gpc238 (
      {stage1_13[29]},
      {stage2_13[15]}
   );
   gpc1_1 gpc239 (
      {stage1_13[30]},
      {stage2_13[16]}
   );
   gpc1_1 gpc240 (
      {stage1_13[31]},
      {stage2_13[17]}
   );
   gpc1_1 gpc241 (
      {stage1_13[32]},
      {stage2_13[18]}
   );
   gpc1_1 gpc242 (
      {stage1_14[12]},
      {stage2_14[11]}
   );
   gpc1_1 gpc243 (
      {stage1_14[13]},
      {stage2_14[12]}
   );
   gpc1_1 gpc244 (
      {stage1_14[14]},
      {stage2_14[13]}
   );
   gpc1_1 gpc245 (
      {stage1_14[15]},
      {stage2_14[14]}
   );
   gpc1_1 gpc246 (
      {stage1_14[16]},
      {stage2_14[15]}
   );
   gpc1_1 gpc247 (
      {stage1_14[17]},
      {stage2_14[16]}
   );
   gpc1_1 gpc248 (
      {stage1_14[18]},
      {stage2_14[17]}
   );
   gpc1_1 gpc249 (
      {stage1_14[19]},
      {stage2_14[18]}
   );
   gpc1_1 gpc250 (
      {stage1_14[20]},
      {stage2_14[19]}
   );
   gpc1_1 gpc251 (
      {stage1_14[21]},
      {stage2_14[20]}
   );
   gpc1_1 gpc252 (
      {stage1_14[22]},
      {stage2_14[21]}
   );
   gpc1_1 gpc253 (
      {stage1_14[23]},
      {stage2_14[22]}
   );
   gpc1_1 gpc254 (
      {stage1_14[24]},
      {stage2_14[23]}
   );
   gpc1_1 gpc255 (
      {stage1_16[12]},
      {stage2_16[6]}
   );
   gpc1_1 gpc256 (
      {stage1_16[13]},
      {stage2_16[7]}
   );
   gpc1_1 gpc257 (
      {stage1_16[14]},
      {stage2_16[8]}
   );
   gpc1_1 gpc258 (
      {stage1_16[15]},
      {stage2_16[9]}
   );
   gpc1_1 gpc259 (
      {stage1_16[16]},
      {stage2_16[10]}
   );
   gpc1_1 gpc260 (
      {stage1_16[17]},
      {stage2_16[11]}
   );
   gpc1_1 gpc261 (
      {stage1_16[18]},
      {stage2_16[12]}
   );
   gpc1163_5 gpc262 (
      {stage2_0[0], stage2_0[1], stage2_0[2]},
      {stage2_1[0], stage2_1[1], stage2_1[2], stage2_1[3], stage2_1[4], stage2_1[5]},
      {stage2_2[0]},
      {stage2_3[0]},
      {stage3_4[0],stage3_3[0],stage3_2[0],stage3_1[0],stage3_0[0]}
   );
   gpc1163_5 gpc263 (
      {stage2_0[3], 1'b0, 1'b0},
      {stage2_1[6], stage2_1[7], stage2_1[8], stage2_1[9], stage2_1[10], stage2_1[11]},
      {stage2_2[1]},
      {stage2_3[1]},
      {stage3_4[1],stage3_3[1],stage3_2[1],stage3_1[1],stage3_0[1]}
   );
   gpc606_5 gpc264 (
      {stage2_1[12], stage2_1[13], stage2_1[14], stage2_1[15], stage2_1[16], stage2_1[17]},
      {stage2_3[2], stage2_3[3], stage2_3[4], stage2_3[5], stage2_3[6], stage2_3[7]},
      {stage3_5[0],stage3_4[2],stage3_3[2],stage3_2[2],stage3_1[2]}
   );
   gpc615_5 gpc265 (
      {stage2_2[2], stage2_2[3], stage2_2[4], stage2_2[5], stage2_2[6]},
      {stage2_3[8]},
      {stage2_4[0], stage2_4[1], stage2_4[2], stage2_4[3], stage2_4[4], stage2_4[5]},
      {stage3_6[0],stage3_5[1],stage3_4[3],stage3_3[3],stage3_2[3]}
   );
   gpc615_5 gpc266 (
      {stage2_4[6], stage2_4[7], stage2_4[8], stage2_4[9], stage2_4[10]},
      {stage2_5[0]},
      {stage2_6[0], stage2_6[1], stage2_6[2], stage2_6[3], stage2_6[4], stage2_6[5]},
      {stage3_8[0],stage3_7[0],stage3_6[1],stage3_5[2],stage3_4[4]}
   );
   gpc615_5 gpc267 (
      {stage2_4[11], stage2_4[12], stage2_4[13], stage2_4[14], stage2_4[15]},
      {stage2_5[1]},
      {stage2_6[6], stage2_6[7], stage2_6[8], stage2_6[9], stage2_6[10], stage2_6[11]},
      {stage3_8[1],stage3_7[1],stage3_6[2],stage3_5[3],stage3_4[5]}
   );
   gpc606_5 gpc268 (
      {stage2_5[2], stage2_5[3], stage2_5[4], stage2_5[5], stage2_5[6], stage2_5[7]},
      {stage2_7[0], stage2_7[1], stage2_7[2], stage2_7[3], stage2_7[4], stage2_7[5]},
      {stage3_9[0],stage3_8[2],stage3_7[2],stage3_6[3],stage3_5[4]}
   );
   gpc606_5 gpc269 (
      {stage2_5[8], stage2_5[9], stage2_5[10], stage2_5[11], stage2_5[12], stage2_5[13]},
      {stage2_7[6], stage2_7[7], stage2_7[8], stage2_7[9], stage2_7[10], stage2_7[11]},
      {stage3_9[1],stage3_8[3],stage3_7[3],stage3_6[4],stage3_5[5]}
   );
   gpc1163_5 gpc270 (
      {stage2_8[0], stage2_8[1], stage2_8[2]},
      {stage2_9[0], stage2_9[1], stage2_9[2], stage2_9[3], stage2_9[4], stage2_9[5]},
      {stage2_10[0]},
      {stage2_11[0]},
      {stage3_12[0],stage3_11[0],stage3_10[0],stage3_9[2],stage3_8[4]}
   );
   gpc606_5 gpc271 (
      {stage2_8[3], stage2_8[4], stage2_8[5], stage2_8[6], stage2_8[7], stage2_8[8]},
      {stage2_10[1], stage2_10[2], stage2_10[3], stage2_10[4], stage2_10[5], stage2_10[6]},
      {stage3_12[1],stage3_11[1],stage3_10[1],stage3_9[3],stage3_8[5]}
   );
   gpc606_5 gpc272 (
      {stage2_8[9], stage2_8[10], stage2_8[11], stage2_8[12], stage2_8[13], stage2_8[14]},
      {stage2_10[7], stage2_10[8], stage2_10[9], stage2_10[10], stage2_10[11], stage2_10[12]},
      {stage3_12[2],stage3_11[2],stage3_10[2],stage3_9[4],stage3_8[6]}
   );
   gpc606_5 gpc273 (
      {stage2_11[1], stage2_11[2], stage2_11[3], stage2_11[4], stage2_11[5], stage2_11[6]},
      {stage2_13[0], stage2_13[1], stage2_13[2], stage2_13[3], stage2_13[4], stage2_13[5]},
      {stage3_15[0],stage3_14[0],stage3_13[0],stage3_12[3],stage3_11[3]}
   );
   gpc615_5 gpc274 (
      {stage2_11[7], stage2_11[8], stage2_11[9], stage2_11[10], stage2_11[11]},
      {stage2_12[0]},
      {stage2_13[6], stage2_13[7], stage2_13[8], stage2_13[9], stage2_13[10], stage2_13[11]},
      {stage3_15[1],stage3_14[1],stage3_13[1],stage3_12[4],stage3_11[4]}
   );
   gpc615_5 gpc275 (
      {stage2_11[12], stage2_11[13], stage2_11[14], stage2_11[15], stage2_11[16]},
      {stage2_12[1]},
      {stage2_13[12], stage2_13[13], stage2_13[14], stage2_13[15], stage2_13[16], stage2_13[17]},
      {stage3_15[2],stage3_14[2],stage3_13[2],stage3_12[5],stage3_11[5]}
   );
   gpc606_5 gpc276 (
      {stage2_12[2], stage2_12[3], stage2_12[4], stage2_12[5], stage2_12[6], stage2_12[7]},
      {stage2_14[0], stage2_14[1], stage2_14[2], stage2_14[3], stage2_14[4], stage2_14[5]},
      {stage3_16[0],stage3_15[3],stage3_14[3],stage3_13[3],stage3_12[6]}
   );
   gpc606_5 gpc277 (
      {stage2_14[6], stage2_14[7], stage2_14[8], stage2_14[9], stage2_14[10], stage2_14[11]},
      {stage2_16[0], stage2_16[1], stage2_16[2], stage2_16[3], stage2_16[4], stage2_16[5]},
      {stage3_18[0],stage3_17[0],stage3_16[1],stage3_15[4],stage3_14[4]}
   );
   gpc615_5 gpc278 (
      {stage2_14[12], stage2_14[13], stage2_14[14], stage2_14[15], stage2_14[16]},
      {stage2_15[0]},
      {stage2_16[6], stage2_16[7], stage2_16[8], stage2_16[9], stage2_16[10], stage2_16[11]},
      {stage3_18[1],stage3_17[1],stage3_16[2],stage3_15[5],stage3_14[5]}
   );
   gpc606_5 gpc279 (
      {stage2_15[1], stage2_15[2], stage2_15[3], stage2_15[4], stage2_15[5], stage2_15[6]},
      {stage2_17[0], stage2_17[1], stage2_17[2], stage2_17[3], stage2_17[4], stage2_17[5]},
      {stage3_19[0],stage3_18[2],stage3_17[2],stage3_16[3],stage3_15[6]}
   );
   gpc1_1 gpc280 (
      {stage2_1[18]},
      {stage3_1[3]}
   );
   gpc1_1 gpc281 (
      {stage2_1[19]},
      {stage3_1[4]}
   );
   gpc1_1 gpc282 (
      {stage2_1[20]},
      {stage3_1[5]}
   );
   gpc1_1 gpc283 (
      {stage2_1[21]},
      {stage3_1[6]}
   );
   gpc1_1 gpc284 (
      {stage2_2[7]},
      {stage3_2[4]}
   );
   gpc1_1 gpc285 (
      {stage2_3[9]},
      {stage3_3[4]}
   );
   gpc1_1 gpc286 (
      {stage2_3[10]},
      {stage3_3[5]}
   );
   gpc1_1 gpc287 (
      {stage2_5[14]},
      {stage3_5[6]}
   );
   gpc1_1 gpc288 (
      {stage2_5[15]},
      {stage3_5[7]}
   );
   gpc1_1 gpc289 (
      {stage2_5[16]},
      {stage3_5[8]}
   );
   gpc1_1 gpc290 (
      {stage2_5[17]},
      {stage3_5[9]}
   );
   gpc1_1 gpc291 (
      {stage2_8[15]},
      {stage3_8[7]}
   );
   gpc1_1 gpc292 (
      {stage2_9[6]},
      {stage3_9[5]}
   );
   gpc1_1 gpc293 (
      {stage2_9[7]},
      {stage3_9[6]}
   );
   gpc1_1 gpc294 (
      {stage2_11[17]},
      {stage3_11[6]}
   );
   gpc1_1 gpc295 (
      {stage2_13[18]},
      {stage3_13[4]}
   );
   gpc1_1 gpc296 (
      {stage2_14[17]},
      {stage3_14[6]}
   );
   gpc1_1 gpc297 (
      {stage2_14[18]},
      {stage3_14[7]}
   );
   gpc1_1 gpc298 (
      {stage2_14[19]},
      {stage3_14[8]}
   );
   gpc1_1 gpc299 (
      {stage2_14[20]},
      {stage3_14[9]}
   );
   gpc1_1 gpc300 (
      {stage2_14[21]},
      {stage3_14[10]}
   );
   gpc1_1 gpc301 (
      {stage2_14[22]},
      {stage3_14[11]}
   );
   gpc1_1 gpc302 (
      {stage2_14[23]},
      {stage3_14[12]}
   );
   gpc1_1 gpc303 (
      {stage2_15[7]},
      {stage3_15[7]}
   );
   gpc1_1 gpc304 (
      {stage2_16[12]},
      {stage3_16[4]}
   );
   gpc1_1 gpc305 (
      {stage2_18[0]},
      {stage3_18[3]}
   );
   gpc1_1 gpc306 (
      {stage2_18[1]},
      {stage3_18[4]}
   );
   gpc1_1 gpc307 (
      {stage2_18[2]},
      {stage3_18[5]}
   );
   gpc1_1 gpc308 (
      {stage2_18[3]},
      {stage3_18[6]}
   );
   gpc1_1 gpc309 (
      {stage2_19[0]},
      {stage3_19[1]}
   );
   gpc1_1 gpc310 (
      {stage2_19[1]},
      {stage3_19[2]}
   );
   gpc606_5 gpc311 (
      {stage3_1[0], stage3_1[1], stage3_1[2], stage3_1[3], stage3_1[4], stage3_1[5]},
      {stage3_3[0], stage3_3[1], stage3_3[2], stage3_3[3], stage3_3[4], stage3_3[5]},
      {stage4_5[0],stage4_4[0],stage4_3[0],stage4_2[0],stage4_1[0]}
   );
   gpc615_5 gpc312 (
      {stage3_2[0], stage3_2[1], stage3_2[2], stage3_2[3], stage3_2[4]},
      {1'b0},
      {stage3_4[0], stage3_4[1], stage3_4[2], stage3_4[3], stage3_4[4], stage3_4[5]},
      {stage4_6[0],stage4_5[1],stage4_4[1],stage4_3[1],stage4_2[1]}
   );
   gpc117_4 gpc313 (
      {stage3_5[0], stage3_5[1], stage3_5[2], stage3_5[3], stage3_5[4], stage3_5[5], stage3_5[6]},
      {stage3_6[0]},
      {stage3_7[0]},
      {stage4_8[0],stage4_7[0],stage4_6[1],stage4_5[2]}
   );
   gpc615_5 gpc314 (
      {stage3_6[1], stage3_6[2], stage3_6[3], stage3_6[4], 1'b0},
      {stage3_7[1]},
      {stage3_8[0], stage3_8[1], stage3_8[2], stage3_8[3], stage3_8[4], stage3_8[5]},
      {stage4_10[0],stage4_9[0],stage4_8[1],stage4_7[1],stage4_6[2]}
   );
   gpc615_5 gpc315 (
      {stage3_9[0], stage3_9[1], stage3_9[2], stage3_9[3], stage3_9[4]},
      {stage3_10[0]},
      {stage3_11[0], stage3_11[1], stage3_11[2], stage3_11[3], stage3_11[4], stage3_11[5]},
      {stage4_13[0],stage4_12[0],stage4_11[0],stage4_10[1],stage4_9[1]}
   );
   gpc606_5 gpc316 (
      {stage3_12[0], stage3_12[1], stage3_12[2], stage3_12[3], stage3_12[4], stage3_12[5]},
      {stage3_14[0], stage3_14[1], stage3_14[2], stage3_14[3], stage3_14[4], stage3_14[5]},
      {stage4_16[0],stage4_15[0],stage4_14[0],stage4_13[1],stage4_12[1]}
   );
   gpc615_5 gpc317 (
      {stage3_13[0], stage3_13[1], stage3_13[2], stage3_13[3], stage3_13[4]},
      {stage3_14[6]},
      {stage3_15[0], stage3_15[1], stage3_15[2], stage3_15[3], stage3_15[4], stage3_15[5]},
      {stage4_17[0],stage4_16[1],stage4_15[1],stage4_14[1],stage4_13[2]}
   );
   gpc615_5 gpc318 (
      {stage3_16[0], stage3_16[1], stage3_16[2], stage3_16[3], stage3_16[4]},
      {stage3_17[0]},
      {stage3_18[0], stage3_18[1], stage3_18[2], stage3_18[3], stage3_18[4], stage3_18[5]},
      {stage4_20[0],stage4_19[0],stage4_18[0],stage4_17[1],stage4_16[2]}
   );
   gpc1_1 gpc319 (
      {stage3_0[0]},
      {stage4_0[0]}
   );
   gpc1_1 gpc320 (
      {stage3_0[1]},
      {stage4_0[1]}
   );
   gpc1_1 gpc321 (
      {stage3_1[6]},
      {stage4_1[1]}
   );
   gpc1_1 gpc322 (
      {stage3_5[7]},
      {stage4_5[3]}
   );
   gpc1_1 gpc323 (
      {stage3_5[8]},
      {stage4_5[4]}
   );
   gpc1_1 gpc324 (
      {stage3_5[9]},
      {stage4_5[5]}
   );
   gpc1_1 gpc325 (
      {stage3_7[2]},
      {stage4_7[2]}
   );
   gpc1_1 gpc326 (
      {stage3_7[3]},
      {stage4_7[3]}
   );
   gpc1_1 gpc327 (
      {stage3_8[6]},
      {stage4_8[2]}
   );
   gpc1_1 gpc328 (
      {stage3_8[7]},
      {stage4_8[3]}
   );
   gpc1_1 gpc329 (
      {stage3_9[5]},
      {stage4_9[2]}
   );
   gpc1_1 gpc330 (
      {stage3_9[6]},
      {stage4_9[3]}
   );
   gpc1_1 gpc331 (
      {stage3_10[1]},
      {stage4_10[2]}
   );
   gpc1_1 gpc332 (
      {stage3_10[2]},
      {stage4_10[3]}
   );
   gpc1_1 gpc333 (
      {stage3_11[6]},
      {stage4_11[1]}
   );
   gpc1_1 gpc334 (
      {stage3_12[6]},
      {stage4_12[2]}
   );
   gpc1_1 gpc335 (
      {stage3_14[7]},
      {stage4_14[2]}
   );
   gpc1_1 gpc336 (
      {stage3_14[8]},
      {stage4_14[3]}
   );
   gpc1_1 gpc337 (
      {stage3_14[9]},
      {stage4_14[4]}
   );
   gpc1_1 gpc338 (
      {stage3_14[10]},
      {stage4_14[5]}
   );
   gpc1_1 gpc339 (
      {stage3_14[11]},
      {stage4_14[6]}
   );
   gpc1_1 gpc340 (
      {stage3_14[12]},
      {stage4_14[7]}
   );
   gpc1_1 gpc341 (
      {stage3_15[6]},
      {stage4_15[2]}
   );
   gpc1_1 gpc342 (
      {stage3_15[7]},
      {stage4_15[3]}
   );
   gpc1_1 gpc343 (
      {stage3_17[1]},
      {stage4_17[2]}
   );
   gpc1_1 gpc344 (
      {stage3_17[2]},
      {stage4_17[3]}
   );
   gpc1_1 gpc345 (
      {stage3_18[6]},
      {stage4_18[1]}
   );
   gpc1_1 gpc346 (
      {stage3_19[0]},
      {stage4_19[1]}
   );
   gpc1_1 gpc347 (
      {stage3_19[1]},
      {stage4_19[2]}
   );
   gpc1_1 gpc348 (
      {stage3_19[2]},
      {stage4_19[3]}
   );
   gpc1325_5 gpc349 (
      {stage4_5[0], stage4_5[1], stage4_5[2], stage4_5[3], stage4_5[4]},
      {stage4_6[0], stage4_6[1]},
      {stage4_7[0], stage4_7[1], stage4_7[2]},
      {stage4_8[0]},
      {stage5_9[0],stage5_8[0],stage5_7[0],stage5_6[0],stage5_5[0]}
   );
   gpc1343_5 gpc350 (
      {stage4_8[1], stage4_8[2], stage4_8[3]},
      {stage4_9[0], stage4_9[1], stage4_9[2], stage4_9[3]},
      {stage4_10[0], stage4_10[1], stage4_10[2]},
      {stage4_11[0]},
      {stage5_12[0],stage5_11[0],stage5_10[0],stage5_9[1],stage5_8[1]}
   );
   gpc623_5 gpc351 (
      {stage4_12[0], stage4_12[1], stage4_12[2]},
      {stage4_13[0], stage4_13[1]},
      {stage4_14[0], stage4_14[1], stage4_14[2], stage4_14[3], stage4_14[4], stage4_14[5]},
      {stage5_16[0],stage5_15[0],stage5_14[0],stage5_13[0],stage5_12[1]}
   );
   gpc1343_5 gpc352 (
      {stage4_14[6], stage4_14[7], 1'b0},
      {stage4_15[0], stage4_15[1], stage4_15[2], stage4_15[3]},
      {stage4_16[0], stage4_16[1], stage4_16[2]},
      {stage4_17[0]},
      {stage5_18[0],stage5_17[0],stage5_16[1],stage5_15[1],stage5_14[1]}
   );
   gpc623_5 gpc353 (
      {stage4_17[1], stage4_17[2], stage4_17[3]},
      {stage4_18[0], stage4_18[1]},
      {stage4_19[0], stage4_19[1], stage4_19[2], stage4_19[3], 1'b0, 1'b0},
      {stage5_21[0],stage5_20[0],stage5_19[0],stage5_18[1],stage5_17[1]}
   );
   gpc1_1 gpc354 (
      {stage4_0[0]},
      {stage5_0[0]}
   );
   gpc1_1 gpc355 (
      {stage4_0[1]},
      {stage5_0[1]}
   );
   gpc1_1 gpc356 (
      {stage4_1[0]},
      {stage5_1[0]}
   );
   gpc1_1 gpc357 (
      {stage4_1[1]},
      {stage5_1[1]}
   );
   gpc1_1 gpc358 (
      {stage4_2[0]},
      {stage5_2[0]}
   );
   gpc1_1 gpc359 (
      {stage4_2[1]},
      {stage5_2[1]}
   );
   gpc1_1 gpc360 (
      {stage4_3[0]},
      {stage5_3[0]}
   );
   gpc1_1 gpc361 (
      {stage4_3[1]},
      {stage5_3[1]}
   );
   gpc1_1 gpc362 (
      {stage4_4[0]},
      {stage5_4[0]}
   );
   gpc1_1 gpc363 (
      {stage4_4[1]},
      {stage5_4[1]}
   );
   gpc1_1 gpc364 (
      {stage4_5[5]},
      {stage5_5[1]}
   );
   gpc1_1 gpc365 (
      {stage4_6[2]},
      {stage5_6[1]}
   );
   gpc1_1 gpc366 (
      {stage4_7[3]},
      {stage5_7[1]}
   );
   gpc1_1 gpc367 (
      {stage4_10[3]},
      {stage5_10[1]}
   );
   gpc1_1 gpc368 (
      {stage4_11[1]},
      {stage5_11[1]}
   );
   gpc1_1 gpc369 (
      {stage4_13[2]},
      {stage5_13[1]}
   );
   gpc1_1 gpc370 (
      {stage4_20[0]},
      {stage5_20[1]}
   );
endmodule
module rowadder2_1_22(input [21:0] src0, input [21:0] src1, output [22:0] dst0);
    wire [21:0] gene;
    wire [21:0] prop;
    wire [23:0] out;
    wire [23:0] carryout;
    LUT2 #(
        .INIT(4'h8)
    ) lut_0_gene (
        .I0(src0[0]),
        .I1(src1[0]),
        .O(gene[0])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_0_prop (
        .I0(src0[0]),
        .I1(src1[0]),
        .O(prop[0])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_1_gene (
        .I0(src0[1]),
        .I1(src1[1]),
        .O(gene[1])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_1_prop (
        .I0(src0[1]),
        .I1(src1[1]),
        .O(prop[1])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_2_gene (
        .I0(src0[2]),
        .I1(src1[2]),
        .O(gene[2])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_2_prop (
        .I0(src0[2]),
        .I1(src1[2]),
        .O(prop[2])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_3_gene (
        .I0(src0[3]),
        .I1(src1[3]),
        .O(gene[3])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_3_prop (
        .I0(src0[3]),
        .I1(src1[3]),
        .O(prop[3])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_4_gene (
        .I0(src0[4]),
        .I1(src1[4]),
        .O(gene[4])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_4_prop (
        .I0(src0[4]),
        .I1(src1[4]),
        .O(prop[4])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_5_gene (
        .I0(src0[5]),
        .I1(src1[5]),
        .O(gene[5])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_5_prop (
        .I0(src0[5]),
        .I1(src1[5]),
        .O(prop[5])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_6_gene (
        .I0(src0[6]),
        .I1(src1[6]),
        .O(gene[6])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_6_prop (
        .I0(src0[6]),
        .I1(src1[6]),
        .O(prop[6])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_7_gene (
        .I0(src0[7]),
        .I1(src1[7]),
        .O(gene[7])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_7_prop (
        .I0(src0[7]),
        .I1(src1[7]),
        .O(prop[7])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_8_gene (
        .I0(src0[8]),
        .I1(src1[8]),
        .O(gene[8])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_8_prop (
        .I0(src0[8]),
        .I1(src1[8]),
        .O(prop[8])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_9_gene (
        .I0(src0[9]),
        .I1(src1[9]),
        .O(gene[9])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_9_prop (
        .I0(src0[9]),
        .I1(src1[9]),
        .O(prop[9])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_10_gene (
        .I0(src0[10]),
        .I1(src1[10]),
        .O(gene[10])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_10_prop (
        .I0(src0[10]),
        .I1(src1[10]),
        .O(prop[10])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_11_gene (
        .I0(src0[11]),
        .I1(src1[11]),
        .O(gene[11])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_11_prop (
        .I0(src0[11]),
        .I1(src1[11]),
        .O(prop[11])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_12_gene (
        .I0(src0[12]),
        .I1(src1[12]),
        .O(gene[12])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_12_prop (
        .I0(src0[12]),
        .I1(src1[12]),
        .O(prop[12])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_13_gene (
        .I0(src0[13]),
        .I1(src1[13]),
        .O(gene[13])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_13_prop (
        .I0(src0[13]),
        .I1(src1[13]),
        .O(prop[13])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_14_gene (
        .I0(src0[14]),
        .I1(src1[14]),
        .O(gene[14])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_14_prop (
        .I0(src0[14]),
        .I1(src1[14]),
        .O(prop[14])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_15_gene (
        .I0(src0[15]),
        .I1(src1[15]),
        .O(gene[15])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_15_prop (
        .I0(src0[15]),
        .I1(src1[15]),
        .O(prop[15])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_16_gene (
        .I0(src0[16]),
        .I1(src1[16]),
        .O(gene[16])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_16_prop (
        .I0(src0[16]),
        .I1(src1[16]),
        .O(prop[16])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_17_gene (
        .I0(src0[17]),
        .I1(src1[17]),
        .O(gene[17])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_17_prop (
        .I0(src0[17]),
        .I1(src1[17]),
        .O(prop[17])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_18_gene (
        .I0(src0[18]),
        .I1(src1[18]),
        .O(gene[18])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_18_prop (
        .I0(src0[18]),
        .I1(src1[18]),
        .O(prop[18])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_19_gene (
        .I0(src0[19]),
        .I1(src1[19]),
        .O(gene[19])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_19_prop (
        .I0(src0[19]),
        .I1(src1[19]),
        .O(prop[19])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_20_gene (
        .I0(src0[20]),
        .I1(src1[20]),
        .O(gene[20])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_20_prop (
        .I0(src0[20]),
        .I1(src1[20]),
        .O(prop[20])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_21_gene (
        .I0(src0[21]),
        .I1(src1[21]),
        .O(gene[21])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_21_prop (
        .I0(src0[21]),
        .I1(src1[21]),
        .O(prop[21])
    );
    CARRY4 carry4_3_0 (
        .CO(carryout[3:0]),
        .O(out[3:0]),
        .CI(1'h0),
        .CYINIT(1'h0),
        .DI(gene[3:0]),
        .S(prop[3:0])
    );
    CARRY4 carry4_7_4 (
        .CO(carryout[7:4]),
        .O(out[7:4]),
        .CI(carryout[3]),
        .CYINIT(1'h0),
        .DI(gene[7:4]),
        .S(prop[7:4])
    );
    CARRY4 carry4_11_8 (
        .CO(carryout[11:8]),
        .O(out[11:8]),
        .CI(carryout[7]),
        .CYINIT(1'h0),
        .DI(gene[11:8]),
        .S(prop[11:8])
    );
    CARRY4 carry4_15_12 (
        .CO(carryout[15:12]),
        .O(out[15:12]),
        .CI(carryout[11]),
        .CYINIT(1'h0),
        .DI(gene[15:12]),
        .S(prop[15:12])
    );
    CARRY4 carry4_19_16 (
        .CO(carryout[19:16]),
        .O(out[19:16]),
        .CI(carryout[15]),
        .CYINIT(1'h0),
        .DI(gene[19:16]),
        .S(prop[19:16])
    );
    CARRY4 carry4_23_20 (
        .CO(carryout[23:20]),
        .O(out[23:20]),
        .CI(carryout[19]),
        .CYINIT(1'h0),
        .DI({2'h0, gene[21:20]}),
        .S({2'h0, prop[21:20]})
    );
    assign dst0 = {carryout[21], out[21:0]};
endmodule


module comp2_1test_64_16();
    reg [15:0] src0;
    reg [15:0] src1;
    reg [15:0] src2;
    reg [15:0] src3;
    reg [15:0] src4;
    reg [15:0] src5;
    reg [15:0] src6;
    reg [15:0] src7;
    reg [15:0] src8;
    reg [15:0] src9;
    reg [15:0] src10;
    reg [15:0] src11;
    reg [15:0] src12;
    reg [15:0] src13;
    reg [15:0] src14;
    reg [15:0] src15;
    reg [15:0] src16;
    reg [15:0] src17;
    reg [15:0] src18;
    reg [15:0] src19;
    reg [15:0] src20;
    reg [15:0] src21;
    reg [15:0] src22;
    reg [15:0] src23;
    reg [15:0] src24;
    reg [15:0] src25;
    reg [15:0] src26;
    reg [15:0] src27;
    reg [15:0] src28;
    reg [15:0] src29;
    reg [15:0] src30;
    reg [15:0] src31;
    reg [15:0] src32;
    reg [15:0] src33;
    reg [15:0] src34;
    reg [15:0] src35;
    reg [15:0] src36;
    reg [15:0] src37;
    reg [15:0] src38;
    reg [15:0] src39;
    reg [15:0] src40;
    reg [15:0] src41;
    reg [15:0] src42;
    reg [15:0] src43;
    reg [15:0] src44;
    reg [15:0] src45;
    reg [15:0] src46;
    reg [15:0] src47;
    reg [15:0] src48;
    reg [15:0] src49;
    reg [15:0] src50;
    reg [15:0] src51;
    reg [15:0] src52;
    reg [15:0] src53;
    reg [15:0] src54;
    reg [15:0] src55;
    reg [15:0] src56;
    reg [15:0] src57;
    reg [15:0] src58;
    reg [15:0] src59;
    reg [15:0] src60;
    reg [15:0] src61;
    reg [15:0] src62;
    reg [15:0] src63;
    reg [21:0] exp;
    wire [21:0] dst;
    assign test = dst == exp;
    compressor2_1_64_16 compressor2_1_64_16_inst(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .src31(src31),
        .src32(src32),
        .src33(src33),
        .src34(src34),
        .src35(src35),
        .src36(src36),
        .src37(src37),
        .src38(src38),
        .src39(src39),
        .src40(src40),
        .src41(src41),
        .src42(src42),
        .src43(src43),
        .src44(src44),
        .src45(src45),
        .src46(src46),
        .src47(src47),
        .src48(src48),
        .src49(src49),
        .src50(src50),
        .src51(src51),
        .src52(src52),
        .src53(src53),
        .src54(src54),
        .src55(src55),
        .src56(src56),
        .src57(src57),
        .src58(src58),
        .src59(src59),
        .src60(src60),
        .src61(src61),
        .src62(src62),
        .src63(src63),
        .dst(dst)
    );
    initial begin
        $monitor("0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x %x", src0, src1, src2, src3, src4, src5, src6, src7, src8, src9, src10, src11, src12, src13, src14, src15, src16, src17, src18, src19, src20, src21, src22, src23, src24, src25, src26, src27, src28, src29, src30, src31, src32, src33, src34, src35, src36, src37, src38, src39, src40, src41, src42, src43, src44, src45, src46, src47, src48, src49, src50, src51, src52, src53, src54, src55, src56, src57, src58, src59, src60, src61, src62, src63, dst, exp, test);
        src0 <= 16'h2c9e;
        src1 <= 16'hca7;
        src2 <= 16'hef9c;
        src3 <= 16'ha6f7;
        src4 <= 16'h7371;
        src5 <= 16'hb0be;
        src6 <= 16'hb2d4;
        src7 <= 16'hec85;
        src8 <= 16'hdc68;
        src9 <= 16'hed01;
        src10 <= 16'h5009;
        src11 <= 16'hf842;
        src12 <= 16'h544;
        src13 <= 16'ha45e;
        src14 <= 16'hf312;
        src15 <= 16'haee8;
        src16 <= 16'h3cf2;
        src17 <= 16'hf097;
        src18 <= 16'hb01c;
        src19 <= 16'hd94e;
        src20 <= 16'hea50;
        src21 <= 16'h5440;
        src22 <= 16'h610f;
        src23 <= 16'h9d36;
        src24 <= 16'h683f;
        src25 <= 16'h4721;
        src26 <= 16'he921;
        src27 <= 16'h41b3;
        src28 <= 16'hf11d;
        src29 <= 16'h23b7;
        src30 <= 16'hfc58;
        src31 <= 16'hf8db;
        src32 <= 16'h94bc;
        src33 <= 16'hdea7;
        src34 <= 16'h5cca;
        src35 <= 16'h4bc9;
        src36 <= 16'ha686;
        src37 <= 16'h415f;
        src38 <= 16'h8bff;
        src39 <= 16'h8de4;
        src40 <= 16'hee84;
        src41 <= 16'h561e;
        src42 <= 16'h935d;
        src43 <= 16'h235b;
        src44 <= 16'hf582;
        src45 <= 16'h4677;
        src46 <= 16'h25d1;
        src47 <= 16'h7c5b;
        src48 <= 16'hebaf;
        src49 <= 16'h5b9;
        src50 <= 16'h74c3;
        src51 <= 16'h8113;
        src52 <= 16'h337;
        src53 <= 16'ha42a;
        src54 <= 16'h703b;
        src55 <= 16'hc1ce;
        src56 <= 16'h50ae;
        src57 <= 16'h3b22;
        src58 <= 16'h7adc;
        src59 <= 16'haaef;
        src60 <= 16'h8385;
        src61 <= 16'h2999;
        src62 <= 16'h7e8d;
        src63 <= 16'h156e;
        exp <= 22'h22734c;
        #1
        src0 <= 16'hfb3b;
        src1 <= 16'h9cad;
        src2 <= 16'h1f89;
        src3 <= 16'h878;
        src4 <= 16'h455c;
        src5 <= 16'h2062;
        src6 <= 16'h4faa;
        src7 <= 16'hdb43;
        src8 <= 16'h380c;
        src9 <= 16'h41df;
        src10 <= 16'h112;
        src11 <= 16'hc17a;
        src12 <= 16'he2f;
        src13 <= 16'hbcc6;
        src14 <= 16'he00a;
        src15 <= 16'hfb6c;
        src16 <= 16'h3ad5;
        src17 <= 16'hec89;
        src18 <= 16'hfd59;
        src19 <= 16'h4486;
        src20 <= 16'hddc7;
        src21 <= 16'hd027;
        src22 <= 16'haf28;
        src23 <= 16'hacbb;
        src24 <= 16'h7b09;
        src25 <= 16'h1ef5;
        src26 <= 16'he6bb;
        src27 <= 16'h6936;
        src28 <= 16'ha8c1;
        src29 <= 16'h98c3;
        src30 <= 16'h5b92;
        src31 <= 16'h49dc;
        src32 <= 16'he1be;
        src33 <= 16'h341f;
        src34 <= 16'h80b3;
        src35 <= 16'h6623;
        src36 <= 16'hd4b3;
        src37 <= 16'h9831;
        src38 <= 16'h2239;
        src39 <= 16'h77ca;
        src40 <= 16'h4eb;
        src41 <= 16'ha157;
        src42 <= 16'hc0a9;
        src43 <= 16'h6671;
        src44 <= 16'h2fda;
        src45 <= 16'hcb86;
        src46 <= 16'ha56a;
        src47 <= 16'h1d53;
        src48 <= 16'hcccf;
        src49 <= 16'h726b;
        src50 <= 16'h54eb;
        src51 <= 16'h24ce;
        src52 <= 16'ha1c8;
        src53 <= 16'hded1;
        src54 <= 16'h5cb3;
        src55 <= 16'h222f;
        src56 <= 16'h4a30;
        src57 <= 16'h3625;
        src58 <= 16'hf67a;
        src59 <= 16'h85de;
        src60 <= 16'heab8;
        src61 <= 16'h1e9d;
        src62 <= 16'h168b;
        src63 <= 16'hbf94;
        exp <= 22'h1f9b07;
        #1
        src0 <= 16'hc8a9;
        src1 <= 16'hd6fd;
        src2 <= 16'h9fe;
        src3 <= 16'h2a27;
        src4 <= 16'h4aae;
        src5 <= 16'hc015;
        src6 <= 16'h399e;
        src7 <= 16'h7030;
        src8 <= 16'h44f2;
        src9 <= 16'h7f66;
        src10 <= 16'h6b73;
        src11 <= 16'h1699;
        src12 <= 16'h9a67;
        src13 <= 16'h3f9b;
        src14 <= 16'ha321;
        src15 <= 16'h678a;
        src16 <= 16'h9d10;
        src17 <= 16'h9fa6;
        src18 <= 16'h98ff;
        src19 <= 16'h56ef;
        src20 <= 16'hbb64;
        src21 <= 16'h6d9c;
        src22 <= 16'h1c8e;
        src23 <= 16'h1ae8;
        src24 <= 16'hbd91;
        src25 <= 16'h3128;
        src26 <= 16'hf386;
        src27 <= 16'hd80c;
        src28 <= 16'h3eda;
        src29 <= 16'he58c;
        src30 <= 16'h74ab;
        src31 <= 16'h8800;
        src32 <= 16'hd72;
        src33 <= 16'he89b;
        src34 <= 16'h37d2;
        src35 <= 16'h68d8;
        src36 <= 16'h8de9;
        src37 <= 16'h51b1;
        src38 <= 16'ha761;
        src39 <= 16'h842d;
        src40 <= 16'ha292;
        src41 <= 16'hd49e;
        src42 <= 16'h344e;
        src43 <= 16'h82c2;
        src44 <= 16'hcbad;
        src45 <= 16'hd430;
        src46 <= 16'h7a1e;
        src47 <= 16'h7f9b;
        src48 <= 16'h47a2;
        src49 <= 16'h4391;
        src50 <= 16'h3f95;
        src51 <= 16'h66ea;
        src52 <= 16'ha72c;
        src53 <= 16'hb7e9;
        src54 <= 16'h4df2;
        src55 <= 16'h809d;
        src56 <= 16'h3767;
        src57 <= 16'h8274;
        src58 <= 16'h1e31;
        src59 <= 16'h4947;
        src60 <= 16'hf6f1;
        src61 <= 16'h8e7b;
        src62 <= 16'hcda2;
        src63 <= 16'h9062;
        exp <= 22'h1ee9b1;
        #1
        src0 <= 16'h36c8;
        src1 <= 16'h17fe;
        src2 <= 16'h7608;
        src3 <= 16'h1c28;
        src4 <= 16'h839f;
        src5 <= 16'hf860;
        src6 <= 16'h3f52;
        src7 <= 16'hba4f;
        src8 <= 16'h2348;
        src9 <= 16'h3bd0;
        src10 <= 16'hd72d;
        src11 <= 16'hb8b0;
        src12 <= 16'hd5d1;
        src13 <= 16'h6d80;
        src14 <= 16'hbb51;
        src15 <= 16'h44af;
        src16 <= 16'h9e5a;
        src17 <= 16'h60aa;
        src18 <= 16'ha5f2;
        src19 <= 16'h6c74;
        src20 <= 16'h7ceb;
        src21 <= 16'h865e;
        src22 <= 16'hd4f4;
        src23 <= 16'h42b;
        src24 <= 16'h22f3;
        src25 <= 16'haf77;
        src26 <= 16'h8d71;
        src27 <= 16'hc142;
        src28 <= 16'hb9b1;
        src29 <= 16'h22d7;
        src30 <= 16'h1a24;
        src31 <= 16'h200c;
        src32 <= 16'h988e;
        src33 <= 16'h18af;
        src34 <= 16'hc64f;
        src35 <= 16'h35c5;
        src36 <= 16'h5be4;
        src37 <= 16'h86ed;
        src38 <= 16'hbf78;
        src39 <= 16'h7f57;
        src40 <= 16'hf08f;
        src41 <= 16'hf395;
        src42 <= 16'hdd34;
        src43 <= 16'hdc1a;
        src44 <= 16'h5e34;
        src45 <= 16'h458c;
        src46 <= 16'h1d2e;
        src47 <= 16'h9182;
        src48 <= 16'h62af;
        src49 <= 16'h1eb1;
        src50 <= 16'hfcad;
        src51 <= 16'hfc21;
        src52 <= 16'h2609;
        src53 <= 16'h9501;
        src54 <= 16'h3fd0;
        src55 <= 16'hc41e;
        src56 <= 16'h85df;
        src57 <= 16'h8db1;
        src58 <= 16'h86f7;
        src59 <= 16'h19a5;
        src60 <= 16'h26e2;
        src61 <= 16'h89ae;
        src62 <= 16'h3023;
        src63 <= 16'he6ea;
        exp <= 22'h1f2245;
        #1
        src0 <= 16'hfa77;
        src1 <= 16'hca47;
        src2 <= 16'h13d1;
        src3 <= 16'hcf18;
        src4 <= 16'he125;
        src5 <= 16'h3b9f;
        src6 <= 16'h8d32;
        src7 <= 16'h78e3;
        src8 <= 16'h75a0;
        src9 <= 16'hfa39;
        src10 <= 16'h802f;
        src11 <= 16'hccbd;
        src12 <= 16'h5211;
        src13 <= 16'hefc5;
        src14 <= 16'h8af0;
        src15 <= 16'h3c7b;
        src16 <= 16'h242f;
        src17 <= 16'h129d;
        src18 <= 16'ha271;
        src19 <= 16'hc36e;
        src20 <= 16'ha018;
        src21 <= 16'h3389;
        src22 <= 16'hb585;
        src23 <= 16'ha555;
        src24 <= 16'had31;
        src25 <= 16'h4995;
        src26 <= 16'h2d59;
        src27 <= 16'hf2a6;
        src28 <= 16'h4986;
        src29 <= 16'h56dc;
        src30 <= 16'h78c1;
        src31 <= 16'hfba0;
        src32 <= 16'h7735;
        src33 <= 16'h6239;
        src34 <= 16'h2ea6;
        src35 <= 16'ha19a;
        src36 <= 16'h2304;
        src37 <= 16'h721;
        src38 <= 16'ha070;
        src39 <= 16'h60e;
        src40 <= 16'hb8c;
        src41 <= 16'h8dfa;
        src42 <= 16'hb40e;
        src43 <= 16'hd2d7;
        src44 <= 16'h2e86;
        src45 <= 16'h75fe;
        src46 <= 16'hf2b5;
        src47 <= 16'h3aeb;
        src48 <= 16'h23a9;
        src49 <= 16'h58b8;
        src50 <= 16'hc468;
        src51 <= 16'hf773;
        src52 <= 16'h7d7c;
        src53 <= 16'h27f5;
        src54 <= 16'hba7f;
        src55 <= 16'h7208;
        src56 <= 16'h6d3a;
        src57 <= 16'h1bdb;
        src58 <= 16'h260f;
        src59 <= 16'hc8e0;
        src60 <= 16'hceb1;
        src61 <= 16'h4711;
        src62 <= 16'hb8ff;
        src63 <= 16'h16ce;
        exp <= 22'h1f5bdb;
        #1
        src0 <= 16'hce3d;
        src1 <= 16'hbe9e;
        src2 <= 16'he45e;
        src3 <= 16'h676b;
        src4 <= 16'he702;
        src5 <= 16'h415e;
        src6 <= 16'h3d23;
        src7 <= 16'hb58c;
        src8 <= 16'hd7c9;
        src9 <= 16'hdb80;
        src10 <= 16'h4686;
        src11 <= 16'h3bd4;
        src12 <= 16'h5eb8;
        src13 <= 16'h536f;
        src14 <= 16'h5408;
        src15 <= 16'h2cc0;
        src16 <= 16'h351c;
        src17 <= 16'h45e6;
        src18 <= 16'he47a;
        src19 <= 16'haa84;
        src20 <= 16'hb6e4;
        src21 <= 16'ha64b;
        src22 <= 16'h54a7;
        src23 <= 16'h2611;
        src24 <= 16'h216f;
        src25 <= 16'h7bb;
        src26 <= 16'hb3de;
        src27 <= 16'hc0ec;
        src28 <= 16'hd029;
        src29 <= 16'h388c;
        src30 <= 16'h7dd0;
        src31 <= 16'hfcd6;
        src32 <= 16'h842a;
        src33 <= 16'h2b67;
        src34 <= 16'h3800;
        src35 <= 16'h2178;
        src36 <= 16'hd72e;
        src37 <= 16'h5539;
        src38 <= 16'h8a01;
        src39 <= 16'hb208;
        src40 <= 16'h7f0d;
        src41 <= 16'h3052;
        src42 <= 16'h8e74;
        src43 <= 16'h46f2;
        src44 <= 16'hb716;
        src45 <= 16'h2e58;
        src46 <= 16'h2a13;
        src47 <= 16'hee9b;
        src48 <= 16'h28ee;
        src49 <= 16'hb56e;
        src50 <= 16'hcee8;
        src51 <= 16'hb51f;
        src52 <= 16'h5fd6;
        src53 <= 16'h15ff;
        src54 <= 16'hccbc;
        src55 <= 16'h44e4;
        src56 <= 16'hbd2f;
        src57 <= 16'he35;
        src58 <= 16'hfbdb;
        src59 <= 16'h3bfb;
        src60 <= 16'h954e;
        src61 <= 16'h9404;
        src62 <= 16'h8344;
        src63 <= 16'hafc5;
        exp <= 22'h1f9d42;
        #1
        src0 <= 16'hb5c;
        src1 <= 16'h29d9;
        src2 <= 16'h8160;
        src3 <= 16'h2d0a;
        src4 <= 16'hea6a;
        src5 <= 16'hd959;
        src6 <= 16'ha653;
        src7 <= 16'ha876;
        src8 <= 16'h62c6;
        src9 <= 16'h6796;
        src10 <= 16'h6ad1;
        src11 <= 16'h2d48;
        src12 <= 16'h3b23;
        src13 <= 16'h7c2;
        src14 <= 16'h5cf9;
        src15 <= 16'hbe49;
        src16 <= 16'h606;
        src17 <= 16'h6bb2;
        src18 <= 16'h1df5;
        src19 <= 16'h2cf6;
        src20 <= 16'h3db8;
        src21 <= 16'h8277;
        src22 <= 16'he049;
        src23 <= 16'he413;
        src24 <= 16'hbd9a;
        src25 <= 16'hbc47;
        src26 <= 16'hb66d;
        src27 <= 16'h9cd1;
        src28 <= 16'h4e4c;
        src29 <= 16'h6998;
        src30 <= 16'ha9f4;
        src31 <= 16'h184e;
        src32 <= 16'he489;
        src33 <= 16'hf95f;
        src34 <= 16'h65ca;
        src35 <= 16'h3423;
        src36 <= 16'h71fd;
        src37 <= 16'h1c1c;
        src38 <= 16'h1ddb;
        src39 <= 16'hbdef;
        src40 <= 16'h9c12;
        src41 <= 16'h68b2;
        src42 <= 16'heee;
        src43 <= 16'h58ea;
        src44 <= 16'hed4;
        src45 <= 16'h6ad0;
        src46 <= 16'h1c37;
        src47 <= 16'hc4a1;
        src48 <= 16'hf534;
        src49 <= 16'h91b2;
        src50 <= 16'hc32d;
        src51 <= 16'h3f82;
        src52 <= 16'hbe5c;
        src53 <= 16'hf223;
        src54 <= 16'ha676;
        src55 <= 16'h2ec;
        src56 <= 16'h314c;
        src57 <= 16'h4d4e;
        src58 <= 16'h4b4c;
        src59 <= 16'had9a;
        src60 <= 16'hef41;
        src61 <= 16'hc787;
        src62 <= 16'h6c4f;
        src63 <= 16'h7d9f;
        exp <= 22'h1de3b6;
        #1
        src0 <= 16'haeb9;
        src1 <= 16'h74dc;
        src2 <= 16'he14f;
        src3 <= 16'hf4f0;
        src4 <= 16'hc3d6;
        src5 <= 16'h9b00;
        src6 <= 16'h9479;
        src7 <= 16'hc231;
        src8 <= 16'h27e9;
        src9 <= 16'h3f2c;
        src10 <= 16'hc290;
        src11 <= 16'h7dea;
        src12 <= 16'h2cf2;
        src13 <= 16'ha4b8;
        src14 <= 16'h132d;
        src15 <= 16'h4f7a;
        src16 <= 16'h4620;
        src17 <= 16'h4348;
        src18 <= 16'h918a;
        src19 <= 16'h5620;
        src20 <= 16'h50c7;
        src21 <= 16'heb87;
        src22 <= 16'hd1ca;
        src23 <= 16'hf7f5;
        src24 <= 16'h435c;
        src25 <= 16'h6fcd;
        src26 <= 16'h2663;
        src27 <= 16'hd8a5;
        src28 <= 16'h6e69;
        src29 <= 16'h68ef;
        src30 <= 16'h3b21;
        src31 <= 16'h4eaf;
        src32 <= 16'h8321;
        src33 <= 16'hcb1e;
        src34 <= 16'hbc07;
        src35 <= 16'ha4ff;
        src36 <= 16'h80e6;
        src37 <= 16'h485d;
        src38 <= 16'h9e1d;
        src39 <= 16'ha9cd;
        src40 <= 16'h67c6;
        src41 <= 16'hedb0;
        src42 <= 16'h495e;
        src43 <= 16'hf525;
        src44 <= 16'hf541;
        src45 <= 16'h3dbc;
        src46 <= 16'he87a;
        src47 <= 16'h9536;
        src48 <= 16'he7a3;
        src49 <= 16'h8f1e;
        src50 <= 16'h7fe5;
        src51 <= 16'hd158;
        src52 <= 16'hee00;
        src53 <= 16'hc1ec;
        src54 <= 16'h9516;
        src55 <= 16'h6dac;
        src56 <= 16'hf024;
        src57 <= 16'hfb28;
        src58 <= 16'hb294;
        src59 <= 16'h1be;
        src60 <= 16'hdb7c;
        src61 <= 16'he5a8;
        src62 <= 16'hf080;
        src63 <= 16'h5a81;
        exp <= 22'h254133;
        #1
        src0 <= 16'hd913;
        src1 <= 16'h80d5;
        src2 <= 16'hb5a3;
        src3 <= 16'hfa9;
        src4 <= 16'h2522;
        src5 <= 16'h79f;
        src6 <= 16'h1890;
        src7 <= 16'h6040;
        src8 <= 16'hdb43;
        src9 <= 16'h57f;
        src10 <= 16'hc7da;
        src11 <= 16'hba65;
        src12 <= 16'hf38e;
        src13 <= 16'hdf86;
        src14 <= 16'h9c95;
        src15 <= 16'hd499;
        src16 <= 16'h2551;
        src17 <= 16'hbce9;
        src18 <= 16'h7f45;
        src19 <= 16'hb9f0;
        src20 <= 16'h27f6;
        src21 <= 16'h986b;
        src22 <= 16'h3995;
        src23 <= 16'h197c;
        src24 <= 16'h8670;
        src25 <= 16'h359e;
        src26 <= 16'h1a6b;
        src27 <= 16'h6b0e;
        src28 <= 16'h5acf;
        src29 <= 16'hf361;
        src30 <= 16'h5548;
        src31 <= 16'ha9ac;
        src32 <= 16'h19f9;
        src33 <= 16'h8d01;
        src34 <= 16'h453;
        src35 <= 16'h3f31;
        src36 <= 16'h958f;
        src37 <= 16'h81d6;
        src38 <= 16'h6171;
        src39 <= 16'h10c;
        src40 <= 16'h4835;
        src41 <= 16'he3df;
        src42 <= 16'h602b;
        src43 <= 16'h5f8b;
        src44 <= 16'h4b64;
        src45 <= 16'h4e85;
        src46 <= 16'h44a1;
        src47 <= 16'haf08;
        src48 <= 16'h1790;
        src49 <= 16'hb658;
        src50 <= 16'h2501;
        src51 <= 16'h1d6f;
        src52 <= 16'h3dd2;
        src53 <= 16'h9835;
        src54 <= 16'hbb7;
        src55 <= 16'h8461;
        src56 <= 16'h7371;
        src57 <= 16'hd80d;
        src58 <= 16'hf504;
        src59 <= 16'he4fe;
        src60 <= 16'h73dd;
        src61 <= 16'hc25e;
        src62 <= 16'he2a9;
        src63 <= 16'h8ad1;
        exp <= 22'h1d46fc;
        #1
        src0 <= 16'h6e21;
        src1 <= 16'he7d6;
        src2 <= 16'hde84;
        src3 <= 16'he9c9;
        src4 <= 16'hb55;
        src5 <= 16'hab6e;
        src6 <= 16'ha738;
        src7 <= 16'h261f;
        src8 <= 16'h5bd7;
        src9 <= 16'h2fae;
        src10 <= 16'hcd49;
        src11 <= 16'h699d;
        src12 <= 16'hdeb;
        src13 <= 16'h5db8;
        src14 <= 16'h9e3d;
        src15 <= 16'h21c2;
        src16 <= 16'ha543;
        src17 <= 16'h9b6d;
        src18 <= 16'h2003;
        src19 <= 16'hf0ba;
        src20 <= 16'he86f;
        src21 <= 16'h74ff;
        src22 <= 16'h2cef;
        src23 <= 16'h1460;
        src24 <= 16'h1c00;
        src25 <= 16'hb1db;
        src26 <= 16'h6a7b;
        src27 <= 16'h8dd7;
        src28 <= 16'h279c;
        src29 <= 16'h2207;
        src30 <= 16'hec1e;
        src31 <= 16'h9196;
        src32 <= 16'h9725;
        src33 <= 16'hd574;
        src34 <= 16'h9e9c;
        src35 <= 16'hed29;
        src36 <= 16'hf93c;
        src37 <= 16'h30f6;
        src38 <= 16'h39ed;
        src39 <= 16'hccfc;
        src40 <= 16'h6113;
        src41 <= 16'h8691;
        src42 <= 16'hdc58;
        src43 <= 16'h417a;
        src44 <= 16'h3f85;
        src45 <= 16'h1f22;
        src46 <= 16'h50d6;
        src47 <= 16'hf526;
        src48 <= 16'ha570;
        src49 <= 16'h8ba0;
        src50 <= 16'h1848;
        src51 <= 16'he604;
        src52 <= 16'h3efd;
        src53 <= 16'h485;
        src54 <= 16'h2f25;
        src55 <= 16'hd23c;
        src56 <= 16'hd850;
        src57 <= 16'ha7fd;
        src58 <= 16'h6647;
        src59 <= 16'hcf24;
        src60 <= 16'h8f75;
        src61 <= 16'hb81d;
        src62 <= 16'hac0a;
        src63 <= 16'ha1f5;
        exp <= 22'h20a133;
        #1
        src0 <= 16'h419;
        src1 <= 16'had1b;
        src2 <= 16'hf272;
        src3 <= 16'h428f;
        src4 <= 16'hf60d;
        src5 <= 16'h8464;
        src6 <= 16'h483c;
        src7 <= 16'h247c;
        src8 <= 16'hb074;
        src9 <= 16'h6b88;
        src10 <= 16'h18b5;
        src11 <= 16'he771;
        src12 <= 16'hd5b1;
        src13 <= 16'hbc27;
        src14 <= 16'h5625;
        src15 <= 16'h81cd;
        src16 <= 16'hf162;
        src17 <= 16'h6de6;
        src18 <= 16'h3fef;
        src19 <= 16'h5cd8;
        src20 <= 16'h66a5;
        src21 <= 16'hff06;
        src22 <= 16'h7a7e;
        src23 <= 16'h2fc2;
        src24 <= 16'hf5d7;
        src25 <= 16'h851f;
        src26 <= 16'hecf6;
        src27 <= 16'hb284;
        src28 <= 16'h388a;
        src29 <= 16'h12eb;
        src30 <= 16'he1cd;
        src31 <= 16'h6a3e;
        src32 <= 16'ha37f;
        src33 <= 16'h99f0;
        src34 <= 16'hb641;
        src35 <= 16'h30ad;
        src36 <= 16'hd876;
        src37 <= 16'hfe55;
        src38 <= 16'hdfe;
        src39 <= 16'h18a3;
        src40 <= 16'h821c;
        src41 <= 16'h8616;
        src42 <= 16'h4a52;
        src43 <= 16'h6c04;
        src44 <= 16'hda0b;
        src45 <= 16'h16ea;
        src46 <= 16'hf595;
        src47 <= 16'h1a85;
        src48 <= 16'h67ed;
        src49 <= 16'h809b;
        src50 <= 16'h250;
        src51 <= 16'h4c7c;
        src52 <= 16'ha35;
        src53 <= 16'hef83;
        src54 <= 16'h8bf9;
        src55 <= 16'h49ec;
        src56 <= 16'h816;
        src57 <= 16'hdddc;
        src58 <= 16'hedda;
        src59 <= 16'h21c8;
        src60 <= 16'h8382;
        src61 <= 16'h1bca;
        src62 <= 16'h15cc;
        src63 <= 16'ha339;
        exp <= 22'h1f476a;
        #1
        src0 <= 16'h8293;
        src1 <= 16'h2a99;
        src2 <= 16'h863a;
        src3 <= 16'hd2f0;
        src4 <= 16'h3b2f;
        src5 <= 16'h27c9;
        src6 <= 16'h9513;
        src7 <= 16'h686;
        src8 <= 16'h2e49;
        src9 <= 16'h1f41;
        src10 <= 16'hd72;
        src11 <= 16'h1a93;
        src12 <= 16'h867b;
        src13 <= 16'ha7b8;
        src14 <= 16'hd001;
        src15 <= 16'h15d0;
        src16 <= 16'h476b;
        src17 <= 16'hfbe5;
        src18 <= 16'h3aaa;
        src19 <= 16'hbdf8;
        src20 <= 16'h5c9f;
        src21 <= 16'h20cf;
        src22 <= 16'h9fce;
        src23 <= 16'hbd92;
        src24 <= 16'hf2dc;
        src25 <= 16'h66a1;
        src26 <= 16'ha2fe;
        src27 <= 16'h3135;
        src28 <= 16'h6a7b;
        src29 <= 16'h85e;
        src30 <= 16'h2186;
        src31 <= 16'he701;
        src32 <= 16'ha677;
        src33 <= 16'h649e;
        src34 <= 16'hf864;
        src35 <= 16'hbfe;
        src36 <= 16'h7dfa;
        src37 <= 16'h7eab;
        src38 <= 16'h8639;
        src39 <= 16'h957e;
        src40 <= 16'h86;
        src41 <= 16'h8d18;
        src42 <= 16'hc03b;
        src43 <= 16'hbaf9;
        src44 <= 16'hf476;
        src45 <= 16'h76f;
        src46 <= 16'h7236;
        src47 <= 16'h9f1c;
        src48 <= 16'haf78;
        src49 <= 16'hd854;
        src50 <= 16'h81ab;
        src51 <= 16'he9ac;
        src52 <= 16'h1168;
        src53 <= 16'h7621;
        src54 <= 16'hf6cc;
        src55 <= 16'h72d9;
        src56 <= 16'h7d48;
        src57 <= 16'hc430;
        src58 <= 16'hffc5;
        src59 <= 16'h61e8;
        src60 <= 16'h1682;
        src61 <= 16'h1311;
        src62 <= 16'h5be9;
        src63 <= 16'h6cf4;
        exp <= 22'h1e060c;
        #1
        src0 <= 16'h992b;
        src1 <= 16'hbb27;
        src2 <= 16'h7b00;
        src3 <= 16'h1d26;
        src4 <= 16'h1e96;
        src5 <= 16'ha222;
        src6 <= 16'h61cd;
        src7 <= 16'h9745;
        src8 <= 16'h2739;
        src9 <= 16'h7fa1;
        src10 <= 16'h21a0;
        src11 <= 16'h96d3;
        src12 <= 16'hae0b;
        src13 <= 16'h7d9;
        src14 <= 16'hc9ad;
        src15 <= 16'h3a20;
        src16 <= 16'hf810;
        src17 <= 16'he50;
        src18 <= 16'h1a62;
        src19 <= 16'h15ba;
        src20 <= 16'h1d4b;
        src21 <= 16'h1116;
        src22 <= 16'h800d;
        src23 <= 16'hc73f;
        src24 <= 16'hd078;
        src25 <= 16'h262e;
        src26 <= 16'h8aa2;
        src27 <= 16'hec74;
        src28 <= 16'h27d2;
        src29 <= 16'hedab;
        src30 <= 16'he3c;
        src31 <= 16'h7ed3;
        src32 <= 16'he47;
        src33 <= 16'ha98c;
        src34 <= 16'h1ad7;
        src35 <= 16'h6862;
        src36 <= 16'hea3;
        src37 <= 16'h6327;
        src38 <= 16'hf63f;
        src39 <= 16'h2bf8;
        src40 <= 16'hfef5;
        src41 <= 16'h562d;
        src42 <= 16'h1b26;
        src43 <= 16'h4815;
        src44 <= 16'hebef;
        src45 <= 16'hd447;
        src46 <= 16'hd808;
        src47 <= 16'hdb40;
        src48 <= 16'h172e;
        src49 <= 16'h2e74;
        src50 <= 16'haf7b;
        src51 <= 16'hc3d1;
        src52 <= 16'h48d1;
        src53 <= 16'h4c0c;
        src54 <= 16'h202b;
        src55 <= 16'hd827;
        src56 <= 16'h9d64;
        src57 <= 16'he88b;
        src58 <= 16'h1352;
        src59 <= 16'h41b1;
        src60 <= 16'h5865;
        src61 <= 16'h2ea;
        src62 <= 16'h121d;
        src63 <= 16'haae8;
        exp <= 22'h1baffc;
        #1
        src0 <= 16'hb14a;
        src1 <= 16'hc31c;
        src2 <= 16'ha0b2;
        src3 <= 16'haf52;
        src4 <= 16'h2f7;
        src5 <= 16'ha255;
        src6 <= 16'h5d1f;
        src7 <= 16'ha837;
        src8 <= 16'hd70a;
        src9 <= 16'hf326;
        src10 <= 16'h7fdc;
        src11 <= 16'hb20e;
        src12 <= 16'h196a;
        src13 <= 16'h231;
        src14 <= 16'hb468;
        src15 <= 16'h1cd;
        src16 <= 16'h16b9;
        src17 <= 16'h335e;
        src18 <= 16'h3627;
        src19 <= 16'h6407;
        src20 <= 16'h759a;
        src21 <= 16'hb8ce;
        src22 <= 16'h6edd;
        src23 <= 16'hec;
        src24 <= 16'hdba7;
        src25 <= 16'h6945;
        src26 <= 16'h7352;
        src27 <= 16'h8546;
        src28 <= 16'h49e8;
        src29 <= 16'ha794;
        src30 <= 16'h14fc;
        src31 <= 16'hbd0;
        src32 <= 16'hf971;
        src33 <= 16'he49f;
        src34 <= 16'h55e6;
        src35 <= 16'hf66e;
        src36 <= 16'hef5d;
        src37 <= 16'h9f76;
        src38 <= 16'h3576;
        src39 <= 16'h50a7;
        src40 <= 16'ha5b3;
        src41 <= 16'hbf69;
        src42 <= 16'h20b2;
        src43 <= 16'hfd36;
        src44 <= 16'hec12;
        src45 <= 16'hea50;
        src46 <= 16'h77ec;
        src47 <= 16'h4370;
        src48 <= 16'hdaae;
        src49 <= 16'h6270;
        src50 <= 16'hb5f4;
        src51 <= 16'hd2b1;
        src52 <= 16'h9a18;
        src53 <= 16'h4bf3;
        src54 <= 16'h9ac0;
        src55 <= 16'he9ec;
        src56 <= 16'ha683;
        src57 <= 16'h289b;
        src58 <= 16'hecd5;
        src59 <= 16'he0da;
        src60 <= 16'hf4a5;
        src61 <= 16'h6387;
        src62 <= 16'h3aa6;
        src63 <= 16'h6ec6;
        exp <= 22'h22322d;
        #1
        src0 <= 16'hde41;
        src1 <= 16'h11fe;
        src2 <= 16'hc16e;
        src3 <= 16'hb343;
        src4 <= 16'h2a6e;
        src5 <= 16'h9894;
        src6 <= 16'h1aea;
        src7 <= 16'h8cea;
        src8 <= 16'h6ab3;
        src9 <= 16'h46b6;
        src10 <= 16'hd8a7;
        src11 <= 16'h193b;
        src12 <= 16'h6644;
        src13 <= 16'h7e3c;
        src14 <= 16'hb0cd;
        src15 <= 16'h6559;
        src16 <= 16'hb97f;
        src17 <= 16'h5f97;
        src18 <= 16'h1d3b;
        src19 <= 16'hd3f0;
        src20 <= 16'hbfca;
        src21 <= 16'h3df4;
        src22 <= 16'h358c;
        src23 <= 16'hca87;
        src24 <= 16'h3161;
        src25 <= 16'he17d;
        src26 <= 16'h449c;
        src27 <= 16'h88c9;
        src28 <= 16'hd443;
        src29 <= 16'hfef6;
        src30 <= 16'h9cdf;
        src31 <= 16'hf119;
        src32 <= 16'h4f89;
        src33 <= 16'h4e87;
        src34 <= 16'h1614;
        src35 <= 16'h8769;
        src36 <= 16'hbfcc;
        src37 <= 16'h2718;
        src38 <= 16'hd0fc;
        src39 <= 16'hcd11;
        src40 <= 16'ha673;
        src41 <= 16'h8810;
        src42 <= 16'hf8f0;
        src43 <= 16'h14f2;
        src44 <= 16'h8393;
        src45 <= 16'hc8cd;
        src46 <= 16'hf36f;
        src47 <= 16'hcc36;
        src48 <= 16'ha604;
        src49 <= 16'he705;
        src50 <= 16'hde67;
        src51 <= 16'h20d3;
        src52 <= 16'h3331;
        src53 <= 16'hda6a;
        src54 <= 16'hbbef;
        src55 <= 16'h1189;
        src56 <= 16'hb7f6;
        src57 <= 16'h88a6;
        src58 <= 16'h508d;
        src59 <= 16'ha4ea;
        src60 <= 16'h12f4;
        src61 <= 16'hfebc;
        src62 <= 16'h9b00;
        src63 <= 16'hef0e;
        exp <= 22'h22f94c;
        #1
        src0 <= 16'h4f84;
        src1 <= 16'h8e28;
        src2 <= 16'h542f;
        src3 <= 16'hcf6b;
        src4 <= 16'ha02a;
        src5 <= 16'h385b;
        src6 <= 16'h6d41;
        src7 <= 16'h3472;
        src8 <= 16'h2175;
        src9 <= 16'hc4b2;
        src10 <= 16'h5ea1;
        src11 <= 16'h31;
        src12 <= 16'h58f7;
        src13 <= 16'hd3bd;
        src14 <= 16'he909;
        src15 <= 16'h79c2;
        src16 <= 16'hd311;
        src17 <= 16'h4236;
        src18 <= 16'hf6d2;
        src19 <= 16'h1863;
        src20 <= 16'h727e;
        src21 <= 16'hdd4a;
        src22 <= 16'h5220;
        src23 <= 16'h853a;
        src24 <= 16'h7c22;
        src25 <= 16'h337f;
        src26 <= 16'hd4a1;
        src27 <= 16'h9ddb;
        src28 <= 16'h8f68;
        src29 <= 16'ha800;
        src30 <= 16'hbfca;
        src31 <= 16'h1218;
        src32 <= 16'hdd10;
        src33 <= 16'h9781;
        src34 <= 16'h578e;
        src35 <= 16'h292c;
        src36 <= 16'hc18d;
        src37 <= 16'h19d0;
        src38 <= 16'h27ab;
        src39 <= 16'hdf3f;
        src40 <= 16'h70c0;
        src41 <= 16'hf083;
        src42 <= 16'hdb1a;
        src43 <= 16'h906a;
        src44 <= 16'hb2b4;
        src45 <= 16'h3c05;
        src46 <= 16'h2fba;
        src47 <= 16'haa82;
        src48 <= 16'h9dc8;
        src49 <= 16'hdda9;
        src50 <= 16'h51f0;
        src51 <= 16'h8dcb;
        src52 <= 16'hd944;
        src53 <= 16'h51cc;
        src54 <= 16'h7887;
        src55 <= 16'hcc23;
        src56 <= 16'hcfe7;
        src57 <= 16'h8064;
        src58 <= 16'h7390;
        src59 <= 16'h2bc4;
        src60 <= 16'ha1b9;
        src61 <= 16'hbe63;
        src62 <= 16'h9cf6;
        src63 <= 16'h3f6a;
        exp <= 22'h212b4a;
        #1
        src0 <= 16'hfee;
        src1 <= 16'he80f;
        src2 <= 16'h24a7;
        src3 <= 16'h5434;
        src4 <= 16'h3765;
        src5 <= 16'he0b7;
        src6 <= 16'he98a;
        src7 <= 16'hf194;
        src8 <= 16'h34af;
        src9 <= 16'h7b1c;
        src10 <= 16'h544d;
        src11 <= 16'hc6bd;
        src12 <= 16'h8f6a;
        src13 <= 16'hd0a4;
        src14 <= 16'h33a;
        src15 <= 16'h2f58;
        src16 <= 16'hd237;
        src17 <= 16'hc952;
        src18 <= 16'h7c1b;
        src19 <= 16'he1ce;
        src20 <= 16'h47ea;
        src21 <= 16'h75e3;
        src22 <= 16'hee8d;
        src23 <= 16'h2a06;
        src24 <= 16'he74c;
        src25 <= 16'h1093;
        src26 <= 16'h38b3;
        src27 <= 16'h118e;
        src28 <= 16'he4ad;
        src29 <= 16'h2378;
        src30 <= 16'h46fc;
        src31 <= 16'h4522;
        src32 <= 16'hdfb;
        src33 <= 16'h16a4;
        src34 <= 16'hc03d;
        src35 <= 16'ha95;
        src36 <= 16'h27fb;
        src37 <= 16'he12f;
        src38 <= 16'h92df;
        src39 <= 16'hae8c;
        src40 <= 16'hd585;
        src41 <= 16'hcadf;
        src42 <= 16'hd32e;
        src43 <= 16'hd978;
        src44 <= 16'h78da;
        src45 <= 16'h19c9;
        src46 <= 16'h9c8;
        src47 <= 16'h9982;
        src48 <= 16'h55e6;
        src49 <= 16'h1b2f;
        src50 <= 16'he5da;
        src51 <= 16'h8d32;
        src52 <= 16'h1560;
        src53 <= 16'h9117;
        src54 <= 16'hd87f;
        src55 <= 16'h860c;
        src56 <= 16'head9;
        src57 <= 16'h43db;
        src58 <= 16'h4ffa;
        src59 <= 16'h3c50;
        src60 <= 16'h3924;
        src61 <= 16'hfe43;
        src62 <= 16'hbb01;
        src63 <= 16'h9269;
        exp <= 22'h1f4dab;
        #1
        src0 <= 16'h6720;
        src1 <= 16'hc2d3;
        src2 <= 16'h6614;
        src3 <= 16'hf59c;
        src4 <= 16'hf719;
        src5 <= 16'hee96;
        src6 <= 16'hf741;
        src7 <= 16'hb2b1;
        src8 <= 16'he32e;
        src9 <= 16'hcb59;
        src10 <= 16'hd61f;
        src11 <= 16'h2ff8;
        src12 <= 16'hdaa3;
        src13 <= 16'ha2f;
        src14 <= 16'hd006;
        src15 <= 16'h79cb;
        src16 <= 16'ha694;
        src17 <= 16'ha971;
        src18 <= 16'h2dc5;
        src19 <= 16'h7947;
        src20 <= 16'hd8df;
        src21 <= 16'h44d9;
        src22 <= 16'hc4c2;
        src23 <= 16'hff4d;
        src24 <= 16'ha912;
        src25 <= 16'h7fb1;
        src26 <= 16'haee3;
        src27 <= 16'hc58b;
        src28 <= 16'haa9b;
        src29 <= 16'h8e2e;
        src30 <= 16'h172e;
        src31 <= 16'hc8f4;
        src32 <= 16'hcb16;
        src33 <= 16'h1e21;
        src34 <= 16'ha10a;
        src35 <= 16'h9fb2;
        src36 <= 16'h8f13;
        src37 <= 16'h9fab;
        src38 <= 16'h1b9f;
        src39 <= 16'h8c1f;
        src40 <= 16'h662d;
        src41 <= 16'he6ab;
        src42 <= 16'h70c;
        src43 <= 16'hee43;
        src44 <= 16'h86ad;
        src45 <= 16'h2841;
        src46 <= 16'h3671;
        src47 <= 16'h6579;
        src48 <= 16'hd9e1;
        src49 <= 16'hc2ed;
        src50 <= 16'h957a;
        src51 <= 16'h9fac;
        src52 <= 16'h6c61;
        src53 <= 16'h739;
        src54 <= 16'hce29;
        src55 <= 16'h20;
        src56 <= 16'ha328;
        src57 <= 16'h41d8;
        src58 <= 16'h7e37;
        src59 <= 16'h3005;
        src60 <= 16'hd06c;
        src61 <= 16'h821e;
        src62 <= 16'h9bb6;
        src63 <= 16'ha990;
        exp <= 22'h2453ca;
        #1
        src0 <= 16'hf661;
        src1 <= 16'h595d;
        src2 <= 16'haef2;
        src3 <= 16'h3641;
        src4 <= 16'h4470;
        src5 <= 16'h7617;
        src6 <= 16'hfe61;
        src7 <= 16'hcae5;
        src8 <= 16'h488b;
        src9 <= 16'h7501;
        src10 <= 16'h44ea;
        src11 <= 16'h5162;
        src12 <= 16'h5956;
        src13 <= 16'hb135;
        src14 <= 16'h24a2;
        src15 <= 16'h6861;
        src16 <= 16'hcde;
        src17 <= 16'h5572;
        src18 <= 16'hc7b5;
        src19 <= 16'habcf;
        src20 <= 16'ha783;
        src21 <= 16'hc95b;
        src22 <= 16'h7c87;
        src23 <= 16'hb9bc;
        src24 <= 16'hda10;
        src25 <= 16'hbd40;
        src26 <= 16'he10c;
        src27 <= 16'h9b16;
        src28 <= 16'hb952;
        src29 <= 16'hadd9;
        src30 <= 16'h93be;
        src31 <= 16'hb37d;
        src32 <= 16'h8681;
        src33 <= 16'h7563;
        src34 <= 16'hf906;
        src35 <= 16'h6d32;
        src36 <= 16'ha829;
        src37 <= 16'h7a15;
        src38 <= 16'ha5b6;
        src39 <= 16'h3752;
        src40 <= 16'hd198;
        src41 <= 16'ha0f2;
        src42 <= 16'hd9c3;
        src43 <= 16'h7319;
        src44 <= 16'h7a67;
        src45 <= 16'h65b2;
        src46 <= 16'h81a0;
        src47 <= 16'h6c91;
        src48 <= 16'h6be3;
        src49 <= 16'h28bf;
        src50 <= 16'he749;
        src51 <= 16'h79f9;
        src52 <= 16'h27d5;
        src53 <= 16'h162f;
        src54 <= 16'heb45;
        src55 <= 16'h3c77;
        src56 <= 16'hb72c;
        src57 <= 16'hda37;
        src58 <= 16'h5e7f;
        src59 <= 16'ha5e5;
        src60 <= 16'h57a1;
        src61 <= 16'h2159;
        src62 <= 16'he844;
        src63 <= 16'hf0e4;
        exp <= 22'h231590;
        #1
        src0 <= 16'h95ee;
        src1 <= 16'he5b5;
        src2 <= 16'hc2d9;
        src3 <= 16'h7363;
        src4 <= 16'hf0f8;
        src5 <= 16'hda8a;
        src6 <= 16'h237;
        src7 <= 16'h7925;
        src8 <= 16'h995a;
        src9 <= 16'hd379;
        src10 <= 16'h6a44;
        src11 <= 16'h905b;
        src12 <= 16'hc090;
        src13 <= 16'h688a;
        src14 <= 16'h648;
        src15 <= 16'hce1e;
        src16 <= 16'h6452;
        src17 <= 16'hc9c3;
        src18 <= 16'h78aa;
        src19 <= 16'h4ab;
        src20 <= 16'h7c95;
        src21 <= 16'h32ea;
        src22 <= 16'h1656;
        src23 <= 16'h5b2f;
        src24 <= 16'h835b;
        src25 <= 16'h62fd;
        src26 <= 16'hc789;
        src27 <= 16'hc0fc;
        src28 <= 16'h2264;
        src29 <= 16'hce37;
        src30 <= 16'h10c9;
        src31 <= 16'he36c;
        src32 <= 16'hddbe;
        src33 <= 16'h2a80;
        src34 <= 16'he1cc;
        src35 <= 16'h3e32;
        src36 <= 16'h3b32;
        src37 <= 16'hc1a9;
        src38 <= 16'hdc87;
        src39 <= 16'h3414;
        src40 <= 16'hc4bf;
        src41 <= 16'h1508;
        src42 <= 16'ha90d;
        src43 <= 16'haa11;
        src44 <= 16'ha05;
        src45 <= 16'hc456;
        src46 <= 16'ha182;
        src47 <= 16'h51de;
        src48 <= 16'h7973;
        src49 <= 16'h7b45;
        src50 <= 16'hb41c;
        src51 <= 16'h9d88;
        src52 <= 16'ha04f;
        src53 <= 16'h902b;
        src54 <= 16'h40d;
        src55 <= 16'h31b1;
        src56 <= 16'hb9ce;
        src57 <= 16'h50f7;
        src58 <= 16'hae9a;
        src59 <= 16'h69e0;
        src60 <= 16'h5103;
        src61 <= 16'h13f1;
        src62 <= 16'h3ba1;
        src63 <= 16'h7097;
        exp <= 22'h1f831b;
        #1
        src0 <= 16'h7d9c;
        src1 <= 16'ha084;
        src2 <= 16'h2e27;
        src3 <= 16'h9fa7;
        src4 <= 16'hd7f0;
        src5 <= 16'h3e53;
        src6 <= 16'h76df;
        src7 <= 16'ha2b7;
        src8 <= 16'h6b3f;
        src9 <= 16'h6b13;
        src10 <= 16'h956c;
        src11 <= 16'h4fe7;
        src12 <= 16'hf2ee;
        src13 <= 16'h8cc4;
        src14 <= 16'h2e31;
        src15 <= 16'hadf;
        src16 <= 16'he2c2;
        src17 <= 16'hfe5f;
        src18 <= 16'hd8b4;
        src19 <= 16'hb024;
        src20 <= 16'ha5e6;
        src21 <= 16'h5a52;
        src22 <= 16'hae53;
        src23 <= 16'h717f;
        src24 <= 16'h1561;
        src25 <= 16'h134c;
        src26 <= 16'he56b;
        src27 <= 16'h1fa9;
        src28 <= 16'h502c;
        src29 <= 16'h811e;
        src30 <= 16'h7067;
        src31 <= 16'hb13a;
        src32 <= 16'h56a4;
        src33 <= 16'hbac0;
        src34 <= 16'h83c2;
        src35 <= 16'hff8f;
        src36 <= 16'h7fe6;
        src37 <= 16'h54e5;
        src38 <= 16'h333a;
        src39 <= 16'hacd6;
        src40 <= 16'hb35;
        src41 <= 16'h338e;
        src42 <= 16'h2a0f;
        src43 <= 16'h6bb8;
        src44 <= 16'h46e2;
        src45 <= 16'h5f57;
        src46 <= 16'h37a4;
        src47 <= 16'h95eb;
        src48 <= 16'hf84e;
        src49 <= 16'h4041;
        src50 <= 16'h9e19;
        src51 <= 16'hb147;
        src52 <= 16'h9af6;
        src53 <= 16'h7688;
        src54 <= 16'h43f3;
        src55 <= 16'h7e89;
        src56 <= 16'hcda7;
        src57 <= 16'hcc22;
        src58 <= 16'hf892;
        src59 <= 16'h85f6;
        src60 <= 16'h77a3;
        src61 <= 16'h34b6;
        src62 <= 16'h5588;
        src63 <= 16'h5818;
        exp <= 22'h1f9af2;
        #1
        src0 <= 16'h28e3;
        src1 <= 16'hf60e;
        src2 <= 16'h47a2;
        src3 <= 16'h3498;
        src4 <= 16'h7335;
        src5 <= 16'hd070;
        src6 <= 16'h28b;
        src7 <= 16'h68bc;
        src8 <= 16'ha31b;
        src9 <= 16'hbc23;
        src10 <= 16'h54ed;
        src11 <= 16'hd00d;
        src12 <= 16'h9b12;
        src13 <= 16'h966b;
        src14 <= 16'h65f5;
        src15 <= 16'h7fdd;
        src16 <= 16'hb910;
        src17 <= 16'h3cb2;
        src18 <= 16'h2435;
        src19 <= 16'haee5;
        src20 <= 16'hffa7;
        src21 <= 16'hcc11;
        src22 <= 16'hae78;
        src23 <= 16'h35ca;
        src24 <= 16'h6cc9;
        src25 <= 16'he0be;
        src26 <= 16'h2086;
        src27 <= 16'h66ce;
        src28 <= 16'hdc5d;
        src29 <= 16'hee7d;
        src30 <= 16'he90f;
        src31 <= 16'h65c7;
        src32 <= 16'h586;
        src33 <= 16'h960;
        src34 <= 16'h81c0;
        src35 <= 16'h1bcd;
        src36 <= 16'h3e1c;
        src37 <= 16'hd60;
        src38 <= 16'h29ad;
        src39 <= 16'h7a89;
        src40 <= 16'h31be;
        src41 <= 16'h8ffb;
        src42 <= 16'hfca2;
        src43 <= 16'h1493;
        src44 <= 16'h309d;
        src45 <= 16'h906;
        src46 <= 16'hffd9;
        src47 <= 16'hd362;
        src48 <= 16'h50b5;
        src49 <= 16'h14b;
        src50 <= 16'h7972;
        src51 <= 16'h1598;
        src52 <= 16'hda20;
        src53 <= 16'hbd89;
        src54 <= 16'hf1b8;
        src55 <= 16'h8dd4;
        src56 <= 16'h8675;
        src57 <= 16'h3d69;
        src58 <= 16'h4b3b;
        src59 <= 16'ha642;
        src60 <= 16'h56e9;
        src61 <= 16'hae86;
        src62 <= 16'hbaa6;
        src63 <= 16'hf0cb;
        exp <= 22'h1f276a;
        #1
        src0 <= 16'hd4e3;
        src1 <= 16'ha702;
        src2 <= 16'h8699;
        src3 <= 16'he684;
        src4 <= 16'h37b5;
        src5 <= 16'h195e;
        src6 <= 16'hfe3e;
        src7 <= 16'hbf30;
        src8 <= 16'ha11f;
        src9 <= 16'h593;
        src10 <= 16'he00b;
        src11 <= 16'h1447;
        src12 <= 16'h18bc;
        src13 <= 16'h8059;
        src14 <= 16'hba11;
        src15 <= 16'h411b;
        src16 <= 16'hc1ee;
        src17 <= 16'h17d3;
        src18 <= 16'he0a0;
        src19 <= 16'he285;
        src20 <= 16'hd737;
        src21 <= 16'hb9e3;
        src22 <= 16'hd84a;
        src23 <= 16'h5b6b;
        src24 <= 16'h4e24;
        src25 <= 16'h8995;
        src26 <= 16'h20e6;
        src27 <= 16'hf48d;
        src28 <= 16'h4f5;
        src29 <= 16'h338f;
        src30 <= 16'h45a3;
        src31 <= 16'he31a;
        src32 <= 16'h8fd9;
        src33 <= 16'ha755;
        src34 <= 16'h5aaf;
        src35 <= 16'hd179;
        src36 <= 16'heb82;
        src37 <= 16'h8c9e;
        src38 <= 16'h57c4;
        src39 <= 16'h5701;
        src40 <= 16'h2a9c;
        src41 <= 16'he2e5;
        src42 <= 16'hf20a;
        src43 <= 16'h4c2c;
        src44 <= 16'haf03;
        src45 <= 16'h4a5f;
        src46 <= 16'hb3f5;
        src47 <= 16'hd38d;
        src48 <= 16'ha440;
        src49 <= 16'h3469;
        src50 <= 16'h1141;
        src51 <= 16'hde77;
        src52 <= 16'h9810;
        src53 <= 16'hcdbf;
        src54 <= 16'h6182;
        src55 <= 16'h125d;
        src56 <= 16'hb1bf;
        src57 <= 16'h611e;
        src58 <= 16'h4cd6;
        src59 <= 16'hbd8e;
        src60 <= 16'heb2d;
        src61 <= 16'h115a;
        src62 <= 16'ha1b1;
        src63 <= 16'h4a9a;
        exp <= 22'h21d5e2;
        #1
        src0 <= 16'h9c41;
        src1 <= 16'h8313;
        src2 <= 16'h39f3;
        src3 <= 16'hc743;
        src4 <= 16'h5c5b;
        src5 <= 16'hf59c;
        src6 <= 16'hbb92;
        src7 <= 16'hb912;
        src8 <= 16'h2b2e;
        src9 <= 16'h65b;
        src10 <= 16'hd87f;
        src11 <= 16'h4a94;
        src12 <= 16'h4d73;
        src13 <= 16'h35f6;
        src14 <= 16'hbe17;
        src15 <= 16'h6bbd;
        src16 <= 16'h3858;
        src17 <= 16'h963;
        src18 <= 16'h76f6;
        src19 <= 16'hf83c;
        src20 <= 16'hfee2;
        src21 <= 16'hfa67;
        src22 <= 16'h1b67;
        src23 <= 16'h6b58;
        src24 <= 16'h9aa1;
        src25 <= 16'h75f1;
        src26 <= 16'hf02;
        src27 <= 16'h7576;
        src28 <= 16'h202c;
        src29 <= 16'h5566;
        src30 <= 16'he2d;
        src31 <= 16'h7506;
        src32 <= 16'h3bb9;
        src33 <= 16'h1027;
        src34 <= 16'h663b;
        src35 <= 16'h7f34;
        src36 <= 16'h6657;
        src37 <= 16'h1725;
        src38 <= 16'hefd8;
        src39 <= 16'he2dc;
        src40 <= 16'h6b42;
        src41 <= 16'h99d1;
        src42 <= 16'h9eb1;
        src43 <= 16'hdd6e;
        src44 <= 16'hf5ae;
        src45 <= 16'ha8a7;
        src46 <= 16'h7cee;
        src47 <= 16'h7148;
        src48 <= 16'h63dd;
        src49 <= 16'h7650;
        src50 <= 16'h25f9;
        src51 <= 16'h5aba;
        src52 <= 16'h65a2;
        src53 <= 16'h4627;
        src54 <= 16'hee95;
        src55 <= 16'h385c;
        src56 <= 16'hfcf3;
        src57 <= 16'h5c44;
        src58 <= 16'h1a2b;
        src59 <= 16'hf289;
        src60 <= 16'hd6a5;
        src61 <= 16'hb486;
        src62 <= 16'h71f9;
        src63 <= 16'he869;
        exp <= 22'h1fb010;
        #1
        src0 <= 16'ha3d2;
        src1 <= 16'h42b0;
        src2 <= 16'hf256;
        src3 <= 16'h8829;
        src4 <= 16'h1ebb;
        src5 <= 16'h7b5a;
        src6 <= 16'haba;
        src7 <= 16'ha281;
        src8 <= 16'h1c4a;
        src9 <= 16'hae69;
        src10 <= 16'hc098;
        src11 <= 16'hb9e0;
        src12 <= 16'h9e8f;
        src13 <= 16'h4c75;
        src14 <= 16'haa5e;
        src15 <= 16'hd37f;
        src16 <= 16'he9a2;
        src17 <= 16'h801b;
        src18 <= 16'hadf0;
        src19 <= 16'h78a3;
        src20 <= 16'hd4f5;
        src21 <= 16'h7f85;
        src22 <= 16'hbaba;
        src23 <= 16'hbcb;
        src24 <= 16'hbffc;
        src25 <= 16'hdf0c;
        src26 <= 16'h1448;
        src27 <= 16'h6669;
        src28 <= 16'h6868;
        src29 <= 16'h5539;
        src30 <= 16'hd14;
        src31 <= 16'h3f6a;
        src32 <= 16'h4202;
        src33 <= 16'h8968;
        src34 <= 16'hde2b;
        src35 <= 16'h823f;
        src36 <= 16'h360e;
        src37 <= 16'h6a7d;
        src38 <= 16'h48f7;
        src39 <= 16'hf89;
        src40 <= 16'hbd23;
        src41 <= 16'hb850;
        src42 <= 16'h49d;
        src43 <= 16'h5065;
        src44 <= 16'h7c26;
        src45 <= 16'hf2e8;
        src46 <= 16'h71b5;
        src47 <= 16'h323e;
        src48 <= 16'ha4da;
        src49 <= 16'h5b8f;
        src50 <= 16'hf532;
        src51 <= 16'hdc62;
        src52 <= 16'hb7b0;
        src53 <= 16'h71f;
        src54 <= 16'hd3f1;
        src55 <= 16'hbde2;
        src56 <= 16'h779a;
        src57 <= 16'h24bc;
        src58 <= 16'h188e;
        src59 <= 16'h8a95;
        src60 <= 16'h2bbb;
        src61 <= 16'hc4e1;
        src62 <= 16'h8bd0;
        src63 <= 16'h5049;
        exp <= 22'h1f56a6;
        #1
        src0 <= 16'h92fd;
        src1 <= 16'h46c3;
        src2 <= 16'ha057;
        src3 <= 16'he180;
        src4 <= 16'he07d;
        src5 <= 16'ha399;
        src6 <= 16'h3b2c;
        src7 <= 16'hd1ad;
        src8 <= 16'h833a;
        src9 <= 16'h96f3;
        src10 <= 16'hfb;
        src11 <= 16'h3059;
        src12 <= 16'h412c;
        src13 <= 16'h86a1;
        src14 <= 16'hebdb;
        src15 <= 16'h25b0;
        src16 <= 16'hd055;
        src17 <= 16'h3e94;
        src18 <= 16'h142f;
        src19 <= 16'h23a1;
        src20 <= 16'h8970;
        src21 <= 16'h1a69;
        src22 <= 16'h2514;
        src23 <= 16'h317;
        src24 <= 16'hb442;
        src25 <= 16'h4ae2;
        src26 <= 16'ha6db;
        src27 <= 16'ha3f1;
        src28 <= 16'h5c93;
        src29 <= 16'hfc7d;
        src30 <= 16'h4a9;
        src31 <= 16'ha26;
        src32 <= 16'hf30f;
        src33 <= 16'h8781;
        src34 <= 16'hbf6e;
        src35 <= 16'h45d5;
        src36 <= 16'h70b9;
        src37 <= 16'h1a98;
        src38 <= 16'h3b57;
        src39 <= 16'h86b5;
        src40 <= 16'h1824;
        src41 <= 16'hffa;
        src42 <= 16'hfc52;
        src43 <= 16'ha7ee;
        src44 <= 16'hacf6;
        src45 <= 16'ha20e;
        src46 <= 16'h9a6f;
        src47 <= 16'hd04b;
        src48 <= 16'h4823;
        src49 <= 16'h8814;
        src50 <= 16'hb64f;
        src51 <= 16'h29f8;
        src52 <= 16'h6f9d;
        src53 <= 16'h9890;
        src54 <= 16'h92b0;
        src55 <= 16'h5c8d;
        src56 <= 16'h292a;
        src57 <= 16'hf825;
        src58 <= 16'h9c27;
        src59 <= 16'h970c;
        src60 <= 16'ha236;
        src61 <= 16'hed1a;
        src62 <= 16'hc29f;
        src63 <= 16'h9b8e;
        exp <= 22'h1f131e;
        #1
        src0 <= 16'ha650;
        src1 <= 16'hf4e9;
        src2 <= 16'h31e9;
        src3 <= 16'h1eb8;
        src4 <= 16'he103;
        src5 <= 16'hafd0;
        src6 <= 16'h9019;
        src7 <= 16'h240d;
        src8 <= 16'h660b;
        src9 <= 16'ha0c9;
        src10 <= 16'he61;
        src11 <= 16'h3164;
        src12 <= 16'h73a5;
        src13 <= 16'h3fba;
        src14 <= 16'hb935;
        src15 <= 16'hd7c1;
        src16 <= 16'h8ecb;
        src17 <= 16'h300a;
        src18 <= 16'h306d;
        src19 <= 16'hd82;
        src20 <= 16'h5590;
        src21 <= 16'h4bfb;
        src22 <= 16'hfbf9;
        src23 <= 16'h2e69;
        src24 <= 16'h215;
        src25 <= 16'h6329;
        src26 <= 16'h230f;
        src27 <= 16'h8f93;
        src28 <= 16'h5394;
        src29 <= 16'ha288;
        src30 <= 16'hf2ab;
        src31 <= 16'h6664;
        src32 <= 16'h8945;
        src33 <= 16'hc340;
        src34 <= 16'h48af;
        src35 <= 16'he7ee;
        src36 <= 16'haa1f;
        src37 <= 16'h144c;
        src38 <= 16'h851e;
        src39 <= 16'h8aa8;
        src40 <= 16'h78fe;
        src41 <= 16'hbbb7;
        src42 <= 16'h8f35;
        src43 <= 16'h3b59;
        src44 <= 16'h43b;
        src45 <= 16'h91f0;
        src46 <= 16'h450a;
        src47 <= 16'hafcf;
        src48 <= 16'h2f33;
        src49 <= 16'hd82a;
        src50 <= 16'haee0;
        src51 <= 16'h4483;
        src52 <= 16'h69ee;
        src53 <= 16'h1eae;
        src54 <= 16'hc51d;
        src55 <= 16'ha1d2;
        src56 <= 16'h2270;
        src57 <= 16'h62f7;
        src58 <= 16'h34ec;
        src59 <= 16'h5575;
        src60 <= 16'ha5a1;
        src61 <= 16'hac19;
        src62 <= 16'h1098;
        src63 <= 16'h7788;
        exp <= 22'h1c9504;
        #1
        src0 <= 16'haeb0;
        src1 <= 16'hb894;
        src2 <= 16'h5fff;
        src3 <= 16'hdfc5;
        src4 <= 16'hf21e;
        src5 <= 16'h3adf;
        src6 <= 16'he3f0;
        src7 <= 16'hed34;
        src8 <= 16'hd0e6;
        src9 <= 16'h35e5;
        src10 <= 16'h15ac;
        src11 <= 16'he5f0;
        src12 <= 16'h3b31;
        src13 <= 16'h7d94;
        src14 <= 16'h8130;
        src15 <= 16'ha24b;
        src16 <= 16'hb5a3;
        src17 <= 16'h2b01;
        src18 <= 16'h39de;
        src19 <= 16'h5e77;
        src20 <= 16'h6a4c;
        src21 <= 16'hc236;
        src22 <= 16'h2c5c;
        src23 <= 16'h4123;
        src24 <= 16'hba89;
        src25 <= 16'h23d3;
        src26 <= 16'h772a;
        src27 <= 16'heeac;
        src28 <= 16'hc704;
        src29 <= 16'he9bc;
        src30 <= 16'hb67c;
        src31 <= 16'he276;
        src32 <= 16'h5c34;
        src33 <= 16'h9933;
        src34 <= 16'h74d3;
        src35 <= 16'h25b5;
        src36 <= 16'he98;
        src37 <= 16'hb679;
        src38 <= 16'h9b66;
        src39 <= 16'h61ed;
        src40 <= 16'hc922;
        src41 <= 16'h8e5a;
        src42 <= 16'he781;
        src43 <= 16'h152b;
        src44 <= 16'hbaeb;
        src45 <= 16'hd54a;
        src46 <= 16'h2fe6;
        src47 <= 16'hbc2d;
        src48 <= 16'h148e;
        src49 <= 16'haef2;
        src50 <= 16'hc47b;
        src51 <= 16'h14ba;
        src52 <= 16'h28fb;
        src53 <= 16'h424b;
        src54 <= 16'h9bfd;
        src55 <= 16'h14e9;
        src56 <= 16'h4086;
        src57 <= 16'h7b75;
        src58 <= 16'hc992;
        src59 <= 16'h2609;
        src60 <= 16'hb9d1;
        src61 <= 16'hec86;
        src62 <= 16'h7be6;
        src63 <= 16'h63d8;
        exp <= 22'h2131fd;
        #1
        src0 <= 16'he772;
        src1 <= 16'hf5fa;
        src2 <= 16'h2e21;
        src3 <= 16'h46d8;
        src4 <= 16'h7986;
        src5 <= 16'h8345;
        src6 <= 16'h312d;
        src7 <= 16'h6bd5;
        src8 <= 16'h8a1e;
        src9 <= 16'hadd4;
        src10 <= 16'h7353;
        src11 <= 16'h3b28;
        src12 <= 16'h9347;
        src13 <= 16'hc14f;
        src14 <= 16'h9ada;
        src15 <= 16'h77b7;
        src16 <= 16'h6fcc;
        src17 <= 16'ha93d;
        src18 <= 16'hf49f;
        src19 <= 16'h9b18;
        src20 <= 16'h58d6;
        src21 <= 16'h30cb;
        src22 <= 16'h6791;
        src23 <= 16'h3fb6;
        src24 <= 16'h583e;
        src25 <= 16'h452e;
        src26 <= 16'ha344;
        src27 <= 16'h90b5;
        src28 <= 16'h9ede;
        src29 <= 16'h5e6b;
        src30 <= 16'h5f5f;
        src31 <= 16'hfb8c;
        src32 <= 16'h10f3;
        src33 <= 16'h5c92;
        src34 <= 16'hb4c8;
        src35 <= 16'h8750;
        src36 <= 16'h29f8;
        src37 <= 16'h728f;
        src38 <= 16'hebc;
        src39 <= 16'h9a62;
        src40 <= 16'he178;
        src41 <= 16'h788f;
        src42 <= 16'h9a66;
        src43 <= 16'hf34;
        src44 <= 16'h5855;
        src45 <= 16'h4beb;
        src46 <= 16'h61be;
        src47 <= 16'h2d4e;
        src48 <= 16'hdd98;
        src49 <= 16'hf603;
        src50 <= 16'h7ce6;
        src51 <= 16'h22bd;
        src52 <= 16'h89aa;
        src53 <= 16'h9bb5;
        src54 <= 16'h5e50;
        src55 <= 16'h8373;
        src56 <= 16'h447c;
        src57 <= 16'hc9a9;
        src58 <= 16'h8fc9;
        src59 <= 16'h49bc;
        src60 <= 16'h119;
        src61 <= 16'h6583;
        src62 <= 16'h7b9a;
        src63 <= 16'h9407;
        exp <= 22'h1e3b7d;
        #1
        src0 <= 16'h5b6b;
        src1 <= 16'hc869;
        src2 <= 16'h2e96;
        src3 <= 16'hdf9d;
        src4 <= 16'h55a;
        src5 <= 16'h6d03;
        src6 <= 16'hb822;
        src7 <= 16'h607a;
        src8 <= 16'h2124;
        src9 <= 16'h101b;
        src10 <= 16'h1c0b;
        src11 <= 16'h8558;
        src12 <= 16'h128d;
        src13 <= 16'hb283;
        src14 <= 16'hd3b;
        src15 <= 16'hd9bb;
        src16 <= 16'h9bb1;
        src17 <= 16'hecce;
        src18 <= 16'hdf05;
        src19 <= 16'h1a52;
        src20 <= 16'h5a56;
        src21 <= 16'he81b;
        src22 <= 16'h717e;
        src23 <= 16'h5ec7;
        src24 <= 16'hc81d;
        src25 <= 16'hb418;
        src26 <= 16'h982d;
        src27 <= 16'h3a93;
        src28 <= 16'hb844;
        src29 <= 16'ha7a6;
        src30 <= 16'h8bf4;
        src31 <= 16'h23e1;
        src32 <= 16'h437b;
        src33 <= 16'hf552;
        src34 <= 16'h3172;
        src35 <= 16'he50c;
        src36 <= 16'hf8d7;
        src37 <= 16'h65fe;
        src38 <= 16'h3bca;
        src39 <= 16'h95bb;
        src40 <= 16'h65fb;
        src41 <= 16'h57cc;
        src42 <= 16'hbb55;
        src43 <= 16'hb47;
        src44 <= 16'h4d01;
        src45 <= 16'h702b;
        src46 <= 16'hc6ec;
        src47 <= 16'hc873;
        src48 <= 16'ha73f;
        src49 <= 16'h371e;
        src50 <= 16'hb472;
        src51 <= 16'hd4c;
        src52 <= 16'hf39d;
        src53 <= 16'hc3c2;
        src54 <= 16'hc3dc;
        src55 <= 16'h25b3;
        src56 <= 16'h1bb6;
        src57 <= 16'h2944;
        src58 <= 16'ha6a9;
        src59 <= 16'h47d4;
        src60 <= 16'h832a;
        src61 <= 16'he04;
        src62 <= 16'hf8cf;
        src63 <= 16'h7ee;
        exp <= 22'h1e85e6;
        #1
        src0 <= 16'h60a8;
        src1 <= 16'h395e;
        src2 <= 16'hcee7;
        src3 <= 16'h9814;
        src4 <= 16'h8b06;
        src5 <= 16'hef65;
        src6 <= 16'h502f;
        src7 <= 16'h4780;
        src8 <= 16'h962c;
        src9 <= 16'hd73e;
        src10 <= 16'h3f3;
        src11 <= 16'hc182;
        src12 <= 16'hdcd1;
        src13 <= 16'h7402;
        src14 <= 16'hd9d2;
        src15 <= 16'h8892;
        src16 <= 16'hd262;
        src17 <= 16'hfc4c;
        src18 <= 16'hda12;
        src19 <= 16'h6895;
        src20 <= 16'he728;
        src21 <= 16'h7512;
        src22 <= 16'h7be3;
        src23 <= 16'haa70;
        src24 <= 16'h24b5;
        src25 <= 16'hf097;
        src26 <= 16'h7a39;
        src27 <= 16'h2cc3;
        src28 <= 16'h7c0d;
        src29 <= 16'hca97;
        src30 <= 16'h683f;
        src31 <= 16'h2e26;
        src32 <= 16'h42c5;
        src33 <= 16'hf92;
        src34 <= 16'h3e4e;
        src35 <= 16'h9527;
        src36 <= 16'h3716;
        src37 <= 16'h58a3;
        src38 <= 16'h947d;
        src39 <= 16'h3abf;
        src40 <= 16'h40d2;
        src41 <= 16'h14c3;
        src42 <= 16'ha62c;
        src43 <= 16'ha873;
        src44 <= 16'h97e7;
        src45 <= 16'hed26;
        src46 <= 16'h144b;
        src47 <= 16'h965d;
        src48 <= 16'h74b1;
        src49 <= 16'h46ed;
        src50 <= 16'h678;
        src51 <= 16'h3971;
        src52 <= 16'h1e89;
        src53 <= 16'hc16f;
        src54 <= 16'h22e;
        src55 <= 16'h7bbd;
        src56 <= 16'h21bb;
        src57 <= 16'h8cab;
        src58 <= 16'ha0fb;
        src59 <= 16'h2030;
        src60 <= 16'hbf5c;
        src61 <= 16'h9210;
        src62 <= 16'h8b4;
        src63 <= 16'h8db4;
        exp <= 22'h1e2fdd;
        #1
        src0 <= 16'he3a0;
        src1 <= 16'h3e90;
        src2 <= 16'h4549;
        src3 <= 16'hd96f;
        src4 <= 16'hf9c3;
        src5 <= 16'ha7a2;
        src6 <= 16'hc0b2;
        src7 <= 16'h3a4f;
        src8 <= 16'h25e4;
        src9 <= 16'hc9c7;
        src10 <= 16'hac0;
        src11 <= 16'h191d;
        src12 <= 16'h4d43;
        src13 <= 16'hf6b3;
        src14 <= 16'h5e41;
        src15 <= 16'h76b0;
        src16 <= 16'hd775;
        src17 <= 16'h23f3;
        src18 <= 16'hdd97;
        src19 <= 16'hfaa3;
        src20 <= 16'h7a5f;
        src21 <= 16'hf35;
        src22 <= 16'h6dad;
        src23 <= 16'h48c0;
        src24 <= 16'he3d7;
        src25 <= 16'hdadf;
        src26 <= 16'ha262;
        src27 <= 16'h3586;
        src28 <= 16'h8a42;
        src29 <= 16'hcd36;
        src30 <= 16'h7fc9;
        src31 <= 16'hd35e;
        src32 <= 16'h61d1;
        src33 <= 16'h573b;
        src34 <= 16'h9a9e;
        src35 <= 16'hc674;
        src36 <= 16'h8cce;
        src37 <= 16'h7da2;
        src38 <= 16'h3dc7;
        src39 <= 16'h4070;
        src40 <= 16'h42bd;
        src41 <= 16'h5915;
        src42 <= 16'h79d3;
        src43 <= 16'ha145;
        src44 <= 16'h5bea;
        src45 <= 16'ha921;
        src46 <= 16'h4dd1;
        src47 <= 16'h7f0e;
        src48 <= 16'hf6e8;
        src49 <= 16'h6509;
        src50 <= 16'h1df9;
        src51 <= 16'h8a4;
        src52 <= 16'hd4a0;
        src53 <= 16'hc142;
        src54 <= 16'h8362;
        src55 <= 16'h2e6;
        src56 <= 16'h53f4;
        src57 <= 16'h6dc4;
        src58 <= 16'hf031;
        src59 <= 16'h150f;
        src60 <= 16'haf36;
        src61 <= 16'h4e60;
        src62 <= 16'h159a;
        src63 <= 16'h7fcf;
        exp <= 22'h1f82e5;
        #1
        src0 <= 16'h3025;
        src1 <= 16'he7bd;
        src2 <= 16'h23f6;
        src3 <= 16'h30f;
        src4 <= 16'ha1bf;
        src5 <= 16'h8ab2;
        src6 <= 16'h4aad;
        src7 <= 16'h2aec;
        src8 <= 16'h4312;
        src9 <= 16'hc35e;
        src10 <= 16'hdb97;
        src11 <= 16'hf3dc;
        src12 <= 16'h1a4b;
        src13 <= 16'hbabc;
        src14 <= 16'hbcbc;
        src15 <= 16'h3c60;
        src16 <= 16'hc00b;
        src17 <= 16'h3d4;
        src18 <= 16'hcc19;
        src19 <= 16'h5213;
        src20 <= 16'h64d0;
        src21 <= 16'hf957;
        src22 <= 16'h8c23;
        src23 <= 16'ha9cd;
        src24 <= 16'h7da9;
        src25 <= 16'h5388;
        src26 <= 16'h4400;
        src27 <= 16'h4ebd;
        src28 <= 16'hf90d;
        src29 <= 16'h14fd;
        src30 <= 16'hd2d;
        src31 <= 16'h8d7d;
        src32 <= 16'h321d;
        src33 <= 16'hda81;
        src34 <= 16'hbcb6;
        src35 <= 16'h98ca;
        src36 <= 16'h8d16;
        src37 <= 16'h6240;
        src38 <= 16'heaaf;
        src39 <= 16'h24f8;
        src40 <= 16'h8a72;
        src41 <= 16'h623e;
        src42 <= 16'h298b;
        src43 <= 16'hada6;
        src44 <= 16'hfa0f;
        src45 <= 16'h9ffd;
        src46 <= 16'hdd73;
        src47 <= 16'hce68;
        src48 <= 16'he46c;
        src49 <= 16'h3458;
        src50 <= 16'hb2c8;
        src51 <= 16'h1428;
        src52 <= 16'hf2ab;
        src53 <= 16'hc593;
        src54 <= 16'hb4ed;
        src55 <= 16'h8d18;
        src56 <= 16'ha212;
        src57 <= 16'h862;
        src58 <= 16'h7d62;
        src59 <= 16'hb45e;
        src60 <= 16'h8ead;
        src61 <= 16'hf057;
        src62 <= 16'h3c9f;
        src63 <= 16'hf8e;
        exp <= 22'h20f3fa;
        #1
        src0 <= 16'h7229;
        src1 <= 16'hbdf4;
        src2 <= 16'h6223;
        src3 <= 16'h151;
        src4 <= 16'he1d3;
        src5 <= 16'hc20f;
        src6 <= 16'hd0bf;
        src7 <= 16'h65ec;
        src8 <= 16'h1891;
        src9 <= 16'hdb5;
        src10 <= 16'h95d9;
        src11 <= 16'h5635;
        src12 <= 16'h9c77;
        src13 <= 16'h1137;
        src14 <= 16'h9e8b;
        src15 <= 16'h6874;
        src16 <= 16'hbc28;
        src17 <= 16'h5054;
        src18 <= 16'h8137;
        src19 <= 16'h3a10;
        src20 <= 16'hae40;
        src21 <= 16'h4726;
        src22 <= 16'h4bd4;
        src23 <= 16'h64de;
        src24 <= 16'h9fb6;
        src25 <= 16'ha28c;
        src26 <= 16'h816b;
        src27 <= 16'h96ee;
        src28 <= 16'hb183;
        src29 <= 16'h1b9f;
        src30 <= 16'h7c79;
        src31 <= 16'hf7cb;
        src32 <= 16'hc42f;
        src33 <= 16'h90f8;
        src34 <= 16'h34f1;
        src35 <= 16'h4449;
        src36 <= 16'h5950;
        src37 <= 16'h24dc;
        src38 <= 16'hf365;
        src39 <= 16'haef3;
        src40 <= 16'hb8a6;
        src41 <= 16'h1138;
        src42 <= 16'h429;
        src43 <= 16'h7a99;
        src44 <= 16'h60cb;
        src45 <= 16'h94e8;
        src46 <= 16'hcac;
        src47 <= 16'hf1f6;
        src48 <= 16'h7b5f;
        src49 <= 16'h775f;
        src50 <= 16'h336b;
        src51 <= 16'h4aff;
        src52 <= 16'hbfd7;
        src53 <= 16'h9b1;
        src54 <= 16'h8654;
        src55 <= 16'h8343;
        src56 <= 16'h44f9;
        src57 <= 16'hba4c;
        src58 <= 16'h6cc6;
        src59 <= 16'h62ef;
        src60 <= 16'h6d41;
        src61 <= 16'he3f6;
        src62 <= 16'h5dfd;
        src63 <= 16'h3cdf;
        exp <= 22'h1d6a29;
        #1
        src0 <= 16'hc110;
        src1 <= 16'h84a0;
        src2 <= 16'hdadc;
        src3 <= 16'h312;
        src4 <= 16'h5b9;
        src5 <= 16'hdd1b;
        src6 <= 16'h71e9;
        src7 <= 16'he9d6;
        src8 <= 16'h5e79;
        src9 <= 16'h17bb;
        src10 <= 16'h27d9;
        src11 <= 16'h1767;
        src12 <= 16'ha3c9;
        src13 <= 16'h49d6;
        src14 <= 16'hb8e8;
        src15 <= 16'h7f2b;
        src16 <= 16'hcebe;
        src17 <= 16'h1e47;
        src18 <= 16'h3675;
        src19 <= 16'h29fe;
        src20 <= 16'h7ae9;
        src21 <= 16'hd504;
        src22 <= 16'h823d;
        src23 <= 16'hfeb1;
        src24 <= 16'h221a;
        src25 <= 16'hde20;
        src26 <= 16'hf43f;
        src27 <= 16'h9a44;
        src28 <= 16'h10c9;
        src29 <= 16'h4bd1;
        src30 <= 16'h66fb;
        src31 <= 16'hfef6;
        src32 <= 16'heaad;
        src33 <= 16'h9b22;
        src34 <= 16'hc95;
        src35 <= 16'h747e;
        src36 <= 16'hd03;
        src37 <= 16'h9b06;
        src38 <= 16'hadce;
        src39 <= 16'h787a;
        src40 <= 16'he225;
        src41 <= 16'h4550;
        src42 <= 16'h522b;
        src43 <= 16'ha95d;
        src44 <= 16'h579a;
        src45 <= 16'h6efc;
        src46 <= 16'ha035;
        src47 <= 16'h8e3a;
        src48 <= 16'hc860;
        src49 <= 16'hc19f;
        src50 <= 16'h2dcc;
        src51 <= 16'hc1ec;
        src52 <= 16'h74cc;
        src53 <= 16'h612d;
        src54 <= 16'h54c9;
        src55 <= 16'h4b79;
        src56 <= 16'he9bd;
        src57 <= 16'h2ee3;
        src58 <= 16'h4426;
        src59 <= 16'h5943;
        src60 <= 16'h676b;
        src61 <= 16'ha125;
        src62 <= 16'ha4d0;
        src63 <= 16'h5e93;
        exp <= 22'h1f4c15;
        #1
        src0 <= 16'h6a62;
        src1 <= 16'h5629;
        src2 <= 16'h7c6b;
        src3 <= 16'h3ec5;
        src4 <= 16'h96a7;
        src5 <= 16'h2df7;
        src6 <= 16'hd6b5;
        src7 <= 16'h6c0f;
        src8 <= 16'h7dc;
        src9 <= 16'h89e5;
        src10 <= 16'h91a8;
        src11 <= 16'h109d;
        src12 <= 16'hff92;
        src13 <= 16'h28b7;
        src14 <= 16'hb20b;
        src15 <= 16'h23c3;
        src16 <= 16'hb89a;
        src17 <= 16'h3c12;
        src18 <= 16'hd77d;
        src19 <= 16'h1943;
        src20 <= 16'h5d6e;
        src21 <= 16'h42ca;
        src22 <= 16'h6ab7;
        src23 <= 16'h74e2;
        src24 <= 16'h17e9;
        src25 <= 16'h9502;
        src26 <= 16'hff5b;
        src27 <= 16'h5b2d;
        src28 <= 16'hf7e4;
        src29 <= 16'hca11;
        src30 <= 16'hb255;
        src31 <= 16'hb030;
        src32 <= 16'h72e8;
        src33 <= 16'h7a6d;
        src34 <= 16'h774;
        src35 <= 16'h2bb8;
        src36 <= 16'ha7fa;
        src37 <= 16'hccbe;
        src38 <= 16'h7b2c;
        src39 <= 16'h580e;
        src40 <= 16'hbfb1;
        src41 <= 16'h882;
        src42 <= 16'h69e3;
        src43 <= 16'hcf64;
        src44 <= 16'h70e7;
        src45 <= 16'hd069;
        src46 <= 16'h8b64;
        src47 <= 16'h12ca;
        src48 <= 16'h4b3c;
        src49 <= 16'hd17;
        src50 <= 16'he3b9;
        src51 <= 16'hc6f7;
        src52 <= 16'h13d4;
        src53 <= 16'hd87a;
        src54 <= 16'hbba2;
        src55 <= 16'h4a19;
        src56 <= 16'hcbdf;
        src57 <= 16'h8e0e;
        src58 <= 16'h5cb6;
        src59 <= 16'h1393;
        src60 <= 16'h28b0;
        src61 <= 16'h3c0f;
        src62 <= 16'h9a0d;
        src63 <= 16'hbba7;
        exp <= 22'h1e0984;
        #1
        src0 <= 16'h1789;
        src1 <= 16'h2947;
        src2 <= 16'hc76f;
        src3 <= 16'h6eec;
        src4 <= 16'h5918;
        src5 <= 16'h971f;
        src6 <= 16'h5192;
        src7 <= 16'h134b;
        src8 <= 16'h7dcb;
        src9 <= 16'hfd2c;
        src10 <= 16'h63ad;
        src11 <= 16'h6ca3;
        src12 <= 16'hde1d;
        src13 <= 16'h51b9;
        src14 <= 16'h7b49;
        src15 <= 16'h342f;
        src16 <= 16'hc40e;
        src17 <= 16'ha098;
        src18 <= 16'h81ed;
        src19 <= 16'h9a11;
        src20 <= 16'h6a78;
        src21 <= 16'hc1d3;
        src22 <= 16'h6a87;
        src23 <= 16'hbae2;
        src24 <= 16'h7150;
        src25 <= 16'h6345;
        src26 <= 16'h5426;
        src27 <= 16'hd34e;
        src28 <= 16'hee60;
        src29 <= 16'ha250;
        src30 <= 16'h279b;
        src31 <= 16'hc289;
        src32 <= 16'hec4c;
        src33 <= 16'hd048;
        src34 <= 16'h690f;
        src35 <= 16'he1f7;
        src36 <= 16'hd6d2;
        src37 <= 16'h5fc7;
        src38 <= 16'h2a94;
        src39 <= 16'h34de;
        src40 <= 16'hbb4a;
        src41 <= 16'h70e6;
        src42 <= 16'h9309;
        src43 <= 16'h4596;
        src44 <= 16'h3bf3;
        src45 <= 16'h7f05;
        src46 <= 16'hfad;
        src47 <= 16'hf81d;
        src48 <= 16'h1e71;
        src49 <= 16'h4613;
        src50 <= 16'hf1f4;
        src51 <= 16'h694e;
        src52 <= 16'h7a37;
        src53 <= 16'h3598;
        src54 <= 16'h41a9;
        src55 <= 16'h94fb;
        src56 <= 16'hc65c;
        src57 <= 16'h87cc;
        src58 <= 16'hf41;
        src59 <= 16'h3c7c;
        src60 <= 16'h55b2;
        src61 <= 16'h2243;
        src62 <= 16'h2412;
        src63 <= 16'h7299;
        exp <= 22'h1e93fd;
        #1
        src0 <= 16'ha47e;
        src1 <= 16'hae5b;
        src2 <= 16'hbfb8;
        src3 <= 16'h464a;
        src4 <= 16'h74dc;
        src5 <= 16'h8ea4;
        src6 <= 16'hcdb0;
        src7 <= 16'hf594;
        src8 <= 16'h2ec9;
        src9 <= 16'h3068;
        src10 <= 16'h74fb;
        src11 <= 16'h12cb;
        src12 <= 16'ha7b9;
        src13 <= 16'hecc5;
        src14 <= 16'h9fe3;
        src15 <= 16'h1785;
        src16 <= 16'hf8d0;
        src17 <= 16'h5082;
        src18 <= 16'hb2f;
        src19 <= 16'h6fc3;
        src20 <= 16'habbf;
        src21 <= 16'hf5f;
        src22 <= 16'h552;
        src23 <= 16'hd0ee;
        src24 <= 16'h7855;
        src25 <= 16'hdea1;
        src26 <= 16'h5f9b;
        src27 <= 16'h3432;
        src28 <= 16'h4999;
        src29 <= 16'h125d;
        src30 <= 16'h953a;
        src31 <= 16'h27d9;
        src32 <= 16'h51a0;
        src33 <= 16'h8330;
        src34 <= 16'hcbfa;
        src35 <= 16'ha08d;
        src36 <= 16'hd1d9;
        src37 <= 16'h7bf2;
        src38 <= 16'hf1f1;
        src39 <= 16'h8bdc;
        src40 <= 16'h7fab;
        src41 <= 16'hb504;
        src42 <= 16'h27e0;
        src43 <= 16'h64ac;
        src44 <= 16'h1595;
        src45 <= 16'h3845;
        src46 <= 16'h300a;
        src47 <= 16'h7bc3;
        src48 <= 16'h4349;
        src49 <= 16'h4829;
        src50 <= 16'ha9da;
        src51 <= 16'hbe5e;
        src52 <= 16'h30cc;
        src53 <= 16'h1d6b;
        src54 <= 16'hf186;
        src55 <= 16'h159d;
        src56 <= 16'ha680;
        src57 <= 16'he11b;
        src58 <= 16'h70b4;
        src59 <= 16'h5444;
        src60 <= 16'ha612;
        src61 <= 16'h4c5d;
        src62 <= 16'hc466;
        src63 <= 16'h77b4;
        exp <= 22'h1e37db;
        #1
        src0 <= 16'h15b0;
        src1 <= 16'hb6a6;
        src2 <= 16'h298e;
        src3 <= 16'hc303;
        src4 <= 16'h9d01;
        src5 <= 16'hb7b9;
        src6 <= 16'he007;
        src7 <= 16'he192;
        src8 <= 16'h9bc2;
        src9 <= 16'he757;
        src10 <= 16'h4d5d;
        src11 <= 16'hf8ed;
        src12 <= 16'hcb1f;
        src13 <= 16'h62f9;
        src14 <= 16'hdfbc;
        src15 <= 16'h3406;
        src16 <= 16'hde5;
        src17 <= 16'hf62d;
        src18 <= 16'h8f15;
        src19 <= 16'h46c7;
        src20 <= 16'h32d4;
        src21 <= 16'he474;
        src22 <= 16'h5661;
        src23 <= 16'hd800;
        src24 <= 16'h7b7a;
        src25 <= 16'h1236;
        src26 <= 16'h8e59;
        src27 <= 16'h3e94;
        src28 <= 16'hd0a5;
        src29 <= 16'h1b30;
        src30 <= 16'h9fb2;
        src31 <= 16'ha539;
        src32 <= 16'h627d;
        src33 <= 16'hd77;
        src34 <= 16'h8397;
        src35 <= 16'hf679;
        src36 <= 16'h402c;
        src37 <= 16'hea27;
        src38 <= 16'h685a;
        src39 <= 16'ha5e0;
        src40 <= 16'h24a8;
        src41 <= 16'h98d5;
        src42 <= 16'hbc9d;
        src43 <= 16'h5378;
        src44 <= 16'h1c9e;
        src45 <= 16'h6a4c;
        src46 <= 16'h10ed;
        src47 <= 16'hc6cf;
        src48 <= 16'h6b33;
        src49 <= 16'hd98c;
        src50 <= 16'h7538;
        src51 <= 16'h67ff;
        src52 <= 16'hd398;
        src53 <= 16'hb80c;
        src54 <= 16'h11e7;
        src55 <= 16'h1430;
        src56 <= 16'h1e49;
        src57 <= 16'h1ce;
        src58 <= 16'hf8c9;
        src59 <= 16'h6c1f;
        src60 <= 16'h12a3;
        src61 <= 16'h606f;
        src62 <= 16'h3ddd;
        src63 <= 16'h4cb4;
        exp <= 22'h1f2a87;
        #1
        src0 <= 16'h521f;
        src1 <= 16'h8f90;
        src2 <= 16'h33df;
        src3 <= 16'h9c08;
        src4 <= 16'h4389;
        src5 <= 16'h75c;
        src6 <= 16'hc0bd;
        src7 <= 16'h434a;
        src8 <= 16'hf1b3;
        src9 <= 16'hfacd;
        src10 <= 16'hb5c;
        src11 <= 16'h3f24;
        src12 <= 16'ha3d9;
        src13 <= 16'h7676;
        src14 <= 16'h3beb;
        src15 <= 16'he4c1;
        src16 <= 16'ha2c7;
        src17 <= 16'h4839;
        src18 <= 16'h5f06;
        src19 <= 16'h3074;
        src20 <= 16'hbd4a;
        src21 <= 16'h379b;
        src22 <= 16'hdde6;
        src23 <= 16'h2966;
        src24 <= 16'hf1ae;
        src25 <= 16'ha2ff;
        src26 <= 16'hd2e3;
        src27 <= 16'h9dbc;
        src28 <= 16'hf313;
        src29 <= 16'ha9c0;
        src30 <= 16'h524e;
        src31 <= 16'h9b8d;
        src32 <= 16'he113;
        src33 <= 16'h43d7;
        src34 <= 16'h8e0d;
        src35 <= 16'haa65;
        src36 <= 16'h8597;
        src37 <= 16'had00;
        src38 <= 16'hbc6f;
        src39 <= 16'hc416;
        src40 <= 16'h1b1d;
        src41 <= 16'h1a9;
        src42 <= 16'h7033;
        src43 <= 16'h21e8;
        src44 <= 16'h9a4a;
        src45 <= 16'hd61a;
        src46 <= 16'h2fcc;
        src47 <= 16'ha69b;
        src48 <= 16'h621;
        src49 <= 16'h77f7;
        src50 <= 16'hc20d;
        src51 <= 16'h319a;
        src52 <= 16'h95d0;
        src53 <= 16'hdd06;
        src54 <= 16'he884;
        src55 <= 16'h4657;
        src56 <= 16'hf6d2;
        src57 <= 16'hde0a;
        src58 <= 16'hc72b;
        src59 <= 16'h15e8;
        src60 <= 16'hfb66;
        src61 <= 16'h3b52;
        src62 <= 16'h3be3;
        src63 <= 16'h3587;
        exp <= 22'h20ecc7;
        #1
        src0 <= 16'hf9ae;
        src1 <= 16'hba1a;
        src2 <= 16'h9b56;
        src3 <= 16'h1d49;
        src4 <= 16'hfd27;
        src5 <= 16'h5c1;
        src6 <= 16'h56c1;
        src7 <= 16'h507c;
        src8 <= 16'hf3e3;
        src9 <= 16'h8d8c;
        src10 <= 16'hedc2;
        src11 <= 16'hae95;
        src12 <= 16'h981e;
        src13 <= 16'hd0c5;
        src14 <= 16'hd478;
        src15 <= 16'h347f;
        src16 <= 16'h1f0f;
        src17 <= 16'he896;
        src18 <= 16'hcc93;
        src19 <= 16'hc3d5;
        src20 <= 16'hee72;
        src21 <= 16'h5d80;
        src22 <= 16'h5b93;
        src23 <= 16'h1449;
        src24 <= 16'h6449;
        src25 <= 16'hd518;
        src26 <= 16'ha86f;
        src27 <= 16'h6f47;
        src28 <= 16'h4251;
        src29 <= 16'hd15;
        src30 <= 16'hdbf3;
        src31 <= 16'h7c3f;
        src32 <= 16'he558;
        src33 <= 16'h4baa;
        src34 <= 16'h9685;
        src35 <= 16'hdbac;
        src36 <= 16'ha11;
        src37 <= 16'he6a7;
        src38 <= 16'h1ef9;
        src39 <= 16'hc437;
        src40 <= 16'hbc51;
        src41 <= 16'h8be5;
        src42 <= 16'hc742;
        src43 <= 16'hd97c;
        src44 <= 16'hce5f;
        src45 <= 16'h1ed2;
        src46 <= 16'hf912;
        src47 <= 16'h8685;
        src48 <= 16'hb318;
        src49 <= 16'hfa1a;
        src50 <= 16'h6ba6;
        src51 <= 16'h4fee;
        src52 <= 16'h320c;
        src53 <= 16'h125a;
        src54 <= 16'h45;
        src55 <= 16'h80b9;
        src56 <= 16'h9f9e;
        src57 <= 16'h27dc;
        src58 <= 16'hc851;
        src59 <= 16'h3e1a;
        src60 <= 16'h6a37;
        src61 <= 16'hb999;
        src62 <= 16'h1e3e;
        src63 <= 16'h4004;
        exp <= 22'h223dae;
        #1
        src0 <= 16'hfb5;
        src1 <= 16'h6679;
        src2 <= 16'h1fbd;
        src3 <= 16'h27a6;
        src4 <= 16'hc18a;
        src5 <= 16'hd7e7;
        src6 <= 16'hddd6;
        src7 <= 16'h8126;
        src8 <= 16'hc72d;
        src9 <= 16'hee0c;
        src10 <= 16'h9634;
        src11 <= 16'haee5;
        src12 <= 16'h71c3;
        src13 <= 16'h7a45;
        src14 <= 16'h8c41;
        src15 <= 16'h8a4d;
        src16 <= 16'h8067;
        src17 <= 16'h9312;
        src18 <= 16'h77ff;
        src19 <= 16'hd0f9;
        src20 <= 16'ha724;
        src21 <= 16'haa4;
        src22 <= 16'hd49;
        src23 <= 16'h2d30;
        src24 <= 16'ha233;
        src25 <= 16'h8f16;
        src26 <= 16'h1378;
        src27 <= 16'h6099;
        src28 <= 16'h3534;
        src29 <= 16'he3d3;
        src30 <= 16'hbe20;
        src31 <= 16'h69f4;
        src32 <= 16'h4ae0;
        src33 <= 16'hb5fa;
        src34 <= 16'hda4d;
        src35 <= 16'hb637;
        src36 <= 16'hf09f;
        src37 <= 16'h63db;
        src38 <= 16'h71b5;
        src39 <= 16'h9c37;
        src40 <= 16'h4120;
        src41 <= 16'h7030;
        src42 <= 16'h112;
        src43 <= 16'hf0ef;
        src44 <= 16'h6540;
        src45 <= 16'hb975;
        src46 <= 16'ha0d9;
        src47 <= 16'hd03c;
        src48 <= 16'h68d5;
        src49 <= 16'h7d69;
        src50 <= 16'hdd61;
        src51 <= 16'hd2c6;
        src52 <= 16'he5b8;
        src53 <= 16'haedf;
        src54 <= 16'h5df1;
        src55 <= 16'h8ebc;
        src56 <= 16'hbccc;
        src57 <= 16'h7fe4;
        src58 <= 16'h2e89;
        src59 <= 16'ha0b2;
        src60 <= 16'hdde1;
        src61 <= 16'hd9be;
        src62 <= 16'h6561;
        src63 <= 16'hce85;
        exp <= 22'h231805;
        #1
        src0 <= 16'hd98f;
        src1 <= 16'h78ec;
        src2 <= 16'hb5c8;
        src3 <= 16'h330;
        src4 <= 16'hf70e;
        src5 <= 16'had00;
        src6 <= 16'he96f;
        src7 <= 16'h124a;
        src8 <= 16'h3856;
        src9 <= 16'h7685;
        src10 <= 16'h3151;
        src11 <= 16'h2d1f;
        src12 <= 16'hb8c3;
        src13 <= 16'hea44;
        src14 <= 16'h1b72;
        src15 <= 16'hb2ea;
        src16 <= 16'hf4f9;
        src17 <= 16'hd0e4;
        src18 <= 16'ha5a6;
        src19 <= 16'h6f41;
        src20 <= 16'hc3d7;
        src21 <= 16'h550f;
        src22 <= 16'h8f55;
        src23 <= 16'h5966;
        src24 <= 16'h2678;
        src25 <= 16'h4fbe;
        src26 <= 16'ha41f;
        src27 <= 16'h57d4;
        src28 <= 16'hc6ba;
        src29 <= 16'hcc55;
        src30 <= 16'h6d89;
        src31 <= 16'hf24;
        src32 <= 16'h5187;
        src33 <= 16'ha97d;
        src34 <= 16'hdcb9;
        src35 <= 16'h8291;
        src36 <= 16'h4a3;
        src37 <= 16'hd832;
        src38 <= 16'h5e6d;
        src39 <= 16'h20bd;
        src40 <= 16'h42a9;
        src41 <= 16'he166;
        src42 <= 16'h7d9e;
        src43 <= 16'h6f66;
        src44 <= 16'h6010;
        src45 <= 16'hdfea;
        src46 <= 16'hfd0d;
        src47 <= 16'h6861;
        src48 <= 16'hb951;
        src49 <= 16'h7be8;
        src50 <= 16'h78c8;
        src51 <= 16'h4b7d;
        src52 <= 16'h2718;
        src53 <= 16'ha9a6;
        src54 <= 16'h6eb0;
        src55 <= 16'hb52b;
        src56 <= 16'hcfcf;
        src57 <= 16'h1925;
        src58 <= 16'h46b3;
        src59 <= 16'hc7b9;
        src60 <= 16'h2514;
        src61 <= 16'h5869;
        src62 <= 16'h5013;
        src63 <= 16'h65c6;
        exp <= 22'h200dc7;
        #1
        src0 <= 16'h83d7;
        src1 <= 16'h9459;
        src2 <= 16'hc098;
        src3 <= 16'hd3e0;
        src4 <= 16'h9694;
        src5 <= 16'haa83;
        src6 <= 16'h3f04;
        src7 <= 16'h88f0;
        src8 <= 16'h8426;
        src9 <= 16'h2967;
        src10 <= 16'h8d3d;
        src11 <= 16'hef0e;
        src12 <= 16'h21e;
        src13 <= 16'h6aa7;
        src14 <= 16'haf4d;
        src15 <= 16'he558;
        src16 <= 16'h6f0f;
        src17 <= 16'h6449;
        src18 <= 16'h6318;
        src19 <= 16'ha7c;
        src20 <= 16'hba41;
        src21 <= 16'hca85;
        src22 <= 16'h46d9;
        src23 <= 16'hf503;
        src24 <= 16'h550d;
        src25 <= 16'h850a;
        src26 <= 16'hee2c;
        src27 <= 16'h8aa7;
        src28 <= 16'h2f96;
        src29 <= 16'h50b4;
        src30 <= 16'h375d;
        src31 <= 16'hb860;
        src32 <= 16'hf843;
        src33 <= 16'hb596;
        src34 <= 16'h1560;
        src35 <= 16'h1ecd;
        src36 <= 16'h4572;
        src37 <= 16'hc7d9;
        src38 <= 16'he271;
        src39 <= 16'heda;
        src40 <= 16'h2c3f;
        src41 <= 16'hb9f9;
        src42 <= 16'h5054;
        src43 <= 16'h69ed;
        src44 <= 16'h44a;
        src45 <= 16'h230f;
        src46 <= 16'hf14a;
        src47 <= 16'h2949;
        src48 <= 16'h9eeb;
        src49 <= 16'h6a4f;
        src50 <= 16'he384;
        src51 <= 16'h9213;
        src52 <= 16'hfc98;
        src53 <= 16'h9202;
        src54 <= 16'h28e1;
        src55 <= 16'he8bc;
        src56 <= 16'h2d6c;
        src57 <= 16'hfbfc;
        src58 <= 16'heb15;
        src59 <= 16'h7e2f;
        src60 <= 16'h30d2;
        src61 <= 16'h7eeb;
        src62 <= 16'h8506;
        src63 <= 16'he5ca;
        exp <= 22'h2134b6;
        #1
        src0 <= 16'h1acc;
        src1 <= 16'hc92c;
        src2 <= 16'haff5;
        src3 <= 16'he51b;
        src4 <= 16'hd4cf;
        src5 <= 16'h59f6;
        src6 <= 16'h8545;
        src7 <= 16'hfd2a;
        src8 <= 16'hc927;
        src9 <= 16'h2465;
        src10 <= 16'h3959;
        src11 <= 16'hbb1;
        src12 <= 16'he40f;
        src13 <= 16'h7c72;
        src14 <= 16'he199;
        src15 <= 16'hdad9;
        src16 <= 16'h32c2;
        src17 <= 16'h8dc3;
        src18 <= 16'he605;
        src19 <= 16'hec98;
        src20 <= 16'h9af9;
        src21 <= 16'h2994;
        src22 <= 16'hbd48;
        src23 <= 16'ha823;
        src24 <= 16'h97da;
        src25 <= 16'he4e4;
        src26 <= 16'h603e;
        src27 <= 16'h36c0;
        src28 <= 16'h7c0c;
        src29 <= 16'h87da;
        src30 <= 16'hf892;
        src31 <= 16'h5035;
        src32 <= 16'he4bb;
        src33 <= 16'hbbda;
        src34 <= 16'hc743;
        src35 <= 16'h466e;
        src36 <= 16'h9d28;
        src37 <= 16'h9e5e;
        src38 <= 16'h5bb5;
        src39 <= 16'hbfeb;
        src40 <= 16'h4ac1;
        src41 <= 16'h876b;
        src42 <= 16'h91c7;
        src43 <= 16'hfb6d;
        src44 <= 16'hdd8e;
        src45 <= 16'h3c23;
        src46 <= 16'h9db3;
        src47 <= 16'hcd7d;
        src48 <= 16'h41c8;
        src49 <= 16'hfbbc;
        src50 <= 16'hfe94;
        src51 <= 16'he794;
        src52 <= 16'h2683;
        src53 <= 16'h44e9;
        src54 <= 16'heaea;
        src55 <= 16'h7362;
        src56 <= 16'h7f39;
        src57 <= 16'h4897;
        src58 <= 16'hb1eb;
        src59 <= 16'h5696;
        src60 <= 16'h5209;
        src61 <= 16'h5790;
        src62 <= 16'hba25;
        src63 <= 16'h43ca;
        exp <= 22'h24e632;
        #1
        src0 <= 16'h8c;
        src1 <= 16'h9b12;
        src2 <= 16'he5d1;
        src3 <= 16'hb236;
        src4 <= 16'h96e7;
        src5 <= 16'h33e8;
        src6 <= 16'h3232;
        src7 <= 16'h88da;
        src8 <= 16'h6650;
        src9 <= 16'hf4d;
        src10 <= 16'h9e52;
        src11 <= 16'hc9b9;
        src12 <= 16'hced5;
        src13 <= 16'h2c38;
        src14 <= 16'h6aa2;
        src15 <= 16'hebcb;
        src16 <= 16'h18a8;
        src17 <= 16'hc41b;
        src18 <= 16'ha6e6;
        src19 <= 16'hbafc;
        src20 <= 16'h3b90;
        src21 <= 16'he7d8;
        src22 <= 16'ha713;
        src23 <= 16'h9d74;
        src24 <= 16'h70c3;
        src25 <= 16'h70dd;
        src26 <= 16'h3212;
        src27 <= 16'hf1cb;
        src28 <= 16'h9335;
        src29 <= 16'h2aeb;
        src30 <= 16'h5e23;
        src31 <= 16'h63fa;
        src32 <= 16'hf3dc;
        src33 <= 16'h703b;
        src34 <= 16'h1067;
        src35 <= 16'h1f9;
        src36 <= 16'h7ab4;
        src37 <= 16'hbd86;
        src38 <= 16'hee8c;
        src39 <= 16'hb2f2;
        src40 <= 16'h3587;
        src41 <= 16'hc205;
        src42 <= 16'hcc36;
        src43 <= 16'h3874;
        src44 <= 16'hbb3f;
        src45 <= 16'h5fa6;
        src46 <= 16'hea97;
        src47 <= 16'h9bd;
        src48 <= 16'he20;
        src49 <= 16'h33b;
        src50 <= 16'h5117;
        src51 <= 16'hb2e8;
        src52 <= 16'h781a;
        src53 <= 16'hefa2;
        src54 <= 16'hf0c1;
        src55 <= 16'h7a45;
        src56 <= 16'h9a2b;
        src57 <= 16'ha0e1;
        src58 <= 16'h8c10;
        src59 <= 16'hd806;
        src60 <= 16'ha3ed;
        src61 <= 16'hb5fc;
        src62 <= 16'hf135;
        src63 <= 16'h87f0;
        exp <= 22'h21cada;
        #1
        src0 <= 16'hc93e;
        src1 <= 16'had2a;
        src2 <= 16'h962;
        src3 <= 16'hea15;
        src4 <= 16'hfd78;
        src5 <= 16'hb1c1;
        src6 <= 16'h1806;
        src7 <= 16'hed97;
        src8 <= 16'h63ce;
        src9 <= 16'he8a1;
        src10 <= 16'hff7;
        src11 <= 16'h84cd;
        src12 <= 16'h83d3;
        src13 <= 16'hb401;
        src14 <= 16'h1f6d;
        src15 <= 16'hb629;
        src16 <= 16'h6a91;
        src17 <= 16'hbf1a;
        src18 <= 16'he809;
        src19 <= 16'hd16a;
        src20 <= 16'ha2db;
        src21 <= 16'hfade;
        src22 <= 16'h7c8e;
        src23 <= 16'h2df;
        src24 <= 16'hf9cb;
        src25 <= 16'h9e90;
        src26 <= 16'hd13d;
        src27 <= 16'hc091;
        src28 <= 16'hcd60;
        src29 <= 16'h400f;
        src30 <= 16'hca74;
        src31 <= 16'h11fa;
        src32 <= 16'h7829;
        src33 <= 16'h1baa;
        src34 <= 16'h9ad0;
        src35 <= 16'h8936;
        src36 <= 16'h23bb;
        src37 <= 16'hc524;
        src38 <= 16'h6cbe;
        src39 <= 16'h3c41;
        src40 <= 16'h2a9d;
        src41 <= 16'h5774;
        src42 <= 16'h8efb;
        src43 <= 16'he3bf;
        src44 <= 16'ha8d9;
        src45 <= 16'h5426;
        src46 <= 16'h71f0;
        src47 <= 16'h800f;
        src48 <= 16'hc813;
        src49 <= 16'h890f;
        src50 <= 16'h117c;
        src51 <= 16'he7e2;
        src52 <= 16'h34e4;
        src53 <= 16'h1696;
        src54 <= 16'h410a;
        src55 <= 16'h96b9;
        src56 <= 16'hfa02;
        src57 <= 16'h96c3;
        src58 <= 16'h2796;
        src59 <= 16'hcd7c;
        src60 <= 16'hae59;
        src61 <= 16'hfb75;
        src62 <= 16'ha85f;
        src63 <= 16'h1f20;
        exp <= 22'h22b3fd;
        #1
        src0 <= 16'h6428;
        src1 <= 16'ha2e1;
        src2 <= 16'hadfe;
        src3 <= 16'hbfa1;
        src4 <= 16'h8ffc;
        src5 <= 16'hee17;
        src6 <= 16'h1246;
        src7 <= 16'ha0a0;
        src8 <= 16'hf4d6;
        src9 <= 16'h858b;
        src10 <= 16'h2b31;
        src11 <= 16'hecc9;
        src12 <= 16'h9b5c;
        src13 <= 16'h17b7;
        src14 <= 16'h10dc;
        src15 <= 16'h8b4c;
        src16 <= 16'h607a;
        src17 <= 16'h9e9c;
        src18 <= 16'hc517;
        src19 <= 16'h926c;
        src20 <= 16'h6d09;
        src21 <= 16'h95d2;
        src22 <= 16'h9daa;
        src23 <= 16'had97;
        src24 <= 16'hfd49;
        src25 <= 16'he172;
        src26 <= 16'heb9b;
        src27 <= 16'ha92a;
        src28 <= 16'h2a3;
        src29 <= 16'h281b;
        src30 <= 16'he526;
        src31 <= 16'h5724;
        src32 <= 16'h3972;
        src33 <= 16'hf324;
        src34 <= 16'hc210;
        src35 <= 16'h4f04;
        src36 <= 16'hd301;
        src37 <= 16'h7ef2;
        src38 <= 16'h691d;
        src39 <= 16'h44d0;
        src40 <= 16'h1637;
        src41 <= 16'hf025;
        src42 <= 16'hfbb1;
        src43 <= 16'h5819;
        src44 <= 16'hc8f8;
        src45 <= 16'hff20;
        src46 <= 16'h9793;
        src47 <= 16'h9234;
        src48 <= 16'hac3;
        src49 <= 16'hdb3c;
        src50 <= 16'h7adb;
        src51 <= 16'h9391;
        src52 <= 16'hfe24;
        src53 <= 16'h19dd;
        src54 <= 16'h951;
        src55 <= 16'h3a37;
        src56 <= 16'h2ec9;
        src57 <= 16'hc40d;
        src58 <= 16'h5e9f;
        src59 <= 16'h264c;
        src60 <= 16'h3e27;
        src61 <= 16'h16c1;
        src62 <= 16'ha615;
        src63 <= 16'h9e9c;
        exp <= 22'h21f151;
        #1
        src0 <= 16'h585f;
        src1 <= 16'hbc8a;
        src2 <= 16'h4da;
        src3 <= 16'ha93e;
        src4 <= 16'h3fe0;
        src5 <= 16'h6acf;
        src6 <= 16'haaca;
        src7 <= 16'hbbca;
        src8 <= 16'h49b5;
        src9 <= 16'hebb8;
        src10 <= 16'ha3d5;
        src11 <= 16'hfb03;
        src12 <= 16'hcee3;
        src13 <= 16'h68cf;
        src14 <= 16'hc64c;
        src15 <= 16'hfec1;
        src16 <= 16'h6543;
        src17 <= 16'he85b;
        src18 <= 16'h8053;
        src19 <= 16'h3e51;
        src20 <= 16'he320;
        src21 <= 16'h7275;
        src22 <= 16'h70a6;
        src23 <= 16'hc318;
        src24 <= 16'hc439;
        src25 <= 16'he12c;
        src26 <= 16'h9467;
        src27 <= 16'h9f7c;
        src28 <= 16'h5fd2;
        src29 <= 16'he291;
        src30 <= 16'hae58;
        src31 <= 16'hc236;
        src32 <= 16'h29c9;
        src33 <= 16'h1e9e;
        src34 <= 16'h4000;
        src35 <= 16'h8a0f;
        src36 <= 16'h7ae5;
        src37 <= 16'hac9;
        src38 <= 16'hceaf;
        src39 <= 16'h97a8;
        src40 <= 16'h5347;
        src41 <= 16'h37de;
        src42 <= 16'h4de;
        src43 <= 16'h329b;
        src44 <= 16'h2485;
        src45 <= 16'h73ae;
        src46 <= 16'h271b;
        src47 <= 16'hedb2;
        src48 <= 16'h9e91;
        src49 <= 16'hbaa3;
        src50 <= 16'h13df;
        src51 <= 16'h6302;
        src52 <= 16'hf34f;
        src53 <= 16'h9a38;
        src54 <= 16'h7953;
        src55 <= 16'hc242;
        src56 <= 16'hb3fb;
        src57 <= 16'h683;
        src58 <= 16'hf4c0;
        src59 <= 16'he037;
        src60 <= 16'hbb30;
        src61 <= 16'h8c46;
        src62 <= 16'h9146;
        src63 <= 16'h2927;
        exp <= 22'h225fb8;
        #1
        src0 <= 16'he763;
        src1 <= 16'h9aba;
        src2 <= 16'hc8c7;
        src3 <= 16'h6a4a;
        src4 <= 16'h65ce;
        src5 <= 16'h6e82;
        src6 <= 16'h802a;
        src7 <= 16'he9ff;
        src8 <= 16'h2ddb;
        src9 <= 16'h2731;
        src10 <= 16'hb0ba;
        src11 <= 16'h5c8d;
        src12 <= 16'h3e4e;
        src13 <= 16'hfd28;
        src14 <= 16'h2ae1;
        src15 <= 16'h95de;
        src16 <= 16'h83de;
        src17 <= 16'h2482;
        src18 <= 16'h7f0d;
        src19 <= 16'h9243;
        src20 <= 16'h12cb;
        src21 <= 16'h9b03;
        src22 <= 16'h4716;
        src23 <= 16'h51a9;
        src24 <= 16'h1ad5;
        src25 <= 16'hcc17;
        src26 <= 16'ha9f1;
        src27 <= 16'h1a79;
        src28 <= 16'h14ce;
        src29 <= 16'h53b7;
        src30 <= 16'hf51d;
        src31 <= 16'h9726;
        src32 <= 16'h65e5;
        src33 <= 16'h572a;
        src34 <= 16'hd412;
        src35 <= 16'h2cca;
        src36 <= 16'hda87;
        src37 <= 16'h3849;
        src38 <= 16'hc9fb;
        src39 <= 16'h5de3;
        src40 <= 16'he74e;
        src41 <= 16'h6b6d;
        src42 <= 16'hf181;
        src43 <= 16'h49ca;
        src44 <= 16'hf925;
        src45 <= 16'h4805;
        src46 <= 16'h47a3;
        src47 <= 16'h79e6;
        src48 <= 16'hfc7a;
        src49 <= 16'h5695;
        src50 <= 16'hd6e4;
        src51 <= 16'h211e;
        src52 <= 16'h4c12;
        src53 <= 16'hf694;
        src54 <= 16'hfbae;
        src55 <= 16'h14d4;
        src56 <= 16'h1cdd;
        src57 <= 16'hb6f7;
        src58 <= 16'h45ee;
        src59 <= 16'haba5;
        src60 <= 16'he2f0;
        src61 <= 16'hae65;
        src62 <= 16'hb6ed;
        src63 <= 16'hef14;
        exp <= 22'h2116d2;
        #1
        src0 <= 16'h305;
        src1 <= 16'hf9a;
        src2 <= 16'h8506;
        src3 <= 16'h3723;
        src4 <= 16'hd011;
        src5 <= 16'h4613;
        src6 <= 16'h972a;
        src7 <= 16'hf576;
        src8 <= 16'hbb61;
        src9 <= 16'haf70;
        src10 <= 16'heff9;
        src11 <= 16'he7ec;
        src12 <= 16'hae64;
        src13 <= 16'h4b0b;
        src14 <= 16'h13c1;
        src15 <= 16'h9d44;
        src16 <= 16'hbc3d;
        src17 <= 16'h544;
        src18 <= 16'h2b2;
        src19 <= 16'h44c9;
        src20 <= 16'hdf61;
        src21 <= 16'h7468;
        src22 <= 16'hdc2e;
        src23 <= 16'h4bd5;
        src24 <= 16'h926b;
        src25 <= 16'h9b37;
        src26 <= 16'hf8b8;
        src27 <= 16'hbc44;
        src28 <= 16'hc893;
        src29 <= 16'hac5c;
        src30 <= 16'ha187;
        src31 <= 16'hcb5;
        src32 <= 16'hdee4;
        src33 <= 16'hef9;
        src34 <= 16'hf737;
        src35 <= 16'h98de;
        src36 <= 16'h1631;
        src37 <= 16'hda7c;
        src38 <= 16'hdff6;
        src39 <= 16'h1312;
        src40 <= 16'h9883;
        src41 <= 16'h303b;
        src42 <= 16'ha155;
        src43 <= 16'hd02a;
        src44 <= 16'h43c9;
        src45 <= 16'h38f0;
        src46 <= 16'h3e9b;
        src47 <= 16'hff6;
        src48 <= 16'h6b6e;
        src49 <= 16'h5efd;
        src50 <= 16'ha5da;
        src51 <= 16'h59e1;
        src52 <= 16'hb93;
        src53 <= 16'h16c3;
        src54 <= 16'ha9eb;
        src55 <= 16'ha37e;
        src56 <= 16'hf295;
        src57 <= 16'h10fa;
        src58 <= 16'hab69;
        src59 <= 16'h83;
        src60 <= 16'hb4f7;
        src61 <= 16'h26c1;
        src62 <= 16'hd05f;
        src63 <= 16'h6d9c;
        exp <= 22'h1f5388;
        #1
        src0 <= 16'h43f0;
        src1 <= 16'h9029;
        src2 <= 16'h320c;
        src3 <= 16'he5d5;
        src4 <= 16'h20bd;
        src5 <= 16'h7199;
        src6 <= 16'hbaa7;
        src7 <= 16'h7ea3;
        src8 <= 16'hb42b;
        src9 <= 16'hbfe;
        src10 <= 16'h87cc;
        src11 <= 16'hda5;
        src12 <= 16'hf6da;
        src13 <= 16'h2591;
        src14 <= 16'hc257;
        src15 <= 16'hb52e;
        src16 <= 16'hd27e;
        src17 <= 16'hca5f;
        src18 <= 16'h9586;
        src19 <= 16'hada8;
        src20 <= 16'h5890;
        src21 <= 16'hcfed;
        src22 <= 16'ha20f;
        src23 <= 16'h13c2;
        src24 <= 16'h728d;
        src25 <= 16'h4f77;
        src26 <= 16'h48c;
        src27 <= 16'hf05b;
        src28 <= 16'hfedb;
        src29 <= 16'h6a28;
        src30 <= 16'hacfe;
        src31 <= 16'h940b;
        src32 <= 16'h8c7c;
        src33 <= 16'h55d9;
        src34 <= 16'he106;
        src35 <= 16'ha7c5;
        src36 <= 16'h1ee8;
        src37 <= 16'h173e;
        src38 <= 16'ha7d2;
        src39 <= 16'hfc00;
        src40 <= 16'h64f4;
        src41 <= 16'h5e08;
        src42 <= 16'h5373;
        src43 <= 16'h776c;
        src44 <= 16'h5f7d;
        src45 <= 16'h3707;
        src46 <= 16'h9a5b;
        src47 <= 16'h933;
        src48 <= 16'ha81f;
        src49 <= 16'hd9bd;
        src50 <= 16'h44d8;
        src51 <= 16'hb73;
        src52 <= 16'ha72f;
        src53 <= 16'h4236;
        src54 <= 16'hee4d;
        src55 <= 16'h85cc;
        src56 <= 16'h9a54;
        src57 <= 16'h95ba;
        src58 <= 16'h8cdc;
        src59 <= 16'hae29;
        src60 <= 16'ha9e3;
        src61 <= 16'h4685;
        src62 <= 16'hff67;
        src63 <= 16'h1b60;
        exp <= 22'h207360;
        #1
        src0 <= 16'h1f53;
        src1 <= 16'hb85b;
        src2 <= 16'h4f97;
        src3 <= 16'he9c2;
        src4 <= 16'hff8c;
        src5 <= 16'hb465;
        src6 <= 16'h6374;
        src7 <= 16'h5cff;
        src8 <= 16'hbd6e;
        src9 <= 16'h3ecb;
        src10 <= 16'h508e;
        src11 <= 16'hcfb3;
        src12 <= 16'h2398;
        src13 <= 16'h6bf8;
        src14 <= 16'h20a9;
        src15 <= 16'h5581;
        src16 <= 16'h534e;
        src17 <= 16'ha0d5;
        src18 <= 16'hb6ef;
        src19 <= 16'h6668;
        src20 <= 16'h712f;
        src21 <= 16'ha22;
        src22 <= 16'h149c;
        src23 <= 16'h47a;
        src24 <= 16'h6a00;
        src25 <= 16'ha03b;
        src26 <= 16'h5322;
        src27 <= 16'hfd8a;
        src28 <= 16'hd58;
        src29 <= 16'h7660;
        src30 <= 16'h4eab;
        src31 <= 16'hf627;
        src32 <= 16'he2ee;
        src33 <= 16'h6c55;
        src34 <= 16'hc821;
        src35 <= 16'h1cd1;
        src36 <= 16'he3e6;
        src37 <= 16'hc3f8;
        src38 <= 16'h2dbf;
        src39 <= 16'h1ee;
        src40 <= 16'ha2a5;
        src41 <= 16'h496f;
        src42 <= 16'hc2a6;
        src43 <= 16'h9d7e;
        src44 <= 16'hddd6;
        src45 <= 16'hbe32;
        src46 <= 16'hca04;
        src47 <= 16'hbb00;
        src48 <= 16'h7a2d;
        src49 <= 16'h9c11;
        src50 <= 16'h278d;
        src51 <= 16'h45d6;
        src52 <= 16'h8cc5;
        src53 <= 16'h7880;
        src54 <= 16'hf19b;
        src55 <= 16'h7c19;
        src56 <= 16'h1b49;
        src57 <= 16'h1e7a;
        src58 <= 16'h81ce;
        src59 <= 16'hf3e4;
        src60 <= 16'hae46;
        src61 <= 16'hffd1;
        src62 <= 16'h447e;
        src63 <= 16'h80c6;
        exp <= 22'h20035f;
        #1
        src0 <= 16'h515d;
        src1 <= 16'hfec;
        src2 <= 16'h85a;
        src3 <= 16'hadba;
        src4 <= 16'hd16c;
        src5 <= 16'h9d25;
        src6 <= 16'h5522;
        src7 <= 16'hb508;
        src8 <= 16'h6973;
        src9 <= 16'hacfb;
        src10 <= 16'hfe08;
        src11 <= 16'h189b;
        src12 <= 16'h8ac;
        src13 <= 16'h9763;
        src14 <= 16'h5790;
        src15 <= 16'h1f9a;
        src16 <= 16'hfb21;
        src17 <= 16'h3c45;
        src18 <= 16'h35ff;
        src19 <= 16'hd642;
        src20 <= 16'hfab0;
        src21 <= 16'h3ca3;
        src22 <= 16'hb6e6;
        src23 <= 16'hf155;
        src24 <= 16'h9456;
        src25 <= 16'he0c8;
        src26 <= 16'hd8cb;
        src27 <= 16'h1c34;
        src28 <= 16'hfae5;
        src29 <= 16'haa8;
        src30 <= 16'h1e93;
        src31 <= 16'h4e63;
        src32 <= 16'h33be;
        src33 <= 16'hfe7d;
        src34 <= 16'hd48e;
        src35 <= 16'h8b7c;
        src36 <= 16'h3579;
        src37 <= 16'h4448;
        src38 <= 16'h49bd;
        src39 <= 16'hc01a;
        src40 <= 16'hd6b;
        src41 <= 16'h63f1;
        src42 <= 16'h3d8a;
        src43 <= 16'hf15d;
        src44 <= 16'h116;
        src45 <= 16'h5614;
        src46 <= 16'h163f;
        src47 <= 16'h1e47;
        src48 <= 16'hcc0e;
        src49 <= 16'h44ad;
        src50 <= 16'h6d5d;
        src51 <= 16'h33b6;
        src52 <= 16'h608e;
        src53 <= 16'ha4b;
        src54 <= 16'h8783;
        src55 <= 16'h9123;
        src56 <= 16'hade3;
        src57 <= 16'hdc3c;
        src58 <= 16'h4a0a;
        src59 <= 16'haa;
        src60 <= 16'h6394;
        src61 <= 16'hfef5;
        src62 <= 16'h20cd;
        src63 <= 16'h3167;
        exp <= 22'h1cd4e4;
        #1
        src0 <= 16'h28c9;
        src1 <= 16'h3f99;
        src2 <= 16'hcb83;
        src3 <= 16'h1b9f;
        src4 <= 16'hd117;
        src5 <= 16'h3ba3;
        src6 <= 16'h59b6;
        src7 <= 16'h2ead;
        src8 <= 16'hab3f;
        src9 <= 16'h8e9e;
        src10 <= 16'h5cd9;
        src11 <= 16'hd7ca;
        src12 <= 16'h1a0a;
        src13 <= 16'hd8eb;
        src14 <= 16'hf748;
        src15 <= 16'ha6a6;
        src16 <= 16'hb7ba;
        src17 <= 16'h9d26;
        src18 <= 16'hcc75;
        src19 <= 16'h787c;
        src20 <= 16'h4864;
        src21 <= 16'h9562;
        src22 <= 16'h25cd;
        src23 <= 16'hfec5;
        src24 <= 16'h4412;
        src25 <= 16'h9660;
        src26 <= 16'h871e;
        src27 <= 16'h2703;
        src28 <= 16'hd33f;
        src29 <= 16'h2021;
        src30 <= 16'h4d53;
        src31 <= 16'h1924;
        src32 <= 16'h2caa;
        src33 <= 16'hf05d;
        src34 <= 16'h37b7;
        src35 <= 16'h3e22;
        src36 <= 16'habc3;
        src37 <= 16'h8134;
        src38 <= 16'h83b;
        src39 <= 16'h11ae;
        src40 <= 16'h3761;
        src41 <= 16'h92df;
        src42 <= 16'he31d;
        src43 <= 16'hbdbd;
        src44 <= 16'h8f65;
        src45 <= 16'ha3bb;
        src46 <= 16'hae13;
        src47 <= 16'hf2e5;
        src48 <= 16'hb294;
        src49 <= 16'heda6;
        src50 <= 16'h1584;
        src51 <= 16'h58b9;
        src52 <= 16'hdde5;
        src53 <= 16'he6d4;
        src54 <= 16'hc8ae;
        src55 <= 16'h435c;
        src56 <= 16'h2e4c;
        src57 <= 16'h3f98;
        src58 <= 16'hda6e;
        src59 <= 16'heedf;
        src60 <= 16'h8e9c;
        src61 <= 16'hae10;
        src62 <= 16'he069;
        src63 <= 16'hcb70;
        exp <= 22'h217a79;
        #1
        src0 <= 16'h84d0;
        src1 <= 16'h3388;
        src2 <= 16'h334e;
        src3 <= 16'h6f16;
        src4 <= 16'hec2f;
        src5 <= 16'h30a8;
        src6 <= 16'h9331;
        src7 <= 16'hb769;
        src8 <= 16'had3;
        src9 <= 16'h9d1d;
        src10 <= 16'h93c7;
        src11 <= 16'h6c8d;
        src12 <= 16'hb3e9;
        src13 <= 16'h59f0;
        src14 <= 16'hcc07;
        src15 <= 16'h98fd;
        src16 <= 16'ha7db;
        src17 <= 16'h58f6;
        src18 <= 16'hdf94;
        src19 <= 16'h1140;
        src20 <= 16'h87e0;
        src21 <= 16'h91f8;
        src22 <= 16'ha054;
        src23 <= 16'h841c;
        src24 <= 16'hcc95;
        src25 <= 16'h73d9;
        src26 <= 16'ha003;
        src27 <= 16'h3726;
        src28 <= 16'hefe5;
        src29 <= 16'h205e;
        src30 <= 16'hdca8;
        src31 <= 16'hed51;
        src32 <= 16'h22d3;
        src33 <= 16'h3c06;
        src34 <= 16'h1b9b;
        src35 <= 16'h2ae;
        src36 <= 16'h7f84;
        src37 <= 16'hef30;
        src38 <= 16'h2356;
        src39 <= 16'hab8e;
        src40 <= 16'hb821;
        src41 <= 16'h4b8c;
        src42 <= 16'h6f0;
        src43 <= 16'h8a17;
        src44 <= 16'hd2d2;
        src45 <= 16'h6a0d;
        src46 <= 16'h69fe;
        src47 <= 16'hbd3;
        src48 <= 16'h26bb;
        src49 <= 16'h44ea;
        src50 <= 16'h7f79;
        src51 <= 16'ha568;
        src52 <= 16'h9dbd;
        src53 <= 16'h403;
        src54 <= 16'h3f87;
        src55 <= 16'h479e;
        src56 <= 16'h74d2;
        src57 <= 16'h459;
        src58 <= 16'hd73b;
        src59 <= 16'hb33;
        src60 <= 16'hd3dc;
        src61 <= 16'h16ad;
        src62 <= 16'hddd0;
        src63 <= 16'h476a;
        exp <= 22'h1d25f3;
        #1
        src0 <= 16'haf28;
        src1 <= 16'h2d11;
        src2 <= 16'h97df;
        src3 <= 16'h41a6;
        src4 <= 16'hf456;
        src5 <= 16'h3b50;
        src6 <= 16'h3b95;
        src7 <= 16'hbf07;
        src8 <= 16'h2bac;
        src9 <= 16'ha662;
        src10 <= 16'ha696;
        src11 <= 16'h9f9f;
        src12 <= 16'h2501;
        src13 <= 16'h3542;
        src14 <= 16'h5435;
        src15 <= 16'hc96f;
        src16 <= 16'h696f;
        src17 <= 16'h2274;
        src18 <= 16'h3e33;
        src19 <= 16'h94c6;
        src20 <= 16'hffc6;
        src21 <= 16'hc72a;
        src22 <= 16'h40f;
        src23 <= 16'h72ad;
        src24 <= 16'hd74f;
        src25 <= 16'ha611;
        src26 <= 16'hb775;
        src27 <= 16'h1321;
        src28 <= 16'h8856;
        src29 <= 16'hacef;
        src30 <= 16'had2d;
        src31 <= 16'hbc80;
        src32 <= 16'h8341;
        src33 <= 16'hf3ac;
        src34 <= 16'h5037;
        src35 <= 16'he526;
        src36 <= 16'h4fa9;
        src37 <= 16'h4c;
        src38 <= 16'h5ad;
        src39 <= 16'hb623;
        src40 <= 16'h6a54;
        src41 <= 16'hf17e;
        src42 <= 16'hfd49;
        src43 <= 16'h417d;
        src44 <= 16'h4b84;
        src45 <= 16'he067;
        src46 <= 16'hbaac;
        src47 <= 16'h885d;
        src48 <= 16'heb0d;
        src49 <= 16'h5ace;
        src50 <= 16'he5ac;
        src51 <= 16'hd812;
        src52 <= 16'ha034;
        src53 <= 16'hd192;
        src54 <= 16'hdb1;
        src55 <= 16'h4de5;
        src56 <= 16'h6060;
        src57 <= 16'hde29;
        src58 <= 16'h8d87;
        src59 <= 16'h36bc;
        src60 <= 16'h1cf6;
        src61 <= 16'h2f55;
        src62 <= 16'h838c;
        src63 <= 16'hb606;
        exp <= 22'h210ed3;
        #1
        src0 <= 16'hae47;
        src1 <= 16'h956f;
        src2 <= 16'hd1fe;
        src3 <= 16'hd35d;
        src4 <= 16'hdd49;
        src5 <= 16'h8879;
        src6 <= 16'hd9d9;
        src7 <= 16'h30e8;
        src8 <= 16'hd367;
        src9 <= 16'h8cc6;
        src10 <= 16'hc64d;
        src11 <= 16'haa65;
        src12 <= 16'hfe0b;
        src13 <= 16'h3952;
        src14 <= 16'ha346;
        src15 <= 16'h4937;
        src16 <= 16'h54b7;
        src17 <= 16'h44c0;
        src18 <= 16'ha130;
        src19 <= 16'h6791;
        src20 <= 16'hea25;
        src21 <= 16'h9561;
        src22 <= 16'h3212;
        src23 <= 16'hd6cb;
        src24 <= 16'he2e8;
        src25 <= 16'haae0;
        src26 <= 16'hca28;
        src27 <= 16'hb206;
        src28 <= 16'h28c4;
        src29 <= 16'h5201;
        src30 <= 16'he420;
        src31 <= 16'hd0ee;
        src32 <= 16'hcdcd;
        src33 <= 16'h8595;
        src34 <= 16'h4f60;
        src35 <= 16'h9ed6;
        src36 <= 16'h4302;
        src37 <= 16'h2b5e;
        src38 <= 16'h63f1;
        src39 <= 16'hc079;
        src40 <= 16'h7d51;
        src41 <= 16'h1ff7;
        src42 <= 16'h43ad;
        src43 <= 16'h252b;
        src44 <= 16'h2689;
        src45 <= 16'hdde5;
        src46 <= 16'h66e1;
        src47 <= 16'h3c85;
        src48 <= 16'hbffc;
        src49 <= 16'h84c7;
        src50 <= 16'h9e2b;
        src51 <= 16'ha8cb;
        src52 <= 16'he9f2;
        src53 <= 16'h1b30;
        src54 <= 16'h2dd5;
        src55 <= 16'h48c7;
        src56 <= 16'hcc9c;
        src57 <= 16'h621b;
        src58 <= 16'h8c96;
        src59 <= 16'hd88f;
        src60 <= 16'hedcd;
        src61 <= 16'h98fb;
        src62 <= 16'h3868;
        src63 <= 16'h5815;
        exp <= 22'h22e79f;
        #1
        src0 <= 16'hbffe;
        src1 <= 16'he8e5;
        src2 <= 16'hfdea;
        src3 <= 16'h3bd0;
        src4 <= 16'hef06;
        src5 <= 16'hcb3f;
        src6 <= 16'h304a;
        src7 <= 16'h7a86;
        src8 <= 16'h54f5;
        src9 <= 16'h5b64;
        src10 <= 16'hc74d;
        src11 <= 16'h6a1;
        src12 <= 16'h257;
        src13 <= 16'he062;
        src14 <= 16'h56e2;
        src15 <= 16'hbc18;
        src16 <= 16'h34ee;
        src17 <= 16'hdc0e;
        src18 <= 16'hb971;
        src19 <= 16'h65e8;
        src20 <= 16'haf9d;
        src21 <= 16'h1b08;
        src22 <= 16'hc4ee;
        src23 <= 16'h1af1;
        src24 <= 16'h7582;
        src25 <= 16'hd2f7;
        src26 <= 16'h6999;
        src27 <= 16'hb068;
        src28 <= 16'hb50;
        src29 <= 16'h3660;
        src30 <= 16'h46db;
        src31 <= 16'h2e0f;
        src32 <= 16'h751c;
        src33 <= 16'h997e;
        src34 <= 16'h2278;
        src35 <= 16'h45eb;
        src36 <= 16'hf9b4;
        src37 <= 16'ha308;
        src38 <= 16'h4a8d;
        src39 <= 16'h3066;
        src40 <= 16'hdea7;
        src41 <= 16'h1459;
        src42 <= 16'h2520;
        src43 <= 16'h5dd0;
        src44 <= 16'hf252;
        src45 <= 16'h5b0a;
        src46 <= 16'hc8db;
        src47 <= 16'h5ceb;
        src48 <= 16'hdeff;
        src49 <= 16'ha1b6;
        src50 <= 16'hc0ad;
        src51 <= 16'hd93a;
        src52 <= 16'hfaf4;
        src53 <= 16'hf4ba;
        src54 <= 16'hf319;
        src55 <= 16'hf47f;
        src56 <= 16'hd1c5;
        src57 <= 16'hcf1;
        src58 <= 16'hff86;
        src59 <= 16'h939;
        src60 <= 16'h7dc8;
        src61 <= 16'h2b77;
        src62 <= 16'he376;
        src63 <= 16'hbbbf;
        exp <= 22'h224922;
        #1
        src0 <= 16'h1ff4;
        src1 <= 16'h6631;
        src2 <= 16'h61e;
        src3 <= 16'hd59f;
        src4 <= 16'h8f7d;
        src5 <= 16'h2da3;
        src6 <= 16'h4cae;
        src7 <= 16'ha69e;
        src8 <= 16'hb610;
        src9 <= 16'hee1b;
        src10 <= 16'h3925;
        src11 <= 16'hb4f3;
        src12 <= 16'ha066;
        src13 <= 16'hc6de;
        src14 <= 16'hed4;
        src15 <= 16'h65cf;
        src16 <= 16'h7095;
        src17 <= 16'h3d91;
        src18 <= 16'hadd2;
        src19 <= 16'hc4d4;
        src20 <= 16'h7105;
        src21 <= 16'hf584;
        src22 <= 16'ha573;
        src23 <= 16'h6b00;
        src24 <= 16'h9fc3;
        src25 <= 16'h7fdb;
        src26 <= 16'h93f7;
        src27 <= 16'hedb;
        src28 <= 16'hc8d5;
        src29 <= 16'h7104;
        src30 <= 16'ha292;
        src31 <= 16'h67c6;
        src32 <= 16'h9b9d;
        src33 <= 16'hd234;
        src34 <= 16'hc7e1;
        src35 <= 16'h6bc0;
        src36 <= 16'h850f;
        src37 <= 16'h9ec6;
        src38 <= 16'hee44;
        src39 <= 16'h4616;
        src40 <= 16'h1d96;
        src41 <= 16'hf1be;
        src42 <= 16'h4063;
        src43 <= 16'h3770;
        src44 <= 16'h1249;
        src45 <= 16'hc5ff;
        src46 <= 16'hff5;
        src47 <= 16'h2a59;
        src48 <= 16'ha3f1;
        src49 <= 16'h4825;
        src50 <= 16'hd2d2;
        src51 <= 16'h380f;
        src52 <= 16'ha29d;
        src53 <= 16'hc140;
        src54 <= 16'h39d6;
        src55 <= 16'hc85d;
        src56 <= 16'hcc52;
        src57 <= 16'h2276;
        src58 <= 16'h18b7;
        src59 <= 16'h302;
        src60 <= 16'h6164;
        src61 <= 16'h5f8e;
        src62 <= 16'he07d;
        src63 <= 16'h86e0;
        exp <= 22'h1f4216;
        #1
        src0 <= 16'h27a4;
        src1 <= 16'h7f37;
        src2 <= 16'he85a;
        src3 <= 16'h54ae;
        src4 <= 16'h51b9;
        src5 <= 16'hebd6;
        src6 <= 16'h1d0f;
        src7 <= 16'h2897;
        src8 <= 16'he927;
        src9 <= 16'h5674;
        src10 <= 16'hc118;
        src11 <= 16'h52e5;
        src12 <= 16'h7b78;
        src13 <= 16'h43a1;
        src14 <= 16'h76d7;
        src15 <= 16'h7a1d;
        src16 <= 16'h13cc;
        src17 <= 16'h34cd;
        src18 <= 16'hbbd3;
        src19 <= 16'h598c;
        src20 <= 16'he439;
        src21 <= 16'hf589;
        src22 <= 16'hfc04;
        src23 <= 16'h975c;
        src24 <= 16'hcbbd;
        src25 <= 16'hc260;
        src26 <= 16'h9021;
        src27 <= 16'hf0b8;
        src28 <= 16'he194;
        src29 <= 16'haf98;
        src30 <= 16'h2f72;
        src31 <= 16'h406f;
        src32 <= 16'hd494;
        src33 <= 16'hbf03;
        src34 <= 16'h70f5;
        src35 <= 16'hb8b6;
        src36 <= 16'h1bbc;
        src37 <= 16'h1583;
        src38 <= 16'hb8ae;
        src39 <= 16'h241c;
        src40 <= 16'hf406;
        src41 <= 16'ha959;
        src42 <= 16'h9b8e;
        src43 <= 16'h30ea;
        src44 <= 16'hef47;
        src45 <= 16'h9ca5;
        src46 <= 16'h5a25;
        src47 <= 16'h79f8;
        src48 <= 16'he214;
        src49 <= 16'ha76c;
        src50 <= 16'hd435;
        src51 <= 16'hd02;
        src52 <= 16'h75;
        src53 <= 16'hd572;
        src54 <= 16'h8f86;
        src55 <= 16'h611f;
        src56 <= 16'h721d;
        src57 <= 16'h34f5;
        src58 <= 16'h23b2;
        src59 <= 16'hda2c;
        src60 <= 16'hf73c;
        src61 <= 16'h7498;
        src62 <= 16'h1076;
        src63 <= 16'h63f6;
        exp <= 22'h219178;
        #1
        src0 <= 16'hcf9f;
        src1 <= 16'hebc8;
        src2 <= 16'h5011;
        src3 <= 16'h5fde;
        src4 <= 16'hbbb1;
        src5 <= 16'h2959;
        src6 <= 16'h3db5;
        src7 <= 16'h63eb;
        src8 <= 16'hbf32;
        src9 <= 16'h9566;
        src10 <= 16'h331d;
        src11 <= 16'h367c;
        src12 <= 16'h57e4;
        src13 <= 16'h28fa;
        src14 <= 16'h7ae0;
        src15 <= 16'hec87;
        src16 <= 16'h3508;
        src17 <= 16'h5dfa;
        src18 <= 16'h833d;
        src19 <= 16'hff10;
        src20 <= 16'h58f1;
        src21 <= 16'hce54;
        src22 <= 16'hed;
        src23 <= 16'hdf43;
        src24 <= 16'hd01a;
        src25 <= 16'hcb61;
        src26 <= 16'hcc6d;
        src27 <= 16'h3e1b;
        src28 <= 16'h2821;
        src29 <= 16'h3d4;
        src30 <= 16'h406;
        src31 <= 16'h7c8d;
        src32 <= 16'h20e8;
        src33 <= 16'hce82;
        src34 <= 16'ha4cb;
        src35 <= 16'h8e21;
        src36 <= 16'he5e0;
        src37 <= 16'h97a8;
        src38 <= 16'h8ff9;
        src39 <= 16'he50f;
        src40 <= 16'hce2;
        src41 <= 16'h1118;
        src42 <= 16'h8975;
        src43 <= 16'h963c;
        src44 <= 16'h851a;
        src45 <= 16'hd41b;
        src46 <= 16'hdc06;
        src47 <= 16'he0cf;
        src48 <= 16'hfcd0;
        src49 <= 16'h6d7f;
        src50 <= 16'h7a74;
        src51 <= 16'h6a71;
        src52 <= 16'hf37a;
        src53 <= 16'h13d0;
        src54 <= 16'h5de3;
        src55 <= 16'hc962;
        src56 <= 16'hfccc;
        src57 <= 16'hd1e0;
        src58 <= 16'h4fbc;
        src59 <= 16'h633e;
        src60 <= 16'ha504;
        src61 <= 16'haf5f;
        src62 <= 16'h358;
        src63 <= 16'ha670;
        exp <= 22'h216df4;
        #1
        src0 <= 16'hd76b;
        src1 <= 16'haf40;
        src2 <= 16'h1b51;
        src3 <= 16'h14b7;
        src4 <= 16'h2ee2;
        src5 <= 16'hef37;
        src6 <= 16'h23a6;
        src7 <= 16'h495f;
        src8 <= 16'heb2b;
        src9 <= 16'h88c2;
        src10 <= 16'hf2e3;
        src11 <= 16'hbb2e;
        src12 <= 16'hb8fe;
        src13 <= 16'he9c0;
        src14 <= 16'h3e5f;
        src15 <= 16'h4358;
        src16 <= 16'hf72c;
        src17 <= 16'hd96b;
        src18 <= 16'h9ab0;
        src19 <= 16'h2e8f;
        src20 <= 16'h6b15;
        src21 <= 16'hf247;
        src22 <= 16'ha9ea;
        src23 <= 16'hf44e;
        src24 <= 16'h23aa;
        src25 <= 16'he43e;
        src26 <= 16'hcf55;
        src27 <= 16'h3ca8;
        src28 <= 16'h78d7;
        src29 <= 16'h50a1;
        src30 <= 16'h97de;
        src31 <= 16'h4e35;
        src32 <= 16'hfad0;
        src33 <= 16'h1f99;
        src34 <= 16'hc53;
        src35 <= 16'h79ec;
        src36 <= 16'h7286;
        src37 <= 16'h4a52;
        src38 <= 16'hf6af;
        src39 <= 16'h45b2;
        src40 <= 16'h7f5d;
        src41 <= 16'hf3ea;
        src42 <= 16'h2ee0;
        src43 <= 16'hf848;
        src44 <= 16'h4e21;
        src45 <= 16'hb044;
        src46 <= 16'hcccf;
        src47 <= 16'h4b92;
        src48 <= 16'he674;
        src49 <= 16'heaf1;
        src50 <= 16'hf9c4;
        src51 <= 16'h3019;
        src52 <= 16'h660a;
        src53 <= 16'h9b11;
        src54 <= 16'hbd57;
        src55 <= 16'hf40d;
        src56 <= 16'h6ba5;
        src57 <= 16'haa7f;
        src58 <= 16'h9778;
        src59 <= 16'ha9d2;
        src60 <= 16'hff1c;
        src61 <= 16'h5dab;
        src62 <= 16'h3792;
        src63 <= 16'hbbaa;
        exp <= 22'h248166;
        #1
        src0 <= 16'hf00f;
        src1 <= 16'h6f;
        src2 <= 16'h9cf6;
        src3 <= 16'h5652;
        src4 <= 16'h8819;
        src5 <= 16'h3fbe;
        src6 <= 16'h1892;
        src7 <= 16'he16c;
        src8 <= 16'h2626;
        src9 <= 16'h2b3;
        src10 <= 16'h70be;
        src11 <= 16'h4f8;
        src12 <= 16'h9194;
        src13 <= 16'hf546;
        src14 <= 16'hafd7;
        src15 <= 16'h9dff;
        src16 <= 16'h4c3e;
        src17 <= 16'he363;
        src18 <= 16'hee5a;
        src19 <= 16'he2e1;
        src20 <= 16'hca8d;
        src21 <= 16'hcfc4;
        src22 <= 16'h6f74;
        src23 <= 16'h7977;
        src24 <= 16'h1bdd;
        src25 <= 16'hffe7;
        src26 <= 16'hd041;
        src27 <= 16'h3460;
        src28 <= 16'h66d4;
        src29 <= 16'he373;
        src30 <= 16'hedba;
        src31 <= 16'hc1a;
        src32 <= 16'h331e;
        src33 <= 16'h2499;
        src34 <= 16'h1756;
        src35 <= 16'h5047;
        src36 <= 16'h95d5;
        src37 <= 16'h39b7;
        src38 <= 16'hda85;
        src39 <= 16'had20;
        src40 <= 16'h6941;
        src41 <= 16'h4766;
        src42 <= 16'h455e;
        src43 <= 16'hcc01;
        src44 <= 16'h863f;
        src45 <= 16'h59c7;
        src46 <= 16'h582d;
        src47 <= 16'h20d7;
        src48 <= 16'hea6f;
        src49 <= 16'hca9c;
        src50 <= 16'he129;
        src51 <= 16'h51c4;
        src52 <= 16'hda2b;
        src53 <= 16'h12eb;
        src54 <= 16'he950;
        src55 <= 16'h6848;
        src56 <= 16'h4a56;
        src57 <= 16'hf1c2;
        src58 <= 16'ha46a;
        src59 <= 16'hacbf;
        src60 <= 16'heef1;
        src61 <= 16'h687b;
        src62 <= 16'h6b3e;
        src63 <= 16'hd5c2;
        exp <= 22'h217f5a;
        #1
        src0 <= 16'h4489;
        src1 <= 16'h4092;
        src2 <= 16'h6b3;
        src3 <= 16'h3bfa;
        src4 <= 16'hce75;
        src5 <= 16'hb3b8;
        src6 <= 16'h3bc0;
        src7 <= 16'h35af;
        src8 <= 16'hb77d;
        src9 <= 16'h2df5;
        src10 <= 16'hb8b9;
        src11 <= 16'h1ba8;
        src12 <= 16'h7c7;
        src13 <= 16'h5532;
        src14 <= 16'h8be3;
        src15 <= 16'hca9d;
        src16 <= 16'hb0ae;
        src17 <= 16'hceed;
        src18 <= 16'h2396;
        src19 <= 16'h27f9;
        src20 <= 16'he71b;
        src21 <= 16'hc144;
        src22 <= 16'h35c2;
        src23 <= 16'h62eb;
        src24 <= 16'h63e3;
        src25 <= 16'h42aa;
        src26 <= 16'h6f04;
        src27 <= 16'ha1df;
        src28 <= 16'h7684;
        src29 <= 16'h7629;
        src30 <= 16'h516c;
        src31 <= 16'h5749;
        src32 <= 16'hec;
        src33 <= 16'hac2e;
        src34 <= 16'h25c7;
        src35 <= 16'hd08b;
        src36 <= 16'hfa33;
        src37 <= 16'h7e4c;
        src38 <= 16'h53fd;
        src39 <= 16'hb8dd;
        src40 <= 16'hed76;
        src41 <= 16'h685f;
        src42 <= 16'h9834;
        src43 <= 16'hfef9;
        src44 <= 16'hbc42;
        src45 <= 16'hd8ab;
        src46 <= 16'hd81f;
        src47 <= 16'hebc0;
        src48 <= 16'hea57;
        src49 <= 16'h89c6;
        src50 <= 16'h2cf3;
        src51 <= 16'hff62;
        src52 <= 16'h6193;
        src53 <= 16'hd8e3;
        src54 <= 16'h6f58;
        src55 <= 16'he989;
        src56 <= 16'h667b;
        src57 <= 16'h3638;
        src58 <= 16'h763c;
        src59 <= 16'hd555;
        src60 <= 16'hce3f;
        src61 <= 16'hfbdb;
        src62 <= 16'h55ce;
        src63 <= 16'h6367;
        exp <= 22'h218fa7;
        #1
        src0 <= 16'hc471;
        src1 <= 16'h4b4a;
        src2 <= 16'hf646;
        src3 <= 16'h95bb;
        src4 <= 16'ha4c7;
        src5 <= 16'h1ff4;
        src6 <= 16'h589e;
        src7 <= 16'h9038;
        src8 <= 16'h9350;
        src9 <= 16'h854d;
        src10 <= 16'hda8b;
        src11 <= 16'haf3f;
        src12 <= 16'h38f8;
        src13 <= 16'hc4b1;
        src14 <= 16'h856a;
        src15 <= 16'h359e;
        src16 <= 16'he838;
        src17 <= 16'h23cd;
        src18 <= 16'hbdd;
        src19 <= 16'h45e6;
        src20 <= 16'he361;
        src21 <= 16'h90c5;
        src22 <= 16'hd96e;
        src23 <= 16'hce9d;
        src24 <= 16'hd547;
        src25 <= 16'h2e2;
        src26 <= 16'h5976;
        src27 <= 16'hfa76;
        src28 <= 16'h204c;
        src29 <= 16'ha879;
        src30 <= 16'h3c12;
        src31 <= 16'hb8;
        src32 <= 16'hfb69;
        src33 <= 16'hc1e6;
        src34 <= 16'hb967;
        src35 <= 16'hafbe;
        src36 <= 16'h71e7;
        src37 <= 16'ha700;
        src38 <= 16'hb161;
        src39 <= 16'he6a6;
        src40 <= 16'hfa93;
        src41 <= 16'hb7b7;
        src42 <= 16'hf442;
        src43 <= 16'hc78f;
        src44 <= 16'hd61c;
        src45 <= 16'hffa2;
        src46 <= 16'h3e47;
        src47 <= 16'h7382;
        src48 <= 16'h66f7;
        src49 <= 16'h1cc6;
        src50 <= 16'h746d;
        src51 <= 16'hae17;
        src52 <= 16'hb201;
        src53 <= 16'ha50;
        src54 <= 16'h6dd;
        src55 <= 16'h71ba;
        src56 <= 16'hf67;
        src57 <= 16'he3e4;
        src58 <= 16'hfd94;
        src59 <= 16'h33ef;
        src60 <= 16'hb72b;
        src61 <= 16'h66f4;
        src62 <= 16'hc2c8;
        src63 <= 16'h87ae;
        exp <= 22'h238592;
        #1
        src0 <= 16'h6435;
        src1 <= 16'hbc6a;
        src2 <= 16'h40b2;
        src3 <= 16'h6959;
        src4 <= 16'h3ff1;
        src5 <= 16'h2b05;
        src6 <= 16'ha06b;
        src7 <= 16'hbaaf;
        src8 <= 16'h1d53;
        src9 <= 16'h772d;
        src10 <= 16'h7c90;
        src11 <= 16'hb3f;
        src12 <= 16'h55e5;
        src13 <= 16'h3c30;
        src14 <= 16'h9f96;
        src15 <= 16'hcc1d;
        src16 <= 16'h529c;
        src17 <= 16'hc2d9;
        src18 <= 16'h63f0;
        src19 <= 16'h304a;
        src20 <= 16'h214e;
        src21 <= 16'h8d6c;
        src22 <= 16'h976;
        src23 <= 16'hfd36;
        src24 <= 16'h8825;
        src25 <= 16'hbb68;
        src26 <= 16'h169f;
        src27 <= 16'h61fe;
        src28 <= 16'he9b6;
        src29 <= 16'h753;
        src30 <= 16'h8e1;
        src31 <= 16'hb17d;
        src32 <= 16'hf880;
        src33 <= 16'ha244;
        src34 <= 16'h4e3f;
        src35 <= 16'h613f;
        src36 <= 16'h4931;
        src37 <= 16'hbf9;
        src38 <= 16'h1500;
        src39 <= 16'h17e2;
        src40 <= 16'h6b7a;
        src41 <= 16'h4bb2;
        src42 <= 16'h89ab;
        src43 <= 16'h56e7;
        src44 <= 16'h40f3;
        src45 <= 16'h9173;
        src46 <= 16'h60;
        src47 <= 16'hbceb;
        src48 <= 16'h3b35;
        src49 <= 16'hec83;
        src50 <= 16'h1ff;
        src51 <= 16'h2ef4;
        src52 <= 16'h34fa;
        src53 <= 16'hdcb9;
        src54 <= 16'had15;
        src55 <= 16'h170f;
        src56 <= 16'h1964;
        src57 <= 16'hee64;
        src58 <= 16'h64be;
        src59 <= 16'hdfff;
        src60 <= 16'h4bc9;
        src61 <= 16'h59b5;
        src62 <= 16'h211f;
        src63 <= 16'hb08;
        exp <= 22'h19b1e0;
        #1
        src0 <= 16'h1eda;
        src1 <= 16'h1520;
        src2 <= 16'h62e5;
        src3 <= 16'h609a;
        src4 <= 16'h20ee;
        src5 <= 16'h9f1;
        src6 <= 16'h1548;
        src7 <= 16'h712a;
        src8 <= 16'h7bf;
        src9 <= 16'h2c35;
        src10 <= 16'hc2d;
        src11 <= 16'h253e;
        src12 <= 16'h1fd0;
        src13 <= 16'h284c;
        src14 <= 16'h23ca;
        src15 <= 16'h817b;
        src16 <= 16'h5b72;
        src17 <= 16'h9227;
        src18 <= 16'hb1bf;
        src19 <= 16'ha544;
        src20 <= 16'h2213;
        src21 <= 16'he700;
        src22 <= 16'h444;
        src23 <= 16'h1fad;
        src24 <= 16'he241;
        src25 <= 16'hdd0a;
        src26 <= 16'h4008;
        src27 <= 16'hd621;
        src28 <= 16'h685c;
        src29 <= 16'h4e1e;
        src30 <= 16'h9929;
        src31 <= 16'h1401;
        src32 <= 16'h6be6;
        src33 <= 16'hd3cd;
        src34 <= 16'h84e9;
        src35 <= 16'h6e4a;
        src36 <= 16'h5890;
        src37 <= 16'hdb01;
        src38 <= 16'h38b9;
        src39 <= 16'hc406;
        src40 <= 16'hba1;
        src41 <= 16'h4bb8;
        src42 <= 16'h15ee;
        src43 <= 16'h9977;
        src44 <= 16'h5ad1;
        src45 <= 16'h877f;
        src46 <= 16'hb6c9;
        src47 <= 16'h9652;
        src48 <= 16'h5103;
        src49 <= 16'ha155;
        src50 <= 16'heefc;
        src51 <= 16'hba50;
        src52 <= 16'h9629;
        src53 <= 16'hfd3d;
        src54 <= 16'h530c;
        src55 <= 16'ha4d6;
        src56 <= 16'h8176;
        src57 <= 16'h3060;
        src58 <= 16'ha8b3;
        src59 <= 16'h292a;
        src60 <= 16'heb3d;
        src61 <= 16'h8027;
        src62 <= 16'hf03b;
        src63 <= 16'ha2b3;
        exp <= 22'h1be892;
        #1
        src0 <= 16'hec35;
        src1 <= 16'h8bf9;
        src2 <= 16'h37d;
        src3 <= 16'hd1fe;
        src4 <= 16'h467c;
        src5 <= 16'haf73;
        src6 <= 16'h8a39;
        src7 <= 16'h1988;
        src8 <= 16'h1a24;
        src9 <= 16'ha0e0;
        src10 <= 16'hcc38;
        src11 <= 16'he7ea;
        src12 <= 16'h6e2c;
        src13 <= 16'hd9ce;
        src14 <= 16'hae92;
        src15 <= 16'heca;
        src16 <= 16'hf41f;
        src17 <= 16'hc9cf;
        src18 <= 16'h7d1a;
        src19 <= 16'h4fc3;
        src20 <= 16'hfa8d;
        src21 <= 16'h26b5;
        src22 <= 16'hbad0;
        src23 <= 16'h9eed;
        src24 <= 16'he28d;
        src25 <= 16'he60c;
        src26 <= 16'h2112;
        src27 <= 16'h5c73;
        src28 <= 16'h7c3f;
        src29 <= 16'h922d;
        src30 <= 16'h250b;
        src31 <= 16'h7170;
        src32 <= 16'ha534;
        src33 <= 16'h8e0f;
        src34 <= 16'h91e2;
        src35 <= 16'h750f;
        src36 <= 16'hd806;
        src37 <= 16'h2dd3;
        src38 <= 16'h5caf;
        src39 <= 16'hab6e;
        src40 <= 16'hbecf;
        src41 <= 16'h659b;
        src42 <= 16'hbe29;
        src43 <= 16'h2cd;
        src44 <= 16'h4685;
        src45 <= 16'he372;
        src46 <= 16'hc8f4;
        src47 <= 16'h393a;
        src48 <= 16'h4124;
        src49 <= 16'heb6a;
        src50 <= 16'h320f;
        src51 <= 16'hce09;
        src52 <= 16'hf8ad;
        src53 <= 16'ha567;
        src54 <= 16'h613d;
        src55 <= 16'hd855;
        src56 <= 16'hc0f5;
        src57 <= 16'h7f53;
        src58 <= 16'he349;
        src59 <= 16'he0ee;
        src60 <= 16'hb755;
        src61 <= 16'hde38;
        src62 <= 16'h2c78;
        src63 <= 16'h887;
        exp <= 22'h2379aa;
        #1
        src0 <= 16'h4ce9;
        src1 <= 16'h32d9;
        src2 <= 16'ha3a0;
        src3 <= 16'hf7;
        src4 <= 16'ha0e1;
        src5 <= 16'h7a33;
        src6 <= 16'he0f7;
        src7 <= 16'h1e8c;
        src8 <= 16'h171f;
        src9 <= 16'hd04;
        src10 <= 16'h46da;
        src11 <= 16'h6973;
        src12 <= 16'hc53a;
        src13 <= 16'hb1a3;
        src14 <= 16'h8bcb;
        src15 <= 16'hca44;
        src16 <= 16'h54f1;
        src17 <= 16'hf535;
        src18 <= 16'h53aa;
        src19 <= 16'h36c0;
        src20 <= 16'h356f;
        src21 <= 16'h3be2;
        src22 <= 16'ha9e4;
        src23 <= 16'h6391;
        src24 <= 16'h4726;
        src25 <= 16'h63ed;
        src26 <= 16'h1cda;
        src27 <= 16'h8e8c;
        src28 <= 16'hca0;
        src29 <= 16'hcf6d;
        src30 <= 16'hceba;
        src31 <= 16'he67;
        src32 <= 16'h56fa;
        src33 <= 16'h3003;
        src34 <= 16'hc3f1;
        src35 <= 16'hfd4b;
        src36 <= 16'hb25d;
        src37 <= 16'h355b;
        src38 <= 16'hb9e5;
        src39 <= 16'he7e8;
        src40 <= 16'h401f;
        src41 <= 16'hba5c;
        src42 <= 16'h518d;
        src43 <= 16'haa8c;
        src44 <= 16'h237f;
        src45 <= 16'ha7d6;
        src46 <= 16'h3423;
        src47 <= 16'h14a5;
        src48 <= 16'h3c0;
        src49 <= 16'he40f;
        src50 <= 16'h2243;
        src51 <= 16'h136f;
        src52 <= 16'hba30;
        src53 <= 16'h28d5;
        src54 <= 16'habe7;
        src55 <= 16'hcfbe;
        src56 <= 16'haf29;
        src57 <= 16'h9bb8;
        src58 <= 16'h3458;
        src59 <= 16'hfe79;
        src60 <= 16'h48ef;
        src61 <= 16'hd735;
        src62 <= 16'hd504;
        src63 <= 16'hb1e8;
        exp <= 22'h1dc0a5;
        #1
        src0 <= 16'h8484;
        src1 <= 16'h57b;
        src2 <= 16'hc6f4;
        src3 <= 16'h9d21;
        src4 <= 16'h121d;
        src5 <= 16'h144e;
        src6 <= 16'hfaf2;
        src7 <= 16'h8951;
        src8 <= 16'h853d;
        src9 <= 16'h7db6;
        src10 <= 16'hdc13;
        src11 <= 16'h9a19;
        src12 <= 16'h8c55;
        src13 <= 16'hae1;
        src14 <= 16'h36f8;
        src15 <= 16'h943d;
        src16 <= 16'h266b;
        src17 <= 16'h660b;
        src18 <= 16'h77ca;
        src19 <= 16'hd6a2;
        src20 <= 16'hf1e6;
        src21 <= 16'he09c;
        src22 <= 16'h33b8;
        src23 <= 16'h1e31;
        src24 <= 16'h5178;
        src25 <= 16'hf288;
        src26 <= 16'hec0b;
        src27 <= 16'h578b;
        src28 <= 16'h20;
        src29 <= 16'he9f0;
        src30 <= 16'h7f80;
        src31 <= 16'h9fdd;
        src32 <= 16'h5437;
        src33 <= 16'h29af;
        src34 <= 16'h2024;
        src35 <= 16'h5678;
        src36 <= 16'h75c;
        src37 <= 16'h27ba;
        src38 <= 16'he72e;
        src39 <= 16'h4129;
        src40 <= 16'h9864;
        src41 <= 16'h5d24;
        src42 <= 16'hfc05;
        src43 <= 16'h93e5;
        src44 <= 16'h6772;
        src45 <= 16'heba0;
        src46 <= 16'h1f5;
        src47 <= 16'h179;
        src48 <= 16'hc7c0;
        src49 <= 16'h1ea3;
        src50 <= 16'hf496;
        src51 <= 16'h1e5c;
        src52 <= 16'heb2e;
        src53 <= 16'h7fe1;
        src54 <= 16'hfc6b;
        src55 <= 16'h81e1;
        src56 <= 16'h5526;
        src57 <= 16'h3774;
        src58 <= 16'h277a;
        src59 <= 16'h8e7b;
        src60 <= 16'h5f4c;
        src61 <= 16'h5d51;
        src62 <= 16'h1cec;
        src63 <= 16'h6aca;
        exp <= 22'h1d960f;
        #1
        src0 <= 16'ha1df;
        src1 <= 16'h1325;
        src2 <= 16'h5d14;
        src3 <= 16'hd5f0;
        src4 <= 16'hcc74;
        src5 <= 16'h62ed;
        src6 <= 16'hda22;
        src7 <= 16'h1b65;
        src8 <= 16'h9ea2;
        src9 <= 16'haa32;
        src10 <= 16'h8e84;
        src11 <= 16'h3269;
        src12 <= 16'h47bf;
        src13 <= 16'h6fa9;
        src14 <= 16'had7;
        src15 <= 16'ha674;
        src16 <= 16'h9a4d;
        src17 <= 16'hc6f7;
        src18 <= 16'h16ff;
        src19 <= 16'h9cef;
        src20 <= 16'h1b11;
        src21 <= 16'hd653;
        src22 <= 16'h379b;
        src23 <= 16'h5a42;
        src24 <= 16'h3350;
        src25 <= 16'h2e28;
        src26 <= 16'h62e0;
        src27 <= 16'h418d;
        src28 <= 16'hd597;
        src29 <= 16'h94e6;
        src30 <= 16'hf227;
        src31 <= 16'h34f1;
        src32 <= 16'hd744;
        src33 <= 16'h9612;
        src34 <= 16'ha32e;
        src35 <= 16'h5269;
        src36 <= 16'he45c;
        src37 <= 16'h9644;
        src38 <= 16'h6705;
        src39 <= 16'h7f33;
        src40 <= 16'ha1cd;
        src41 <= 16'hbd2c;
        src42 <= 16'h17d7;
        src43 <= 16'h270b;
        src44 <= 16'h2657;
        src45 <= 16'hbda3;
        src46 <= 16'hdc08;
        src47 <= 16'hd94;
        src48 <= 16'hf73b;
        src49 <= 16'hbf33;
        src50 <= 16'h8d18;
        src51 <= 16'hfdc3;
        src52 <= 16'h6d48;
        src53 <= 16'h3125;
        src54 <= 16'h2c7d;
        src55 <= 16'hcc8d;
        src56 <= 16'h52e4;
        src57 <= 16'h7064;
        src58 <= 16'h437e;
        src59 <= 16'hdae7;
        src60 <= 16'ha9cb;
        src61 <= 16'h5562;
        src62 <= 16'h26e2;
        src63 <= 16'h7825;
        exp <= 22'h1f3728;
        #1
        src0 <= 16'h14a6;
        src1 <= 16'h2de4;
        src2 <= 16'h9abb;
        src3 <= 16'h78a;
        src4 <= 16'hf1ea;
        src5 <= 16'h520f;
        src6 <= 16'h8698;
        src7 <= 16'h506;
        src8 <= 16'h987f;
        src9 <= 16'h69d0;
        src10 <= 16'h593b;
        src11 <= 16'h78fc;
        src12 <= 16'he236;
        src13 <= 16'h45fd;
        src14 <= 16'hfc90;
        src15 <= 16'hfcab;
        src16 <= 16'h8a19;
        src17 <= 16'h6095;
        src18 <= 16'had99;
        src19 <= 16'h4c5b;
        src20 <= 16'h7d83;
        src21 <= 16'hd023;
        src22 <= 16'h1d7f;
        src23 <= 16'h7f;
        src24 <= 16'h5f90;
        src25 <= 16'hcd8c;
        src26 <= 16'h28ea;
        src27 <= 16'hae0d;
        src28 <= 16'heed3;
        src29 <= 16'he736;
        src30 <= 16'h4971;
        src31 <= 16'h177a;
        src32 <= 16'h3fa5;
        src33 <= 16'h89d2;
        src34 <= 16'h2932;
        src35 <= 16'hfa1d;
        src36 <= 16'he340;
        src37 <= 16'h46ca;
        src38 <= 16'h465;
        src39 <= 16'hb9d;
        src40 <= 16'h8b18;
        src41 <= 16'h8853;
        src42 <= 16'hc71f;
        src43 <= 16'h6588;
        src44 <= 16'h1a1c;
        src45 <= 16'h5f6b;
        src46 <= 16'hb33f;
        src47 <= 16'hdd63;
        src48 <= 16'h4f25;
        src49 <= 16'h98b6;
        src50 <= 16'h6dc0;
        src51 <= 16'h5678;
        src52 <= 16'hfe07;
        src53 <= 16'hd7a8;
        src54 <= 16'haeea;
        src55 <= 16'hc06a;
        src56 <= 16'h251e;
        src57 <= 16'h360a;
        src58 <= 16'h39f7;
        src59 <= 16'hdfaf;
        src60 <= 16'h25ba;
        src61 <= 16'h1926;
        src62 <= 16'h2064;
        src63 <= 16'haa5e;
        exp <= 22'h1e163a;
        #1
        src0 <= 16'h21d3;
        src1 <= 16'hb2b4;
        src2 <= 16'hf152;
        src3 <= 16'ha6e8;
        src4 <= 16'h26a4;
        src5 <= 16'h2f42;
        src6 <= 16'hc8f8;
        src7 <= 16'h8cd6;
        src8 <= 16'h333e;
        src9 <= 16'h9e93;
        src10 <= 16'h1f0;
        src11 <= 16'he7eb;
        src12 <= 16'haecc;
        src13 <= 16'h9e08;
        src14 <= 16'h7b42;
        src15 <= 16'h8bcc;
        src16 <= 16'h3b06;
        src17 <= 16'he983;
        src18 <= 16'h9e84;
        src19 <= 16'h323f;
        src20 <= 16'h5582;
        src21 <= 16'h9505;
        src22 <= 16'h9c94;
        src23 <= 16'h9f9b;
        src24 <= 16'hd25;
        src25 <= 16'h5521;
        src26 <= 16'h36ce;
        src27 <= 16'hfd0b;
        src28 <= 16'hb2b7;
        src29 <= 16'h3f4a;
        src30 <= 16'h1de9;
        src31 <= 16'h40e4;
        src32 <= 16'h5208;
        src33 <= 16'h1d9d;
        src34 <= 16'h2e59;
        src35 <= 16'h1782;
        src36 <= 16'hc755;
        src37 <= 16'h1c17;
        src38 <= 16'h1c94;
        src39 <= 16'ha5a2;
        src40 <= 16'hfe3b;
        src41 <= 16'h7eb1;
        src42 <= 16'h173e;
        src43 <= 16'h371a;
        src44 <= 16'h267f;
        src45 <= 16'hd2d7;
        src46 <= 16'h3a65;
        src47 <= 16'h223f;
        src48 <= 16'hb6ab;
        src49 <= 16'h403e;
        src50 <= 16'h3890;
        src51 <= 16'h5140;
        src52 <= 16'hd6f7;
        src53 <= 16'hb38d;
        src54 <= 16'h1cfa;
        src55 <= 16'h4a10;
        src56 <= 16'h2536;
        src57 <= 16'h983b;
        src58 <= 16'h5e65;
        src59 <= 16'hb520;
        src60 <= 16'h953e;
        src61 <= 16'hf39b;
        src62 <= 16'h9ea6;
        src63 <= 16'h5157;
        exp <= 22'h1c6365;
        #1
        src0 <= 16'hee0d;
        src1 <= 16'h1453;
        src2 <= 16'hd08;
        src3 <= 16'h7ae4;
        src4 <= 16'h76ce;
        src5 <= 16'hb226;
        src6 <= 16'h6a48;
        src7 <= 16'hfff2;
        src8 <= 16'h5600;
        src9 <= 16'ha517;
        src10 <= 16'h7f43;
        src11 <= 16'h196c;
        src12 <= 16'ha30c;
        src13 <= 16'h32bd;
        src14 <= 16'he92c;
        src15 <= 16'hd1b0;
        src16 <= 16'h6ee5;
        src17 <= 16'ha701;
        src18 <= 16'h59d6;
        src19 <= 16'h3dd0;
        src20 <= 16'h978e;
        src21 <= 16'h3fb9;
        src22 <= 16'hd719;
        src23 <= 16'h35c;
        src24 <= 16'h548f;
        src25 <= 16'h649d;
        src26 <= 16'h19fb;
        src27 <= 16'h7416;
        src28 <= 16'h3798;
        src29 <= 16'h1606;
        src30 <= 16'h680e;
        src31 <= 16'hb966;
        src32 <= 16'h102;
        src33 <= 16'hedc2;
        src34 <= 16'h3c41;
        src35 <= 16'h5d2c;
        src36 <= 16'hdaf6;
        src37 <= 16'hed1;
        src38 <= 16'h7b58;
        src39 <= 16'hc088;
        src40 <= 16'h1616;
        src41 <= 16'h5d1d;
        src42 <= 16'ha980;
        src43 <= 16'h2967;
        src44 <= 16'h76e8;
        src45 <= 16'h80f0;
        src46 <= 16'hd66a;
        src47 <= 16'hd60c;
        src48 <= 16'h86b6;
        src49 <= 16'h2f85;
        src50 <= 16'h66b5;
        src51 <= 16'hd97e;
        src52 <= 16'h84aa;
        src53 <= 16'h7d7d;
        src54 <= 16'hb402;
        src55 <= 16'h6c0c;
        src56 <= 16'hbdf;
        src57 <= 16'h25d1;
        src58 <= 16'h55cd;
        src59 <= 16'hdc75;
        src60 <= 16'hface;
        src61 <= 16'h8afd;
        src62 <= 16'h4dc6;
        src63 <= 16'h53bb;
        exp <= 22'h1d939d;
        #1
        src0 <= 16'h58ee;
        src1 <= 16'h466e;
        src2 <= 16'h78fa;
        src3 <= 16'he3f1;
        src4 <= 16'h50d1;
        src5 <= 16'h293d;
        src6 <= 16'h44c2;
        src7 <= 16'hc392;
        src8 <= 16'h11eb;
        src9 <= 16'hc0c0;
        src10 <= 16'h6091;
        src11 <= 16'hdfe6;
        src12 <= 16'h422b;
        src13 <= 16'ha59d;
        src14 <= 16'hf4f1;
        src15 <= 16'h5897;
        src16 <= 16'hfc60;
        src17 <= 16'h8cfa;
        src18 <= 16'h8674;
        src19 <= 16'hf42;
        src20 <= 16'h36c7;
        src21 <= 16'h93d7;
        src22 <= 16'h1d0e;
        src23 <= 16'he2ec;
        src24 <= 16'h53f9;
        src25 <= 16'h1cee;
        src26 <= 16'hab8c;
        src27 <= 16'h989b;
        src28 <= 16'h907;
        src29 <= 16'h7e1;
        src30 <= 16'he6b7;
        src31 <= 16'hb82f;
        src32 <= 16'h2d7a;
        src33 <= 16'h631a;
        src34 <= 16'h38f7;
        src35 <= 16'hb76d;
        src36 <= 16'h981d;
        src37 <= 16'hff84;
        src38 <= 16'hd5fa;
        src39 <= 16'hfda;
        src40 <= 16'hbe6d;
        src41 <= 16'hc18f;
        src42 <= 16'ha5e8;
        src43 <= 16'ha1ca;
        src44 <= 16'hce5d;
        src45 <= 16'hda94;
        src46 <= 16'h7ee2;
        src47 <= 16'had42;
        src48 <= 16'h3beb;
        src49 <= 16'h3277;
        src50 <= 16'h70f6;
        src51 <= 16'hc1ad;
        src52 <= 16'h2a48;
        src53 <= 16'hbb0d;
        src54 <= 16'h1f69;
        src55 <= 16'h4c8a;
        src56 <= 16'h3d1a;
        src57 <= 16'hb1b8;
        src58 <= 16'hb89b;
        src59 <= 16'h1f44;
        src60 <= 16'h6751;
        src61 <= 16'hc228;
        src62 <= 16'hed5a;
        src63 <= 16'h6d18;
        exp <= 22'h1fedb8;
        #1
        src0 <= 16'hed75;
        src1 <= 16'ha8ac;
        src2 <= 16'h2cb;
        src3 <= 16'hbc53;
        src4 <= 16'hfd2c;
        src5 <= 16'h81dd;
        src6 <= 16'h9adf;
        src7 <= 16'h3b94;
        src8 <= 16'hf9d7;
        src9 <= 16'h5148;
        src10 <= 16'h8d66;
        src11 <= 16'hbf48;
        src12 <= 16'hd339;
        src13 <= 16'h21ff;
        src14 <= 16'h4a42;
        src15 <= 16'hf8ae;
        src16 <= 16'h44d3;
        src17 <= 16'hf321;
        src18 <= 16'hbf0c;
        src19 <= 16'heb0a;
        src20 <= 16'ha429;
        src21 <= 16'hc35d;
        src22 <= 16'hddde;
        src23 <= 16'hb869;
        src24 <= 16'h986a;
        src25 <= 16'h714c;
        src26 <= 16'h98e0;
        src27 <= 16'h8f37;
        src28 <= 16'h2d4;
        src29 <= 16'he78d;
        src30 <= 16'h190f;
        src31 <= 16'hef09;
        src32 <= 16'hb4d1;
        src33 <= 16'hd01f;
        src34 <= 16'h1dec;
        src35 <= 16'h4f99;
        src36 <= 16'h84a5;
        src37 <= 16'h43fb;
        src38 <= 16'h17ae;
        src39 <= 16'h64b;
        src40 <= 16'h3928;
        src41 <= 16'h3ce9;
        src42 <= 16'h5cd4;
        src43 <= 16'hceff;
        src44 <= 16'he90d;
        src45 <= 16'h581a;
        src46 <= 16'h64c4;
        src47 <= 16'h94b9;
        src48 <= 16'h375f;
        src49 <= 16'ha8a2;
        src50 <= 16'h8729;
        src51 <= 16'hd0cc;
        src52 <= 16'he0fb;
        src53 <= 16'hed1c;
        src54 <= 16'h7db0;
        src55 <= 16'hd84b;
        src56 <= 16'h427b;
        src57 <= 16'hec02;
        src58 <= 16'h77ef;
        src59 <= 16'h3e5c;
        src60 <= 16'h6016;
        src61 <= 16'h8bf7;
        src62 <= 16'h5e47;
        src63 <= 16'h4e40;
        exp <= 22'h230dc7;
        #1
        src0 <= 16'h9c1b;
        src1 <= 16'h368b;
        src2 <= 16'h6c71;
        src3 <= 16'h8b05;
        src4 <= 16'h7c18;
        src5 <= 16'h3463;
        src6 <= 16'h6def;
        src7 <= 16'ha8ed;
        src8 <= 16'hda65;
        src9 <= 16'h48f8;
        src10 <= 16'hdd72;
        src11 <= 16'h4012;
        src12 <= 16'hcdeb;
        src13 <= 16'h2a6a;
        src14 <= 16'hd6a8;
        src15 <= 16'h8b89;
        src16 <= 16'hd24c;
        src17 <= 16'h35f5;
        src18 <= 16'hb1a8;
        src19 <= 16'h917;
        src20 <= 16'hd3bc;
        src21 <= 16'haf9;
        src22 <= 16'hcf6e;
        src23 <= 16'h493b;
        src24 <= 16'h45bd;
        src25 <= 16'h8515;
        src26 <= 16'habfa;
        src27 <= 16'h5683;
        src28 <= 16'he3bb;
        src29 <= 16'h983c;
        src30 <= 16'h786;
        src31 <= 16'hed46;
        src32 <= 16'h8930;
        src33 <= 16'h3415;
        src34 <= 16'h3d1b;
        src35 <= 16'hb53a;
        src36 <= 16'h5ee0;
        src37 <= 16'hc1a1;
        src38 <= 16'h9a58;
        src39 <= 16'h637e;
        src40 <= 16'hf6fd;
        src41 <= 16'h3aba;
        src42 <= 16'h3ee8;
        src43 <= 16'h8e86;
        src44 <= 16'h5991;
        src45 <= 16'hd66b;
        src46 <= 16'h696a;
        src47 <= 16'h6505;
        src48 <= 16'hed5c;
        src49 <= 16'h3b6d;
        src50 <= 16'hb287;
        src51 <= 16'ha43e;
        src52 <= 16'hcadd;
        src53 <= 16'h8e7d;
        src54 <= 16'h682a;
        src55 <= 16'h6000;
        src56 <= 16'hdf97;
        src57 <= 16'h9cc1;
        src58 <= 16'h91aa;
        src59 <= 16'h53e4;
        src60 <= 16'hf3dc;
        src61 <= 16'hb297;
        src62 <= 16'h1808;
        src63 <= 16'h775f;
        exp <= 22'h21299d;
        #1
        src0 <= 16'h2a4b;
        src1 <= 16'hebc;
        src2 <= 16'hf33b;
        src3 <= 16'he311;
        src4 <= 16'ha033;
        src5 <= 16'h666b;
        src6 <= 16'hda3;
        src7 <= 16'h4fd0;
        src8 <= 16'hefbf;
        src9 <= 16'h14de;
        src10 <= 16'hd2d8;
        src11 <= 16'h3749;
        src12 <= 16'h67b0;
        src13 <= 16'h8b78;
        src14 <= 16'h1c19;
        src15 <= 16'hab30;
        src16 <= 16'hd2c1;
        src17 <= 16'h92f5;
        src18 <= 16'h45f3;
        src19 <= 16'h3d20;
        src20 <= 16'h1d51;
        src21 <= 16'h684;
        src22 <= 16'he522;
        src23 <= 16'he887;
        src24 <= 16'h4769;
        src25 <= 16'hac08;
        src26 <= 16'hdb4d;
        src27 <= 16'h924b;
        src28 <= 16'h662c;
        src29 <= 16'h17b2;
        src30 <= 16'hb706;
        src31 <= 16'hb640;
        src32 <= 16'h3da2;
        src33 <= 16'he158;
        src34 <= 16'h2aa6;
        src35 <= 16'h7797;
        src36 <= 16'h8496;
        src37 <= 16'h7ff;
        src38 <= 16'h22a8;
        src39 <= 16'heba2;
        src40 <= 16'he91c;
        src41 <= 16'h39ee;
        src42 <= 16'hdca;
        src43 <= 16'hb94e;
        src44 <= 16'h2ec7;
        src45 <= 16'hfb99;
        src46 <= 16'hd9fe;
        src47 <= 16'hd420;
        src48 <= 16'hc116;
        src49 <= 16'h7649;
        src50 <= 16'h2060;
        src51 <= 16'he23b;
        src52 <= 16'h4d09;
        src53 <= 16'h19c2;
        src54 <= 16'h1cf8;
        src55 <= 16'he281;
        src56 <= 16'ha350;
        src57 <= 16'he2a4;
        src58 <= 16'hfc7d;
        src59 <= 16'hb2f5;
        src60 <= 16'hb72d;
        src61 <= 16'hbdda;
        src62 <= 16'h84ac;
        src63 <= 16'hc799;
        exp <= 22'h2118ad;
        #1
        src0 <= 16'hb859;
        src1 <= 16'h2510;
        src2 <= 16'hc0e4;
        src3 <= 16'hb150;
        src4 <= 16'h3b0b;
        src5 <= 16'hd0d8;
        src6 <= 16'h7a19;
        src7 <= 16'hfe7c;
        src8 <= 16'h630d;
        src9 <= 16'hff9d;
        src10 <= 16'hc8e3;
        src11 <= 16'hcc94;
        src12 <= 16'h5ef9;
        src13 <= 16'haf32;
        src14 <= 16'h37f;
        src15 <= 16'hb520;
        src16 <= 16'hebc5;
        src17 <= 16'h213c;
        src18 <= 16'h22e2;
        src19 <= 16'hed7b;
        src20 <= 16'h2a1;
        src21 <= 16'hd669;
        src22 <= 16'h1ab5;
        src23 <= 16'h3728;
        src24 <= 16'hc721;
        src25 <= 16'hb9c0;
        src26 <= 16'ha2ad;
        src27 <= 16'h3477;
        src28 <= 16'h8786;
        src29 <= 16'h1e1e;
        src30 <= 16'hb87b;
        src31 <= 16'heb3e;
        src32 <= 16'hc0e5;
        src33 <= 16'hc878;
        src34 <= 16'h3058;
        src35 <= 16'h4e5;
        src36 <= 16'h2a86;
        src37 <= 16'h4074;
        src38 <= 16'h8375;
        src39 <= 16'h9330;
        src40 <= 16'ha7e0;
        src41 <= 16'h7a5c;
        src42 <= 16'ha315;
        src43 <= 16'hc510;
        src44 <= 16'hf89d;
        src45 <= 16'hfe49;
        src46 <= 16'h9e31;
        src47 <= 16'h26;
        src48 <= 16'h6824;
        src49 <= 16'h47f1;
        src50 <= 16'hab79;
        src51 <= 16'h2346;
        src52 <= 16'ha77d;
        src53 <= 16'h6184;
        src54 <= 16'h78a9;
        src55 <= 16'h4d3f;
        src56 <= 16'hb773;
        src57 <= 16'hed17;
        src58 <= 16'h189b;
        src59 <= 16'h95bc;
        src60 <= 16'he336;
        src61 <= 16'he107;
        src62 <= 16'h18bd;
        src63 <= 16'h6512;
        exp <= 22'h21bf28;
        #1
        src0 <= 16'hd33b;
        src1 <= 16'h8edf;
        src2 <= 16'h7111;
        src3 <= 16'hee00;
        src4 <= 16'h11f1;
        src5 <= 16'h8423;
        src6 <= 16'hf0bd;
        src7 <= 16'hf311;
        src8 <= 16'h6187;
        src9 <= 16'h7159;
        src10 <= 16'hbeb5;
        src11 <= 16'h8e7;
        src12 <= 16'hde56;
        src13 <= 16'h8670;
        src14 <= 16'h8c1d;
        src15 <= 16'he05d;
        src16 <= 16'hce33;
        src17 <= 16'h363d;
        src18 <= 16'hc834;
        src19 <= 16'hb665;
        src20 <= 16'h89b0;
        src21 <= 16'h8805;
        src22 <= 16'h5638;
        src23 <= 16'h13b0;
        src24 <= 16'h3a50;
        src25 <= 16'hc6d2;
        src26 <= 16'hb1f8;
        src27 <= 16'h8787;
        src28 <= 16'h9aa;
        src29 <= 16'h7f30;
        src30 <= 16'h79d6;
        src31 <= 16'h70e9;
        src32 <= 16'ha62;
        src33 <= 16'h945d;
        src34 <= 16'he184;
        src35 <= 16'hb77c;
        src36 <= 16'had00;
        src37 <= 16'hc22a;
        src38 <= 16'h53b7;
        src39 <= 16'ha925;
        src40 <= 16'hbea6;
        src41 <= 16'h76b8;
        src42 <= 16'h7a07;
        src43 <= 16'h9acd;
        src44 <= 16'hdd05;
        src45 <= 16'h5297;
        src46 <= 16'h7417;
        src47 <= 16'h8e28;
        src48 <= 16'ha1c;
        src49 <= 16'ha621;
        src50 <= 16'ha459;
        src51 <= 16'h147f;
        src52 <= 16'hfdb9;
        src53 <= 16'hcb5a;
        src54 <= 16'hc198;
        src55 <= 16'h6f77;
        src56 <= 16'h57b4;
        src57 <= 16'ha1e3;
        src58 <= 16'h9caa;
        src59 <= 16'he80f;
        src60 <= 16'hae0d;
        src61 <= 16'ha464;
        src62 <= 16'h48ce;
        src63 <= 16'h2043;
        exp <= 22'h231084;
        #1
        src0 <= 16'hccb5;
        src1 <= 16'h9211;
        src2 <= 16'h8774;
        src3 <= 16'h9ddd;
        src4 <= 16'h875d;
        src5 <= 16'hccdc;
        src6 <= 16'h3d92;
        src7 <= 16'h5fb0;
        src8 <= 16'h1587;
        src9 <= 16'h6282;
        src10 <= 16'h475b;
        src11 <= 16'h1305;
        src12 <= 16'h26c9;
        src13 <= 16'hdf0;
        src14 <= 16'h1ce9;
        src15 <= 16'h6616;
        src16 <= 16'h5b35;
        src17 <= 16'h2d21;
        src18 <= 16'h4c33;
        src19 <= 16'hbe8;
        src20 <= 16'h316e;
        src21 <= 16'hc045;
        src22 <= 16'h86d;
        src23 <= 16'hf76f;
        src24 <= 16'h9aba;
        src25 <= 16'hafd4;
        src26 <= 16'hcd14;
        src27 <= 16'h22df;
        src28 <= 16'h3284;
        src29 <= 16'hfd65;
        src30 <= 16'hdd36;
        src31 <= 16'hdaed;
        src32 <= 16'hddb3;
        src33 <= 16'hba65;
        src34 <= 16'hcd7f;
        src35 <= 16'h9cb4;
        src36 <= 16'h41e6;
        src37 <= 16'h737c;
        src38 <= 16'hf4f9;
        src39 <= 16'hcabd;
        src40 <= 16'hee9a;
        src41 <= 16'hf41a;
        src42 <= 16'h10b;
        src43 <= 16'ha6eb;
        src44 <= 16'h527c;
        src45 <= 16'hb197;
        src46 <= 16'h3cf2;
        src47 <= 16'hd4c9;
        src48 <= 16'h712f;
        src49 <= 16'he097;
        src50 <= 16'h570f;
        src51 <= 16'h77a9;
        src52 <= 16'h5dfa;
        src53 <= 16'hf47c;
        src54 <= 16'hd3fe;
        src55 <= 16'ha0f;
        src56 <= 16'hb9b9;
        src57 <= 16'hbab0;
        src58 <= 16'h13b5;
        src59 <= 16'hab6b;
        src60 <= 16'h7160;
        src61 <= 16'hdaf;
        src62 <= 16'h8aa1;
        src63 <= 16'h577b;
        exp <= 22'h1ff1d0;
        #1
        src0 <= 16'h1a7d;
        src1 <= 16'h7418;
        src2 <= 16'h234c;
        src3 <= 16'h9db9;
        src4 <= 16'hff5d;
        src5 <= 16'hdaae;
        src6 <= 16'ha1b1;
        src7 <= 16'h40a7;
        src8 <= 16'h496d;
        src9 <= 16'h5369;
        src10 <= 16'h2c5a;
        src11 <= 16'ha46d;
        src12 <= 16'h8d6e;
        src13 <= 16'h2704;
        src14 <= 16'hbcd5;
        src15 <= 16'hcb1a;
        src16 <= 16'h953c;
        src17 <= 16'h49f6;
        src18 <= 16'h78c0;
        src19 <= 16'he0b4;
        src20 <= 16'h990a;
        src21 <= 16'hb197;
        src22 <= 16'hed4e;
        src23 <= 16'h990e;
        src24 <= 16'h8cc8;
        src25 <= 16'hb49f;
        src26 <= 16'h1e67;
        src27 <= 16'h3260;
        src28 <= 16'ha17a;
        src29 <= 16'ha8ef;
        src30 <= 16'h76dc;
        src31 <= 16'hf6d1;
        src32 <= 16'h1;
        src33 <= 16'he38b;
        src34 <= 16'hfd89;
        src35 <= 16'h1852;
        src36 <= 16'hff82;
        src37 <= 16'hb376;
        src38 <= 16'h2e6e;
        src39 <= 16'hcec6;
        src40 <= 16'h13e3;
        src41 <= 16'h1630;
        src42 <= 16'hc68;
        src43 <= 16'h8832;
        src44 <= 16'hfaf9;
        src45 <= 16'h8ad1;
        src46 <= 16'h3b8b;
        src47 <= 16'h5c7e;
        src48 <= 16'h87ec;
        src49 <= 16'hdeed;
        src50 <= 16'h4d3a;
        src51 <= 16'hc049;
        src52 <= 16'h3b9c;
        src53 <= 16'hcaf;
        src54 <= 16'h6806;
        src55 <= 16'h4fba;
        src56 <= 16'hfdf0;
        src57 <= 16'h13c;
        src58 <= 16'h7c8b;
        src59 <= 16'hed5e;
        src60 <= 16'h5141;
        src61 <= 16'h5908;
        src62 <= 16'he07c;
        src63 <= 16'hb9f4;
        exp <= 22'h20b22a;
        #1
        src0 <= 16'hb0f4;
        src1 <= 16'hde1f;
        src2 <= 16'h14a9;
        src3 <= 16'h3ec7;
        src4 <= 16'h112f;
        src5 <= 16'he369;
        src6 <= 16'hee67;
        src7 <= 16'h46a3;
        src8 <= 16'h99a1;
        src9 <= 16'hcbc3;
        src10 <= 16'h4ccc;
        src11 <= 16'hb7c3;
        src12 <= 16'h6978;
        src13 <= 16'hfa7b;
        src14 <= 16'ha5b5;
        src15 <= 16'h734b;
        src16 <= 16'hcca8;
        src17 <= 16'h968e;
        src18 <= 16'h38ec;
        src19 <= 16'h7287;
        src20 <= 16'h424b;
        src21 <= 16'h7d37;
        src22 <= 16'hd205;
        src23 <= 16'h54fa;
        src24 <= 16'hcfd8;
        src25 <= 16'h94e2;
        src26 <= 16'h2d85;
        src27 <= 16'hada9;
        src28 <= 16'hb5f6;
        src29 <= 16'haa69;
        src30 <= 16'hb0cb;
        src31 <= 16'h1840;
        src32 <= 16'h9616;
        src33 <= 16'h44a5;
        src34 <= 16'h76d8;
        src35 <= 16'h3c41;
        src36 <= 16'h744a;
        src37 <= 16'hf05c;
        src38 <= 16'hd404;
        src39 <= 16'h675c;
        src40 <= 16'h3ee;
        src41 <= 16'h9ad4;
        src42 <= 16'hc890;
        src43 <= 16'hc979;
        src44 <= 16'hb976;
        src45 <= 16'h79f9;
        src46 <= 16'hcb76;
        src47 <= 16'h80a1;
        src48 <= 16'h3e07;
        src49 <= 16'hc9cd;
        src50 <= 16'hb06b;
        src51 <= 16'h7c7a;
        src52 <= 16'h23c4;
        src53 <= 16'hd871;
        src54 <= 16'h8d6c;
        src55 <= 16'he852;
        src56 <= 16'hff93;
        src57 <= 16'hb5c8;
        src58 <= 16'h11e3;
        src59 <= 16'h264e;
        src60 <= 16'h8946;
        src61 <= 16'h2fc0;
        src62 <= 16'h5a2a;
        src63 <= 16'h317;
        exp <= 22'h21da31;
        #1
        src0 <= 16'h2eff;
        src1 <= 16'hafe3;
        src2 <= 16'h9d54;
        src3 <= 16'h7d4f;
        src4 <= 16'h6671;
        src5 <= 16'hbc77;
        src6 <= 16'hef45;
        src7 <= 16'h6e8a;
        src8 <= 16'h34d8;
        src9 <= 16'ha529;
        src10 <= 16'ha4ad;
        src11 <= 16'h5337;
        src12 <= 16'he8db;
        src13 <= 16'hcb99;
        src14 <= 16'h4508;
        src15 <= 16'h3a57;
        src16 <= 16'h1590;
        src17 <= 16'hf469;
        src18 <= 16'hbdd8;
        src19 <= 16'h8eaf;
        src20 <= 16'hd46f;
        src21 <= 16'he004;
        src22 <= 16'h754b;
        src23 <= 16'hd369;
        src24 <= 16'h2001;
        src25 <= 16'h2e56;
        src26 <= 16'h714c;
        src27 <= 16'had5e;
        src28 <= 16'ha0f9;
        src29 <= 16'hfbf0;
        src30 <= 16'h662a;
        src31 <= 16'hbd3d;
        src32 <= 16'h6f89;
        src33 <= 16'h84e2;
        src34 <= 16'h9736;
        src35 <= 16'hdeed;
        src36 <= 16'heb7;
        src37 <= 16'hbc9b;
        src38 <= 16'he2cc;
        src39 <= 16'hbbb9;
        src40 <= 16'h50f9;
        src41 <= 16'h63ca;
        src42 <= 16'h3177;
        src43 <= 16'h6209;
        src44 <= 16'hbe58;
        src45 <= 16'hb36;
        src46 <= 16'h7ffe;
        src47 <= 16'he4f2;
        src48 <= 16'h578a;
        src49 <= 16'hea5f;
        src50 <= 16'h25b3;
        src51 <= 16'h285b;
        src52 <= 16'h192;
        src53 <= 16'h42a;
        src54 <= 16'h405a;
        src55 <= 16'h7ae8;
        src56 <= 16'hd89e;
        src57 <= 16'h22a6;
        src58 <= 16'h53b2;
        src59 <= 16'hfb0f;
        src60 <= 16'hadd0;
        src61 <= 16'hc208;
        src62 <= 16'hc1ad;
        src63 <= 16'h7c36;
        exp <= 22'h2194c7;
        #1
        src0 <= 16'hb4c8;
        src1 <= 16'h9a5f;
        src2 <= 16'he538;
        src3 <= 16'hbae;
        src4 <= 16'h943a;
        src5 <= 16'h5308;
        src6 <= 16'h3bf3;
        src7 <= 16'hac00;
        src8 <= 16'h70fd;
        src9 <= 16'hab00;
        src10 <= 16'h168;
        src11 <= 16'hf1b8;
        src12 <= 16'habc4;
        src13 <= 16'h1a38;
        src14 <= 16'h1fe4;
        src15 <= 16'h45f2;
        src16 <= 16'h8c87;
        src17 <= 16'hc4fe;
        src18 <= 16'h7abe;
        src19 <= 16'h94c0;
        src20 <= 16'h6cc9;
        src21 <= 16'he099;
        src22 <= 16'hc725;
        src23 <= 16'hf8e3;
        src24 <= 16'h8027;
        src25 <= 16'hfbd6;
        src26 <= 16'h881e;
        src27 <= 16'he4dc;
        src28 <= 16'h50db;
        src29 <= 16'h7981;
        src30 <= 16'h6c52;
        src31 <= 16'h832d;
        src32 <= 16'h97c5;
        src33 <= 16'hce18;
        src34 <= 16'hef64;
        src35 <= 16'h8e6b;
        src36 <= 16'hec1e;
        src37 <= 16'hbdc3;
        src38 <= 16'h9362;
        src39 <= 16'h60d3;
        src40 <= 16'h7f1c;
        src41 <= 16'h20b8;
        src42 <= 16'h2d60;
        src43 <= 16'h54e;
        src44 <= 16'hb63;
        src45 <= 16'h9855;
        src46 <= 16'h3e7;
        src47 <= 16'he0b3;
        src48 <= 16'h2493;
        src49 <= 16'h5acf;
        src50 <= 16'h128b;
        src51 <= 16'h9a88;
        src52 <= 16'h4da9;
        src53 <= 16'ha873;
        src54 <= 16'h6f2f;
        src55 <= 16'h618a;
        src56 <= 16'hea28;
        src57 <= 16'hfa74;
        src58 <= 16'h1f76;
        src59 <= 16'hc410;
        src60 <= 16'hda76;
        src61 <= 16'h6839;
        src62 <= 16'h27b;
        src63 <= 16'h9734;
        exp <= 22'h20cfd0;
        #1
        src0 <= 16'he2cc;
        src1 <= 16'h62d0;
        src2 <= 16'hc8ce;
        src3 <= 16'h52a2;
        src4 <= 16'h1455;
        src5 <= 16'hf0c2;
        src6 <= 16'hc772;
        src7 <= 16'hf3df;
        src8 <= 16'h37be;
        src9 <= 16'h7939;
        src10 <= 16'h3266;
        src11 <= 16'h2f59;
        src12 <= 16'haeff;
        src13 <= 16'h5a63;
        src14 <= 16'h3996;
        src15 <= 16'hf249;
        src16 <= 16'h8263;
        src17 <= 16'h4c93;
        src18 <= 16'h8fdd;
        src19 <= 16'h394d;
        src20 <= 16'hc7a0;
        src21 <= 16'h4576;
        src22 <= 16'h4889;
        src23 <= 16'h3ed;
        src24 <= 16'h9b91;
        src25 <= 16'hf737;
        src26 <= 16'h3aeb;
        src27 <= 16'hcc09;
        src28 <= 16'h4448;
        src29 <= 16'h3f1e;
        src30 <= 16'h48ca;
        src31 <= 16'h5e87;
        src32 <= 16'h3803;
        src33 <= 16'hbd8;
        src34 <= 16'hb132;
        src35 <= 16'h8da5;
        src36 <= 16'h2496;
        src37 <= 16'h3563;
        src38 <= 16'h9a90;
        src39 <= 16'hdbbf;
        src40 <= 16'hb106;
        src41 <= 16'h8d2e;
        src42 <= 16'h99c7;
        src43 <= 16'h3bac;
        src44 <= 16'h176;
        src45 <= 16'h972b;
        src46 <= 16'hf54e;
        src47 <= 16'hf639;
        src48 <= 16'h735;
        src49 <= 16'hcc27;
        src50 <= 16'hd94f;
        src51 <= 16'h26b;
        src52 <= 16'h63c1;
        src53 <= 16'h55bc;
        src54 <= 16'h721c;
        src55 <= 16'h4ede;
        src56 <= 16'h1f79;
        src57 <= 16'hafe;
        src58 <= 16'hc8e;
        src59 <= 16'h6a70;
        src60 <= 16'h47ba;
        src61 <= 16'h9e6c;
        src62 <= 16'h417;
        src63 <= 16'h66c2;
        exp <= 22'h1c2654;
        #1
        src0 <= 16'h86f2;
        src1 <= 16'hcccb;
        src2 <= 16'h9cb0;
        src3 <= 16'h8231;
        src4 <= 16'hf2ef;
        src5 <= 16'ha578;
        src6 <= 16'h8e2b;
        src7 <= 16'he07d;
        src8 <= 16'h33e8;
        src9 <= 16'h6579;
        src10 <= 16'h4d63;
        src11 <= 16'h2288;
        src12 <= 16'h39d1;
        src13 <= 16'h8de8;
        src14 <= 16'h576;
        src15 <= 16'he075;
        src16 <= 16'h7849;
        src17 <= 16'h2bf8;
        src18 <= 16'h1b09;
        src19 <= 16'h2cdd;
        src20 <= 16'he666;
        src21 <= 16'h4b39;
        src22 <= 16'hdc95;
        src23 <= 16'hc24;
        src24 <= 16'he6d4;
        src25 <= 16'ha939;
        src26 <= 16'h1d98;
        src27 <= 16'h2e3e;
        src28 <= 16'ha1dc;
        src29 <= 16'h771d;
        src30 <= 16'h4c3e;
        src31 <= 16'h31da;
        src32 <= 16'hc9e8;
        src33 <= 16'h6c32;
        src34 <= 16'he599;
        src35 <= 16'hc224;
        src36 <= 16'hc3cc;
        src37 <= 16'h25df;
        src38 <= 16'h2a65;
        src39 <= 16'hb300;
        src40 <= 16'h1dc2;
        src41 <= 16'h8ec3;
        src42 <= 16'hd400;
        src43 <= 16'hb0e1;
        src44 <= 16'h174e;
        src45 <= 16'h6652;
        src46 <= 16'h38c;
        src47 <= 16'hde69;
        src48 <= 16'hd0b6;
        src49 <= 16'h61a6;
        src50 <= 16'hd7a4;
        src51 <= 16'h1800;
        src52 <= 16'h4ad8;
        src53 <= 16'he25c;
        src54 <= 16'hfa7f;
        src55 <= 16'h4baf;
        src56 <= 16'h94a2;
        src57 <= 16'h3cc2;
        src58 <= 16'h8175;
        src59 <= 16'hdff8;
        src60 <= 16'h49db;
        src61 <= 16'h4a1c;
        src62 <= 16'h9770;
        src63 <= 16'h6268;
        exp <= 22'h1f35f4;
        #1
        src0 <= 16'hb58;
        src1 <= 16'hef6e;
        src2 <= 16'h62af;
        src3 <= 16'h5403;
        src4 <= 16'h8136;
        src5 <= 16'h2be;
        src6 <= 16'hee4c;
        src7 <= 16'hff32;
        src8 <= 16'h3403;
        src9 <= 16'h95df;
        src10 <= 16'h6b8a;
        src11 <= 16'h1596;
        src12 <= 16'hc747;
        src13 <= 16'hde47;
        src14 <= 16'h2dbd;
        src15 <= 16'h9954;
        src16 <= 16'hd6bb;
        src17 <= 16'hb41c;
        src18 <= 16'h50f4;
        src19 <= 16'h9ea1;
        src20 <= 16'hf0a9;
        src21 <= 16'h5ae2;
        src22 <= 16'h44c6;
        src23 <= 16'h13da;
        src24 <= 16'h980e;
        src25 <= 16'h9e88;
        src26 <= 16'hf717;
        src27 <= 16'h12d3;
        src28 <= 16'h47f2;
        src29 <= 16'h6d0d;
        src30 <= 16'h2a93;
        src31 <= 16'hb70b;
        src32 <= 16'hc196;
        src33 <= 16'hf2e5;
        src34 <= 16'h65f;
        src35 <= 16'h5939;
        src36 <= 16'h54dc;
        src37 <= 16'h2be0;
        src38 <= 16'h9f8c;
        src39 <= 16'hb459;
        src40 <= 16'h501c;
        src41 <= 16'h2201;
        src42 <= 16'h4dfb;
        src43 <= 16'h77ce;
        src44 <= 16'ha281;
        src45 <= 16'h571b;
        src46 <= 16'h6b8d;
        src47 <= 16'h64f8;
        src48 <= 16'h7e17;
        src49 <= 16'h34c7;
        src50 <= 16'h6c29;
        src51 <= 16'h432b;
        src52 <= 16'h65ab;
        src53 <= 16'h833c;
        src54 <= 16'h1934;
        src55 <= 16'h7e09;
        src56 <= 16'h494c;
        src57 <= 16'hedef;
        src58 <= 16'hb9;
        src59 <= 16'h21bd;
        src60 <= 16'hec0f;
        src61 <= 16'h761c;
        src62 <= 16'h8ce7;
        src63 <= 16'haaab;
        exp <= 22'h1d90be;
        #1
        src0 <= 16'hc763;
        src1 <= 16'h23e9;
        src2 <= 16'h88d6;
        src3 <= 16'h1123;
        src4 <= 16'hacdd;
        src5 <= 16'h8d5d;
        src6 <= 16'he6d5;
        src7 <= 16'hf685;
        src8 <= 16'had58;
        src9 <= 16'h1067;
        src10 <= 16'h4e4b;
        src11 <= 16'h1453;
        src12 <= 16'hdb3d;
        src13 <= 16'h89b8;
        src14 <= 16'h4715;
        src15 <= 16'hf160;
        src16 <= 16'h1d80;
        src17 <= 16'h7adc;
        src18 <= 16'h5849;
        src19 <= 16'hcfdc;
        src20 <= 16'hcdec;
        src21 <= 16'h2f74;
        src22 <= 16'h7505;
        src23 <= 16'h2e52;
        src24 <= 16'h5137;
        src25 <= 16'hce9c;
        src26 <= 16'haa2a;
        src27 <= 16'hb690;
        src28 <= 16'h57f7;
        src29 <= 16'hc3c;
        src30 <= 16'hf589;
        src31 <= 16'h3597;
        src32 <= 16'h60c8;
        src33 <= 16'hc954;
        src34 <= 16'h9091;
        src35 <= 16'h7188;
        src36 <= 16'heac;
        src37 <= 16'ha0be;
        src38 <= 16'h4b06;
        src39 <= 16'hb802;
        src40 <= 16'hda1a;
        src41 <= 16'h8fd2;
        src42 <= 16'h205b;
        src43 <= 16'haaf3;
        src44 <= 16'hde4;
        src45 <= 16'h4639;
        src46 <= 16'h2366;
        src47 <= 16'hddc1;
        src48 <= 16'h7fb6;
        src49 <= 16'hda3f;
        src50 <= 16'h7bad;
        src51 <= 16'hd5c5;
        src52 <= 16'h3cfa;
        src53 <= 16'ha844;
        src54 <= 16'hfa4c;
        src55 <= 16'h5dc0;
        src56 <= 16'h8019;
        src57 <= 16'he50a;
        src58 <= 16'ha1b3;
        src59 <= 16'h14a9;
        src60 <= 16'ha16b;
        src61 <= 16'h41fc;
        src62 <= 16'h7baf;
        src63 <= 16'hbfb7;
        exp <= 22'h2057da;
        #1
        src0 <= 16'h5b32;
        src1 <= 16'hbac1;
        src2 <= 16'h8a50;
        src3 <= 16'hb57b;
        src4 <= 16'hbf39;
        src5 <= 16'he286;
        src6 <= 16'h9347;
        src7 <= 16'hd958;
        src8 <= 16'h7b9;
        src9 <= 16'h45cb;
        src10 <= 16'h19a6;
        src11 <= 16'hacd1;
        src12 <= 16'hc271;
        src13 <= 16'h6943;
        src14 <= 16'hbadb;
        src15 <= 16'h48d4;
        src16 <= 16'hc341;
        src17 <= 16'h13d7;
        src18 <= 16'hd3dd;
        src19 <= 16'hda42;
        src20 <= 16'h1f06;
        src21 <= 16'hc2e9;
        src22 <= 16'hccfd;
        src23 <= 16'hadee;
        src24 <= 16'hc7c0;
        src25 <= 16'h5a9;
        src26 <= 16'h4719;
        src27 <= 16'h5cca;
        src28 <= 16'h2674;
        src29 <= 16'h1e00;
        src30 <= 16'h4429;
        src31 <= 16'hf861;
        src32 <= 16'h90df;
        src33 <= 16'h389a;
        src34 <= 16'h9aa9;
        src35 <= 16'he57;
        src36 <= 16'h2a21;
        src37 <= 16'h2c51;
        src38 <= 16'h3fc9;
        src39 <= 16'h41b2;
        src40 <= 16'hde65;
        src41 <= 16'h4b6a;
        src42 <= 16'hae5a;
        src43 <= 16'h5cee;
        src44 <= 16'ha015;
        src45 <= 16'h1c4f;
        src46 <= 16'hdf92;
        src47 <= 16'h275e;
        src48 <= 16'hcb90;
        src49 <= 16'h1250;
        src50 <= 16'h841;
        src51 <= 16'h2f11;
        src52 <= 16'hf974;
        src53 <= 16'h1c77;
        src54 <= 16'h6d69;
        src55 <= 16'hac05;
        src56 <= 16'ha745;
        src57 <= 16'h9a13;
        src58 <= 16'hc015;
        src59 <= 16'hcbe;
        src60 <= 16'hb357;
        src61 <= 16'hb46e;
        src62 <= 16'ha073;
        src63 <= 16'h1d92;
        exp <= 22'h1e3726;
        #1
        src0 <= 16'hc03e;
        src1 <= 16'h7706;
        src2 <= 16'hbd8d;
        src3 <= 16'hbe87;
        src4 <= 16'hfd7e;
        src5 <= 16'hd482;
        src6 <= 16'heb1a;
        src7 <= 16'h6da2;
        src8 <= 16'h1bf6;
        src9 <= 16'h814;
        src10 <= 16'h7f7;
        src11 <= 16'h17b8;
        src12 <= 16'hb6d2;
        src13 <= 16'hcd0f;
        src14 <= 16'h2d3a;
        src15 <= 16'h278b;
        src16 <= 16'h217b;
        src17 <= 16'ha7ea;
        src18 <= 16'h7ade;
        src19 <= 16'hf16b;
        src20 <= 16'h52f4;
        src21 <= 16'haad9;
        src22 <= 16'h93c5;
        src23 <= 16'h7bba;
        src24 <= 16'h2e1;
        src25 <= 16'h8d98;
        src26 <= 16'h45f5;
        src27 <= 16'h6301;
        src28 <= 16'h22db;
        src29 <= 16'h7728;
        src30 <= 16'hfc95;
        src31 <= 16'h7d14;
        src32 <= 16'ha396;
        src33 <= 16'h6982;
        src34 <= 16'heea5;
        src35 <= 16'he01c;
        src36 <= 16'ha86c;
        src37 <= 16'h99a1;
        src38 <= 16'hdd41;
        src39 <= 16'hc6a7;
        src40 <= 16'h16f;
        src41 <= 16'hc88;
        src42 <= 16'heff5;
        src43 <= 16'h903a;
        src44 <= 16'hf559;
        src45 <= 16'h45a5;
        src46 <= 16'h32ca;
        src47 <= 16'hc0dc;
        src48 <= 16'hf37c;
        src49 <= 16'h6aab;
        src50 <= 16'h9997;
        src51 <= 16'h9934;
        src52 <= 16'h4659;
        src53 <= 16'hca6a;
        src54 <= 16'h8fed;
        src55 <= 16'h9665;
        src56 <= 16'hbb73;
        src57 <= 16'h74fd;
        src58 <= 16'h83ee;
        src59 <= 16'h3a51;
        src60 <= 16'hbb88;
        src61 <= 16'ha61b;
        src62 <= 16'h7e;
        src63 <= 16'h7c8b;
        exp <= 22'h219e82;
        #1
        src0 <= 16'hbf43;
        src1 <= 16'hb63e;
        src2 <= 16'h9ceb;
        src3 <= 16'h6a45;
        src4 <= 16'hac2a;
        src5 <= 16'h2d74;
        src6 <= 16'h1359;
        src7 <= 16'h1489;
        src8 <= 16'hd087;
        src9 <= 16'h866b;
        src10 <= 16'h76c9;
        src11 <= 16'h327e;
        src12 <= 16'hb1c8;
        src13 <= 16'h5bbb;
        src14 <= 16'hfd03;
        src15 <= 16'h9a40;
        src16 <= 16'h810;
        src17 <= 16'hfb46;
        src18 <= 16'hc845;
        src19 <= 16'h798d;
        src20 <= 16'h3378;
        src21 <= 16'hba95;
        src22 <= 16'hd8d7;
        src23 <= 16'h61eb;
        src24 <= 16'h4538;
        src25 <= 16'hdcd3;
        src26 <= 16'h86c2;
        src27 <= 16'h188f;
        src28 <= 16'h7d64;
        src29 <= 16'hab75;
        src30 <= 16'h8c26;
        src31 <= 16'hc615;
        src32 <= 16'h916e;
        src33 <= 16'h2f9c;
        src34 <= 16'h57d3;
        src35 <= 16'h1690;
        src36 <= 16'h42d7;
        src37 <= 16'hd80c;
        src38 <= 16'h5c6b;
        src39 <= 16'h1790;
        src40 <= 16'ha378;
        src41 <= 16'h84aa;
        src42 <= 16'h1ae;
        src43 <= 16'h8e1d;
        src44 <= 16'h134e;
        src45 <= 16'h8010;
        src46 <= 16'hef9;
        src47 <= 16'h6474;
        src48 <= 16'h1ef7;
        src49 <= 16'h2bab;
        src50 <= 16'h3597;
        src51 <= 16'h54ff;
        src52 <= 16'he6df;
        src53 <= 16'h1fc7;
        src54 <= 16'h70a2;
        src55 <= 16'h8748;
        src56 <= 16'h22e8;
        src57 <= 16'h637f;
        src58 <= 16'he32b;
        src59 <= 16'h18f1;
        src60 <= 16'hea55;
        src61 <= 16'h37d6;
        src62 <= 16'hb2e5;
        src63 <= 16'h13e9;
        exp <= 22'h1c89de;
        #1
        src0 <= 16'he68f;
        src1 <= 16'h2099;
        src2 <= 16'hb635;
        src3 <= 16'hbdc;
        src4 <= 16'h2c4d;
        src5 <= 16'h2c1f;
        src6 <= 16'h1d05;
        src7 <= 16'h9490;
        src8 <= 16'h8f38;
        src9 <= 16'h569b;
        src10 <= 16'h416c;
        src11 <= 16'hf830;
        src12 <= 16'he234;
        src13 <= 16'h4b3;
        src14 <= 16'hc065;
        src15 <= 16'hea79;
        src16 <= 16'h176e;
        src17 <= 16'h57c8;
        src18 <= 16'h128c;
        src19 <= 16'h143c;
        src20 <= 16'h961c;
        src21 <= 16'h94dd;
        src22 <= 16'h49e9;
        src23 <= 16'h7d4e;
        src24 <= 16'h77cc;
        src25 <= 16'h9c68;
        src26 <= 16'h534b;
        src27 <= 16'h4910;
        src28 <= 16'hb4c5;
        src29 <= 16'heb55;
        src30 <= 16'h2996;
        src31 <= 16'had10;
        src32 <= 16'hde0e;
        src33 <= 16'hffb;
        src34 <= 16'h2bd4;
        src35 <= 16'h3a5a;
        src36 <= 16'h3992;
        src37 <= 16'h2327;
        src38 <= 16'h6c80;
        src39 <= 16'h247e;
        src40 <= 16'hcc47;
        src41 <= 16'h20db;
        src42 <= 16'hd515;
        src43 <= 16'h7ef2;
        src44 <= 16'hc758;
        src45 <= 16'h2d04;
        src46 <= 16'h60bb;
        src47 <= 16'h1ad3;
        src48 <= 16'h4db8;
        src49 <= 16'h4a5b;
        src50 <= 16'h773;
        src51 <= 16'h2668;
        src52 <= 16'h4628;
        src53 <= 16'h2fff;
        src54 <= 16'hd5ac;
        src55 <= 16'hf19e;
        src56 <= 16'h8bb0;
        src57 <= 16'hced5;
        src58 <= 16'h72ef;
        src59 <= 16'h4674;
        src60 <= 16'h426e;
        src61 <= 16'h44ef;
        src62 <= 16'h4e84;
        src63 <= 16'h7826;
        exp <= 22'h1a8c3a;
        #1
        src0 <= 16'hc9dd;
        src1 <= 16'h6984;
        src2 <= 16'h2107;
        src3 <= 16'hb3f7;
        src4 <= 16'h1c84;
        src5 <= 16'h81bc;
        src6 <= 16'h4feb;
        src7 <= 16'h156b;
        src8 <= 16'h60d2;
        src9 <= 16'h49a2;
        src10 <= 16'hc889;
        src11 <= 16'h8711;
        src12 <= 16'h1fc0;
        src13 <= 16'h63ec;
        src14 <= 16'h438b;
        src15 <= 16'hcb58;
        src16 <= 16'hc49;
        src17 <= 16'hbd56;
        src18 <= 16'h41cc;
        src19 <= 16'h2123;
        src20 <= 16'hb6e2;
        src21 <= 16'h6c4;
        src22 <= 16'hb272;
        src23 <= 16'h12f9;
        src24 <= 16'heb90;
        src25 <= 16'h47e5;
        src26 <= 16'h890c;
        src27 <= 16'hb087;
        src28 <= 16'h20c6;
        src29 <= 16'h9c4c;
        src30 <= 16'h4ec7;
        src31 <= 16'hf25f;
        src32 <= 16'hf1e9;
        src33 <= 16'hbdba;
        src34 <= 16'hec84;
        src35 <= 16'h8659;
        src36 <= 16'hc552;
        src37 <= 16'hf866;
        src38 <= 16'h17af;
        src39 <= 16'h343e;
        src40 <= 16'hc683;
        src41 <= 16'h1417;
        src42 <= 16'h502b;
        src43 <= 16'h2fbe;
        src44 <= 16'h3319;
        src45 <= 16'h93a1;
        src46 <= 16'ha810;
        src47 <= 16'hd48d;
        src48 <= 16'h2a16;
        src49 <= 16'hffaa;
        src50 <= 16'h6ce1;
        src51 <= 16'h1210;
        src52 <= 16'hcd0b;
        src53 <= 16'h143d;
        src54 <= 16'h2607;
        src55 <= 16'hb493;
        src56 <= 16'ha61a;
        src57 <= 16'h2919;
        src58 <= 16'habc2;
        src59 <= 16'h44ef;
        src60 <= 16'h4ed2;
        src61 <= 16'hbcfb;
        src62 <= 16'hb468;
        src63 <= 16'hecb9;
        exp <= 22'h1e4ed5;
        #1
        src0 <= 16'h2af7;
        src1 <= 16'he375;
        src2 <= 16'h124b;
        src3 <= 16'hc45c;
        src4 <= 16'h43f7;
        src5 <= 16'h1a0d;
        src6 <= 16'h3d4e;
        src7 <= 16'h9b27;
        src8 <= 16'h14c7;
        src9 <= 16'hf73d;
        src10 <= 16'ha1d8;
        src11 <= 16'h344;
        src12 <= 16'hf153;
        src13 <= 16'h549d;
        src14 <= 16'hd04b;
        src15 <= 16'h9487;
        src16 <= 16'h1b1e;
        src17 <= 16'h5817;
        src18 <= 16'ha5cc;
        src19 <= 16'h9fb2;
        src20 <= 16'hfd07;
        src21 <= 16'h4737;
        src22 <= 16'h2486;
        src23 <= 16'hd953;
        src24 <= 16'hb34;
        src25 <= 16'h127e;
        src26 <= 16'he45e;
        src27 <= 16'h66f;
        src28 <= 16'h608b;
        src29 <= 16'ha1d;
        src30 <= 16'h144d;
        src31 <= 16'hfa8b;
        src32 <= 16'h2201;
        src33 <= 16'h9fc0;
        src34 <= 16'h9cc7;
        src35 <= 16'hc6d;
        src36 <= 16'hd935;
        src37 <= 16'hb6d3;
        src38 <= 16'h865f;
        src39 <= 16'hfce1;
        src40 <= 16'h6555;
        src41 <= 16'hbbf0;
        src42 <= 16'hc9f6;
        src43 <= 16'hf211;
        src44 <= 16'h9cf8;
        src45 <= 16'h4c57;
        src46 <= 16'hd040;
        src47 <= 16'h7980;
        src48 <= 16'h6a7c;
        src49 <= 16'h66b;
        src50 <= 16'h6391;
        src51 <= 16'hfe88;
        src52 <= 16'ha486;
        src53 <= 16'h53c8;
        src54 <= 16'h5700;
        src55 <= 16'hb56a;
        src56 <= 16'h830c;
        src57 <= 16'h6b40;
        src58 <= 16'ha335;
        src59 <= 16'hb9e4;
        src60 <= 16'hdac3;
        src61 <= 16'h92bc;
        src62 <= 16'he452;
        src63 <= 16'hcce;
        exp <= 22'h20048b;
        #1
        src0 <= 16'hf785;
        src1 <= 16'h2f38;
        src2 <= 16'h61bc;
        src3 <= 16'h2a2d;
        src4 <= 16'h715f;
        src5 <= 16'h76c5;
        src6 <= 16'h72fe;
        src7 <= 16'h512;
        src8 <= 16'h8903;
        src9 <= 16'h8e93;
        src10 <= 16'h7edd;
        src11 <= 16'h11fb;
        src12 <= 16'ha069;
        src13 <= 16'hfbcd;
        src14 <= 16'h1223;
        src15 <= 16'hef8d;
        src16 <= 16'h9522;
        src17 <= 16'h3430;
        src18 <= 16'h81ac;
        src19 <= 16'he28a;
        src20 <= 16'h134d;
        src21 <= 16'hc7d6;
        src22 <= 16'ha5f5;
        src23 <= 16'he89d;
        src24 <= 16'h4f97;
        src25 <= 16'h9f8d;
        src26 <= 16'h60d5;
        src27 <= 16'h87f6;
        src28 <= 16'hddfa;
        src29 <= 16'h4e79;
        src30 <= 16'h7622;
        src31 <= 16'h3f49;
        src32 <= 16'ha3db;
        src33 <= 16'hd3cc;
        src34 <= 16'hd748;
        src35 <= 16'h3f75;
        src36 <= 16'hcc02;
        src37 <= 16'h1079;
        src38 <= 16'h72b;
        src39 <= 16'h55f2;
        src40 <= 16'h3fa0;
        src41 <= 16'h16c1;
        src42 <= 16'h8836;
        src43 <= 16'hc4d7;
        src44 <= 16'h3a52;
        src45 <= 16'h3e4;
        src46 <= 16'hda42;
        src47 <= 16'h550f;
        src48 <= 16'h31f4;
        src49 <= 16'hb1f5;
        src50 <= 16'h422;
        src51 <= 16'ha45e;
        src52 <= 16'hac55;
        src53 <= 16'h2b2f;
        src54 <= 16'h8fe8;
        src55 <= 16'hdbfb;
        src56 <= 16'hdc;
        src57 <= 16'h955a;
        src58 <= 16'hfc7b;
        src59 <= 16'ha297;
        src60 <= 16'hb137;
        src61 <= 16'h2a47;
        src62 <= 16'h5a94;
        src63 <= 16'h45d8;
        exp <= 22'h1e042b;
        #1
        src0 <= 16'he104;
        src1 <= 16'h9b1a;
        src2 <= 16'hc06f;
        src3 <= 16'hdc82;
        src4 <= 16'hc626;
        src5 <= 16'he023;
        src6 <= 16'h2376;
        src7 <= 16'h803e;
        src8 <= 16'hc151;
        src9 <= 16'hc0ad;
        src10 <= 16'h52d6;
        src11 <= 16'h702d;
        src12 <= 16'hb6e6;
        src13 <= 16'h9c5b;
        src14 <= 16'h1214;
        src15 <= 16'h9841;
        src16 <= 16'hd2e8;
        src17 <= 16'h22e0;
        src18 <= 16'h56e5;
        src19 <= 16'hb7ef;
        src20 <= 16'ha8;
        src21 <= 16'h2cbe;
        src22 <= 16'h1eba;
        src23 <= 16'h5280;
        src24 <= 16'hd1cc;
        src25 <= 16'h2754;
        src26 <= 16'h8a13;
        src27 <= 16'h5da;
        src28 <= 16'hfd74;
        src29 <= 16'h27ec;
        src30 <= 16'hf17e;
        src31 <= 16'h879e;
        src32 <= 16'he631;
        src33 <= 16'h88e7;
        src34 <= 16'h4dd1;
        src35 <= 16'hfef0;
        src36 <= 16'hbb8c;
        src37 <= 16'h3743;
        src38 <= 16'h9e8;
        src39 <= 16'h3a62;
        src40 <= 16'hc2a9;
        src41 <= 16'hc577;
        src42 <= 16'hc415;
        src43 <= 16'h3504;
        src44 <= 16'h10b1;
        src45 <= 16'h23b7;
        src46 <= 16'hfd31;
        src47 <= 16'hea1e;
        src48 <= 16'h1dd;
        src49 <= 16'h5d0b;
        src50 <= 16'h668e;
        src51 <= 16'h439d;
        src52 <= 16'h8234;
        src53 <= 16'h47b2;
        src54 <= 16'h42f4;
        src55 <= 16'h9e97;
        src56 <= 16'h2c88;
        src57 <= 16'hf59a;
        src58 <= 16'h8f73;
        src59 <= 16'h42ed;
        src60 <= 16'h2013;
        src61 <= 16'heff;
        src62 <= 16'hb98b;
        src63 <= 16'h7c34;
        exp <= 22'h1f0e21;
        #1
        src0 <= 16'h8e71;
        src1 <= 16'he6;
        src2 <= 16'hf2a9;
        src3 <= 16'he83;
        src4 <= 16'hedc5;
        src5 <= 16'hd2af;
        src6 <= 16'h8a01;
        src7 <= 16'h4490;
        src8 <= 16'h5afe;
        src9 <= 16'hf17d;
        src10 <= 16'hbdaf;
        src11 <= 16'h7d7c;
        src12 <= 16'hdfc7;
        src13 <= 16'h1b30;
        src14 <= 16'h8926;
        src15 <= 16'ha185;
        src16 <= 16'hd4ec;
        src17 <= 16'heacd;
        src18 <= 16'hd15e;
        src19 <= 16'h818e;
        src20 <= 16'h84a7;
        src21 <= 16'h421e;
        src22 <= 16'h55f2;
        src23 <= 16'hef63;
        src24 <= 16'hf290;
        src25 <= 16'h653;
        src26 <= 16'hf785;
        src27 <= 16'h6b34;
        src28 <= 16'h1cfa;
        src29 <= 16'he188;
        src30 <= 16'hbd54;
        src31 <= 16'h49e6;
        src32 <= 16'h632c;
        src33 <= 16'h34a7;
        src34 <= 16'hf941;
        src35 <= 16'hc3e1;
        src36 <= 16'h8772;
        src37 <= 16'h226f;
        src38 <= 16'hbcc2;
        src39 <= 16'hee83;
        src40 <= 16'hb1fd;
        src41 <= 16'h297c;
        src42 <= 16'h2bee;
        src43 <= 16'h9485;
        src44 <= 16'he4b6;
        src45 <= 16'h7fdd;
        src46 <= 16'h29f7;
        src47 <= 16'h7c5a;
        src48 <= 16'hb68b;
        src49 <= 16'hb2cb;
        src50 <= 16'hd687;
        src51 <= 16'h9527;
        src52 <= 16'h6a96;
        src53 <= 16'hbb9a;
        src54 <= 16'h4f92;
        src55 <= 16'h2545;
        src56 <= 16'h20f7;
        src57 <= 16'h3a06;
        src58 <= 16'had39;
        src59 <= 16'hc28;
        src60 <= 16'h7ff2;
        src61 <= 16'h81e;
        src62 <= 16'h959d;
        src63 <= 16'h8dec;
        exp <= 22'h21cdd4;
        #1
        src0 <= 16'hcdee;
        src1 <= 16'h5cfd;
        src2 <= 16'h9648;
        src3 <= 16'h849b;
        src4 <= 16'h16dd;
        src5 <= 16'h17b9;
        src6 <= 16'h76ca;
        src7 <= 16'h9d93;
        src8 <= 16'h4e40;
        src9 <= 16'h5cb7;
        src10 <= 16'h5668;
        src11 <= 16'h1340;
        src12 <= 16'h262f;
        src13 <= 16'hc141;
        src14 <= 16'hddc5;
        src15 <= 16'h208b;
        src16 <= 16'hebfe;
        src17 <= 16'h515e;
        src18 <= 16'h1724;
        src19 <= 16'h2028;
        src20 <= 16'h42ba;
        src21 <= 16'h6cfa;
        src22 <= 16'h9dcc;
        src23 <= 16'h9b32;
        src24 <= 16'h673f;
        src25 <= 16'h2865;
        src26 <= 16'hd615;
        src27 <= 16'h3629;
        src28 <= 16'h3e;
        src29 <= 16'h97f1;
        src30 <= 16'hac06;
        src31 <= 16'h6e41;
        src32 <= 16'ha205;
        src33 <= 16'h7d39;
        src34 <= 16'hf200;
        src35 <= 16'h1b9;
        src36 <= 16'ha639;
        src37 <= 16'hcc2f;
        src38 <= 16'h9413;
        src39 <= 16'hd146;
        src40 <= 16'h5bc;
        src41 <= 16'habcd;
        src42 <= 16'h8a3e;
        src43 <= 16'h9ad6;
        src44 <= 16'h8a84;
        src45 <= 16'h7756;
        src46 <= 16'h10db;
        src47 <= 16'h94b2;
        src48 <= 16'h46f0;
        src49 <= 16'ha86e;
        src50 <= 16'hbd29;
        src51 <= 16'ha596;
        src52 <= 16'h42c5;
        src53 <= 16'ha433;
        src54 <= 16'h44c8;
        src55 <= 16'h96ee;
        src56 <= 16'h3a41;
        src57 <= 16'h1748;
        src58 <= 16'h1fee;
        src59 <= 16'hc8e3;
        src60 <= 16'hc6f2;
        src61 <= 16'hc26d;
        src62 <= 16'hc742;
        src63 <= 16'hd252;
        exp <= 22'h1e09a6;
        #1
        $finish;
    end
endmodule

