module testbench();
    reg [14:0] src0;
    reg [14:0] src1;
    reg [14:0] src2;
    reg [14:0] src3;
    reg [14:0] src4;
    reg [14:0] src5;
    reg [14:0] src6;
    reg [14:0] src7;
    reg [14:0] src8;
    reg [14:0] src9;
    reg [14:0] src10;
    reg [14:0] src11;
    reg [14:0] src12;
    reg [14:0] src13;
    reg [14:0] src14;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [18:0] srcsum;
    wire [18:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13] + src0[14])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13] + src1[14])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13] + src2[14])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13] + src3[14])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13] + src4[14])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13] + src5[14])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13] + src6[14])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13] + src7[14])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13] + src8[14])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13] + src9[14])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13] + src10[14])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13] + src11[14])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12] + src12[13] + src12[14])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13] + src13[14])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14])<<14);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1ffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h19e357cd6167640c8c165a8a47aeaa645797680672b720d8cfc5acae3;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1cebea1ba8b4609f336ad6e56833593be1c39b77a0690fa14126e2cb1;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h10b85d284f0bb97cf0eda758d0b2285a41f10b9b3f12362a8e8171cf0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1faadad0ac3d1775240a0d6109d2c3a6e83341681c34714948819146f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h7e76fa6d94d478a8ce685cf3273a7a9becdc4d978a9dd2e98242661e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h311e33968536d084286565669ea0fce042ccbeaafebf6d16d9f602a0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h154ca55da8ab796704eec6b721778f32d2e6ec2de5d3c7b63248e5ab;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h6d468cc9ba0051cea255b44cbef7816db4d71cfdf30bd976c22f023f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h191d3c91836e2664948698fff975dc7705be7df886617b937fa245817;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1258e834aeb7c2994e8142da675d4f7fe63fd8d61720108c9c1ae9a5e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h65fc79313218b9f733de15b9caafe0c65c3bb817a1367776bdf141a4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1d4e82ff5258b794ca4fe60173dbaa88080d0f85606c61a74e406b72a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1690ff9a74ade307165774395e9dce2a19ca8f47036d08879864f1fe8;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hef39f410eb63681a513aebf773843441c23a962447fb24e5b224364a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1d1d7375bf739bf8a2b7d5a598a579175ab9f5288fb1f201ea9ced87d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1a0cead006873212b0abaf540039cd120dbabeafd28c424273fdb0400;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hc4fe7a6d145c601da3f67759cc664d133eed2544d0e1df864b083b58;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h47e2ccd30e9f19a5fe33e3b0d85600c98583491e8b97020df8fc5cb6;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hd56555181ebcd2e3c340694e1027d9f51b78127c7fd8f570f511defa;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hb611cae079b1335b6f33c710b94ec0424a571f643820a3d2299d1832;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h102c94218e34b662c5028ee227b29761b22c0223731e0e7ffbafe5f8b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h843ce34fe6e4035d920521deecf99b32ca803a0e761eb0eb84c51d7;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h169f88814698c8e5d7a9dd5d2bf65bd1b1997c416f8530239e1f3e1b3;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h138f9e1daf440231720b7cc93196b0e2f41f63d7f3c24ff1801b043d5;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h5d5acd454e37082d99532388307c60a1f4c3950ed7cdd1afe00c6c73;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1ce52c9ec069de8c045f02c3f7f69ebaa3248833410e63f2eccea5d8;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h19960209d92e099f991d738f9d4bd4b9e1bdf633e077196729d35c535;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1a0551678407dd90d05d6b3abd80278aec7007d79c9dc4dc4e47ef2b8;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1dd6b97919a51a61aa318c3bc31757fe821cf9df17127402e89be48fc;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h10b63c9feef23e0fa1d31f2e52eafab53b526d9c624fe9582a6a97d99;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h10e68a34e9baa2e50c6f950f33ac86b0fa1ef96a42e009aa736cdbea;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'ha0e1a5d115e72291a2dbe0b36315d0dfad4ca8a9138b394f766a9efc;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h9b02cb3d263a56425c3306aab611fb2998a3a0eb1ffbfe745c2fa024;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1063d75f73eabd8ec881c58ee45b51e9d2d1712cdd155e92c18100abd;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h17d4e3b61e6aa9efc635f12b3c20febcba38bedd718ffd7b16a17d699;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hbed527aef868439ade80186666c0fcda4ff1e94eadb8650b1f3ecfb2;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'haf27cff46a1f32a70d4fa0fbff3787665a2bae63e2e5fdc052689127;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h155f5cb35de650e67d349f92d94055b7c62bfd138cc8ad13bafa2ba6d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h107965976b728ffaecc8ea318e9afc28b11a6f002dfb2848d4d97ad07;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h18fb2a9198eb723864192cf43152d9f9943a1b1d20a8eaa5f98ed08ca;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hc8e3518206644d06bf5cdf297b2e38100cfd6bc29b0dfb096d55142c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h9f81ac25b3a2d8871c9aa0ddee05a906a65a4d0602a5d15e782608d6;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hb97c352eb252a9016f8f6ab056e81a6224d45ae883f724f0a5c507f5;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h120d143abaebe3a92a8ac9366996f9e95d83966b012fb7b7addef5067;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1dace9b8c9f3e72229abf70f370b0ca17545ba19695ad9d837b049211;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hc23e151729722b36d6878c4319aaf79d88380f5ae541e994db83c4ad;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1e491d2af49bf502ef281289d19d7576f1581700a742e089ec3df6411;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h13d9915fd2e0aa367a0210a85deede1858a5cf84a3c11774b0bb7aa2f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hf3146f5497b5c2b4c5293b12c68c8ceba64941bf3ecf51268ae59155;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h6d7fa2111f2c1e37c092d2c3051d0050daa64e8750469b52c049fa02;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h93d08b7947163d893d445b4479550a81c72e7049ab2ce9773df2be67;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1d055a11fedbb0ab59f5005eb8a3bb3b507a368c54496d69119f69266;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'ha48e3a55234e2682ee8c130726932e06f99c08c22bcc5e7bb58f6732;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'ha4a1e792b2561e74108b710abd66812e26675f3460725b9a7766d312;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1c91024a315845deb84256b4b8a2b1569126c1aca59cc41541c4c97a5;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1c0ae992c189d592495e1df59bcbdc8b26bf16c848592fc00ef96a7e4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h12ed2c06991d7e48de6b0307593982b43d8739e669f8da23919814b63;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1fac181dacd00e35310670ba90322bda29a7d6c3364d3f9951d5bba96;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1f81d84be4cd29c62c63f0acad95eafc6f1a874e0d825e46a550b68b4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1a435764044d739b749f61b08726184cdb36fccf5a81f82198148c44;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h12b259ebeb4951e3e0f5c416b9ed911e4c28c043a25924c31498054a3;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h15f52b78569ebabcb093695362e6da130408a0772ffded7b5f1581149;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1adb94985651c1b2aa4e4449156f85d518e633e700f5d8352bd3f561c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h18d2ab34dfe383a52303d46b979ebd179fc4e111e3e915f468d1d2138;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h6a822c278ce8a401c7b5bec85fc9adf60bb5e00921285df23fb7ddd6;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hf2c7a6f906b177ecf9b03e4664ae7b5dc9b987bc49e785a63b8bce05;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1820dd5816c544150dc94346aabedcdd99c58770ff402d8c26a09ca5b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1470cf08e16d363a12f979d278c86491e2e2d112a3c3bbef152085730;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1e1fc6724d3a7d411934ba4d0d5470117b86077b5d88f63411bc9462d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h6a56ad0eb6f797fc8a17f118cb681b0dc0fe51c7907b95d1c64edca3;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h2dcbde52f36cee8a14d9012f30075a30f3fb26b88b36390b79635216;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h21760e79e44592f6bbae26e76cb3b2ed0ea3fb8dc648a6d9ce17b5d9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hb86b131c782df4f3963b1d3a488a79cd93c9d791af9ee49f44c07bdd;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h45c7a9927e6c8924e33fdfec32c94598f8fdd5c4118376095ceca25b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h5a2f4a7f1d8263b72022b74da9b67720cd6f293f65345ca1d04ac85d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1345e7342e0d1746885fef68d8c4f02154dbd9607a5abae3fd50ebe16;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h146a79f15956e042e29ebaee814edbf8c5d7bef246f7ce06ae01ddd7c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h19d71c68939bc8ce3e479417daecc46969ecb2c70d203dfa713b1439e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h10423352094787da676aa2d83758c77712356b3453de3d1b43b532b54;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hd359b381b598b578d2e5000622eaa835e4ebf41a3df31610f2e47dca;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1abdac7d9db19abc46011d12aa61830ba63154780d832939de3e00a91;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1f7f705763d8920c5b47524454e355ba6018f644f6f2afec788e25002;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hf8eaa8ef0ac33cff21e536185d1ea21a6f5118a26a5fc14572e5be89;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h3b801055def8fffecf9b9aaf86c7c05d13b51dc7bd0deac286d4f2f0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h557fe12df951707310b05f8036490050508ef6ac9999d331cc72c9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1476a2e5845cab51fdd2a121a47ede0b0a49be999a5a05f99e325aa65;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1a92e3f70a4abcb9a9a8bd8a97209b0c9dc732b85bc72b16025440921;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1225606810ca1520b87c4a62b9b0349ff69943eea9ed6e0f365e117f4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h190a34a439fc96f8c086ded0e437501ccf71d46909a253b0cc0eac19a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h14f91abf8df5d3bfef46e14dc7eb12d1dd6a2c5fa83d745b6367ee6eb;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1ff613043a42beee48b8868a9b06426c7cd81f844fdfaf2c09efec215;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h126c63d9a9563c20c41fa56c9f26a891c088c24078740b82bb1f72316;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1351e77086e3c894590c42f307cd52e2bcb24878e2411f942df6f18aa;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hddf9fcbb4b8c4ed9af6e3c24241897e9c20a517c4ea5f6f440d8e402;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1f211ea39fc985e6893601565300155d7f18b6926d8bd124e90719dc5;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'haf4c1695ce63425452111171d2f6fa4846cb74d7cf17decf6d71ec42;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hfcded88fd87ae412ec00413443fae2ba04d4463e5c5b9524c44296c6;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h31d1ee14d2d71d6f407e41229c09276b5be202dbcf117e33402f569d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h13fdb971b108ad456ff092b35c8908b2557ef607911f9d9f829a68bfd;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hb152e52eb7396180343ca03e3e8847d894ac2f78d53236e5689579ed;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h102a8b229242b2ebc3829ef8f1ad608721a67a2e2fb2f18c5f281d4f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h9dd37bbc203db0a1c138c9e02747c7e42787765a3b1c8308e2d4a108;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h9c059262bab448cbfe114132338fb0f124ec78102f7b0e6ec24feea4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1147521e4108944c5f838b899b511c1fc2bd39dbd6af947c34cc364fd;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h2f4684c6e621e82f08f2e0df5f1f5cbfec6aba9389580f7522cde10e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h43ca6e25b5ab007ab6475cb5da56a09e61ab7ce9ca67407c06dd85ed;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h821468345ffd2f2ed2d9f8285ea614ea896b3262c8d72788a08affa;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h74c9fffb3d595849119c08452bf1018dc8f28e4984dde8313b3ede6d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h12527bbc91a28e3080072d31b698d5663e696e07d57b76cf112e89dbe;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h197f15790a32dc711dd6dcb33a102c9bcef87029ec2bc6f3d7d6ef1f6;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h12b8ceefd39fa7325863b4f65fa235ed34808a30e61f17a91018b09c8;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h6ceae7f0b1c6d616ddd3299d23d69af7756719094eaae07e34d7c9de;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hfa24bb397d79870e88322c0da4815eb97cdeaecc71bef47b903f6ea6;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1307126f1be1ce4a7b409a989d285c36dd272c6f21352621d8e941f5c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h125e6da42fb4fbb1b193970d7b0bf5f87857e4e70572dd3b760c2c33d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1dd7278d46de9fcd01ea9efd8c72217bd595d4525420d85c82c5ef122;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'ha31ec1e61bee25b3d7cfcd4f7cc3bf45f392979793d7ec8d6a6c5153;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h8381b878d710d44ba0e3e1d37a36ad929b2f60dd9a5b9314c6c336e4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hd6474fc740ef3214e6c339eb8a0e134c0fb6d74bd3d867f1c292f02d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h129265fc0dab21d3dcb610ab1d31fe5da39e00ff7c715cf90e7d55341;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h602b8df1e303f6899de02a605b2deb9276be4d9b97cc3830a292a1c7;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1f77c6b1bbe0edb4a4ba1e262477c08174991c303f95373adf089b38f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1aa6aff7cc1be8b58ecea63236d04eb24dbdc2386fc824dc14e2f855f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1eafceb44d2e63a32f7f130c0579f2807ce6d97b122cefb2680cfd5ac;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'he319b921d243d23e1bcc650b54bd3497e2dac13a24adb7fb539a64f3;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h762e83f2a02c93c9d5af0c1d447364b9b5231e0d54133382c06ea265;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hcd73adfdb5fa5a035e0399c777fb5da6e261969a79ba7a3494a3c0a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1959a833deaedacdd912250d0515b76ff325280c6e1ea50d5ba00685d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'ha3f54f5f5a4ff0d78da7c05fcf02e90e0856421b0a6b9040dcc27df0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h80c1066ca9a0cac87548953da5d2eabe486e3dddc953204163653eea;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h7deb00c6a71505823d4070e839bd17c83a3a4bcc1948f2c7d2a6382a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h181c9ac61d382ea5b92750a9377a281c7ab2e98182369ccddfed0c4e0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1511dbb709ca08b0a166e8cd9bf44e139aeda0754922d3ae2709a2ef1;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1aa51122af706563a3188598bad744edd4c91b18b1ab251d9d9a72283;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1a0f580ae782187ae854c9ac866fba9a458cd5927d43d60958407d696;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1aa8bebef651e05d1aa6d674d09a7a5d051bdaaeef3cbf27994e895a9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h677e76a116bdce2731f6b3810a5c21efa0b9321288cadf71f9840a4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1db1f02048cb98868f6a6b4cce2b9af887cf4773f9fd73d3971b52b91;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1dd2fc95c67fca713f4e46b877c78e7d2028a7242ca284d1f37613060;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1107fd8e630704e28ebd3a8465ccd627b323f342d6e3635c9d66ff195;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h982e2a634a0a6d9637b96cfa40cc73a8038e19cd110b8e0778329f14;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h11d528e237aca6d4c91f547a4d79ae0976727068c276fba8097443f5e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1c0c079bd6acd078f30883f281acacdb9b1e9c7b58a91cfb2014bd4f1;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1bbf6878a6aae674c4fae1fad501a0e4cb1201226f5e64b5d24674afe;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h178fbb9cdffe5d4d913271b4460c21ce2a80f8aa9457790f1a98ad221;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hde15a11d25f155a39cefa7e20a486853ead3176c4daccf2d7da3ff9b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h8ec7605ef2758f1b4fd4055818a0218fd4d91996e090d349dad36c88;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hfabbee385911ccb4be78c5024aaed798b2bb2465598ce2cdcc4e1065;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h193572811b62c865c827d7854a6f771261c429c32c1c6b9336b4b5ca4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h32c7f9b0ae6442b5197774ad93d9a6695ff7bb805b3cbc40b7df6d8a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h17ed93a6f6de082b6116d6dc02d8397fa33a6d928a7da5e88810b99d7;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hfe7df774d2c6f6eb3981aec314c3151dc4f61b11beb353fb7174f0d5;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h16ec75adaca62cb76373cf04fae0b0c469b4a05ac5a96b1dd8fece01b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h10730684bc2fc527bd4eec357e30e78669d941529f7130c7bea70238d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1bad65d23c9b879028ff7011b62a40d7dc2b5b7e0a0d5f9a8a4c0b660;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hffbc4cc44fc15deb8f5b18d4a90f6f103fc6fb66a6aad0131a946cf1;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h89595f27fadf4e259755e1e4a281671ac861fce0c2f2faaa058dab3e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h2790e6e0710987dafcaa3e3b88c36b09ed7e0ae2e55794f93587eb0e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h100d3a5c939efa99f037e9ed310bcd3a995f10d672456ebafb9669b22;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1138d8c2fea31a6d9766b3c90d7a8e6d2d9b46040f138190b29253308;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h13f2256d459d9236f9ddbf565bc96347df0d3344e846645f941e1ac03;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h84b10ed100fe48a092c70ecb163fd46ce2696e8d023e468350bc869c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hd2f7f86ad28f2758af0fcb031392074ba714bc11e1651957b1e2b8a5;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1e26edf74159b08792ced551dd7bd3115f017472687c67ab25d0fc166;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h11ad8204c5852d0a6aff26cd9cb6f564b5791599166359a7410954c39;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h18e561e45030635adb023d596f2470370963db902bf1805c33d857f6c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h4523bf0e2deb5b783ed285ad7f63c84a2d0e251078e2eb78dea19278;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h19e741a9e9ae59bcf7ad91a9d275099106b83cb26c7f5825d4b4b2cfb;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1f457110e7e6fb7d22315241827d9c4c0a2777ba8139fd07c75ee416e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h3c3c17be83ea877021f643645c7e9aedca6c065940b2e91fc56a8252;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h115694ed03dc7732d927ae972fe2f5ed36453396c797b3fdc27c77a7d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h475cf49535c3eee84696dabd736d4b913731b55456c154bd4d91fed7;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1cf3cf3517daeaee515abe3eeae231239e11557025bc34ade413d279d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1ab414a84b52c32c7f78778b8a3771b33ba0d7b5f1ecbd8a50674ca6a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h9520f99e69620c76678e3559967e72eb48798b314280f8f4aa3a4ea9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1c43255f1511b78aa2084d0b5f21df248902bdee0aa8c7af82372173a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hc0601dbc86d395e0a0511b006446314fe0162ec1d9fcd06778049c18;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1b0b413d61b010ba276f5d312404e1ff6d0f8beec38bf302912cbd347;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1b477db160e106e61609a4b3f4dce67ff7d018e4a9218fbaef8a12d0c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h10ba53c6b5b7309a9becd5fd7200aa12dc7845fabb29137d83a312f3c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1e35f27dfb7cd5952738a51898b7224071f06909d4360c480aa35613f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1642069b4b0f39c0f8e7004b705b4b75f5bd07fd312ac0d675134efcb;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'ha283fc63b57c9adc8df5f044314e85fc2a3d7418eb2c904cff49c387;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h2973cea2c3945e5499aaf53c0eb8967a65a9255a19359466955d308e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h7e562d71147f8d87e7e0628b4d6df7c6f8ec40e699a73030bc61c056;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h135df826cb18a2bd3c0692a32dc3f4ee7402337f2c418eca11d539a23;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'he5ed5d7bda532048354ee7e747ad259295ede1129c14891f7e1eed3a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h813f4333c2347073a459e725cd0ba200fb96abcb6a14c862b1f9650c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h78490ae8e1608abba97df77624a724ee524a3ffa7d373cf91c6f1d13;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hb644a24dc4d40e6b1010d1cd4c5b39dd1e3cfe2339005e4baaa4c689;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h9c29ac7c8ebb01728d7420257b434a76164501db17d412e6aa13e270;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h9fa3ad0feb14457bb1f4f080e2b42dc4bbf6bcefd1e3113ae5789868;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hef9b0fbb02c51f55e364c0d14ae79d7b570267b1ced83259804aaa8e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h17080d30eed3b5db602e2abb7d617f6f65746bcf641e44c31252e0b43;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1e7563b89f2c713dc60e4e34696d3454ce8b612cb0b09637283698bf0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1ef62ed95f9981db726a0d8a3e73a3d72d64d2bcb1790b52467a9b636;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h137dc071713b4979476aa5a9bf34ed77fb7fc193bcc6e0154ae80bbce;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h82befe243c226a911de3d16c876e32eca99e5103b8115848dff1b1b3;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h3cf09d5a6866b2a31b646ff41d564e32a11a2e6567a9aaf53a49aee5;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hbaaf779a80de40a1c3179d815e22ccfa41f6399dc24ef680611cf9ae;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h12296a7196fe6ce0dc66c9423269f416a094d178df6ecb109186fef90;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h149d25ff7f009a66213f1383d472792a7b7d4ab9a07dcaa03ac844479;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h858ed85cd6767a9b95eba7d9993ff8112e5ed345c15282edc01549ab;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1d9971cc1edd7229f9bcd0d365ac97d0cd4d9c842d055c124ffa518c4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1a642df59ce764e0387a66a7b7b54790b0714ff163f5f7772a863a1d5;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h156cbc14d1e404d90a45131b347f599dd1616101d199403b408782f78;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1ee15c4368972b5cf2c23c30a310910b31677bfdd767b4f71e870ba2e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h13c9f521c2c04e231f6fd18b3cdcb686bc3000c2d24d0f324b8a6c082;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h186e57038452c4ec17523cd9f884ad8c97d33a05d955587ec965e5988;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hc7b7188cae410b1fe7f6986f73c8a060748318c2e157279697b8ec80;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h134bc598c5f7a828c42916d5127cc5f302aa9f932b6277a1a1dfb6660;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'he37fdb21b06aaf616f1dc7b777aef5c1e2c68685f7d04c6c8ea300f0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h5ae3a53158ee95912eb18c66b4462a0d291030f15d4a885823598c20;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h177449650a30f75695d70065395d2d2a9fa196e367f763864ae4f0cba;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h34bba369fdb92e6f87bb6855141db4dc21cfaab5699d000c5c625eb7;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1b77122ed4e2dbbd5952646dc9fb3a0c1c303dccfc697a7c3c9d9707;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h139df4e50e545e0b161174de0ff61b55ecda6a2c3b7320853d0b37308;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h70e20f25c3fe15e904648a5bf033ce7cfac5bd4d855fde27e3c62e8c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h176ec69a9ba814004c9349275949456d85ca5f04acc35795f1f34247;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'ha587ebc099f3f1a7e9bd54f9f275aca212dbd125cfdea5aaf2760808;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h15a791bf02ac1cf8ee1bc694baf4ca17a0f5bf3e7800ba4e437a0ea47;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h83ebc1f97f69cd6e4d2e3b7e81c13bda76fd1d43a9f17ced9c12ddb6;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1fd012fe80b31516302b56aa2b98b4ceda18b809b25b5574150578d96;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hd92eefd997c2a0e7ed55c6448338422c7a6e8043b3285e890fde79b7;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1bb76ef3e85fdaf27e5897be7f8ff0a4d0235723c21b3aec526291ff1;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'ha7f929b62decf562776a5505e4e4bf11201cb2cd9e10435153f01de0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hef5748ec9fecda7b3b6ddcf46b7a7cbbfd701281a697b93a33a7504d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h15f779e90c19c413054162b2f34c5523a7903d5f0a72c666ad91b462f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hfefd0f63483c31088fa6e90963e47c0154555edd55f1ca3f1e074fff;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h11160824447dc6645941e1146fcbc2ffab4999b13aeff1d90edcd6959;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h2743e15c248283fcc64444c8e1ccb6f8ef74660eec56e4e384425098;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h167b926a38bfe7ecd0dbdfed4a5aac85f2432eae41f7c7e665f6857c4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h14a303a2416b0c27ad93f382688928b61b808ed0a795d38e0ab748aa7;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h213cd08648e7a809dc5c170aecc1fac1aa3155c482b29c3921d8676e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h2ed6a81460acc15ae8d87b1710f2bd86dd64b36e692105d3d9578de7;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h178f2659157344dbc6f0dfe9aee1237387aaab545bc2f6cc88f348dda;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'ha9beaa21885a4a377c3754eaebe8f1926b2f238ef7f804cec49c5079;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h85ec7a61ac20af470a0e8d2dd6a21667acbfd85b44cc13b70563bd14;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1043da113c2580c14e977ccc1070d41bfd5c79f0d48719c05a4e54449;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hfa53313967498d1c0cdfc66434d9c64f427faf0270667b6c80671e85;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h9579aa4bbdd6487cd36e62035ec994b129792565713d3ecd212f3566;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1aeb5de0aba7f52861557292b9daa576cd1f87714e3efe4c36f95b06d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h30ab2d0c25de56dbbcd4666d69fcdec7a27bd1bfc7899caee4835577;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1023b57f16a7bef3bb1ba7d2b7b3a17f9f82ef74ea2341f204480d565;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h175a587222d327854461547b5dd4b18382f1a427736bfa41ae499871a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h130dcd0978fa477d970161b00b231dc8ded17dd66e0f9e04a2ae8d73c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hd4e2e5accf9871f37f5bfb91d21e71f0485a869d06dc6cb7d5cf1b81;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h18fb17e401b1736df11c654a7a5570aa5ab7c7c966a4e153fa7f3dfbe;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1a10f9c51b4b60b134ec30155dd424a2f39509c4b0dd238bfa0aa3a24;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h6bb451dc772f07abcb8e6a5f2d6a13e73c871a2845bad8864c489dde;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hd8b6fc60e0060abff5d7f7e0985be2f2ab064f11c82f9d4bd5e84447;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h71969940a72c4de3abc84c1c83c04d11419bdffbd138e357d19c9585;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1ee0d6a8226b47988fc359c818335797a5a3c596c0af6b374bbe2facd;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h16054e93ef9d21fc9dd452048084253282aebf9f7a835f7c93ef103f5;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h8d4d5a22100b8eeb830cc810f0d3579d709e4671a341ed6b660e6460;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hb53ba15ee784b09fd7e1bd5bb7d4b511fdaecf1d2e19e0a29a4b10ea;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1e5553164efd695359dd7f4d6157c8320b5b3d92b8416e25c941e423f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h171b2a2e5423c797651d8e8c37c85d2458a5611c137cca4fbba3c58c8;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1d8f7fa84622a71fe3f3714c70dcd5232f7bd7997cec4b9e1dc285084;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h2c0d6fb55d091ab81e4a6f355c82c87ef66e17cc408ef5842708c81;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1a92b52f448695e85ec2288987b514ef03c8f4dc096d29e4dd3b40557;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h136586de60800451a51c905c8c17b75877d092dae57b12c1f09902598;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hc089e889f5c298fb0099b5c97ad8cfd2c2097f3625d494ad03cffce7;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1cbf7a7e7305e30f262995b3f4532fb50ddd1d0cbb3eed2e00076e33f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hbacdeb32e414e9e3cfee0bed37a54c515b2a4fbd4aab403961f44940;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h80a26bfedf8f1400f30b0728b87cdbfaa2ff1caee065bcbd2fd3c3b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1db015562c01bc597e79652fff9e8761da74eba5d1efff1f0097c627e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hdf98e879c4b79541b9a3b0a33d6769c7e9a1d51a69ec67556b2b2b05;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h6bb535aea0b2d328d529cfc55ee2547031727cf1e233c7a811ffa8f2;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h30b631fe47e4f0c22bcede4fbc0c97f6c32b852dae726fafb683d709;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h210e445342fd0f8484066abfc1447c1dd96cfac8281a5a42264dbd01;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'ha4b966bfd69b400f9e55c5ab8e27e7e37eec353cada4e4d7240a4df3;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'had1f156e66bb343c5a96880f6f3dda902b0bb8268ad28ab291429958;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h968eecc39c93bcc84a71e36c4b9fada14f2dc679bf683e864483fd12;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h14657cfc19b2a021da7d83b84057ea40d921e125051c68e13a2a508b0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h14a43b33b962d5240b5d856260f29c2a7577cd3843160c04c1d272415;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hd5b17f55887b49521ffb90fbb563b34f7cae7213a2d8a22f4080b4b0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h3c40d4315563a272d6d9c09aa4249f53d4e66f92dab675ce45aee4a6;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h69061f86553aa66d67947959fa4ae96aa2108b970efffe1329816250;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h114b492ab1857ca651585af789b2fd334a849ca500814232aa03f11c7;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h114858a0bedfb86faf9f6aee7ba78aab1d42a15146074332273b265bf;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1f58c7dd25e9465e907ef99e83ae4aad267aa4d1d50b047333f75547;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hdb4c45d709d6420546b630d454b7c11054944b76a0c62448ba7ac54b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h9bddd9b4a963b1bcd8785b48961e47eda9664c8eaff6a41f03abb50d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1eb0a21f00cfc6533a78f85442c7b0c460c178ae771c1cc3093213815;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h66f4249eed219e8caaca9d904a855a294f8a4bebc79fd44df742bb6f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1c5172770a3d1a213bfa32a7e3dc1ff9182d2a46d5fe255a56a915173;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1f2ebb14f77a393cab5091f312e7cbd886b9ce1bb69bd7f732cda72c6;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1cc3be21ae28ad7664e151a78d7d9654309b07c3dc07a50e0ab71c28c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h5da07b3c913be123805b8ad987e48e0e893e3ce800e3cb8e76196bc7;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h8425dbb0f222dc3e99525322a57003570d17b922c0e72c4389621940;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h53d836580c55fd34f616910423851bfa9679c1e74b7cef18a8f1b916;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h18b12f2d2d023831df6ecc44bc48881235a0ca9393c1167b67d0c9394;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hdc3ab5d94790db1af99d993b60a83acb892b403e61fed83afb60326d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hfe898bd0c3fa2dbb621f8e9abbe9f1ebe003418e82fa63dd802ab201;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h16dc5063f88ab69c88ede27b3c5356f7819aff4f55e1d2165da36773a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h694ca04a48c263a60fc44065af1952b0f9fad220b46e3ba4997e0ff4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h2ea814c64c9aae72a8c2b2fa50a53947a20dc22649ccf588dfba5ec2;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1711322f1d897fc9addd65d396700457c9fdfe2d5623f6aa8a13c0c4c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h11948f5bdb9328d414ab8f6a96caa4d09e79172d7a9fb4d42c7db3349;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h12c3d4bef7184f89fa2954725ad744206a02ffce7faf2774460db6893;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h8fc8c91983fb75bca7c08ecf6c04b1d5d19fbf2b65ae8380dede2140;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hbc96ffde1e72fc370b64b00c2bc8860f0591d51b22ad9a3b88f597fc;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1d4de8830a4e5aad2169dbf0856ff2f6299541128da285e7b220b6bff;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h5e4b4db5de850ca0b62fece5fe11c45968ecdf593c2596fa5a8d3b22;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h8ed55a5efe0f1cce251b0d63cdc975cd426f10dbc4d3e6af78baf37f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h94a3a0124d0640b2d81172c7c543239a0e09a522addd1c365007079d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h47180f44e7293c15f4a23ddeb9da279ee6f99ab791815e28cc373c2b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h10dec74fc8e57023be950ca9ed0fe008bc886cc7a83cefc546314d3b2;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hbd2e750c27c29b4be5508cb07b4c20b3d0d179805c51b98e3f5f741e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1f334a719cbb1fcc53aa0a8a541e210271a0826d84a9169753bc4eadb;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h73c0099566fdf5d45e469325615a2c4adce4d47570420dd7fc93d7c1;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1947bc2c26fa9939449518b56d8ce7b987419ea28f4a5d7f6a0b825e1;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h13b285d28727fe25811d1e83bc263180c0ba957a6d7e700b210da680d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h11009f9224386336030eaf3ec2691c1d2c5ecd47018a315c73b59ef44;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h5014656577a536a8631afbb2c071f49b56646591d974fec3f6475a3;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h6df7e133f790b3549b0305b3d8fc2a576b0731cf9bbe44f35fbb7c29;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hf390fa42cd64893f3e9e49085d6747acb145390ebfe2e6011442ca42;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1dcb1c03daee9c0f954ac3793c642651b1257b05508d3450e6b790bd9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h17ada062a60d5c1a0187125b8435b1fee59744a5db9c9c3e5e453b312;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1a08ccbdc39a0e4538e70df883e59575bffe8ea6c8f09cffe68a93deb;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'he8091291ffbe3a5751cb5598451dc4836f3329c87fdabf35c413e0f7;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1fd5785b8b978fe448f2a85315b8c2bc78d22d374e0d93e69ad7a6cc3;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'ha7dd8c491e3fc99d811268cc128535947a78ed3802bb8201a586a522;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h182c2e1451d098dbf5ba807f4613329577cbff75591ac1b4b8523a489;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hdf2f8b6313b8d3ef3b1802e7ae633e027caf483f4c822ae17d30d7f1;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h184d656b54f0ad6c666478b6848c736710c82ff607c64a1ca699c2d1;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h34d65489af9f8e30b24fe0dd243a1c77ef71461c960b26ad14141fc6;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1c5e9e30f81630e39b4910267c556b611593401a92d28f4920921aded;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h172330204d6cad15ae28ae230b76dcb959cb3abb0abd49a8c20e5261d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h707f2ade90c7249b257119659944930c48f430ecf515554fe9111685;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h5c451abf2e86e5402c78a216d1fc7c601d92445a92ab1168bd9948fd;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h127b3bd7f6aa31d69eebc3c6f948b70fcb419a3db478bf08574b470dc;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h7c0e7214004db450ff31ceea79f90df1d3f3e0c4ece64a0dd8cc7443;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1bc859ca9a6d41fe443445afd148f883b61a238260de243a922c16a3c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hcc63c4578e1b607318752e5757794f0c1604e4374511b7ee0f50b214;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hc084f4f328f3bbc704af7f0ba437515222fa23beb3499ce226635100;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'heb15d86ae13365c3f48782c047247529c45060979b3ac9de4144abdb;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1d3bac0df0c5556dd206d324cef3c91f49c90b01a53aa31c034ae4791;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h10df731c8fce81b4d01c4d25f70050cc08e1147c5177b6409e40d709a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h6ba2f586426a37b3102e29c9ee9fe56a9a2adb2cbaf8a156d13f06ee;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h17017a95e9cd56405cfc609c9331c3b2f6e46affe7c234d9f02099d8b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1f878c749fc4871d52ec37b546c246efe9396d73562dbc875bdb6390d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h2f8b17b5546c32941e950681841287af3c7a101bc889a1a4db1a6bb9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hcbce069ae12a8eb3094980fb3b668f482b4d239049619c58b13a7f1e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h230816384e17bdd6809d15cf82b1f0814553908a2b62fde38e89ba3b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1ba725a85b367ceee215b37677c1e3adb71601b7cd4c350d5396a2d92;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hb2c04e3a6ffefd456af3d3fffef3263db7e6029f27f1ca0e5de940b9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h79f22a7d5caf038aea6e6f7ff688fc7db3605bcf7868b5efeff54d2f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h505b2fad2f9b81f1240ed958ff043ba65ccfb6850e32189f6793f334;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h191da661bc7736128769001739d0cacd0f7e8eafdb3803c5c9c1e4c73;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1250490c99036224bb78c1e4d99a633edceeeeae336c4b2e1435db737;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hff0d41c8d383aa9fe293e6cc801acd851bc885559dd7e0d0788fb2f6;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h11775eb614e571d7c61f60b1978c6a0c1cdd1b62054e85f0ebbba5562;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1b3e57ceb97c3d5e45d189a121a8ce16ffa22ef335207a9ff0d19bdd0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1fc034667e90a36d364b8637e2f45a847aa080951a7e724f5ff36bca8;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hab90d9526f4e4ec69a9c5ccac1d18b9a133aa4b676c30e8723627c4b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hbe2beed703b38c49bfa4880cea7105a570d682ffc433c3391ae64ae4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1fff0a0773bbf5633c1b6d5c0928ef9b8d6d63416ee2d221d544bb73e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1982875c13257d712bfc95201c52823b6e505491c56b084291732c783;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h158c60a47771a2400a14713eaf23938e896e00ba7852b131d75df89f3;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h74134187491ee8f3a32d80ec0d8605eee450811a125c4bfdc14cc143;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h18a995754236ee50b91969fedd6c834334051c3b93a24656d63260075;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h576b61dcc8db8a4db5bd7e4abd4908de5e4854e557069fa568c0e539;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h12ac42c09f0010f5ac3481db9a86c7b5f47b57836252bc3843f246b75;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h139f960eb5cc42a79e9f173e4336a4cd1d155ba1eccfceb1bf3084d2;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h77903d6899358c3a21c483419621f3f64e945f39fe93e5bfc0413b42;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h33593d9d8de155d393ab9aa7877b0c54ec2f6047f13410e600f8feca;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hc05c1d2d603f152ddf78f2b7f84f7e92c8640ae054394d5777e8f66f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hc9359cef0efdf474d3e789ba890eb9452d76a98323c395b5145dff14;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h115c499253d29b4c4fa7682deb2ddba8e9ba7be1e79e51cc9caa9d3a1;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1eea18f5f432a1c9f817850280ca31aca477eb3a670e20f1f2d74326;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1abce41903e0e44336c9d29b85ad60e9caca82dd99f979828722a113c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h13607b1ee68c86aaa72b1fb41bcd71d434eb549cbe7375a8a74b24deb;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1755183c9ee13c9c3824dfdce385f6e5ce6d014319e80d5b14994a611;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1b7266dbf0de2c82be1417ccfa2b5018c27068a9553d385c8438ab28d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h129b16e3a1338a0b62c93c5c968af0a0a371a84c100f09be57110e95f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h68c9a3d8b04c7afb0472091bc1784db030da16123bcab5a5561e0d39;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h59d9398fc6309416197a0d14d3e2d24fe8f2275c559c3a522e6850c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h13b0898fb813a044e3c789709a426f5fc6f19766d1fb4827c5e8380a3;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1b1c7d394b9db1961128f07bd42117f0c480d8eb09176c5395267cfbc;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hb2b56902fd5d329892b2d14cfa45801d59ce7b16ba08eb42b01b73b0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1b119175b43121f0f7b128e73814e99a58cd292740433227781dcdc81;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hda7049fdf0ba8136615f20d45e69d3be59836a884bdbb632deb0d663;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1d6bc4ba2844e642a0f7abb5d235803ba8acd2b4f5bc651a02f7afb9e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h18cc50e6fa66f6a47ff9431f5d65b2d42def4c5e6dc794d24db9ad016;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h2cff5d9a49a3814fad1aabe203337f0f16b9c0975d4f7ddc87cb4fda;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hc1ee32d9ab1956a8b28ff6efb887f80ad7563d54a009bbc9ff9a1080;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'heaa384999390060d391c80ee29e4199e9d6fccd736ff3f1c5feafe58;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h11e570b452f6895c9c2916d8500b356ac48964ef5fa7c439c961123e3;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1171aa1b75c770f04ffeca9bd1c8271ae32fd8c70634eb820c4cb6ccb;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h163714baff1dcf01f3a92a9352d7c77f295999708c62c3b960019f384;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1ebd230f0b91a0f49d815ad94df1820c1a1c88627915fda8edd1e6865;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h190fdb52f88b77e766d8cc0a296c05de4c31b738c5431856f96520aa3;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h62fae1827638452b5a6c644fcea03a2306cf52e9b4d44104be03ff06;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h15c5a2516be189918903f5009460b8b3a0d04ffdc8d12ae7308deff1f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hf1d26777a0c9ccff399c6f8eabf900429cd7dd43b1c0b4974e65d723;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h300f0c39a1c4447d98bcd72944b89bc2b85e19d475a9fdc5d01b668c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h174018b763482bb7521307a878ce81efd9f5abb8fb411b6e7b70a6eb8;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1c2248e448ed7028391a2a61ca30f4f73d26185f12ca025388dc8a963;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hd0624a412371662a74c793d06f2f0b833c4b3849d975d958c764b525;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h414dbf9f74e06d258afbae45eb58e0ca32d073f9db24f6a619ae7b1d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h11a4b77fa3d44a087a9ebc85cd53ab6c0bd838d30b00c5771adfed584;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h16645132ad3fe323250367256d08528b2830c0b9a44db148f5410677c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h11fbc9895b60dc8bf9ccef801cc35fc50e255d981c3323b60ee2704c0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hced5cbfe6f5956694f9d6796618f90c9989c91c0037cc041c8b2409e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h2403bf3e7a4e88ca8a930ecd494709f979edc9e20ef2543d8c124234;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hdfbb9468d5d25cafb2f3a28f34d5f5a4732a7b804026296951c099db;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h16786bcdeea2cbf6e58b91f1f5067db86bf72c2a4116bf4b0b472646d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'heeace6f13d752111fe04b66284d6decd4338facdd1661f3fdd1a5dc2;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h19de7584ade69daf72a01ae9634821c9f9d858af3e81e3d256bb84cd5;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1c6893295860c2ad724011aa29a7aad800962c43ac94b2858142e334e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1578cf5a89d43669fd72ac35efb0aa794f8efd4453986294ea2071bbf;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hdd1c78b68043a793fcd87d35b6ea155755b5bfc1c0bb73f94182483f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hffeeb03bf10963927608e4e791d0f790757b843666f83c7d2c787450;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h115af13ddf45dab64c6a6b9ce66e72f195a08b3f688d78feaf8354cac;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hb65a1b52af6f2f7bfd7dd24b5ec30a764fc55d2e7f08a259a4d0b957;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h66cdfe267130d249cb8ee89bc780d781c365fe4844c7eebc4f8df5fa;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hdf0e1d51de742ba67c167775207e088cfb7b64ad5c51675fe3f314be;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h910c97be474431e36dc05b7ec962632055fe531536d4213f81635790;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h104d8d387e004ca52dc3847ab2fb127de9a32bf386688fda9997a4191;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h16333576889a95c79ef9700cb900cdebc52bc690c78e94c70ae0beaad;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1e8eedba8c16ecd042d260c3c614f1b58773ac5e66812de0401008387;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1284afffc155d917ee394418acbe9fec9c2c153bec3547afeb2421e69;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h123eb04ccb0015c241933afc7b8e6992cae6c6dc3a10a42954f4d5095;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1aeae7396dc13cd5254de3cb5bbcfa513fe1da7c3f9ee6b97d77bb3ed;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h3c0b07f5d6b9b4733e0610ffd6ef0f7d4ec1fc19985a93a10f2840a4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hd8f46ac6b78518db53a307d6273da5d700f3506852442a2d7061b5ad;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h11b09a52b6089fadfcdde1fb97c3d5217906832ba28bea43e0a1339d7;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1b72cd398a995f7e04b07723ad23f3ec62b6ca844fa24da2c11b7dc52;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1d335009ccdd2a118d7ba5419627b16a15189cf4e44aa29c9ae309f70;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1bb8609e6295a57328949f2ae6f1198aadadab7dd580cb9cdb15e342b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1d4d7594fedf16fc975e3ee7eb42797cd8fab68dae063e9d47a2c990f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h189967a2a9ce116b4e612d3813bc992acd064df95777d707d4ed7bfc2;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h4d32622e0c2e825f65531fc37fc213b8d8e16d08a0a43a016b5b55ba;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1b248f36a776898189529c242f6d483ffce45f93498f0b24c4d74a6b1;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hdc3a590fe717252395765a0702e903680018c94bbf99ede39fdfdedf;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1ae7bdf30b34b48395f1f4cfc3f2ef4edd0cca2f5d113638a50c7f5b8;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h839266ac0a0193475cd6a8cd0bb553f8cac1e2dd53d0a3fb651119ff;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1cb6c98ecebd8f1fad7050a43ed124ab7bf6ff461f0e898c160eea0ce;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h8f59a8646e05f77151dd63d7b31d15c48b8a9d88e9f7d1ab1065c018;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1677da5fb82a2aac71bc77a7158e4276b1160e3164c28aba7cc829fd0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h18fd6c23822530871fb9c6a856b2e61062405b06b427e5a14074442ce;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h194ec2a99a308c9fbb9c1e0e0711f7e3ac65ff2f8ac18d9cbd9344cab;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1d9e6eeda6ccf531c176dece735d02cef66122bf5b8583e59ee280c4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hf6c40102e87f94d2c8dbfaa6636c6c8482058c7c2a293331b3893464;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1b439ddb1f1f00b4d0a7d9822b3a3d9db837d90316235da1be363c67c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hc2f5ab62d75d4bf7beba66629550022085e4dfefc6c4077db9138cbb;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h89647da9a2c6dd703ed24bd4137f4a723767e705b96d4e60e11b9760;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1d2f3e42ca5b701610f5a4c4e4553a14af15c6e208d25c69fe3ad2ed7;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h852d638b19d364e03829de2cc1c109e23f2b3a69c9f1bf3399d3c843;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h11ffc0c31d8c30c25b06ce703aeb79a0d37c1d257eadaff969d722a14;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h151164f4ff973819e5a2440b9eeef107be128b20b16e643b80816a9aa;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h19fa9e980faee4815e9be246b85151013c358de39411e6581fb0079f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h155199a2dc6c590fa49fdec3f4d96dbebadd83000dd282a4f783e8a1f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h6c99b3f0d96cee479f3cadbb9493a1e41d1e2e0332df05d8606bbffa;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h187ea1253e6d58181831f57ae3946ec463eb1efe78fc2e85788f0acd9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h578be0eb35e2a4868e655a0204385144229ac39ee59378a7f82ff73b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1ecf0012592452fe4163e21c07c2d36f891dbddd1064a994ea97afa78;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'he3448ad2cdf2619f0716125cfe2d94fcab28e377ee6acb14339ebb91;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1f93aa504c46a9bebdefb5e2965f777331444d0612591137d65561c67;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h6a793df20daae0910b7a884fff4256c7d93a4c9a53fdca5f48aba2f9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1b7260040b32b16f6671c2735017a034a5a9aff2d6f8f115fd78a9fae;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h3efa97069297d8f7f0800cb032e7e8055c7e453f55a45780b65855a0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hf207946cc2b5b5b332d03f8911a633c0f848901acd4706892c59d772;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1d4a0d6ee263e32f759f58b455311cb5bd9c470d771e0f81fff924850;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h119cc7925bd7e04bde55effc1e8df53f917e8c97a30ed1e4871e951a1;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h673d6b5a487317023b9b2a0e3caa2e0d3f5a51bd272233f49d77294e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h15265dba7d67c17c82efdd4baa7259af9c69d424ce9cfed64c2d79c45;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1f6d9ff20131492920e8f441e068fed8e322cf7c0e645ad9692dc654d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h12a765aaaf7a49c4ef9a0870e59519abc770637f3305cfa4572779d25;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h188de9b68acf9188f0c9c4626913fff0acb7d8f7188ecf8a87051e225;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hda9c27d50e663c8b13a6ae5458d67597b34a6050e102032f095d03a1;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h17e91b234a1cd42b5def2963a7c338603b3043f7694891a1e11d44260;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1f3213a8f0d38443272e82974a2198ca44d2ec29b40916a230e5defd2;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1728a4f505cb0118b175b60333f1fcba8be7d46d6ff043d0bb3d4f2c2;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h957b1034a993591cbd204414c9d09c1977429a196dd922ec6f5e825f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h62f272d7b2ebf736ca18b0e504086b70350b08bf755980f9435d3523;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hf1a0aa16512dab6b5aae7270d27f23365402a13c3e30261318f92d95;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1734891a9fa52c86ee3061fa3b3547753d37b940767f0ede0ee3d3973;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1c66b7f438f8df4b3784f515a9e0c7c148c1daa71ddf6ee5c30c872d4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h8a764f15c964f9ace634eb728bc2355da04bab7d4474bc3741d56eb5;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1e816782ba569d2bc9e051a61e7211e32152e2cb5265c8ea3908fc2db;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h16b80c4992f00af392265a379ef01dc39b854e663f063b9e30af387fd;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h9650e9610727a18e8763045366b36aec1505c2199e8568ccaf08e53e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h954bbe94d3019bce1ffe0870ecb1095f3b830d1a617174d796827bd0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h40633d77020a382987e8118e7d038bf9a665a4d59c43fbf100f1933f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1f141d160c58790a0433df08a708cc51877fa6d9b2dd45030507f969b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1fe3f28e50cbaf609751cd871bfe1e2ce75d1154f8385e2f31982b11d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1ed3252fe97095eb40081eb584ad655268b570bee4381daf879013ed3;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hd9f44fe8ab7a26704c57a1144c986411d45960d1e2240b755a487a5;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h178e78d4e402d4795c6c59ac79fb98068d2edf8983fe9cc99ac7a7622;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hc7ab9a14a335d2bb11daeb6323fb2b48ed9b4b03d0529c78e741b8eb;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h30c02241cbc546cc406daa1895548543682fbee26d73e8cad8ce14d3;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'he8785955528c2b268c2d60b95150aac4947820854d2435db924b2175;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1a11a5858c7a1c602825253f35330347394ee2084317c26baeb2474a8;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h793c47f988b2876bc27e8605740f6f4e5b980337a8487f29a1bcf1c6;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1ffe0fa55179453135ef592e8ab6748418d2f1123dc41cb4c68244671;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h23c683eb118d1bcff0e268414af9ff620eb43da01e03c1c51eaad748;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1717cc0645df1eb4055c851f7d0c480360f86ecd5cc8cd7626f6804f6;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h15dd1fa7e2f06635c767fadb08beed16e417f58480f2ffb3f46b1d2a6;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h8e3f67c1e36e8afad36a6b2c056acc2b40479ad76c45f33dc79205c3;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hd9892096509405e75a86c40a94e6b9dcfbd8d33782120cdca9bc664;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1a02e195d3e9a25cc0d80b5f7b37a792247c6732de6f7e0e4f715b191;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h12c4687d55c25e03261cc056e3a2d4566ead4e12de07af574080b3694;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1e0daef2ed45e7e5c8cce3312f61c4b228f8b5adb87a97c9d5b7dd28a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1876829705db3567a0a97f3e68dca8228c24057c7da74de5dcd49b3b7;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h18735ebdbb6a0835720dce9ff1e293ec958652c150b6f02c79e67593b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h3f0fa84fa67736386d64f8cc4231df148ab543233c025689919017dc;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1b8f84c7341a5ed01228f98261d26cf6772075c1e7c550ef26f73e3da;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1807855e7f5f50bb9a288cf8779327fd7aec969ef0c66423d876d7dc5;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h469c60d348e7d749b770ba5079aa76501d7538d72fdf6cd964cf7799;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h155568bfefda0153651735bfdf427123124aebc84c45da7eef484a5f9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1e1654bf9e4fee98e8522932f4997951ee14cebae99e90da35ef69429;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h3ab70d4cbe5f400331a69eb44c461bbbe8c8c9b50a11f2c617ae8f97;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h5426cb879b83c1d9f9bad5ee5a69f98d18f555341c93f588c2c91f92;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1770bd8a36247c3d1770aba9d4045d2c981b486b212cc9fb9af334bdc;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h14c9ff41e4a892b97012691277e1eb7002777f7a5dfe3a245059ce5b9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h3a6523cf194bbd553cba28f8a9bf0ed76c3234b107e5896782a32869;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h5e35853b1f0508adccf87ddef1a08bfd81dd1368dd5d7135fa074e5e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hd56f05a7713eb4a6ae0f85965ebfde8ac5bbdd08d202fd041653491a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h18b4cd0da1da91e3af0f38e529dfc15b42ce2df2f82b0e20caff8621b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h180a1e1f0b70efd470935aaf9717431f9a90f996cd283c874169e5fa2;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h163b339fedc67592cb4927631f4accede8ef5ca7bb3b8f7cc09e9271b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hf4cc659f8ee3f0fe401818255630177730e0dad7a9d2a4796a74b3b5;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h66161817c433f4bbb6cab91f47fdcac614511495a0a38777170ea750;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'he3cb8577cdd0de9d98fc86bdbef546b75154d9d2b7bb68c1b2b7e09;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1b552ebc969234f69eb3b9e56d575dca407024677a96ae670a15dd90e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h13e8f1191605c304b83f915d19f777f8138c4081ba756560f590c83c5;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1bdc08248b2de8a51382330801b91d7048824f632c3f0bf32b9f2ae65;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h9dc78f5c36ddcf855284d2ab647162b82720bca86ee27a5f4997b898;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1771d2286134b447932eb4350fe9cb776df493b0fb79b123494382426;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h131f05b105af3c638c03efa19bf86747eb0354282536baf4c67076840;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h10e85bf953b4bd7ed177b19f1c8f16d992442bc58a35e940dcd2da37f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h829463a0b148a910e31e99d0555af6c4da61c50e6e173e54f12b7acb;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h169e74ea5e32511a0cdfe8e9b5ac893e3b8096f6317fcb85d9c4539eb;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1099865299fac32e48ed98097e741fc890bee9e1919766b8abbd2eea7;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hbd0aeb84044f1490a69d60e52bcdd241e3c80dc41478165838ddb60a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h48d271b4e2f32e56cf2b5ad9e7d7d14680de6e591b658944cf1fcf1e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h92928aa6f5fefb778147da46b7edc7ae895460d0fba91dd8ea0af8fd;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1f6d1a05fac86256b14acfba56791c9157f5ca4963c4fcee32fce2f50;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1034ac74863b0f75c4b4c2ad2d5ddbf6ce520a7b233a9bc363325b7b7;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h173ce88be577ecc98d3497a5d223abef328933ba5e8013edddab3252;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h139981751e4357e7cbd61a6a8f6e7d7f22725b974d87d1562965ad0f9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h801808e413ec4984de3568a8f3d8d305ff81c6318d368b1356508304;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h8350ca41224f03a2d908d39a0748f70ed879e9cb86de5153982d6711;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hc7fcda79cfd52de513428fe6c09b7cd923a8a83885319c4e8b5fa938;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1abbab4dcb99c435e4d0bd20f4f34884b17af820b7e679d3443e09452;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h19377affdb240d8f71f83f0fc4078d09f86bfec349327a27b4756aa16;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h8982f17eb91bbde3fb21c6e8309909e91c08194c5c9d314e046658a0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1c9faec7e927961cf9f2a0ae94092b1bfef991cb2f71d485be03d0be1;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hd35f558f21dd5e51cabd9fba49d44d7045f0f835c8fea148defc5fd8;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hadd7038219e34bef7b88584ce995113fbcb4671dccf309502acb7061;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1d0811ca3bada875207c2b19d79ceacca55990e242f611c2b36c776b2;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hd34817dc2287f643250bdd14b27cd957c44ecabae238e58d9cdfe781;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1875c67ff4f5729714185bda09256d1995827c75b135d0d7e90a47dcf;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1f7322f9af2421bf670563b1820d1bd7a80247ef861eec197920183f1;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1a9641ed97851bb45b469bf556df8839a7cfb7fb9ec689933346b7153;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hd1b272224b7c98fb857472fda069c64f341442e8eb8663408a668fd4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h7e63d9ac51085c7c2a7a20a0c6e7a16cb7ffb0f4621cd69fedada60a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1f5cae8ac916539dd8438cad626009e921a4462c7d9a2450455478596;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h53d5122c15f9932a75d9c7f1424eb5225881e9b85f1dd9100bb53327;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h154a2e3568b1fd9b0767d306a7c5546c35e02eea4b023234b719a24d5;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h10821e85d172712e43540d1e59541c61d6f54ca4efce2f8f84b8fabfd;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h134c5988b293ccf0d9719904188fc8da3d06dd94f0783599775bc60ad;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1bcbf0f651bbbb4b7039d3484b4975a98305e9daee33112ff81cd35ed;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hac80222ec0719d880efb160c980ec24ce1a0779fc1a9d702e06a76c8;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h4aa06548ffc2462dc51639f9b64edbb63c6e1cda93595e87254525da;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h50a030c4f3b4c117e5edb06e3f26bde1edcb01026589cc4feedd327b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h19f832b592f360654f0edd02b2499576b3754eea86359ec8a22810c0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hc0c57c0106018aa95db38d4b99f2f4b23926fa8b85025d0aa4e85096;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h34649444cf5c6c954a8d1e5792a73b1f0ae40ea6c688804c0c06474c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1e8c65df7450b2943a3db94ff0442c9d6a437b732cf7d2362b1bb5c31;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1fe95fb7ae6b159a20db491c1c078806b1e2b966b8e1ea12f4197f03f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1167736f6a20d6f2a74a62322465278aed1df4764b290a9d0ab32a393;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1fcd17c0fab48e1f4091f25a76baeb088a49c386bc1da743a8a475c3f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h145267ffdebb281d69bd5f07fd2a6bb62eaec7be79cf206c38645b99a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h16d9c1683f3c1e5ca5bb871c883bf4f24090d7a23e5f8ca4717667022;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h627260c4ece8c3ef07c3d4ff4c96cbe62c6592348b6d57f5a4630a05;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h16f97e83f24a9c426c6fd29503c3737c86930f8f49a002e9c49376236;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h19c7b974a100cca82461c6677d579ded7653c4318f684ddf4074e4401;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1742a6de492c794718d6bee2bc2b6e40203cb77e5e5d243b44a45e94e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hb34e41a36436a8ced8265053de6687d6f1b4f87e27e626e9b9f2ea4c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h16f663358e64050e8e9f91b7b22f617390ec125fd1632a6b81062c247;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1f96eb1280298fcdd149ef1ff17a8f4fdb2e5764d173d5996ae30a3f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h13e0a3e40b069cec3678f30cb91f874ead0f145fbd62ba1101333431c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h18c27c81e510317380e8fd0ed7d45e2ff122eb4553a862d046da0e1a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hc53339934b492adb10e5237a2c5938875b26b00f302140766049a1e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1a0cc54399a2894960c89e8631876b9008e8ae4351fec20ff1294bf7d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hd2d75a0288676e4fed3be595e033f4cb00e245e6eea7c32cf2c40525;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1265130deaf2aeeb54fdad52437c2991cdc3456fc049c93b1b2c2d3ed;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1d6997d381b1113aab5f678aeb5af6ecb2ec2d49d72b916d1ab7a79e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h74adb036a2858bd19c61d7bf9f6f36d6327498d39f6b57ea2babf04f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1ea856c20328d021d3a8dedb2ce76dfd06c4282d5afca848b3fd41d29;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h6f021418ed10aa5d8ac6815ef27804e897892f8074ee886a0f320984;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h15da3fa89429c3d86ead16e3403f9a10392519d7b94e3f5c300ea7b36;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hfcbde95f59c6572cf667d578358a36f9826d7bf54f81300dc565febd;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h28e3e164a8f444c103740e20cbf10077e4c6647f69ceaa42f573dc19;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h192152c866da61f8fa9b397130850f28eccd3b8c8f50aac83c72caeb8;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'ha9a06c83b2d1c5d8abd5fb417acbde0c509a731f42740f69c2efb002;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h13ba25c04188962afdb70cec400a09e181dd2012b9b2fc67cfc1a3993;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h19d757f0dab30272c70ea32f7dd11ee9c44eec7f492b8c120738fc07d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h3d911ffb1b53351668717319c01065f228af928ac07462a8e15947cc;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h9382b82f25d3c8ec42b683955308d6eb17ae503d78521dec73621933;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h804eac51b329c5ace3a39e3119a96d39b45cae9a5168277919bfa6c2;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h86d1b8269b15bce9c556c287a8b3c63d24fcecc209b5fb9ea3698dd0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h12e69eb36afa51bf145967a47c08eca83e0ffe5aea8509bf7a22a32ba;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h12ee92e7c69b6353b1bbdbfba37d65fa7d479c74eee25d47ade5e3f0b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h772645ccd0ba0ce60af3b0809b38f9f0f8b77dbfac4261bbfcefd084;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h4636b9201841440c4aa0f9c0e07218373c31d21e96e06ab6bbd2377;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h10f55a1668202e478a59e9271c4dc5d9d3228a8958d2757bd4230859c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hde1cba6dd141530bfefed15f78553a1c926a02767bb20ac286f0a886;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hf87913a143d50823b72f2f25422c7822bb01b9cc1934e7c7cc59f29a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h194272d992bf6020aacba1d994c75c8f71272aedd1e5f5d57582abf33;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1b281704de92f21878100e6f7b416a70b1ab4b533ae612c386fe75d71;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1e0b3a3caee296f53ed099e2b5ab55a43057b120e1198a2ae98720262;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h119728adb5d22c73eb3f2b0adb521cdbbf600779fe1969aa9baa3da81;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h16271cd9fed7eb5b4484085515f925ecd6646e8a218896124219b3094;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hb2d2f1c32235e132dd64fa13b6f2fe3e9bdd64b48fce8c6de5a984a1;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h2afaf6fdcea0b36af4f7ddc11de4ea52a77b970b13b82692770f9bf2;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h5de4b46f0bc9634a57708f6dd3da9a7210044bfca4959cc315f6e23f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h123ea2a4584b7bbc9b828a5a030e9c81f25d9ffc42932fd58b97ff4a5;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1f15c60f443068c3555f0fc577039208a4355c7ecb491e6a9538c1f69;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hd590c6a08ce2afdca14c6b4c62bf4996f2bc505668d5a7e565c18486;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1b0f237ac617d72fc93fa1f10b47f535654dac933a015a880d4ff212d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h108706b1d4f3e544a40a889973a27e1b5250a2bfcf14ff5634e51f2ef;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h119d1111fddfad7539081ba2bd777c39b0cba837389b891c7a4dfa325;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h74015b4836ceb090d19d850cd3de5ba6a6eba62f6b8fa4526836b6e1;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h17e0e780732688dc35559060875eae3d3fa906fd9fd5dac622d7a79de;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h11b755f26c996a97720384cc85b7b2829b5798297a3660a6c2e7625ac;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h19db10bfa72ae7f6b6de36254c5513faf6fe23817428a682bb1fab46a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1dee0ad843ae5c633f9bd063dd2fedb00ab2328f3448331b49a7be6c1;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h6bda552f71275eb4ace7c1874d650f71dd3c34fa60b61a44a4949802;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h5f67dc7badafc22845f7143cbb5cd39d9938b5347fd3d755f6ba4df0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1a3e2676aaa15933ecca68faaa74c268fce975493c9aede96e61654d1;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h19587aa23d5b3a55bb0be24322fecbad943db007bcd13d3be2995b97e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h119f13914faaeb2c241db8f1c738790ee30934545810284d95a085472;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h14d7eef3d5f5e91949d14aa9c881a396a60e4dc1a61ffdfc5274614f3;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h95e1afe2e57d40c52c3b6953286a747a742b41d2fa9fc9449186b31b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h8f1ddab9556be4588237b295a5da18c3e4937e2b78553bd14eadd3b8;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1b23835ae5e3343a9f5c23819a64270620cc8b24dd868fd29ff6b625c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1eb20912ef43615e3fce99111ae22793d2459a51032410e1a7ab4d205;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h2181ad0a1a21f2a18c67e44579f19621b0c1b3e8f4ed8a4a5408081;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h13fc209da44787712ddb9a9e925ebc08a3e6516c633f506d84064b40;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h6a2af2473818dc5ab66ad821551c2e2a5eb941539c5068e72c09b2d9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hb36369bd5e23c8327cfd9befb499f7182717d6aa819b113375b4815e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h37e92666af6cc71ba744285ad41e3c71f2e7434775756aae47ced638;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'he928c01b8905f5550a6f261bb209a40d8838577708d2413acc8a250a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'he87f8f6e1e3e7e62b59a27b63cb5351ddf5a7c6918e2678adea84616;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'he53ea20348d7ffdfc11f9ac69246f8f6e8fba1f74bedbe1ac96901d0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hee9a49b3976e67fdd8483bbde204879fc0b9bfacce4defed4a323728;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h6e79ab09fcfc3c9370a14560210d9122ba7214dae5057952fcb9c01;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h132436a70156f7c7f5e6def2aa659fb884dd3f4063840819651132e18;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1eb7d0b72b4bf955921c649a2a7a33c0fa91356148de39c7c07f95c16;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h613c237dd53d0d63e70cfb66c81a048d179dd1cb0516589f0e5bbc39;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h7c16411bae58df227472fe78d69cac6d216b46e280abf7709ac3de77;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h93035d7d47d96120a2f891ace94937b83f0581e28f264e5ee58bb537;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h10b62b7e66d3e4d91d955ca32adcdad39f2e6317000851059206312ca;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hfed782f0d71dee080d9c944666888656f2466f48d420ce08289b0475;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hfc248f8389e6c04426a0e4a2aef88c814f6a92041622d5f4ab7b11a2;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'ha512122d8ebfb933cdcdd83a56659a69988ce1dedf694d2a06187d8c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h10d0903a231b99bd166988a89c4bfc9ec350a4f0dd8bf6fb0db3ac821;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h19128ae924e82c7ace9923404d1499858ae14d6255b944fe0a2c2d0c4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1b4845f00c26fc3955ed3d2352dad63b34fc2333b7bf317f1eef70425;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hc76991b7444069e20bcfa63679fa1ae82ca1617907ff058990bd2bce;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hf0c9eda9ac89d0ae6117a3ac6c37db5b232fd908ba193d1d5d35c592;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h17b86e4ae7ab6e374cdc5eef769359372ee5d92dec1acbf1d8f76f261;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1bbd3f1f28e0377efd3d3c0d7d772c37b32f0a926c54ede16b09883cb;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h33bcbfee9f969db394830a920b21ae429eec144ed44bae07eae11300;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h10b53f3cecf5afae520abeb9cf1b5cdccb7ccedc4c683eccc15013654;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1c7857cf1a74197d2e4edbdea7a09f1c6cfa2b909b984caa294b9bcb5;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h312d6fe3ae109dcf97376f0c3ab3285b472fd9cf76fcc0a60258f44e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1bf340a2355a01ea97415626477f8e14dd322ac4445cd504b510cf9fd;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hf530e9fac40c60fecbba0d4ac416c6c7dc708c26a2ba663f90317846;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h364732e62e19a27f28b4003527ca88d9c51febad0afabbb8a6e6a89f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h18154d99a3e30a46841b905bbac4218966a8300da06b777ed3bd6da7d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1cc7303debb5335ad65bda228f389dc6de751ea4fd43d87419451f6c5;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h6e8dea4849f94f529575e00e8d786834e4fce19a824955ee9bb4d2b4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1d78a90852b8f4c99cba44805a5ecd1063e4d63c770ac32ec5d4dcd4f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'he35ba7ff49847070204ac465047daca1060861a5255becddf55e870d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h11a2e20aad116d10209561ccae432baf438b812c2b7da17f79ed7fc76;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h20009e7336e4c7b69c7117dc38e318311359aec785170e76c2e9cad7;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1a7824f1c2633d4b3f97edc61cec92f021cfef320a4acc76909a514cb;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1258b162e881415983651dd39f82a394dbe1b1aa12cd83620ce399b1e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h3eae8eec359d2682c6757fb6dc877c45be83dbad7afb7a3c47c60a62;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h18442924b1f73bedf1155170d15585a2feb0cfa4a7e8383a1bc5e84a7;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h17577b0f964a221662cbed7a92e659f2fab3167f7f503908b55b8273a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hefa231bfa28eca85f2b1ae373ca2e6fcc2b36f92016d77b6968d39a2;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'he9a73a05298b5f7bb90505b22dc4221e634aa145f947ab6bf8b4cce2;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h135b1e439d1858d2da3285ae3f2c6167309bca50509b0af8afe36c13c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h17dc6af2c8680e451970ab34e9c4c54fa252eb5d7915c97ce8967113b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'heaf30e13a42afc5d2713d2cc0726b22c166cb52ef1d6caf9a8cd303;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h10a8299b38ad9769afff620a66bd0dab658162b518376117adb7a703e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h193c31ac67ddccc0e724e970977998679a3062f35b402a84b7eedbf90;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h29abe67e95de201cbe90e1688e666e2714e499772a3c0f92d88d56ce;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1e1a763dbdc0adf066bae74732fd2b9fa6fb41724b77a3f23e2943de4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1079c10d8f8b0e07a8b13428d833bcd685bfbbdb6930f58020d00cc0c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h6894735108dd1dfacac79de9dcceeb3652c213dd96bc30163372349b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hc3980d90461a44514a3e6ae660fe1fa91921b7b905214fb54868fca5;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h839123067ed8e8c76e35ed3d586fac3150d97a3d735b2c8e2875431e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h198000a0a0120b463697e97fe371582e1d05e8604237597745b4b89b4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h8bb425db22348759ef163b74373634c494322d697de5f4813f8ef56f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h14b85000a14bd161feb417e4c2f6ac6477f5640afd03e55259f750a0c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1459d15c835fc28eab92f30c8c9e4d8e19f56f6318e7f26decf17e342;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1f7385022f9972a7ef511f42069010bc3cf14b92d65ca264a362a9a92;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h75a748800c0c7d5e7ca79a635a165339d4d78802cffc0d2d2d860a49;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hc7f6f07af670995e23e9c1ad21dea60594717a6b2bc9c1a082c7ed96;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1dc46f0faeea96074a832e100c0ded5612d9c73eb60f5bfe855f720d4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h142ce38d96cccc35edce501d155876fec8b4c49c1d5f6642985962aef;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hfdfd5cac9994dc03777b4d7201ae7e3db127713f7c9701bc32bf660b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h221905f5362a79ae2fc7c72b7c009302975ee9817f0f8f6b1f83e74c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h18bec0a572e9bdf8448aff63c278b5969bce27dc64bf1a0dedce7dc9e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h10f11a2d029c8e3dc8ffa8431c4548079c618b14cea500d44cac61047;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h92df59518df9b4d842bce0df6b04464b9eeae0e98f2f22e4945f5dfa;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1fb15445d11aea6a1132d5088439dc7777564e9c72f47d0ef7f671008;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'ha0d34c85dbd2fa2ea30a39ddde3d07e197a812e77b0dde079aa4a030;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'habd9ae2a60eeb50563832e53a52ff9802e5fe29680d23595441d6c2e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hc7d298d1cbe3ea4dfff5ac108c6f84b63674ade4701f38a8a9b8575c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h14ad6601275db7f745143d77d0c9862409fcc5ce6779d933a02085508;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1499f5c89fb92672e3b91e13d69985004ee86c6d418211a26d8cd845a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1bbd2435fc9b6f40ce16a57d0fd61344a5efc11e29f291842ae4ad2b6;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h15fc84dcc1a13027cd30a61968638bb6b12e3e34097b339ade7ef5255;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hf15c17a3cc2a5cd0631a9d6e451f063057870817f087438caed80153;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h372af2482a3e43b6869f6ac09e36544051caad769db28370e203f5a8;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h14cf9a80cfaff71013f60f5f8b834cfe14506f9192eb31fde0eeeba7a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1c74ba6c8a4500492cfcab9d42f5f634f8905f6a9ab910e5efe1f866;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h4848517f3601f9595fe8fd10f5a99a117259b1a8fd209111e2809f6e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h506b616d8162003b8aa85089bdb24a790b6c6f84a76d5babef596388;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1c5d95b10054a73395530e054a1fdbbd16c2b104b8d8b3cb8d27b08b5;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h75d10fd27e65fa6e01d0fbed9ba9ff703e41522e8fb8f53fa605bfc3;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hcc6bffa3fa015b636ba98a4b9c57f7984056f50a61149d5043950212;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hacbaa3ea31b5f31c1768806acfc9087c9ce53a6243291a9af784ecc7;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1abb4120504245f33816a38ee6678cf6bbe6753dbaa25ff1fc2948160;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h12f630e87df59a66fa256ee788f8dc7c1e107a3c83f27ec2e730d9df7;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h19571d0f7426474b198368a605f47cab92fcd8a4b490a132acea49eef;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h19fb3fb08c865ceefe6f7ea1ee8be30efbebfe40ad9dfa97248176929;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1b9c4fd5009fa8c171380f93e16759bfc6498c7d739377d73f76981d0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h184b09cfbb16e440f259dafb28c326b0c48691e42aefacc54cfdffab0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hdebbe29e46c557c760913905af1a23eb0c1852aa0d168b42ecfa6a7;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h17d0476c5ec9d51b6a67188ba9c7f545baecfae5e3ffeec9973d75137;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1efb52e85f12f871c523ba4b63ce5663f5548d3370f3cf31cf2c067ba;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hd2dafd180083e16de6fd31c834c018de6d1b66539329345a7a302a7b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h6b155164d9c207135c611ab0350dde745c768286949195ea0b549122;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'ha5208ae03e7ff7f89f32e98f3bc3369f6a9cb9895f69e2d7050d79a6;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h15654b02bc206e82a775c9462f952e5318bf3e34f8ad9e7662fe2dffe;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h134f1f1ba418f15dfa155a34c32b775b1a878330980936e510d4dbf2a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1adcfe66f064034b7e38f2453b11999c471c2a5d8a8b6287da06c1019;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1a4b1caead731fce9563c05a7be2f7626ada848e178c7d5b82da1130a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h58c3d4ca96d2adbcd14583260490f4c38fc6737407d66e1356d498bf;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1f2ead62d0b6b772f6214230ded384bb52459d077705939b8e9c437a8;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h6177372c58bef824e1946e5213b6f8fe84a6580a869355f222a031f2;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'he9ceb21e06ece525c6d218b26cddb57611e41203a25def8faf11cf1c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1c8c0fcde9fe92ca6ce24b021c9d90b1e761c921b4b65a77d39f6f24;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h2f3b3102f2190582d0374973430cb85ae5f07db13476608e795f30b0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hbb30c1d1685d2f7a8ea3a632472e19b99b8eb37f944d24c6c69e71f0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h13427d6e421c491a3bcca00c611741a7491ace7a35935898fe10e8854;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hd1a93a154c42bab6c007f2f7605d0be1f6efbcb6321b276a8b77e67;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1c4b7356006d304dc041c43cc486d39d637892c8fc76eeb5e5d6d298;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h118cc1104f9575fd3fe5a9ff3000f8df2aa2b30a95dd53b21fe34798a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h2347cb943b4346a8c05e0aaf7b4e661a7922dd9e176972450b471c60;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h321f62e04352f588d41fce1239fc6363d9bf117dafa327efbff7574;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hd60f3f3442f5b840bc05882fe8fba273b947252d1c0edf67034d3524;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h7e7d9c081798df3fb32c8c87976e4f5bb12a774a3d3be1e083faa730;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1695b4c992eb6f4d9528246f08876e72863cebb66ac88a17d35dfb5a0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'he1dec43c5edf1fb3476482c82a46303de636c5acaeb690d41abcf0cc;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hfbd5f3550f37790c32e8a1d06cce2f893956a44ab0bc4ba5eec8c380;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h14b6d9efa26816423d866ba3d6c7885b3c56a39abe7135732b57533cd;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h18a07f6129c5b030480217d9345a197127cd57740ed0f634fb65348ac;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h34446b36480a1c5722eab1f867022b72681e1e0f655a56ac411dd9f2;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h15d1f86ce66b2c365c8732fd7a74ec4cf006b9ba82ec655c9bf3f86a6;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hb12ef58f0044f85c19472c7ebf05a213ea7806689b2fd708bfec5ce6;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'ha8bf1784d979ca9b35826a259242ee59fae90af3228a6d961905ba26;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1afdf92bd0a70572ff6baf63b8502c1a4cef1eed0783a9da0defa4c65;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'he197ddea4038f4dd87640a55e97c5ebb193948b2bf134b0ee6801c80;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h110076381d62e91d87bc3f023b45692ba2fd813df5333106cea1865c4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hde1cb0b16e934580c8f6e71761fee58a6a66c3e610fdd74112598697;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h6563dd596d1846eef8c1d056672bd668cc659a71321167aa27dc42bc;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h126c40129ea8960fe2797a441f62b1b7da5d8043a676a2924590e566d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h16778bd03ee643b900d54e1cec9f12c9d91d4599075f9c82ff971ef5a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h7b0192f40ee198f474b1f7020742829a521f25a9ce156b56701efa70;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hc9550c889a732a53b24ea6b554393c85c61407c347443c5a82b4eb8;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h699e54bc86f2812998597b0b37cb8145e796a04de1e23e185fb53624;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h12a739850723ab7f15c620abd140cb9cb206fb732d5311971d0e85bd3;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1a329a3acc8b446aeaecd56bacf2587b8d3193d84eef957fe3b96cbe5;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1b7191d39b354b3def86326dac01e43cef061e4a9bfc764bba5acdd9a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1e28b4e52e8fa30f6b8670b6ac128658fcaeb22a86d2c22c8a9770934;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h8954372b352db53b878b78150ee17b8df22d60466b84382a407e6624;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h122cd9cccfab157e41274bea334f4c46ea5436f0f2a12494957e440a9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1ceb25ac6f846e9125bf52531b05a41029987480bfacff90ea02076f8;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hb89fc58959e1b5b99951cc7f143ffe5d240681a50fe203d9739706e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1dede7c23d646b4ffcce908c217a5afc036bd3f03c083265bbd09fa0b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1f132d99bc3423dadbc567380e665bbc6db9979200508afbf053f7d7a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h83f75fc09222c2b6fc9b8f0037a7ccc8248e3847ea2b768915593cfb;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h52dc474164d897e6551d5d125e148190158c7490e2dc67ad125c022;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1062cd17104578562096b1ed305919c609a56d26e1a5af0aab542beb6;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h13b3d4326f365ebd82f830110a5c78b46bba16c45f1ff0095bf3b55e5;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h16038890d71be8d73f1b3a5f65390810c54afec8aea988352d5b8e6a5;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h16a10e6a430cd6f8ff9872ebf1b0f444d88b0ee82432000003dc66a83;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h14f8b9c25844709f763acbe800083ab2103e7b2f40cd313980fab4dd5;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h52991985f5523c4b0ff1e8093015e0291584eaea559c936bd76e94a1;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1016f2f4e2c1c675501a722bf516f60a6f8544a554174ce5c7ea8bc39;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1001758b925513f497deadfb21c3d6fcd8f25b9043d39c44d62832c3b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'he1c8320bca4c331721b43823d5fd56a72810fc426da266d31fa7d54d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1730f069c620ac10b5525636d792ba6f4161c03c2d0c01732405aec50;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1cdaf9b32b92f874b39679d206b87e2606e91a9cde03090e6e57b269e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hcdea7032ddf10ec2f296dd99815d396ef18c119fc30d13cd4ba18c99;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h133865ada0cc4bd768273a902acc7f597e115d76700fb7e96db97be91;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1d99e661b45d335003602a8462bde9d18e9df3fd0d28de74510abe660;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h17c1855a56d4cd985312b7176fb0f1cb8f641dfff364da237a3670756;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1515bcbb22359ce3dbee3ba5a950e744425517e2d2eec6c0a1df13e41;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h157d2c4e92cd95e27174e3d31f7cde4b93d1a58a8be5fe9d00cbe608;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1a56ea2a7b9351588eb6c05bf7e9cfbde89ecfea97a95161a8e20726f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h72224dc493ee902da3a6fce1c9a660b4e4e922951f158fadd1536450;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h82bba073e5486509b1000fce3c326780bcdf384872d2d5a1ebc65a98;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'ha33d0b2a581e4271a20c64a2d95eb445429847e7e06b525bb150a6b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h8a069fe97e4fce590540b5175c340d426a2745db3e3f96e2fb50e513;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1e52a1f58ca11667cf56a7b6fb986c9d0bbc31a95059fde7452964e2d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h5f142d699c5928293faadc7093d56c9542bd0e2a7d17a845ce5c7c7b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1062a060e3c4debbf1621713a5ff0bb7cd647ee24863b27baf861b155;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h8127527c036d21e2a79bc1ce8b2defc6ffca18ba1764d31a842af027;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h139278eac81b542c3b56c3073c5a9653daf999ecac15f7cd95dc6aa9e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h8e85b011e465cccbac7b88d687aadb4cbc420c68602e717ac9c7eec2;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h16a0d2f9222dde4f2db89de9d72781d50af5c78bc0bd755a678a2064f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h3baf18435587e834d3cc74e932371962832e610d5be1a37386f3e6f2;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hbbeca4cb02673e2b73650a7556517f29439ea47193749d7708c7c0e7;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1e2a6b44a44ff3a1249402b02987527654b524c474a620c56e57c2576;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h15fede5f27dfdda335ddce85ed795599426c901422d6082aede0bdc39;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1b136eedee16fe54d9ed526c570a5f4024c43ca6bae5a73f9ebfd5563;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h5776649f0cdad67588fb5f8775c72eee136e3e454bd6bbf05926d9b1;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h125aa671e63ad946443e04ec2abe044eee577ae898fe62a4b2aa10827;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h103e89ae87f15dac2324fcbd7fb837452b5810aaf35fed508ab4599af;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h17ae7ece697d4efedf0cc7a587b171b5a1242eb2d606b79c8c0e3f523;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hcc851bb821871b2fa2365929d8024782f581d9cbcf10cd0d9f3b0685;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h620cb3235dad5f8f2c224a99c125492fcb58d3cd94ec429b6cc6c908;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h75697c77c8bd6366240edc3e818eac8cecd800c8ff785fc052b509af;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hb87cd91c9a8b69819f53d5609274043efd229c6613af8de046224725;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hca8f2d77d4e240f6557ef319c8b00bac30756369142b79b03b6e01fc;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h158ec579f790a18ddfa5c2226a16af63a2c1ff5880b38daa62f20bec0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hbcc7bc3ba232f46f04f59d0fac31232fec965c89f147f10621054552;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hc5d3587044a368c8f7696452321dea9e94fa26f632959dd00f81cf26;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h6180fd21079b9895e14715af0b2209ab09f39fc57978175540d39aae;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hbfc5b13ccb389d59529dc463f41452f16fbeb38f3ae63720d68c0305;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1c81b3ea0fe75bdce5efdf5a0a803d584aaecd44bdebd41c140b450f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h14fc41fa252e8d3193d5496eb0d4a05d0d9b5e4ce6d45411805efe101;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h15911d38c1d3b6c8fe0b2f90a7d76a5156fad99083f849e5925751af9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h38ac333d4edc2668ea39e5508e47b6cd25e7f90c50485528955f4467;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h8ebf7f2c45a6ac5df953c8c0d889315b00eb1914a7771cfe93b7c618;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h10fc6808727a546708c8dfdf5ffb68c418b54eb2a804a63ae8937f6a7;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1e3290138a44529f6d560bb5c36efcf3fbc55e19a5f4cfd9d21911b0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'haef22f9ac0864041ec1bdcba114877a7227278e4b5970c337dac8f65;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h11845e1ffe1aa0ab17e5bc747bf4d6aa33ad930534775c607dca9ebdd;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h733b1f081d14376b18a02e046969ad226e39a2aeb3df9669bd203260;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hef9c611ec89931f71d6b0ee5281c0bad7e37da99507d0c38791731cc;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hb7b060ce327b163e1fb1dc8e82a06efabea2762ded9d0f3411fd0b3e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'habd7422e79a273b83d4d0e093e936d324866c57990714af2bc207e4b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h88b698d1cacc0b832a3992ed443afef6fb8cdd47db0cbc3af0bdec8a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1dee5d35d30bb107b0f6d10e9cb669e030cb6a939b9efd3c1aef9d374;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h794035a5abfa7cb5ab7624dec1d0670ce013b479b7dccc8ed79df34e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h5665cee6ab34645c4b1607e84abe7874355b9548148420b173dbee17;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'he6fbd742c04aa8524eeae48dcacea265582bd76dec4596584938a05;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1cd1905ffb1c4fc82aa7265a9cc27b3e4f59b0c5e2a4f1f8a0eff0635;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h72bb5dd803a8573dd55a9acf9050af90fcf7d8a4f7cffc383ad6ad84;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h122102bbde59e620b913d589e9458f0106cfea186dcaa7638e7ff8921;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1079cc16dc80fe1df37fa7f2dd3aabd62cd6fe2ad2092024cc26de2cb;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hec93c678f17b6f7efbd8c525905065c7d37e37680495ee40458ccb5a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h16cb998b768380a02d9e95423d9f45ed726670580c435a9d360169f66;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h3fe8ae95b9b325f1841b0aef38e6810c23da4b418606563db6aaf363;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h2b699e13056bc45aa14bb81f8d51c6168f811ba285dd2fa915f9a181;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h416becdaadd1d548597c5257ed1637431cd9e4028be2afc019e00406;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h5deec29ee2e9f917c367b34b9f81a031e98900da7b6ee050f3e97d6a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1ad7649fdb8602794971de7e73e040da6e4b5c8d3cb3b4c3dec885c97;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h176a606c8d17538fca7fa847271ba368fd61c74995c29b360e00f2621;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h3f88811836aeb6eebf70b2de1b15ecd463cc49a85b3db2a5832130a1;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1462686b57a2173149777c4bd42d2fbd8755ee17cfa230f8089a0e9a2;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h163a1c05188f915b964156a548c1c042a53122732741a44e51b4df94e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1ee66e8d6f6866d585809cd4ba51560ea7ddfb50f3e0b5e9a8a211d66;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h41cf216da7af65c5b81a31ed6351e6873761d6d88785067758d9ef3e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1b5428d845f4a59402669ec7c3fb202b9c6495f988dfb2a122ec74667;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h591390ae9beb3bab8ff19bb4494ed38e893246eb12fbd311d8410fc7;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1675dd4f0cd2449811eae52332bd22fb4d326bc9d0eb6aeae5fdf6c88;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'ha3e905b74b7997cba5453858d8a05da6ed23b88f22edf437b8aa2325;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1b3354ef47f8140845008b282764807d3d5ea4d0c6b05310fe2b9eb8b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'he966dd8d606abff72a504ce5f214f4446989efc7d00e7b1dd282439c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'haec5c53ef05b81ba7aede291f4b27710ce7876ac35eb39a75673b779;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h163b5c986e9b1de77635e714e1b18b82cc4a55e00957e5d81eafac0b6;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h12713ff13106b40704954dd4718f20fe51886b1c96c40c465f6329fa1;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1b6941356d828dd8f899c08ad2fb831af2f3c2ea0e8f124a138cfb3bd;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h5fc721fa906d9e29ad89daba333f544ae53b56de6eef4129f3cf4abf;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h117bbf5c5df59aedca38254544a67d673931b080f09a9e5c615162824;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1ed1a3952aed4fc7802e80ea59c82fa12b173be96cd5db50536548e28;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h30c1a9a398829778c5eebd480a0412eb5363d44ef3a074018188bcad;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1bf8cb5d29d8fad55bdd897564ca4aad65caeaada2f501b260c8a30de;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h882704b142111f2fe4f10eb117e174820644e3cc53d784a87488a2a3;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1454f5acd27577eddfafe21eb5856de27a3afc1739a3b5490d1f8f284;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h13a9f5ecf2f9c5eefcf713e2a4af764e5611b317e442195c89b4d2209;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1b2ee1dfdc9018116b4e435a52943773ed4b892bfa9fef311cc769e80;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1baff061b4f4ac444b528a2a728545cc97c760138c9e52e89e5a65107;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hb8eef4940e9c67d49594d92c2ae0d55154ed3d45a379e5ab2dafbda5;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1fcc9d402b74643ba07b1da0ea54b7da04b0b5e2f758e52effa6a56d3;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1b9f45224faaac5a0d7fbbc4ff6e53ccad08506372cb64e3bbe526e22;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1442e73d70f92befc272344884e7fec839f497dcd0ce831654e7bfdce;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h687cb2bb57cc4d299cf5c226b63fe5f652b256ba4ad06ca590ed185c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'ha760202ea6e8ea37c7eac578dd4787a4155f06a6a705ce0d5c7107b7;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1b896a2708f8eb4c7756bd463a170874b1a8b7ced108df77958d4aeee;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h3e0a22bf8922e2a70ad2656d9dc0f977c48de1480e8024a7d202841b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1dba4f1475e22d15144ce1d01b01293be8f8f552f1b04ed28d58131c3;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1b1c6c736e6b080071cbcab3d17725d395dc5d557645920addecb6826;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h7605fca55bd90192098fbc12611956343e296d04302178242c67a11d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h141e3e1c7465ae80bdab7ecceddd71ec4a374724f122433707455afcf;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1cb9be3808c1bb176e5f52ad967a1dac230084619960dbc7bab2782da;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h17d408d278f7293264c0f9460d6029a69343a2d9598d1821e9f1ddfc6;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h39f30ae7be93852b120b7a0fdff93c5343a0d9c4c8f2b211b32eb98e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hddc507fde94a3e483b3514896c67afef899c3bdf27448f132362a61e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1fa09cf7ac98e4a6a9a8f33ce8b76d942677b10631588276edbd7b412;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1addd9c21e5a8afa7948359823b4a628c7c7d5ca3cadc12b51e725fd8;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hdfe121769908f671a852f22d18d38657fe876dbf5e8520cc9061f41;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h4158926ccbc350978582cb9bb7bf9fc5c8a7ddd6bca429076e6d32bc;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h14f24bfebc5a493d60b225d25e62fe7c4db8e12d43e459a9f0e1cf2ae;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1c677a4144c2f2255328c4ca57cc3e75fbac1e630262c310c252e5b9e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h10a0ab548218a3a3868c1ca91545f0bc59e02fbe108fef9a5ce074c72;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h116c15a424829a58843265be6412406ce5f8c7027e6430657e8c91a50;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h306adb400ab4244162a95d32a4066f0f57af9fcbb340cbd0ba6fea88;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hb87dacef9af89e1198aef3ad328697095fa43768168bdcf7cfce59da;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h15432210af597ba48a37003af7cbb4c865e43538c6fd1db4d0e2d835f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h168731e893359020b522ba8a5832a81dbd77f055a96f45c2d6e75574a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h16ee8d393ecf642de7001f422519c1256c7e88db167cabd2656e2281c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h2572eafca390e88bfa3e1ad6ad589ad98c66408c94769d3771faea4a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1958a51564821748c67c5823243d34d762a68651a982e8e619b68962c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h108fd82eaeda18b7ea1603f469467c63464468bcc50c5847b8cef26e3;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h14e1b0f7838bb07757fe88aae65b90eedf1b267fcba971ad14b270229;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h2873e27ba8bf751e6c3180b57927e43c0717b38a2559b418e1a33fbe;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h138642451f2e0407db12f9e2eb57671aa1ff5590bdcca43d05c1cee73;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hfa75a256a81d4cd20c9433f8e9bc1d55685af4b6d18064ab9320b896;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h84a113cf89e351ac6e0fbbb3437271450ca8d60e00a2005c720c663d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1a7fd2560e9972ff0f1bce2c7145bd375ec7879545870a42861288d46;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hfd19162c72512da539e1b5bb4decb8f8aa1f94e67d090db45d03c9a8;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h164fbc7b0d4d68f82e82fce6cdb49895807d28776a48b65a77c490626;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hd6076cf35ac874ea2e4db77b4f1e4dc9ab3a46a68ff2a604fbd848ae;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hc21106cb6487d88a262ff1e4e41ad97c603d338290f8b2ff5ebf0bdb;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h8e83d118585bc1e6c59564269899287638c7cbf36a9ea0b8651d0c34;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h6ffd93de54c97b6980233b89824ae64fd8465d69caef5f8724bd7afd;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h5c79763cd84f16e71b4ae43897885d99f39f961243c74deb3ffcbf6d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h5936e7a774b327a8f32ede9b2eb48ab2c3a88ffdb80c8be05276b05;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1170689b9a658cfcd2c2d0bbf39b59a285a79f9ae02698509a98958de;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h39143654c70ef6d0d1266f3fa17b2113ac004bfeb314f48c6cd75cbc;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h66dbce04a4e0cb309c61c9d0a1b5adfc32e6cacd9f5ccd7d74c5ebe1;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1ca4d204569974612662b733e2a89ea5791aedc331af3e6bcdb135b77;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h10dc9780e8392e846a381549d077544d76ea36d24c97244e5386abb7c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h116d4a19625d2e67c57f45d81d3882bc35780bd5b693f91796b205002;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h12a2d03d52891745924b1bef74e6988b5574e40849dd7768a19e0f770;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h146cb86459b85e35e764976d31541695d812e0ec7254c0070b8199c99;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hac7105c0f294809a27eda27a70a7f4c585cbe5d47d7463504d65522e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h417af2df1539f1dd7075fdf02a1e1c6a1e8f6dbf6ffe1da24acf8816;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h769324bdd331dac95de601bd965ef1ac9e35d3ce3e5ca9c778f50864;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1fe42eff27b02399d930f1ef5b620b3cca4803da0dd8ff8014619166b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h3c9c9a1264e7e81cbe7245552b995cbbbcf72a72893774077ca98132;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h15f63de4bb1bde6d0cbce7c759e8c66b1d1ab182f601b284f048fa47f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1722224c50a9589212e815769c27cedbe21a389060039ba7e7ed6ec63;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h162e4d6e90772db97444ea917b376bfdd4921652aac74936186e7d9df;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hef631b10cdb0e359e69dc637fe063e825a26e171f105a5bcef8f7241;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hefe8c2e5b66bac2cfb37b97f31e027d2932a08fcf75e8ec788186948;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1fd9a459a957e13af93654c149764ecf501e830f54256ce9d2d2e92f4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h858a1f0d60feb4f41fbc009f26e30919a563ddf30b20110eef41d096;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h4d695b079edf17d88a17214057a0e3d6fa9a80418a9ab8aca54f581d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h686c25b7cb36bf9da13b715baf163b3c1d4672eecdf35aec9f0aa9b3;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h66a822cfa8d59e09eafd2a75219d47131b55f325185598e07c53af4a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'ha3614fa99a228164a3c133ec13f24da68e3bd8248f8ad79ac78f7767;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h14818c31a50d33721607a49a075f24d7715d99f45a8b287e067e244a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h54c12c12c7b797c57b822724b36cb8e91bcfe633c97a83380d6a8ad3;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1c8d43e4500660e7817dacc7d88e0441af9027e0ebfd0ecaef6750ff9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h16f91ef53b53a8e61bf49795cf2790558a75c900927e1367adf43d4f4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h319e5255516a0b95beb33142988d6d6e6efa2ca37ed2242205287ed6;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h141da19add7d185c8360a1f60558550c6421be6d553853bf1ffed8b2c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hff00ef194364f91a4cb8d963628bd81ee3a4227a7150354006e3846;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hd1003894f37a631a39e7a12cdbf4b673fb3cdd4895b1556d3c9056b1;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'ha01950e483d7b1fd578d6e26d5cce166cb5f4f5006234261d5c5cf78;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1b118f93cebdc7ed74d6da9324db42f0a1cf99fde9edc889a82b97173;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'haa0532fa016f6e6ae957035e8263b8537ddcd43ee40c51b679c1af0f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h41b67717a9d4e6f414463d322a8bb08674c8ac777d02ff4c899ba99;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1fcbfd94be907cfa408fc0b321b4eb9a5c1d79c37d84d7c07e3b4eb59;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hbdaf77226e398546ab88b90623bd1e58a08597ecfe184682a448455f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1e565b9d1c342c864e62ebe07e52c7fc5b5996b1c55aab19f062d9c9d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'he5a01cd12223960d32690f2a409720c202b252176abd7a663e6a9408;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h2d873649008d231e34e5ead0ae468d14b0e8283e0c28eb94d6c47d67;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1c0bcdc2929132110fa5d6ec62c391bc45aef37a2c0adde3e8f216c17;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h133f82bb759a11e90f3aeae1fd5fb575f31b494a8effece6cc55b766d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h11eb2a57459937deb4a8ac76a74f603ae4bebad8210c7db657a34171c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h49b0dcea36d0fbe92e656aa1c96f64df75bc3ab31081ba02aa8b8d3f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h2cd355f12bd7ff87cd0b9bfbea92335b0b4e45b6b810bd61c57166ba;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h820ecb3774b19c65baae78b035065ac2ec85af0c7b41346ca01b47d1;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h19d8b25763c77e6b5b818050811ba8b7a6b7576efb56caae184e9cb1;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1f54b1d2bd74c89bd16311ee6c03d14f04abd3e546334066464f29713;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1c6c9f89448d8cdb7eaec031e70e25e2305c3c6019f2d691dde6dd7a5;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h105868077251e09b53178fb52a260b1b75a56b0ac25829fb05a59ef4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h921985e525694404e1c2d0a6afc3629997102581d310d16ca994b7da;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h12f8b5596a9fecc0c34b4940e8fbe6d73d12bbaa352e9eb912533eaa9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1d9a24dafe2c97ba36af072bdd56989f74d2e76b9ae303f46a24e29df;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h18b677117d7b5bf5b27e307b670cf17dbffb57d33b6b8ae4c8dc55fda;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h9510e0d7424b92e198c6add7c85eb039e20cc89a90a8d3261b31dcbe;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hb5be0eaf4bd635571f829ebab60a2f39a2d3ce584eaf0ac7930d17ec;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h38a767a2e94e7307da36f00ad35c507b3881170f979a8f68ab3cea0d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h20104c0e3993475905ad8373b17567b6b1618c12d9254f50aaa172f0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h16a37ae32fb6ff338892418deb74d4cdac528a39b75a8209448f2f4e8;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hbf6fa4b22278bbdf00627b03f30e4c803b2444815f3e6ddd7df7d1ec;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'he519bd080aee0c50d04cb7df2c85e3e1671b7031e7e73cf63fdf3a2c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hcbd86ab40ac889702644889eeb0dc0bd01bd4824698ce9b35dac2374;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h2ae8c659d2173345c59854bc0e50408ecfb7a385112cb056f6c18424;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h12941d920cdcc6de32245224e35bd9d30dbf1be1c42ef9399d14e31a2;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h20c957523a3affb51754d7d80f310b084662a4ac8a66ace39bc55838;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h2e660cae1843b0c665cba10b27d18a0c56708e33a8be154a18f2fd35;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hc6d488be76e6585ee2259f1d85f4d538fd424c15b8ecbea51111bf4d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1c64f98a186a5adb7b29de86d1ce6b723167a1f410d345710e64de7a7;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hf7f76b03bbb4454863e906edbadb0c233d663476a6843120709059f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h16906ea51e6071d3a54f931ea5bc37743b2136f548d1bd103192ef236;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h17d49dda824d838e9ecb7fb2f923a0faf91ddbfc7a9c24e67c9f996c2;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h8f79261860d0bcd8ffc9fd55c3e1e611dae2147a3e14f6aeb964ade3;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h5a146869244dd1e92f04ca66a4ce54d413140dce816c5449fdc91ec2;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1f7e7e4bf234ec9756ed52f44e61efde06f568c63aaf28a80f9d0e47d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h13d93386ac6e8e59506820d1488eef39f43ddafcb38c85e28961c082d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hc72680aedc8dc69037dc1b26e3fb1a1bb03e0e0f8e6bb859490dc64c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h139437a46a8f2a7c08c6dc7b8bb30a65649cbe2ba7e932085ee362522;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h149dd3b0540dc37ffeeaa7d36a46f2b845152476684df36d2179afba;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h6512d3e9afe3d644cc168e798078b1d7e3aa425c49b9f5d50022db6b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h3fe6d70d73aa0ccf84a2e02d7a26b9a232e3d967f38c0b81c1a636f2;
        #1
        $finish();
    end
endmodule
