module testbench();
    reg [0:0] src0;
    reg [1:0] src1;
    reg [2:0] src2;
    reg [3:0] src3;
    reg [4:0] src4;
    reg [5:0] src5;
    reg [6:0] src6;
    reg [7:0] src7;
    reg [8:0] src8;
    reg [9:0] src9;
    reg [10:0] src10;
    reg [11:0] src11;
    reg [12:0] src12;
    reg [13:0] src13;
    reg [14:0] src14;
    reg [15:0] src15;
    reg [16:0] src16;
    reg [17:0] src17;
    reg [18:0] src18;
    reg [19:0] src19;
    reg [20:0] src20;
    reg [21:0] src21;
    reg [22:0] src22;
    reg [23:0] src23;
    reg [24:0] src24;
    reg [25:0] src25;
    reg [26:0] src26;
    reg [27:0] src27;
    reg [26:0] src28;
    reg [25:0] src29;
    reg [24:0] src30;
    reg [23:0] src31;
    reg [22:0] src32;
    reg [21:0] src33;
    reg [20:0] src34;
    reg [19:0] src35;
    reg [18:0] src36;
    reg [17:0] src37;
    reg [16:0] src38;
    reg [15:0] src39;
    reg [14:0] src40;
    reg [13:0] src41;
    reg [12:0] src42;
    reg [11:0] src43;
    reg [10:0] src44;
    reg [9:0] src45;
    reg [8:0] src46;
    reg [7:0] src47;
    reg [6:0] src48;
    reg [5:0] src49;
    reg [4:0] src50;
    reg [3:0] src51;
    reg [2:0] src52;
    reg [1:0] src53;
    reg [0:0] src54;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [0:0] dst26;
    wire [0:0] dst27;
    wire [0:0] dst28;
    wire [0:0] dst29;
    wire [0:0] dst30;
    wire [0:0] dst31;
    wire [0:0] dst32;
    wire [0:0] dst33;
    wire [0:0] dst34;
    wire [0:0] dst35;
    wire [0:0] dst36;
    wire [0:0] dst37;
    wire [0:0] dst38;
    wire [0:0] dst39;
    wire [0:0] dst40;
    wire [0:0] dst41;
    wire [0:0] dst42;
    wire [0:0] dst43;
    wire [0:0] dst44;
    wire [0:0] dst45;
    wire [0:0] dst46;
    wire [0:0] dst47;
    wire [0:0] dst48;
    wire [0:0] dst49;
    wire [0:0] dst50;
    wire [0:0] dst51;
    wire [0:0] dst52;
    wire [0:0] dst53;
    wire [0:0] dst54;
    wire [0:0] dst55;
    wire [55:0] srcsum;
    wire [55:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .src31(src31),
        .src32(src32),
        .src33(src33),
        .src34(src34),
        .src35(src35),
        .src36(src36),
        .src37(src37),
        .src38(src38),
        .src39(src39),
        .src40(src40),
        .src41(src41),
        .src42(src42),
        .src43(src43),
        .src44(src44),
        .src45(src45),
        .src46(src46),
        .src47(src47),
        .src48(src48),
        .src49(src49),
        .src50(src50),
        .src51(src51),
        .src52(src52),
        .src53(src53),
        .src54(src54),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25),
        .dst26(dst26),
        .dst27(dst27),
        .dst28(dst28),
        .dst29(dst29),
        .dst30(dst30),
        .dst31(dst31),
        .dst32(dst32),
        .dst33(dst33),
        .dst34(dst34),
        .dst35(dst35),
        .dst36(dst36),
        .dst37(dst37),
        .dst38(dst38),
        .dst39(dst39),
        .dst40(dst40),
        .dst41(dst41),
        .dst42(dst42),
        .dst43(dst43),
        .dst44(dst44),
        .dst45(dst45),
        .dst46(dst46),
        .dst47(dst47),
        .dst48(dst48),
        .dst49(dst49),
        .dst50(dst50),
        .dst51(dst51),
        .dst52(dst52),
        .dst53(dst53),
        .dst54(dst54),
        .dst55(dst55));
    assign srcsum = ((src0[0])<<0) + ((src1[0] + src1[1])<<1) + ((src2[0] + src2[1] + src2[2])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15] + src18[16] + src18[17] + src18[18])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13] + src19[14] + src19[15] + src19[16] + src19[17] + src19[18] + src19[19])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6] + src20[7] + src20[8] + src20[9] + src20[10] + src20[11] + src20[12] + src20[13] + src20[14] + src20[15] + src20[16] + src20[17] + src20[18] + src20[19] + src20[20])<<20) + ((src21[0] + src21[1] + src21[2] + src21[3] + src21[4] + src21[5] + src21[6] + src21[7] + src21[8] + src21[9] + src21[10] + src21[11] + src21[12] + src21[13] + src21[14] + src21[15] + src21[16] + src21[17] + src21[18] + src21[19] + src21[20] + src21[21])<<21) + ((src22[0] + src22[1] + src22[2] + src22[3] + src22[4] + src22[5] + src22[6] + src22[7] + src22[8] + src22[9] + src22[10] + src22[11] + src22[12] + src22[13] + src22[14] + src22[15] + src22[16] + src22[17] + src22[18] + src22[19] + src22[20] + src22[21] + src22[22])<<22) + ((src23[0] + src23[1] + src23[2] + src23[3] + src23[4] + src23[5] + src23[6] + src23[7] + src23[8] + src23[9] + src23[10] + src23[11] + src23[12] + src23[13] + src23[14] + src23[15] + src23[16] + src23[17] + src23[18] + src23[19] + src23[20] + src23[21] + src23[22] + src23[23])<<23) + ((src24[0] + src24[1] + src24[2] + src24[3] + src24[4] + src24[5] + src24[6] + src24[7] + src24[8] + src24[9] + src24[10] + src24[11] + src24[12] + src24[13] + src24[14] + src24[15] + src24[16] + src24[17] + src24[18] + src24[19] + src24[20] + src24[21] + src24[22] + src24[23] + src24[24])<<24) + ((src25[0] + src25[1] + src25[2] + src25[3] + src25[4] + src25[5] + src25[6] + src25[7] + src25[8] + src25[9] + src25[10] + src25[11] + src25[12] + src25[13] + src25[14] + src25[15] + src25[16] + src25[17] + src25[18] + src25[19] + src25[20] + src25[21] + src25[22] + src25[23] + src25[24] + src25[25])<<25) + ((src26[0] + src26[1] + src26[2] + src26[3] + src26[4] + src26[5] + src26[6] + src26[7] + src26[8] + src26[9] + src26[10] + src26[11] + src26[12] + src26[13] + src26[14] + src26[15] + src26[16] + src26[17] + src26[18] + src26[19] + src26[20] + src26[21] + src26[22] + src26[23] + src26[24] + src26[25] + src26[26])<<26) + ((src27[0] + src27[1] + src27[2] + src27[3] + src27[4] + src27[5] + src27[6] + src27[7] + src27[8] + src27[9] + src27[10] + src27[11] + src27[12] + src27[13] + src27[14] + src27[15] + src27[16] + src27[17] + src27[18] + src27[19] + src27[20] + src27[21] + src27[22] + src27[23] + src27[24] + src27[25] + src27[26] + src27[27])<<27) + ((src28[0] + src28[1] + src28[2] + src28[3] + src28[4] + src28[5] + src28[6] + src28[7] + src28[8] + src28[9] + src28[10] + src28[11] + src28[12] + src28[13] + src28[14] + src28[15] + src28[16] + src28[17] + src28[18] + src28[19] + src28[20] + src28[21] + src28[22] + src28[23] + src28[24] + src28[25] + src28[26])<<28) + ((src29[0] + src29[1] + src29[2] + src29[3] + src29[4] + src29[5] + src29[6] + src29[7] + src29[8] + src29[9] + src29[10] + src29[11] + src29[12] + src29[13] + src29[14] + src29[15] + src29[16] + src29[17] + src29[18] + src29[19] + src29[20] + src29[21] + src29[22] + src29[23] + src29[24] + src29[25])<<29) + ((src30[0] + src30[1] + src30[2] + src30[3] + src30[4] + src30[5] + src30[6] + src30[7] + src30[8] + src30[9] + src30[10] + src30[11] + src30[12] + src30[13] + src30[14] + src30[15] + src30[16] + src30[17] + src30[18] + src30[19] + src30[20] + src30[21] + src30[22] + src30[23] + src30[24])<<30) + ((src31[0] + src31[1] + src31[2] + src31[3] + src31[4] + src31[5] + src31[6] + src31[7] + src31[8] + src31[9] + src31[10] + src31[11] + src31[12] + src31[13] + src31[14] + src31[15] + src31[16] + src31[17] + src31[18] + src31[19] + src31[20] + src31[21] + src31[22] + src31[23])<<31) + ((src32[0] + src32[1] + src32[2] + src32[3] + src32[4] + src32[5] + src32[6] + src32[7] + src32[8] + src32[9] + src32[10] + src32[11] + src32[12] + src32[13] + src32[14] + src32[15] + src32[16] + src32[17] + src32[18] + src32[19] + src32[20] + src32[21] + src32[22])<<32) + ((src33[0] + src33[1] + src33[2] + src33[3] + src33[4] + src33[5] + src33[6] + src33[7] + src33[8] + src33[9] + src33[10] + src33[11] + src33[12] + src33[13] + src33[14] + src33[15] + src33[16] + src33[17] + src33[18] + src33[19] + src33[20] + src33[21])<<33) + ((src34[0] + src34[1] + src34[2] + src34[3] + src34[4] + src34[5] + src34[6] + src34[7] + src34[8] + src34[9] + src34[10] + src34[11] + src34[12] + src34[13] + src34[14] + src34[15] + src34[16] + src34[17] + src34[18] + src34[19] + src34[20])<<34) + ((src35[0] + src35[1] + src35[2] + src35[3] + src35[4] + src35[5] + src35[6] + src35[7] + src35[8] + src35[9] + src35[10] + src35[11] + src35[12] + src35[13] + src35[14] + src35[15] + src35[16] + src35[17] + src35[18] + src35[19])<<35) + ((src36[0] + src36[1] + src36[2] + src36[3] + src36[4] + src36[5] + src36[6] + src36[7] + src36[8] + src36[9] + src36[10] + src36[11] + src36[12] + src36[13] + src36[14] + src36[15] + src36[16] + src36[17] + src36[18])<<36) + ((src37[0] + src37[1] + src37[2] + src37[3] + src37[4] + src37[5] + src37[6] + src37[7] + src37[8] + src37[9] + src37[10] + src37[11] + src37[12] + src37[13] + src37[14] + src37[15] + src37[16] + src37[17])<<37) + ((src38[0] + src38[1] + src38[2] + src38[3] + src38[4] + src38[5] + src38[6] + src38[7] + src38[8] + src38[9] + src38[10] + src38[11] + src38[12] + src38[13] + src38[14] + src38[15] + src38[16])<<38) + ((src39[0] + src39[1] + src39[2] + src39[3] + src39[4] + src39[5] + src39[6] + src39[7] + src39[8] + src39[9] + src39[10] + src39[11] + src39[12] + src39[13] + src39[14] + src39[15])<<39) + ((src40[0] + src40[1] + src40[2] + src40[3] + src40[4] + src40[5] + src40[6] + src40[7] + src40[8] + src40[9] + src40[10] + src40[11] + src40[12] + src40[13] + src40[14])<<40) + ((src41[0] + src41[1] + src41[2] + src41[3] + src41[4] + src41[5] + src41[6] + src41[7] + src41[8] + src41[9] + src41[10] + src41[11] + src41[12] + src41[13])<<41) + ((src42[0] + src42[1] + src42[2] + src42[3] + src42[4] + src42[5] + src42[6] + src42[7] + src42[8] + src42[9] + src42[10] + src42[11] + src42[12])<<42) + ((src43[0] + src43[1] + src43[2] + src43[3] + src43[4] + src43[5] + src43[6] + src43[7] + src43[8] + src43[9] + src43[10] + src43[11])<<43) + ((src44[0] + src44[1] + src44[2] + src44[3] + src44[4] + src44[5] + src44[6] + src44[7] + src44[8] + src44[9] + src44[10])<<44) + ((src45[0] + src45[1] + src45[2] + src45[3] + src45[4] + src45[5] + src45[6] + src45[7] + src45[8] + src45[9])<<45) + ((src46[0] + src46[1] + src46[2] + src46[3] + src46[4] + src46[5] + src46[6] + src46[7] + src46[8])<<46) + ((src47[0] + src47[1] + src47[2] + src47[3] + src47[4] + src47[5] + src47[6] + src47[7])<<47) + ((src48[0] + src48[1] + src48[2] + src48[3] + src48[4] + src48[5] + src48[6])<<48) + ((src49[0] + src49[1] + src49[2] + src49[3] + src49[4] + src49[5])<<49) + ((src50[0] + src50[1] + src50[2] + src50[3] + src50[4])<<50) + ((src51[0] + src51[1] + src51[2] + src51[3])<<51) + ((src52[0] + src52[1] + src52[2])<<52) + ((src53[0] + src53[1])<<53) + ((src54[0])<<54);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25) + ((dst26[0])<<26) + ((dst27[0])<<27) + ((dst28[0])<<28) + ((dst29[0])<<29) + ((dst30[0])<<30) + ((dst31[0])<<31) + ((dst32[0])<<32) + ((dst33[0])<<33) + ((dst34[0])<<34) + ((dst35[0])<<35) + ((dst36[0])<<36) + ((dst37[0])<<37) + ((dst38[0])<<38) + ((dst39[0])<<39) + ((dst40[0])<<40) + ((dst41[0])<<41) + ((dst42[0])<<42) + ((dst43[0])<<43) + ((dst44[0])<<44) + ((dst45[0])<<45) + ((dst46[0])<<46) + ((dst47[0])<<47) + ((dst48[0])<<48) + ((dst49[0])<<49) + ((dst50[0])<<50) + ((dst51[0])<<51) + ((dst52[0])<<52) + ((dst53[0])<<53) + ((dst54[0])<<54) + ((dst55[0])<<55);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h0;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8d204e51c67150be004dcaba10bb8a0d16ab3127fe5bd2dbf5fe81959667252e573314ec301bfadb69463bced5cd8a3c2c2b6824fc48b7cd57520277dc9fe53bc336949778dba6c7970f04c22fb6a805b093ea276ed1224d2f0fa900a93ec5c351ff;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1f5c269f62558ab0c02ed1366af20b276a1e9f3dc0b7a0385fe204bd260894ecf8866e166d898a76e5cbf3b39ea2fd5bf2203c715b83ef8686cf9925427e20c409e315b2373215afcdfc45d89d82b79ecc4dfe4e87cb883ac0c75cf712e8b16ddd85;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h81326cca8d273bc7d44ec90c84abeff42c988d40eaaad91f56e899972162e53bdada11542d73c01ff877d545e75714e705afef586ef6b7be3582b3e789be504d1aabc340e97ff273d30040dd5f93acce028968031915db94f8fc8fd0b98a74c3e904;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbfb56544f466129193f397585a0949a808c9fe675c37e14b03dfbceabe59cd3fad91a1322781a321450c60e8ab008be7363207c1bdd0b57bbcad9dd5345689a550a334cd1f8fc07f4701b22be0731775758b31dde2515f6038f3ea745d7de555866b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h42d92d3b2b6ca31f541420978ede671c2205580e866e0e7a0ef670f88f1a0da7c1e7cb857b98b0013ecbcec773f4712577e87dd60eeb6bd6c3cc7ea7d2786e5bbb1646e658ba8cd0628779b1fd6452f8e8bd76cee82cb09203d63575502a122ba101;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9f58e49c0619f3aa63c0864579209d2394f08215be7fb4d84489a23b48b64ca04fbfbaef1d353d818935788dba9b01c0028ba94e1019f2d5ab316a4b642e0e1f0fd8ff157dfe3ca10cb66f0577ad166da44de82ac7c0bea4502f7913cc62820b90e3;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdfd792d456ae0858f6a5de17f1f83e71f0ed982dbe36a61d49b073fdccda4f29e8a9d74804750521749a38a1874f8ef42d25e09ac9cee1c23c156480c4670b62d48104a44d800f028bd3de2333c007b08e3eecbdd5455d157070ba77eb9818ee3496;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h332fbbe6831ff76d66e579cbba3097d10670e2f1901ba037d44f63fae53d059a3739e18a75e30132787ded500885f8862c7ae6ccaf83b49cfb434f8bbd854fbe2039f4b92513644ece591242c31d85a02e6f03c54e913909160192d0ff49b8edd4f0;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'haee73060f43ef40d84c3a12d40378302f1e58c41a8524a219a62f4afa27fe78963c5e0369e77265cce8242982217448b29f56fc24185c9c0d612c1ac9ad63faaa64cf5a740ea955732a145666b3eebd1940d838930c0219cdce2ed46ceafaadf4b11;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h75509e64184055a1612ac2040d010f6b1ce16ccbe89325c71dec1c06ca0abe4ea17e3af19e2eba0d92350331e5f9bb3e0688e17e8a673a7b2d45fc000f27ef6381b3c1e7534302848383042a89f50fb80af01c51852f3929b5cbb3e85aca12b85e19;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1500bc44ef9d13f60bd72dc953f81bfd87000b5a46cda71bc5c817aaf94defe5d3d372c0b50246305e37a3f4f24c7d5f2ad7e0b78de3a0620e83d6cdc448ef2ea3b3c399b59c1c7503a499e5061472b24cd8b767bd9841093566d38f913ad633f3aa;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2776cfc19c6f6a9a0654881bbfedaff3dffe54076e3734a5f136ba887304de7332bd10bcd6101fb96e2a1397ebce7a55103fab44273ca2ed371b2eccdf50d2c082e4682831965a37618649a2b544c408cd041d3a6ae555b6e2cebb78b7050a84b9cb;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbc770167c2894a44eb07f6d6e5f540c814cae44063858ff8ca9ee682085b3b5201cec2dd51f9bb8764d0e7bb135fb9f6c09bfcd8c8553dad3d395b2884927899abd196bd10e62a00279f2ce21da16ba75c274741fe192497f2386e3df36271198983;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7967e0b306d315a175f1d507e9cbcef5a0535f2d34d16c119e4feae93737f9872f6e97362aa785da01787873732ee70a86fc7c277f900711b165d98fde56f0afed07b2b76b214b0fb2f70a4103d9cd82af14926730c408b24f82046b263b75f41908;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1a408881aaf006c8165a276ddd5c062ce9598ce0c88d69654107db1014145baa55ebd5e77f78311ff44998680155a4d1620d8d7b34c814ff2bdcf98954dd2423e420edc6a948498a12fe59c5ce3512d06508aede50d1c5aa56a50021f3bf27a5d50b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb284af1a090f94a2ba201f84b59b43764404c311c2ea5ee2fb3aa23be6931d495f9524645288bc1bbd8f59e5a550eb6fdf13688aed0719f563b12dc19989564269543dbe1d9e8a6002bc5045d085a1aa3da44ebf22f01db140c98b3f43fce27b5918;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha411345255a050a478d76c27f6bdd8b5f2cfae93edb83435284b3d9f3501d46eed3a30af157656c0e9e0b9747a18c2fbb9719d16c751db3dd526814e8ae6c164489c61463be8bb84b71a73fb015b9d21d61f1147188e8b472bd2a536703a2d986981;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7a77bff21a19c80520da65665e01ad1761f56fb32120f9db67dd4bfc92ef495310f7d964ddba290861d5038a73db21c62103a80b052982426362ffefdf0fc078267365c1108ae3ba214c3cb61bb964e882ee8ca459e00d9fa5cb0a0007ce62d1bcb8;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbfea62b85fb515b835b8d401fe9d80901fff9334974c01120b8ebbce3e930dcddfe9685d6cf489442bf6b9ee555984cc73040c15f1d69a81c74283fc0dbd9e05fbcd2ebfce6702c7320ea8dd285fac7cc302092241b9d3b6ab3fef9f36e628480f93;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfbcd3964b2051668a04cdbaa449e279e4dd4bc6a6ec7d402c134210ccc28fa11c07d5daba479fda31cb6c420c11edd07bf042ad124af6d18bb4715b29a3e8887e69f82c24c5acc76f96d3ca176be687fce2faa5aaaaff1e1692c4ef71071bb3c82aa;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h259948863c069e1be3edded5c2c5bfa944094da4f953ef4382df0e42ed75b1e696825bac04462b026715529a36943ab3fa6c2dda4f69d96603b0f8e762775a5866ac4079838c65e9f47b0ec113b79f04631ceecc54bed1c1bd0d2f3a54ed1c96092d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb176e8e8895f1b1e2503cab84a3ed0515e2fa8e86c2edc3be252bb923ba5e61359abf21555b5d75fb683194b330c46411a7f47268ffaf54e489afcc956df4432eb1af33720af02af1e59d6c0e133664a2408e17a931221937f1333f77074d4eb2e35;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'haa8d1c86aaea60c498bb8b09ee88347c7617d5ac6dd57734414c0f68b888667b24d52f0791339d1323b9c99ebac4362d0d16a458d180061693cb496ad284d950b65336571318d4f50d6e6af5ed396ab2bc83513e4843348fe60eaab2ac05ce232689;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4062a588b3ded75fae1c8b42742a81e8ee1fc4cbecd4a1e669eeffe9e2659a5c4fbe4c658c4e94b715d89e4208e5527c832b8c794d8a4ee4ad17e2e9f6d655aa9bbeec138f6e9fed16159498cbc8ec2e05d5cf28b837b77566d639303f04f777d3aa;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf1794a7b09b6076dac19171954b86d28511195ccb2e5f21a2b85e247dbc8a917178a98657c5ef4058bbf81924e15a4660c7a152e8b0dfdc4e33d900c4cd9e34a40b225f6c48a2218b1877836edac0260d3d0b90ff77b2a1efcf708f8cbcc786e1fe4;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf15fb47e3e36b3dc68d70e85b9f2fa62e65202efe1347a5b3bb0b7b158ee63fecfa798a956528626af16a12c8146b6f0544e04a16c2fe7fa352b91aaf82274fae9b28534ab9c0f0dbe62bcf67f82ed4dfd9d990cc55696604f4b714742b492d236f0;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he81e52d009e652a6dfed3b1d4d5619e5e88175bb2576748f27f2b158d6e15e60fb75bd1354c3b53107438408c2ca9ab13edf6ea5916f44667f05f0330db292436fa859f19d624ccdfd673cd1bfa69d42c180420cedca07dca7b59899c944522e9d82;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h34c2e8eec90b90b1a75703a768bb513da3ff3cd983f8a9e0bfe72d6a3de522b3e0a49476b17c6db2e1feea1f9dfc876637798320247df60d4c5e816a934afda75fcd3484941f9a5122113e5c517c8551dff6d0833715f56e762d7a63126a4beb97aa;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5fe25fb4c9d162fd4d4b8e92445a9e4e4364da3feb1c6e4766b727026b1d6de855eb80b1be7c05a4b08305c0df3f062ff509ef6131656fbb7f1b85b602d12c8d3d9370128273905c9c825d50ab30a1f92e09ae291f5a48234e291198fa30169c0f88;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he24d0bdd35816258d41faab8cc880a71468808624a796ef0440163073b291cbe5b8c87a87f693a4c84f8d17714cd1c20bab2e59d5e72e049fd1462b240e6f0286678859828905b9b8bb0f6a4ffba628f2fc3afeff6efa74dbc288ac87021b67ded8;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5a1f7854b19fb660735a24db15ca7eb76e5a13b927fe054fa2cfe69102cfabdaad19757e57c5b6fcac5eebdd441bb8a8b4cdf4bf645e8823a0c5209780ceac35d116cca1ba4b255e6b0c41a7fa2a8d79689cbf41add566d60483d4f4caa8d2fc4e10;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h372a5c5bab0a0cdf0d2cb5fe18e317662b006925f4913a7bd67ed85da061b97d63e303b7f81aa0fac0d57369883389ac44968219e7acbf444e7a9002dbdb828334b5f2de34121fc4ec1dff9c5427ca739d3b2f1992b192b86ec80d8da81fccf24c6e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hde71aa47fa5809559570f47493fe48e9b54617e85da8cc4d56a65c79c0ff3b26c0d3ca4d401ac2677432344daae4470ada9c36e5bc92366e0e9a65266d023108bf6f94ab58c2a667fd3fa605f9fc05fbc36de9e02f1935da69dcc758539ed0bf0819;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h37bc9837edf4b0d10164b397c6807decdaf3d7af780fd74a6349f429aee985e1e2760376e1aeb454e861f648eb2ff73e538a1c54c79a21ac8ab5a1dcfd8d0c4563d9b0287a2e30671bbe3eadcdd2d7406f8797d5797354209a22b96b6d2d1277ebca;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h36e6da0231a09159c78dc65e2f5dcfd65ec81bea4582280a7c6e66e4945895c9aa8512e766bbac512230dae944f750c428ff774fdbd27e8c7bdc73d268638fce7a4e49e00ab2abfffe32d3cb706a807f2abfc89272ab6e651ace55f768a535010124;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hed3329bc523200b00a97df3d6fbb7e16e1b076ff73dfcbccbeba90026c14024ddc33e4c6526528de4622cdb86f1b03e4785de6d9445b665d0d0b175154e464e3237995ed776927468556ec1c21170e0312bcf3dfcea57528cc8718f81138469cc874;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h773a5744193657c96e5a97b5ce1369b8b0f452880328988033df3b0d21aa4a21e2e9e7cc01f86ae51b64bab80bd16acb5686a343110e2d9a7e43e6529ee1768ff20daa59862e56d881c4c5d173d28e99042665b0e41e0188723a97db8128bc01be74;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6843c0ea15c891c66bf66f138d5af1b8ea130120ba1c4781dc077ce3029e6794e0b072ef99020b7dc66793964cc3564a177865bae2d8ebc0b4ea2cab555398d4643bf345e550e954e2c4f9b734cfefbd149817bfc8aa8f4ec14217e147d277fa7586;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h659b31bfbd3ebdbfffe8d2febf81b8772b6dbd18db4b4802a19e25fc7a290150bfb680978efb7a7aeeec3bb84e3ca542b56f2fb4e67e7a3b28ada757d8bf6f8d97e2db75b34fbd2a8c9ab168b73df5612452492beac05488868a5806fb497fbf3f25;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha9e86e138d3875ff043056bfb79ae334ed618440dde5880f93f4478b23da2021d607ea3674cb02cd3e6bc1f1a5a216052eff73d56afc3e36808a1a9b71f05fcce04fd4d0a5f30fb1c44bf8e9f15d02d68277a86d9aae2e371dadf96d9fbb1e9bd233;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4c2a4fb1e6fe79b29355d0e4a3dab6261a676996d8339b4db7be5f6d14e81f7921b51a7f2b62b21c3a722196e2bb745cf94943ffdcb8e45027455a6d460187618565c616e347b2b6ba26ce0e42b334b0b62e0ee4016f086318968506acefbf3c71ed;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd6e104b8ad06b2752c994020c36784e5b85670cb9454365d640d9ebddc5131b35453312fc15a985edb297e6f283f46d44d7a50c14cad4c0630a59945d09a257b9f2fa4d11abe89a28f725873c980fde30741f2964f035e19cfbcdea99fdc10abd378;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb30bf5add0022a501e865506f53c68f63631c059c83800ffe75f3c2bc7f6190b9e9b526d0c26eb695706aa57f8693d0b359ff330b6181ed2f543dc441a7344f0fba340c43a85820ae6698d286e00a9172afe45ddaf946bd735e5b7b42c0ec7879c9d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h58f68ca6aee22028a838b2a70d1821fb0479a992d6817a6fd20f4a9274c4473522361bb46d2e56f556850ab3658606c3446496fc78445210fd67a0da266e2c52926701e57532f4880ce7e6964bd535d5c27659295da79bb407f0e29c66a0f6301191;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h768c1f760de41111e8199a44324d93b9ff44c86634af2e4dd6e06e3797fdb55007605e7794991236b9ff7c3780eec1245fa38a33a9d2ad8684300ec08938e0197678b1ee7fdd3a8c5bb24a993e7a2716cc265c52cde91ac224e23c45738dde80458e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h43dcd0ce86ce3f4d2736a0a12254e0c422861146da78edd1339bab618c0141eb85a34e0303e91f5f13d575ff4956c91597495d1a4d1022d7f49cd2eba6594d5489639d0247bebcfba0227e854bcc9422493c735e5dad1010dae7ef4b6e185b88060e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4589d34bc8189b77aa6e067921c4218053a53f206acc87dfe2a7bbafd69e98268432b684220af2e7179956310d4fecb9e886063f022abae10bff40cf1209eb2e7c66bb18560a7fcc7d3c03cebe549e0838e1753f5500787d4015d6a2fd256c14fb25;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb041c045874e297001947575c81e716459ebc453b659f4c5fe1f92cf04a748ed5534c0e4843c0df98f67b0b9cab7578698ca5bb060fc651d16bea3c6b210aaad8d8017ec971da03dcd2b2d2a735d692df688000c01d7059e69d2e39091ce47b5a710;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7487a7132e8b054e4e3c7da114157fcfbaa0276cca28074020dc89acb0a380e36162772c3712ef5ce195275b51a6e95bd14d2948e0b2cdfb4c26e0025097184a2750091d2f9caca4c184ba87ca6e18c930307c8b7a7eb99d243cb39e51452189bb29;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he79e17f9233a322e859ba60b58b1c17bffd0b3794d36614a777917dc2e77061c0b4b425e416b3c851ad2d02cdd54c120f0bff4291961b29c798c224343bfc2321e270887416288c929f71fd6e1916ddabf0c395a37f372656c37c9fb10a37d619e39;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h93694874b67c5c18fd3481a7de85afc3015d485f3a1c97c5690f79d6247faeb24eb3fb85611a48eb6d29c824a6f6e24b869bcce16879946434a494ff5099a967a9e5a4ee245058d11cb74aeab52755008d54fec877a24f476929440139acf9e45f59;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9c57d3f4c6f40989f07ef64bf884d38b1fbb88d1bbfebde3a6a449bbd288ad80859972e7b5461fe349f58aa6826a656cb4d9702d0297eac1add9dd0895a49531a36102d92905a484f0bf5eddd8d67363d3da810a251d11d7202c7bf7db21c9071ce2;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdd23de3f95f7800cc078f7b0455e34c881d11283f7010de5a77d798de4d40ecd7879b5e4ea6845fea0afe122685c28dc664de6e83eccc86531cbe42d2ff8f55824cf05df8f2991cfa466b345e56410fc88192ca5489dfb2b41b0e318ab32377df67f;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc4046f5a482215b95a184eabfe4f620659a83da7d57206ed7f60b8558d9bcdec6ebfc63075485625406e844e3e32db1b7deef51ea3eb149b1e4aa70c077fa373c455951aee4824cfc308abb810643a2985a8665a3bae5929d5f79b121b69138d1226;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbdacc38aa4cd28805a99da0fe889b92f64628092d61240f4af6362a7a6893f6a54466eba7377ecb0213108b2d913b986f493b9f1b3b4f5320d341c205b5f701530018bb08e1340d4d6e6aefa0ed54afb78727806e95586951ae8257c75eb37e35fa5;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1b4d53252f148a8184181d42a3c0ab06dc304ca95605f9dad494e85909fee743a2f02f2c2076f0c0978850e7d392c2aa7b8abad2840907b674e7572b803c97d96d8e3320d1b7f6f9224cb568836788c9a676732deb1a2bd6f5a188b4e31fa9998f16;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd39595aec6f6b608043bff100db94d041a23b0f383b31fb65b4adaeea55deeeacb2f534ef688d9effa7b53557b227a6c5b17fda5131f35c0ba45cce72c7f92189b4d6975481f8cadbf9f8ca8e2c0fac5e6e2b201707d60621533f03c0f735a4cc6f6;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfcce907060afdd222cdc43fa0737741205870f9326b584efdb13412471e6479de1fe3d8a9ea06b9448a2bd2c04c3d775b0ff1622c0b8a37a2304c8729ef4219594491591106f08ede40e840a964ab9b603bab408631ccb2f20e285f9152c093f2ea5;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1246248df9c303500575935ae8f6903e4103cfc48a6280c8dc718fd33b0fdca4947a8325040fcc8eb2e4dcb9608eb77e9c74f741756c1ac6d0a86c85e8c92684b8881ae4a41dda4c2d16b4f2b9052e1199b5ff41a7a29a90718fea6a083f26de88de;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf64f1ec27520a1ec38452bb20b6761dcae3290df9d4377e5258d74141b8c7029d5523b7dc606973f4ca3e4cc74f6cedcc4a32879b8dec2120495289649ca55282dbf8f1ea57491c0be79c5938f62324d103ccdd4a60edbbb92bb53792de07dccdf8a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd4495cd14064284a2959a84956075b1610e3a06b3bf70ace1346e92fc2a5e56d0fbb6faf3cd9eb2c219c8a9e6ea816975d7098e1ca7107ee7edf3eb0b0e944b544ec84482be04a88006a5e028187782a056c382270e3d17cbfb4ae788765279172d0;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7cf8aacc5c13b8f798fa3bf7f19c714d9f111e4476f97b87b5f4c68ed488ed4062e63d880274372e96e3ab8dcd09b7b37b4672e9fbebe5e49ade66d741546d38fa6eb7ade660ac093b867a6cef0875b9a9148b41b5e426d3f98cbc959b19b1e1d5d2;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h18acb1fa7cfd5c106b119786d5dfeac7626a2d6584223661b564930c6992247a112cdd39a64de5a784d7e20f1866f530e68ab520d8e6e6be699ff447999bead245ced53e2ff31dc1ad72e7b33ea4d0b2900e802ffd68dea3ad59b472b16c72f8bd0;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he39b4bc2c7117e1c24e7588035e1d3b4dced8b333417ed50df7ac857544d404acbccd8a8f8086cbdc72be2de635b515a7e006fcaef0be29c5597e0b02f08fe93ad76bb3932b5ba6ef39b425d863d3dd48999f953adc6848b2d9a546d3491c8136313;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc4a4a6995ae9c1cc3a208bc160cfe7066265e2f11c36a33ad2a9d154509008176ebfbef83155f8669bd1698d7fbf3b457e32fbc914e32203200ad92c87832da03864f33e3cda6e624fde8f9c7e99834bf6275f557dd46909dbc3d9acb72c637f4c30;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he28dbf7580cc7c170aa1dc47c2ab5eca9b38ec7acf53f040bfe3a78527ca25d4e0abeceb7e08014abb3cc4925d8b3a684c3c98c51b558e380b19c2fc36af64d5bc3e24fa081dfa384afb998378b17ab2af616ef5a13236ffe49c257f8031238bd628;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hce8e3a2b079749eeaf24e74b2462884a494750b74fd3824b843de6d223de0f3131d6c4a4763a5ba202e96bbfc9680b0d78bf621a69253c1e8aed24bbd89790b5ee619bb9d82bfb7adb763eaffea9545b3bcff657d289b49c237f5caabb634ee99d27;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc9c959f0b86f6949e8dbfc665396d944b751c2b3a3cf7f5f2159900a370a24960ab5b8992838b1b0ff56a0cf42b54b055df386e3070583607921264b9a07150a6fc397b3b64db44b215468be9e648a46f49902811b8b5133eb8dbb1e5d88b822ac55;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfe3f375f16e2ace4e14da9e8c771b276a079fe9dd712573617dbc762cc5ba170014c6c3539f6562f76d8734005017280bc3a851c43a71cdecabd009432c67db26648da611b0f92a2b01baa54860b8fd0f11673c836dcdcb8f05bb401c806168fe4b6;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h981bcfae24278df00d50092833f93a256b371d4b0d87be99309a755c1bb583f71e9d2082fd41c8fcb2fc91bd78d47f852648afc78ca0e248cec2622e4489e3a523e323410113c2a603c11936141e60049502d461d20308dc66c995032ed08d5d60aa;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h619ca09aada6c7bf73dc969fc142e7ec82517c2102719101c9c63963091af781d1e41ffc2c0158a94d892282c6e1702e939d6ca4e26d763074bc65a48727d140a922a17a0bd8f6dcf4174be918cc4e0288032a4c8a167f3ebdeba059917b198ce5a8;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h73fbd6bf4c92fc532e3fe561dac6cde51ba991775454b22f2e1ec47ae5956191acac3c8e70bb9c1d353bc81a46b7a1447ff111753c7fb5047124590f0a1a9cf472c3737e74bc1e170532c10b7c24dcf7ed6dd69abd5188d3829e9a26cc26014bbc9e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf9746203dd7afc8cdf87c9dead6ec27b0ffeab0cdba4a859861f79c352684cf90e1f0bf1b46b5006bd7d1cfb4514c4dc1094053544fccc06f1ccab2de80e1422853415951e4513dea964c12d4c575e258dcc1b3517fda977802a6a1c26074925eb0d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h65a2391446bee26c68d6021f28c298dee9e7e8e8940d1182d22826a43daf84c52b9261ea32586bf3d6e0d3e8934c65dd1bf748cb0d21efd47d1d408b4e0a58339eedd198d4e5bea35a089c9db6990712dcda40695593ccfd7914b872ea188a07beb1;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha1645966c11cdaad18630dc1a2240b41559ae40d593fd294e5feeb72432c68f39c8ec731a715e8f12153d14036b8b5f54e2ec7614229d6fe1ac4c843ec220c6718bb90ff824eca02f1f5b7027e524d9d42ce7b18a578b8000c8d139c8fca2c671e98;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1c1f04e6810d1bf82277f808ef92cc5d3f69a182440737dbf13618ec06551ea1b5ead04028c06c310255307c520e7e5295989e253ab6f5d4171b7c51214825430d033e4eebaf9b47328a079eaf451bc6dd8cda99f7c35a92eb3c2fee13052b88e299;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd2d38c36e6fcf898b01e3b160878a7b9ce2efb9dd14a7bd32bca74adc0940202d39f85d08c49aecf9cc66d5f53f6a4b802629e6e1377413a033fec9e5ae42ae60d0e3de78eaac78fd20fd9bde580ab8eda5dac74ce51e6bf2588ec1b478832418020;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd4b346f34077de84a751494f3c36720a48fd3334cf3fb941e2f398e4bfe30b2c90940e447f1f3e464bb75262fd8af2c1a8c456677e7dcb34888bf1d781d01f838730923c1e40cb06a05b6eb85b109ec8af481293e08586d2b9af6520e26f4fe4c95;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf3ccdd3c32b8847a960e77b4ee969df3a35dad9982e268c82492f0845944c3b540e74435378feff23290b7b46b109a4ac8610c39e6ea7ab32406d47bc04fff28ec652368a1d07c3c2169a3f5f94027dabb237fbe94301de291f422f68d350edccf4b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h795b0f4bca0b279f56510a11e71d33d5f48633abab2f07bf69fe07a37a1fa9e0748959f5c1237404fd9fbbf8310f907d9c4daeacb883f5e5c4c97a98ea446096dff8dc935452b9f5ddb4dc0df2a97896465d7874bbc81ce095cb209257192739b9b3;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h36f6e35d744a35a06084b719d6a7510651e3350a27b1289219b94ea800e922feb8aefc00f09f7482ede9778fe56690255bc73f61c47c938280877d526b23029c8f275c53e94da22ac3efb6d50da2d9eef7f84e19a115aa2bf4a85d153aa7a088361;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h209a150ad1d9c409677086ee68b62b0bad48c22208f0e5931473781da074e9d783695ee5056369227268aa89a9d1efdfc7b266f6fdb382bce9e5c0f8cfc96dc05802f56b7654edceaf7af23d8f18f68d0c93b56dcdd8df29bfca0cb8727afbd6ff3c;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3a7348dc68b4b201a970862ff48ef2a80fc74dd7a23278c8f61f1f6436ffd995a3d4dd256ea89291b9d5a3f72a5b740d9188ad6143b9511d2331a246d7aba8371a75f66b27b9af78b125a08de425872f7171036876434570d7330ef828203e6a218f;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3d95dcc62d305f82c1d1e70677546b2d05fbd910ea5db98a0e806fb1c312c49af53eb8db710110d8446931fa9ada2f802f50fd8145c06b76718e33d7696e51ff697a418ce6be07178df10ffd1cd998c321b9dbfa8dd4813b819ec5617f820c2b7335;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h93817c2d954c298a441a69ae225ace40583b4492d40440bdbf8dcb9681691c2c3f21cd72ac7b2f8e1f29f9594a74b05077b4b838e388d04f1bd2e04fe14a3090defb5a2baf37b5467d1ecfbfdfb3c4d1050d266b601f7e643c19de1eb09aab68321b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9cbf63910624f9130237f29fde06fd7781ea669fcf470fd191459291104cac6b6913d464d5eb21f3f5ca7dc18b4749acdfc291caedf95f3ffb250802d7ab718130e5de42489716c2996bd452cf5efceac35503e6fe146bb6ea447019535391e3dc57;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h76baece9468d0ac615db0b784ce72232c1df1c608db43f13452176f9eb6eb13a1f9563f9ef21323edd8e2f18ae6dfe1b9a5e06b7d68ecc4060ac76cebf3356bdabe1af41f61a855c591f483fe7f11e08d3275aef99ce9b603e686d83fb4958dad2b7;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha4a491c951b9a20f11a7b527ad5b9c0e42f58dc33180984e9279966e71597298e9fe94f11b9a6f2d0083c738cf4b6d0a52f32804eb63ff7607ec9c175c088bb14ddc0f98bded715375a1762b463c0c6b0bd43bac54a48a20d348314f53dcb545cd50;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hede30fd9daa40bd3d9edd6b7e2c436a03fa5930138e9077495a441944c0404ec32722b47589b127e2c2137817ec80e0d8090d9c734f2dd1645f3cae76f5a72ab1a4aa9149886f15049eedbc9d9aa5a117824ac497fb5d998cfa81876a92335fbc7c;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hff7f3ce3bdc1fc4631ea579c9297b2b9d34af47df077ff682fa7b49252b457a8410beeaac3f806772942fe145ff7e779b225853a90a70fbee9a9b523a91808a7c785ba1b618f61903d32dc399d8fb8b6014491d9d7525120fd5d6fdbe218c5161ec1;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5d3d4a4633483ebb1ad32bf07e99770c8633f005a353796ef3d4b422874e19b2f1eda9e274f36e7862f24f9a678dc70fcebc3d7158d9329a22f4a34c3b57192904567c08a14682387047af310fa5c10f0ca0ed526ff9c644475b76c6a5c0be16d6bf;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h573ec8ae644c31609dc356787dfb55f0db47cb0fbb593b54ae108951fc4bc4e3c864d7161e1ccfb2026486eefba823c653bc24fe59e840cbec25bb33154105eb0f7d63a40416613df2e8d06bee13cbc1ec1571d0cff89532d3069dc26feb70d717fc;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h363de9d474c749ffe71dcc61c3f164eb62f67cbb3e35b37acd80ffb06edd4ca7b3e97670f9b47cb7124e3d059f5169c042ce2721254b5f74c1bdff99dcdf685bf97b22e491256e29b0df47a192548ada9a1ed771fef87cf2612ca778a914192ccd29;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9af4ca6bc6441353e28b3b34211920982a1b07cf3193ad0a597e4f7dfb2edc3bdd9bdee77c72974d1af8329f25073c3872c0b2a463a2d2e719eba26ee70c10d10a403768e4b540b227ea7f72158179a7b50123d149aec8de9e20245b1697c2ac85d0;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc0beaa73541ad1b892e385fc1e8068d99fddf720c661edbda1be37aa6fd2b4a36c84c0945f589bc52a54b66ad27e610af8ebbe489a65da4d8ddf263141b16cebac05b4c0fd47e39e541680167918265ff51672a27052804bbc14a1e04a32ed165453;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb4f1c7e1f90c1be6c83d44607aa989a221920c6b9904c4e0bbacb9135a5ff674fba02a5793717ccc219054a4b1b60732c032ab275e95cab4a0284357a9d28cbdb4468e2f4a47141a454ac65721ef922e4ba6fa39b098076a4ebc3fd64e4d09ce1e97;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h64e682fcd8b189a5b2c1acd44579b3102194187c2249b3e9c10a84bf4487d139b76f1c4ff3f53885e99407ef8cef272499f676ec8deece0ab731dbf8ad13eef0a868fd321f89db4690470c99f174ac0edd7b6a5d9e83374e0df4166680e4b26d26;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h156d26c4596e1a74762b024813f29e3020a2ee9d25a3cba7b750948dbc565801fdc8fc402157a32eee1317973ca32fbb344766333febe8cb4ca139408c2eadc59e806f1c084683dabf4173cf6d8fb48ac490a516fc77988f0ac330540a6585a0745c;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6e95193cd2a01d47d1e46718ae1e993550f91defd289b3f796c4f652242f3f8e0407a3c21769bf43750b0a38dd2191b21819cef9e367ad144b659ac443709da22b82479266afcc0484c641bcf05f9fbf1e16749e9743ffc968519592363499441575;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h24b0c1b91f24cee274c166b119ef54066088fe4b269eab94e3a04036dd0a5e430bb46ff486ebdfdfb8ec1d20527da189069c58720c29539a9a83c49fee63c35bb146d18fddf9f2733341032f65e3a2e42bd6a3d37320754188349c98d67e2043299e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h32bf5e3794a6f645fd35c3b0ee5432ea590be9fa689ddbff231499b21b5b9af6c1bc467e0ecf76ba8860fa8f34879bc3ae9da0a1041381c30e38bb82e95c3c39c38ff31d38d96ca7eb38095b9c4636e26340fb03e41e53b5c3edcd083c349a6aad0d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc39ad87853bc4274a334af796d19ab40a0b895ef4535f1a3437992379de2b549f9a0e7650eb594beeb5575e599c54b15569a3e271da71c0c37e337ca2e6781e7b5d24e772b8ed76b5c968b4f0f77c25be71b11874c2b430ae203e3a7bc607e517222;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4aab30684798a16009803b1e9816ae860ad45f772795b3f4002b338878d45556e7284c40a26c4f3bce6fa7dea55cefaaf175ea1b2eaeb47cd094821ff6574f0d10f5e0b94691ff387bd6c1e5ffbdbd5023708e5dd8153c31e0e016fca1b9b57b6c4b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbff879b7a730baf60b96243ca63e588b94524cb719487bad5ed7be05fb7804b0fdd05ff1ff645c0c6e264996ad74ba97ab6c54a10728a854b80c76ff9f672a2d04e88a885788a510d405fc8c7e859bd8c48c57cffaa5daa513d234c9629f53324d5a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h70d6c5e139525cf0e28d5ae5a71a75757b91cf8e6e5bf5275b727455e9be8bb55a022c836a7a8dde8c4b51e718d3d9a85809db97ace51e1de330d1695fa30ee81f5e10b3c68eea32cb522a4bc2498a875404ab522cddeb3d731fca57fc7156413c94;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3341b8d3cb23f859c84b5bbe707133544f12e2705748eb2a854525178fea809e6e78225a2e4cbef00f83ef7632739125aae881ac707e41874664d2bf7b2ec29df7db7cd33ba49bccb925ab9d47f3e13abfe26f36b8edf4d5d4b153840b0d2469f609;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd42b1dfb56afa1a7b846fa653454888893a2133d6ef9632e35c77a7ed82673d34a1e245b61f2adadedb54caf9348469738f1006523d71fa3279373d95835db3f5ee5fc40b0228e7d613acc83a7a4673bdc42f30d3f7c3fdad8c44fd7d11fb4fb0991;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2b9352f71cce851656267e47da1b71e99aa915a8b379217e1db4b50990a3531c59fcfc3e6826278aa9680220e7ad223fb88a57026bc810524510e6900bcb7aa521c1996445f4cabf4aefd28f03cbb29ab6f76f70915676dc1cdc6576bf34326fe19b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdeac3fdde0dda87438ba7bc308c2c6f2058117ccb367ec0e0c90419691e25b99b5bb51a625df1ec7754dcadae248d5dc5ed20340b892b3f5480d554d0583b63f50f76d545ad0410fd0b97b5f4d25e2db8e17ffd3b8ded9fce17be64b4cc7ec794dc0;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8f10dbec16b3fe1f7ff2935d42d2ccc19d176178a77f3461f3c63481ad4bf6554e48b375e73ab9884968474a52a7efaf0c0103c613bdcbf492e1f94e1e4fbc2e25acad4cd7dd75cabe4317b1c3b56a4efc87c8a7b13780675a601b4ce35996b5be89;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h61643362194bebccf57a9bb2a1c71b2eaa0a07c7d157a83d1631bb3f45ddfff6db4cbc463a6d2db559819eb505e9ac3de9e46af166e21e7bf27f4b81687a6a561dbe9c22155820eb1a1b70ebb2d28f77274ca34d47832a73fb1e47ae51acd8c2e081;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'haef3722dfcfc732530cbe340ffd4a420c0a507743d759608492468c7f7953f1bcff37699edaeffddd574ed546bcc087ac09b911a4107eb6627b59d2ee149a080a4307d52bf8e0f9f5183eac644f0aed8e41a6c18911f99bdf15fd0b21282acd1854a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h109bc6586b30c3ce587070b1a8323197b3a270d8c446d8023d45b51d246c57746a3da933b15c47e21ce307b387baf0279523affd6d43438711d6918e78dc09a808dd9047f0c366c84d4d3a94ec825a4e8088616bfa6e578fbdcb27b07d653fd4f14d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbe41933932f751d8c4ca05d8de3949958cfdae504d7e0a6eb5d2833294ee6b5dcc70adaf9e371b305e13aa9f9780ed17b603d4b6cdb314ba5379985549e361b9c665214768532200bb6a64aa638493bb1c0fb5acd7c66340d0d2352cd7f2a8f6b49a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h13993daeb15ee9987a5d50049229bc7d6dfbc6a85f74514f6a52a7cbea169ec61964f38d55b9a593b71c483562388bb9ff0dc880a7ca4a55768e34779d0ab480da1edd3cbb6348a1b90a30f82e3b72cb97d652cef258d0abf65bde18b3e5613f5ce5;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h987d82f7395681788ed82f03b55985d0755567bf93278dcb613f2ce39b037283d7675308f0bebe8f524054cbd560c033fb6095cbe4088a5eb2315687050d322aefd0f82716fd64160b116721ed2affe1ac4462e59c966d76669a6105d903700f79c6;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h153ea762a0e1c60327d104a1ddf74287430a6722d1fed44224d35528e580d440cfcd10bb5285ac4c5fdcda3feeae0a6d128443a413b6aa1ee91867fe352e13bb87c7cc27ece0509958c589bd8f0c17c9d66ab1e2723f96be6c23e136fc8f982cb511;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbb4b9d7025929af67f54d7205331a5ad81101b9d8ca9f499a0278020a4eeba8a1fe945bce4818e9a37dae83648b34058a38ea3c901aea5d0e7c2a68009ede8369d50a719d644347c95efa962cdc1109336b207390dfb42fac10f5f3464811677792e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he8bc4cb02076b0901d5adf7f3635df6c6a721e929fd2f6ca6d6b1f257a292c4310e6631cf60c8483ee473957baee548de6d716791620bd2407e7a64f6ea7d068ddf339c183f1dc03a153a575e24c51da6ead39ec24b05b69c8b6168ac6f94a3e7c0e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h85f2229a693adfd40aaf2dbc7af13fa97efa493d20bcb19d8ebf85f3061e2829aa0f12ad74c1f078d64ae0947b9c938a7007ddfb5009e86ba209f81763d726de30044d7704164702382a5f7f87fef62d9b430608e9110bd344b890828fabdcb19454;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hec71ff3d4333328bb914afe3cdb0de37ba88d903f85b74b744e8ff22867c9f49124e3c13698cee74256ea89900225523cecd2cfbde961cd8b4051794ad40fe62b1f08aba88af678811f262aaf430413a83371f10bd5e9afb0c4bc87cda495be09cb6;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'heeb944a2fb89f4631e2b06124e8628aef3fae83d63269027340bea504d51ef5cc78e54d5aaa1ad5c0eb8f44bba037e3bb7c6368a2302cec62fdadfa8b36afa7e5f0ddf0b1fccba3943f5acacc19e40626a4d9770e0e4432ecc4a9d42c7ee04425e04;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb7bc7f9744f22809da05e48e7628a4d3aae3b32b0ccead9e104940f1c8b2fbb3e4fcffa3389a4d160df62da7abccb0b679dcc96d70151eeacd52810ca0269292eefaf9a1232e1d6956673eeafe0ecfd886af3f6beb684275d8b5ad968ed8879eb191;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'heb5c59b98fb29f693dec1af769e4e5c36a10640f96ea06040809b1e5dc285168793f702080ac7a281245c1dacd71a125d765cbe280ec6adc74624beac9f9d013127e2312bd40800116e436ed8b7485265ec83ae1e301f0f6b3ba5d4cfab3276a80d2;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf9abb2f76f0e42c37f684a6431206653402b6797288ea0ded36fa58d7727c34bae8af981c3136da49a54f30c3f0ecc468ca3649b55f3d791cd84480d0bae46490bd65f25357e499317097f58fe6cee26d46f94916cb9e942cf56014341c7090c976d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2b7b4401aac113c1c59832f427f5f5b84807e511762c85b7ce23e0875ab8d3261c68d5e8a842bd827d3d0d45c2c15c75f828d3fe559d581b13a19dfee7d78acfab353c8dac82b28b7ae12c8c4b0a9ae1fc055dcbb52446ac84c7d30059f33f4f4b06;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5d1024e4f463b22cc2aef242c9f9f78b4eff865e6b5b7c3fee85cabad745b9fe2f6a8a00bf99413e7c59ee84c5dcbd7e96b24824ce96a922d62af85caebed821e772e45708e67fb3736f8e114db8862cd47b43fdb7670593325135e214023980b0f4;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1e53888f8f7ee9cb23cb0635c68a088d48a9b2f58225152c5d7f15fc7d7fe67ad3681c7470a28959f49f6497e9411b80a0edec15964cd9b71e270b65d7175b2f7c97537bc7ebd604acc1cf8d6e6c6fb8493d34f6cbde7f35663cee7e32b1f4ad4533;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he3d0dc30cf6821605e78eecfa54a894f7053fb22d5663f160c80e24d50ee0c5aff662f011160937bfc59b2959f04aa00e59aa052995d7c14a780bbd97671bd4d22038b7c38fcaec5fb6c6f591534321533baf8a530eb656d0311648ec38217b47417;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdf75041e1f0ebc902337bba4620e129391f1788abdafa966ee6f44ace36d95ab12656823e9a889bae3f92768dbd96f730ba0b7a35ed46bb781891362947c7aad38df242514f4ee8c5d65fb35721a90c58b26b00e1d2b93d3204b122bb8080b428f88;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2e817998839363147c43a3f4335a2cb1bd10fc5e58a094f1e598db2f80e21ae5877013e26e82053f2312f4d9b3fc855b33846dfecb504cc40aa7f4b649a087f1454598f3d2e0697cc792a5d50a2c9e9b2d5602d64680e8e78f2557ed620db0bfd9eb;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha4345ea40b8ef048cb4b76b720d9a4dfe92385cc1120a8697e4a10c6fb590d37255c7da2cfa4b5832fa99cfeadb79bb4a2a66acd3728a27a5d8233a8ddf6e47c986fd174a4e027c0e5f4c20c022dd0a28e66fa8bfc37fa49e500bc256d27b9c706e0;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6b5c1242f80ae23e8c892d32d8b2524e0173d5c4d5d989843f0ec6851e3d60aae90146d7c97f110310766ff428cd1064440bfc76373c0b27e989ce114fc4aaa8cb0e06e31f854c3ab0138a5ab0cf14aa31dfe066fee542646f109e2ed2f55f645d43;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6c353843cec0738296d8609d9862092825b60a09f5fa3c597bd0e8d2f586ece62704bc65bad98d4189a7d70ebe0cbb92724d88d1eb77596888487d7ad1f0ee247f3e3d7a1efff391accde13f6f42fdaecc8086fb0cb45337282d19ad93082dde28c4;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5349b72b1f8556d0c03558f8f37e0407bdc216ad5e72f09ad0f14aedb89f6fbeb55edb72785fac1582e489ea3b1fa92835492693fa147b8a2114430ad0dcaa3cd119a599b6bc43e36ea6c011283c6af4060879251ca7db55d4fc0e15b569547b93ee;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h174db11d9f117570cf9c8be539d93b1c202299938e51154035472f03b8236749651d9434fcfeae5a7bd85ba02610f295dec747329528355ec15280a675449fb175cfec44ae6abe2d854220e405ad561e717f6598fa092fb6749ed4c392db435c050f;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc995b2ed9200697819a7fab5bb6b69ff89569d96c855ae7c22fc67ce817714827edc186ff6d5f1c95fde3014f50fc048958bb0794b3f730ff69ed272b79cf9677e4aeb60378eb987a739091efc2fdf70fdc61adeb97114f7203de353b69e80e81705;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h165d6850b51ce713859ef75149910b933b41d0112222b48d07eeab56674dedb0a3217670884196299d254286c517f8e41c1033573ee3a0d08425b43d4a65e563a3762a202a2b20e1123eb458684649525c0a9f5f1f3c651526c745870fef339d1999;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h93d9801411b80d1919ed59e019e8592c00712af0b39d6b859fce1980f68e1a595719fd239b9583fd11c5c0a49139d4c70692281c8a7945f2335fade717161fc5e62ce4ee68e2e5ce0fcec0915d6e8815715ff1e027c4372584598e2705d4b7fbb537;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb1340fd177800e6b468c237b6026be3eacfa2746606d5f743f886f10338af57ab5388a57c04203d7afe2e5ef0008cbb0b930ad9c19625e14e9e3d2befc510f6382dda930d0b563a9cab7b7406398b7ab5aee0fdc9c01bd41543c907d75e4258ef214;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb252b7491906970bceb2021204224e0d6d94cb104aad56df06afe30e806be0bcea9cc07696c909809f0cd261a73b62a39424e36be3500f619ba982fdbe5fd769035c6111e28242fb14c21b1eeefed9d238664a6bed889bf13d3f8d8402abd8d799df;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfad0f733d78aedff04f10cab7a0ff27dc896006e0275ea63c8f668c5d6e5907bc2e8c0222154789ab9d574dac8c6bd7ebd56f3e121fa0a47b0d335c1f1662499b84429b5cf98d4e4a6909e9443aac5e3e1f04fc77cc82f5e1f5401871e673003d721;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6fb80c5e65fe3ac67806a38911bb8781d525756d3bfadacd4c0772d2df13f2de6115acef1b882c83efd28868bdb111aba3bc30ef260b9ce7f502fc3e9ad22ef369e42479255570e495a9690dd329069ad7d178beaa39ba2dbcc999304d24c7497db5;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h496b23aa9ea138654c7b8217f23f532cdc333a1ca12efcf01a0b707903154ca19144bc0e47734fb0a110fea577ff431fcf8d22a51cf3561853ae686f14c96f82f8c8881aac1499c97d2cc193a6133c6f4d7dc6dc996e5468df77f9a98584dec3c26e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h63122530b530deac8694884f6c7c807407a4c85b0cab5837ae289bede8c52360ccaec8362cca3c28e6d7265bb7bcdd75581fa5cc5180b0560abcb53805baa396507fd9a955ac0c2eadfe5bfc195e6392148a559da102b5ab4ff35ac805934241120c;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h61c926ec593d1f4443bae468cef76a21521360cd61ad6223b8cbb094d2a52419e31d4e1472e817814c706555cb73c1252fa3f49c23162298cfe0372f0e14c94546c4919bb7361e18c50fa512a1412ac6f0f597157963462fb95bb02417af55d91e86;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7afe0c49cf39bd94272d4856626a3f187d4ee56f70debfefa9406de0355dcff64ae868bb351f315c7fd447d19deabe35c97e6e238925e18581e56f322d1d154fc60a5758ea10b52b636e69e1f89818e66d58e3dc6aa1c7b9a9df9294b3c7c6994d58;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3e3c90b8532d196cb90bf7c0cf391d35e1ac3332eb403be8e8efdcd7a03a26ce66a237504c6f4ad0437581c5b0a11f081d42d2ed50084d178240b7e4409acf36f1d43de45d8db4fdd4d37a3c3f40bc4a884da7b95d091b4e6b81c4df83230e1a4fb0;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'habc2e2b6156f03a70b05f2d4621abee5a408bdfae54d32f960c2d74f2843afb20cdd84890dd03cb4ba71bbb7efa21cf59db11fdf6213bc99a77d6493680a0a0294ba3ebf399d29776f82f5375f970c1bd417141b62a49ebc2f290899ffc8617f7e0e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hefceb16e146bf400104737b0bf7a788fff662e15002b14521a198d48c4cfaed5ffa3011a3f5d7eaadf4f3f179246903dee48b143f5910da492425a36db702ab536531db18e72029558539dcba56ac720433cd61a90245175cdf486ebfeb03e3cb13f;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h491a0a29bc5b4d7d964530fda63cc324187f8e00bb2ae656725ac6febe03027ae03668b67000adcb7466e862edcee35d2747aec0c123fefa88ee25af41ebb6302f6b46144d4991b95ae31dea08f70bd5efc01d868ebab8174478e6a2a0abec5c80a2;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h440cf98d8d2b55c2366bd146ff8d7fb6be1aaedd11fb5d5fb9b179bc03a004b0db204547a7242c08ef18f996e4e30a2748f0c1f43a990a7f44bc4d88e441e9c71ba96e6c11dbc993e2d2afed453f8111cf767c6e87d659934b4d734e2e4d18738167;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h97526c4b9153b3e6a2056d654558b21fb5d894418057c9034b8e04f2ac9e42ae32475f4b0c4942de8b22428948e84e45aacb9723c10b732de6c62fa9b5fe80eac91f83af293e7eb4b05b2cac41ec448a0590da33020f68e754689e15ae91414b8307;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h734a2b9f2d90231f91f970228e30da02653319ba3cde543b104da72e659c5f648fce0fee92343213ca58e66889635ffd48e88ce6b03ab0c38bd25684b3823a8c1cc5bca1ef91f05a15aea5af5aacf47ce77a2f7bab8ea3649d4440cf825c1c05ce75;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdfdb3228728fa4c9cb06cd74e5e3942b9e06fa2f9e89b29c908e832df45e425f4eb7b08b5f5ce21a20a5fca3c334ede2a2ce34f651c1b6699c33c222c304a8d6f4d79a73e747774fdc9aef7d47779273e916a93cc6bc7b5b6c69aa1927db7e4d176b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h63d59d5e0884d2bd7ae96325a7baf05ba5eed278fff310214201847e812a115296bfc5a37444346c55f9c9a8fa7f4eb67009f5247ceaa43b13ddcdb37b718b3ea1eec637f109e8151e795dd1f1ba09f7a729cef2f1abda47a569d4481cd612eb6ad1;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfac233c9dd9cc712585f3c495428750a875ef3207986c77ff811524a41508908fcc437aea8fb7b573497b627889adf37d670c9d78b74c675ab9a415e809af22b56a1e23e75e6aef84f69e0ca7f1d8c1498d56d7efb37a47c39f8d1bc154a6dfb7197;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8511756d4e7471def0d6cb05025bde934ac860ccf04fbf9c0da3b7d8f5e353f51c1a0e579610822929976eec9fe0f7ee877a3116ecae85ae7c6d20dbc017ce06a0f27c25badbb256fc3ac3843f018ca94003d3b812156bf617225c650104e6ac4cba;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he4c106786d879df4f882eaa1ea59f97eb93ba6988c6c3d6951bcc5a791c753c856c41adc25b97b5df1f0aaef90c03f7299477c3c949dd57059c424a709bb66c4800ffeecd65daffc1b47ae8a329fafdec354b2b8cc1a4685e773efc91d63d0caaa6f;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9cb7106df16fcedf62cd6ec3831e4b77aa8f4f58c1f6b758509d32a08d21cd0f8334c30300a6deae6bb203475fe9a11f4264955c7b16ed7a836ab7cf4f48d2f4869ea4ccfe145680dcdf4715c7e37238d47ab30511bb46d959f83436dd9ad484261e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h63f46db3a731489860be146412e816be700e1a7eaccce3ca5fd70898b4177e8a51c80da7b847d8d75ff2b11026bf03a08c9de9e781318a33118acf37d5d074642aada14a73df4f4e9ac21b3b8f7796bdb7de7fc41317d8b70cc6faa8fdcf3e36cf2a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he7a94b26db3bf04f170b9e9670b24e17b63a564543e65435fd69d1bcd4b040773d07847480002df4a006a44c4eea8041d919e712e7537ac2e401e4502baf6ad445706caf025f82f0f08acf94ce147cd47d181e12a6c50f448a5dc8ec1a32c6e3074f;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h573fa3ea525145d83eb5f696ba26a08a71f757538b83cee8d21367d149924b97a573ccd318e6a5713b2385a40487c02e7d8ab393416fa7501c4816ac1c6d1608d3cc164391b6b2ea13909ca1713ccfef887ff4300fa3fedcd087d7fe416a5fa85f63;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdb2631973ca88a260d24bbdb74d71652fe55d2c38ba6774aaafebe1884dcd26446e38632f948772b680bd093167fc789546e84c9464ce067896421c965193c92a2d834bc0e5851dd19711d1967f5c4a5af3ae8faac6a0c3116019a4151999137ed74;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hffbea02bc6a6b5a39cba2c4736535158c96a772a8db6c3cd6506042dc68aa03dffde760febaa8648fb0c9c38bed80d53f23e6c6d5eb8884b01bcf65f64ef01bfc2b1f5e5d88ecbd51a579dcd9518f7efbdc21a3b74c929a37a4a6f0650e7c49b6121;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd984e522fe21e003d482bf3ccdef36f87647a42297b92420c60b48278ea455bc700f2d502e8b6b76663ab1d28c9bdd04106882ea1986da741c2544d3dbbce2c5bc29437034230992a8a57cf716c7fabf817bc0b73bd0c1062edcde4eb7558636d093;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf631674c549eb5b116fd9a619289c1047e377c6feff5a2a32f0d3b586579caab2d39379be817a41d026280777f6abcec38ecd74efd899bd5e553da01ab3a45e5ddb52b3c4ef9208318e9b7be406dc9b098632cab8b523d529cffd2c799b38b113097;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5a3824e68ae2b7fb066078040b5f1da78ce7c65072322a5b42397bf4765f4e7beee8f9ce24d0bbbf531a365a3897c4090a0b11a3579918b9d470714d6d36f99cb2b1bfc2534fa26cb62f4617a4cf7b4b1860b74dc73dcf2257dc9466523d2e040220;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h750114d12f833a2136673c25886d16a6f21f4bbe2edaf9e5b31b30d6b3e037260f92275284762888d651f73e3756e8e3ed652357bf7f93ad92a83e3ceacd0bb2e9c1a1662c2d52f75c9655f01cb41c0c3f724fe05c5fdd1b937c4a921983cf68b077;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hab880aa38e3da1404c04038a9e3b16d05ba95af777cdff8a80e5f91a1c0216e82e30e0ba20d0135f2e06d15d4ba19de9b3487bdd76b0084f5373e82845fdf741246263e670c1a85f6b6b45ee88f4217a9771e6be187c9c211d80670f05e1842a9f5b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h415fd74a3ec08227f0ee0e347ccc1737ccf1b979ec8033294c4f3563bca22fe47e1a76cfa3ebe010c03b5ef42e08856c71e80ecb18340feff307aaef41791d4eb01f7249653872c562929b23c3bc3f5cae04c5b1399554fcd09ba48e6934e4371712;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'haeb9445304b192fdd68adc635e040e738362dc0e8316f8dd6f962398d9316f53fd1fc7283aa0e7ec0703eb276515a4a72d4bea6e2ff808fd358cc201a5682cf90cb42387a72e2cba97b527a80399b54d5a28b768fe9c6c055363e1e95c236eb9bfcb;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7237e8ca40a2cd3f10af07ff9869cd766f039634d6ee385c6465331505683310c2d74cd7402cc622e6f7cbe69c094eacf8cd9f386283370c190c9556a0f485e342b8958171e46cf29fb9c1c793dc0b6e17d4518c973f1876c7486154f93f91a843be;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h69dcd6242ebf8bd8f542e6cc13bd0c234e2a2d05338ef5a7ae3929671432c370a9f5b8bef5e938ce9e64873d42fc67409560aae80ade14968538c97fa7ea9ca76b6636f3a09a4ad3838246dc21b867da6152d5316998770493f1e515f54cd2ffe3dd;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1634740c86fc7a313f90d019ee3a1ccc239a876dcdc37aee5d34c4b945071cb6b66e21078344e8de9ebbe8639bfbecdffabee380d143435291964b3a78f1c34c06961183beff754ede9f285716b05a177b7f21fac157abdfe9e92cdc32d0a736144a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd22e44a911a515d4653b73cb052c7d14da1a8ffae74ee6d58cd1f6796eb3d269d568f952caf7b8e9f4583b23426e8d71ec8299fd40de3da8031141727ef365641fd780e9c3a864aeadd4372bf3812f913c5a9b20467716fadfc6a3032ece432b1bdf;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdc59201c148daa02d91526dab7b348375f7a371377e10b2113277b6bb34d180080b687a172e96c8571c195155c1e2089e71dfcd4c36d18655ea2b9bce1a07f16b8049234a09a3f80c04ced4b4f86f5c8e14a388275c4e038ab8c185a3b4f077d4486;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8fc550867cfa1d62c7fc9f61ccc2f9f58583b704bf6e28d65b39acb8eecc809ccf23676dd28415593c3d273f794cea1fd27ccfdb0ca255763f105d40fc164e0de61e0a1c71fec03f5ba2f1c3bbdfe1ec49fc9e17311e65c366f25665a688f41c23cc;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbbed1adefd0907863ce5220a05d83029d87be3ec25914615244f7477e9791c357a874613164dc1c9d7c0d5e0213c997b12bc074b2a596095e7a37d5f913db046c2e971f15110b1a72e6a34664717d4b3ec09bb504cd7a70c972a9a628b4ff99a7f6e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6186a070412ab4e12936bd9fce5fd1cf1bc0e1c1cfce6dae098c64c7a174159dce50f8f7c4bd8cf03b587d7e8affcad4f875275325e4bb7541e507f47941bbcd905eb066eaae1d90499a2191dd68b7f6c4d14d909eafe398dc563db3e9c1cd614fc8;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hff977c99f0fc5f73714b04ea8cb8082f0a54a60d88bd6454a2e35e0395afc54c0e8b42da59a5ff31004786ea17679edebfa82049c1d2105c8a34f6d528df821288bc66e37c5a12e5445c922d6ab27b25c5dd0c7df11ccbe291968e16a28e7a0c95e2;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h98a863a17edac64df04e20e38dc9b5f1484845447f87863c9f172f533f47435969552d0415af72a3c8ee4da7c3fae9b79712edf96151699a6a708c82dd19079e3d4c18006e2f6fc1de03c8f19a4c732afbbf623714f7b78a4c92d369936a75efab3d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf2429a2b3cdfa21cf19b85359d36abbeffad471c2ad4f54a0434a5a13d3b36ce62c6d4932b753ce7305a5ba0d1a373234a086a247892b5ef8d639480876edd5f6b44da050b2dd921d8d4a5b8ca17fc24b832f7071be4fd243b87cd85c32f2fd79aed;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha16b2e6dd4ee800ea08cd9adf0e66bab7574837aa6af8029bb20cbb46f4f9bda4a21b27b1cc2c165758ddd4be3ccf3006d88b628d1208d0adbac0dff098dc6c75fa181ec26d7fc49a35389f5d676c6c5507d8fd9f983178e112ba3ea45df81b3cf43;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hcb1a41cacb70b8edcd2007e98c6dc36d6e43aaa508d91c52ad1cd19048a6b0cff4c555e505d7b20657918d4a8c7ad7c46fd09b82b2dc77cc8bd6b3e227717e9f5c2a55e3ba2fe75deb3383878c5c632335684822bb0bb4c6b495a050c8706225d6e7;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2c2352d22285cb74f96fc86326745392e23c5d480ea9aa4336160697a19eff17fcca937ad515e4e3032e2758eab9a265cd2a58e0648e591de1dd8cb258ad43b250d5962207c255c28444c5a07c0fdc2a9c8741079afef34edd34ecb1c54d25f72071;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb36dadfdaa05b8d9a5021cf0dcd84196019c9abf7cd74668f586ac1fbfc07bd758ef2e1a757017efe0c343d0d849e3fa1997f7ea7de51287308719bcb4865a9b415f27dd4a3da90f040434e6e0eaf326c4c3fd4aee70b2852b1433e9e6a6d5ae5e78;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc4c4b5a84c63eb7fab34af90d9c23b843828307ac328f488f5566c0a5eacfeecc7b34d359227477be5b1700f745f8c87e419f27ea4df830025535bf351215eab150628a895d047250fa46ea43612227c033cb37b5a0b4af0f48fc8dbe04420f48d32;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h54f6e69efa287f711cc74ccdcd3801b6112db5a9033ea11a466c6d7429db277d88532246299510c58ba84c9963a99619566348e00b0ee2299bcecc6a8e727b7955656c6ab993c464794a6bd5bfb504ad4ee0a327c03f03c6d5abe915f231078c3039;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he4a0aed6ad0d44b881c840cfeb27e8cf95edd10f0f8f6df5e29c8d528fdbda63e25622a1f80d79e09696c2a779b211ee94d76b3acaa61346f37042b4bf970ec8796cf7b46cff8d97ab5f1311e883b9e228587f9304eb3b79504d41b641cc7a01b565;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h229cdcacbea7c22a96668d4d603417f6141ccce0e9fea57546bbf8c758582e8071589c5ec5f256709a916889352c17aa625dc791f57d8c82efc1acabf883a2402a92aeb0001275ffe2869932038f701a7c46bc0266a29a414c6d0946d14bfe5fc19f;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h18be88ce45d2ef13ac122f6eee148eeb2d892a4165da2313555296823e3df2884b017f367f6f7afd6b105fc37fa72e3b141c74cd5a5f056259dda408c5657cd1cca1db0ccc4c4f51a4820de9ebf2a04cf40147f70c8121ade4b934a036b3ab327ea8;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h63f01d1487b46e976aaa24a4cc089c6e86afa8b4e304418642ec60103bf6a5f810689ba12d8873dd9628cc0ccaedcbf044c36bafb25dd2775c06ea6b50b36b51ac0654993e9fdf1e4389d5046366aac4db63ea70fdad7f0ad55ba9ceded53523521d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5d892c70d2da1dcffb5dc7639bd1ffe6f0025baca24a78d29eaef652d1e9120f214b05c66cd416a844c3f9cd4046acb6a5895379b8a0cc76811c5dea45e8097039b17b80eb5d9004bb57ea27aaff9b47549be04b524dcee1b7ff2e67a1be52d2cdb8;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8e301546e1af2078ec7b789c7a80fe367e7cffb0aac61d89bc60175d2954d864eb96fb9477783bafbc709850ce318791d6ec1cfca42791fffd7e8f97dbb40104381771bef6413581004184a82c4b3d591cbac037b22eab21612571a0908080cfaafc;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc7c2925b780c986ce0dde16c5d0404d90e377aa53331e2fa6895560c20c40a78f6df4d53779a8b74b96b8c60d176af221c8a0bac3dcb3364a5a4e09842061befc48985d557ea56a0b6342a415ee52f620a55781005260ff02647341279978787cbe1;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbf40b2be90a55f65e91b8efc43b838264f8c73572af6a1dcdbdf773bee7c235c2e29dfbf17091e8522e091a84947427819344d9b20262bd9aa6b453ebd87ec9472c4017a86983d5b8707bc034b8a4252ca11d1845598208f8ba465cbfebee42396c3;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hed825773138cbb079941b1accd476ef4aa8cb67621118ec2a70b4e420b2b35e6d5b26d1e9ef7921fe98dfda0a5d06294eff4da5808a5df8b755d5d979db3045621bffac8bb02e1525ef96bfc2eb5b4035a5e4ce7809ddc88d194c2da7f8a54b29463;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h95cddaa5a61c75af50a501591445138cfd99d19d5a0171a90d98f35513b45644d31dff08b8b55a4afaedbb2ca31fab7c489012a5ffddb84c697d46fd082fdbf6892147f01e3b7388682d954725ae36c3f117242c4ec553229d82467d88c03e94cff1;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h19ec6c625441a4f9c0c0e42cc1ff9c7a6fd8bf1c223931a2b8d44983a0977f321c69cb1f13c006ddb4384abd07d661b0b6e5eb156e900ebeed4a40315f8d9684d0990bfc50407910c8fe1b76d7484a963845bc224de5f905d42e1ef44a13ab08ae76;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4f1a0e74aeaa1455b42e0ed6e85ed441619ef8e461cb1da6cac144cabc5e01ae40679257375f193818055a5f75d69810a29dd5fa5889a9013a00666d4a7c046433df39942d7d76b89c16882656babda31054f6de2bbc8fc0aeb50d71b2cfddaa3a92;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8b52718b89f47b7df710aad1578b378c9a635345afcfdf75d3d4979f621404fef8803cf2d380c90f4fe5978e09a4244ac69370e557de34a292a9e9967613c140f4a9e627cb4a4a48d2cbf5562da3e8885d692137b7b548f186ab1908582be7d96f3b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h306785fdaa13878cd0f6745cae10c461ee869672610551066974be65e9bb76b363680fcc8b4d768cc03b25f190b1332ec47016801e83326f12eae31c45876c1ae0be581188627e744cbe6668d2b9d0578518f89572863d50e169c0c4fbdc40e67681;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8226067451c87fc80295ad97ba2f2fb6f4a8acbeec735483aa21dc2abcecb18c92cbeeef03f565ea509fa3571241824147593390fe36688a258a037683b363359deeca9eefcf5439df3ecd49146a1b0fd8338897d530fc5115c2d4e02d9540f1a53c;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdd52a295c99b9bf0ddb1741a81c62867e092773575c2871e2dac4d08b07e3faa2cc5ac816b15fa919f4ba1c88ca2fbcd1d02a4f2a60ce5e3cbf324ab7c5abddfa7ea410f6b7319e0cccbf001ad82c21582206642be99f9015dfee0d10311ce00e8ef;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha347ce059a28c9887e2c3014b8048f9b6ab4e571ec81793fca4f1460b0cc49b0b02171c11342e67298c3039ac16f6c2903775a25b3cabcd47cc94dc03cc2d0095b481851cc773d82cd6d9d75d1e777dc77f2915756bc1b32c26fb7d87580e6393dae;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7701dcdb16377deaf464af00bc1898b21c13c55ebc36c7834ad1e08979f8e68543279f46daa7d93085786daa090fa5cab48fec1b2ff2c0a46cbd8647c9368b3bda367437647719387dc4200b2997553a5769b38f48cb2c467a0514cf639f3e464434;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf7a2a75dd7bd6cc6cda8e745b1b6615ee0fea49ef818faf5dc9e3577bca344b59b60b87c248be1396e0879dbb1b827b0a219f186ac9c471ebdc3f6e24e776772436446597855ae769c1dcf2270d9d068115912475796981a565f88412ca8678a80b5;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h53114f3f4eb904d819e08d2bd7ab8b608da3a2a054c8165180936242c639543e20e1d64a8f547f23ff4e9487da0173b95ee29402e16dfdb840132aea38bc5c828ef0a233f01296d29e1dfa842887f12b460db2460c081644a3aac96629f30fd3336f;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h553bb10ef4a9cf8db10e096aaf4f562ace86dbf83b0b3d85d93a2a8b316d40a690f610ef9a5240ee718ccb9456e774b67110852267d2ee20b3f280f52efe9700400d8fde8ff470e6513be8d1cb1e05b44974180075d38cb20fd087f3dbf7f990af5d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8d6f43f0301ac47328d9bcd08002e5e72628443bd41ccdbd99d53c1b6098b50aa35a03a7ee4ede7c753f5c6680139be719e74f0bee1eedbef3a64b4172a02a6ca4f01976a733adfa421048841ac08367b03c082d60746910ca0c2a4416ca9dda5937;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h727e5ea883c7f89c32025220c30f9b5c954debe86ae9b5e5338c92963d6b497bf4774ec23056ec1a86ac24fdad01d26827497f71de2643740b45836c1702e3ce1d264dfecaf6d8031e8cc9030d802a2fb7c6b871867205c319eabe389fcb36f849d1;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd490da4304e4605cd8579d199011944964a9e375a1db6e6b421015a363ce0696d6d975918e2c47f6176c5f1d0bfe82cf709b981948d2fda6338b9a51cc22d26e4205edc76f8d71d436be0a5b63f93f6438c53329eddc48a242cb661801d6bfba5d76;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbd2153997948ccca5c70488fbe708fddb0e9053bbc7ff77ca9936b3cc1546f8532fe283033bbe89253ca0cbc855ac001a33993f37fc0ac7192cf423afb56f891b30813104a384556dce5952c71b1717316a8fd7c09c3c2212e3267123b70cb431b0;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2dd9cf7495f932989b62399cc30640248013b47493adba33b13e6e156e06c0ef94d85dbad20515847c11a7085c8e327526ce12579ab46f28be81f1eee769af15144106bd9e1f933dea5ca59a9795c3a14411ad30c9983e033b9b92df9b6b43904f91;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4d85360a180778ae9e1e148e5c6b40b3de8cdc2df861bcd2ee04a2e09f8aee8baa2e2f7619438abf5bb8ba32aa5f6cc60bc9d104737104b8cee0a59a0eb9a86e9654f30c3e5a1fd1c245eba5a21d50599144e3e18c1536dfaf3bb28f0ecf4a0d10a3;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf327d559a4a26bd13c66de2ad46d4ddb71705e3201763def04636c6c034269bf750c19526de062f85585e6f986412ee6bc268e52ecb70c0420c056d4d28d6e66cebb5e09c3d284ff41c52ec62deefe6deaf28c1cef95b351ba3a76a1472cada42da2;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h25fae89afa7fc72a71829dcb37d297be0921ac44c0a9a6218b3159e87bb5b4bd644ba7c7dfc34d20d593b0cb8f21219c13076d0703872821e8c32e33b57cd2995733149b66cb196bff61b6b10ec9d1e8f4ddda1e959d3f606436447dccaf9c4633e7;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h62a43ca58e9eedd42d669b670cc8bb009512932e3b139d3a3fee5a07ad68cb885d0cc4ce6a34edc819be4d1044a98d10ef8f8a7032a6867123c98ff706470f47f1949f88f6d0690c0c7bc8ba73e1a9c366868b66a7674f63c19b21b22a5ad95a0c72;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hacae88adef21429602b651be5d0ba925903b2fda39344baefbb5074c4c890f3079aa3aa0fead8dd0242cb29c838bf00681d58adf15abcc9641b72ef5ddf2aa6ac5f5a2b89a0d8169026beebb9b6e57e15f563e49dd09deac2386be73516644262a83;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8ae926f7d0abd92e7183ba438d4ac4130c8c923ec929e59f9366b758de135077d2adf0c6750eb1a1716fb0e33fbe6466c1e0926592882592000d61ae1f7b99c29f37e4574a986bdc1116c95a337fbdbe2725b5e09871c699bdabead8c597911fbdab;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd43b6392cbbc2b6dfee8b5125f31299e12f8c17ff90d63627cd10da7843044e256da379395a96455a4f3add634564ab1545535624cefc83b96b094d32c350c67ea64c9644c150b394692c16fa0672f79c0cb06485ef6360edfb1d87df467e4069633;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hcb99f1f4224cd8bcf203f25d9c6e0e850c24cf65fa1d57c2a2b204bbce968845a03c66868c2225e5aed932e8c9e928b5bfbc30d9bf8d8a10dffe17ec9fc8934105938c2a8d1d4116e2cf83bda4a8028ba9350a612bae70efb1004ee872f94b4146;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2aa04210ca08a21e4d3b8ecfc5896fed20ecb867dce52f315470b9d8ae7b3abf924c414eae8857cf3eafa70ec5db8eb114f790070602d004f29d4a26a4eaa48a4292f33ee703bf7e3acabf4ed635d3afff401a01898e6d6fc00a20e488196ab0dbd6;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9fb98bc69c6bdefa077cd0dd0e195e8cddc70d050c3c02177a065d302f0ae4ae8d1095196c14f00d5a74b9cf4d8f44879b4c2d07bd73b88464270341debd54dcb816c06c8aebb0c400390de683605c41ad31629da0d8f50aa0afe24aba14e10d6cdc;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h46db0e69fdf98077c047bcbe893b69c9c9bae62ed928cc94b0f27c807015852cf357bd8f738feee867189d939f7d4db7c366905eb0303d1ad48226ac406a9b1a0e7574437b5b0ee4e450f50ed39b098c3d1e90f0eff9ae153b3069570a57429e61fc;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd5441b205487818b8043986d74c4e5fd228d363c86a899f18216390a52434b383aa959aca2d877b06658b3723203c2b74b5104b2089d9d4022e00d18ffd929a50193018783460112109fb99a78a1ad2646d182a724b1fc8ab1892fda3643264dc26e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h37a5329438bb1efebc0b15d5d2a49aafdca03db11e38c56f70bcd44988149fc1661e4dc3c3bc669c704b0a1670f6eb1e920e033aef2e514cc9302ea48a69ad09a24772c95a439a7a81eca4899802d500f3eb8adf8b8e8a6163addb74ecdf13de657;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha7cee5cce8501fa021e8c717dea19b55770bdccb7594463eea767b90a3de99754ae6583db122fa59db8081ac5e695d590290a572765e62a3005c4e2d5780495d130b5280a9338827b5c1c7b9caa9684824a9f47b1315224a2aa37bfcc9088e1fba69;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he7974d3ae0a6dffc4c54b0192e619d5935df9d418c3c4d8c980ffaad0a95ecad29ca5bdb092dba7a37c84a558273acff144a5d49cbe2527d0c8a362a0315eb7cc89d3ef9debb5f8699d15d51ed24255bbb85fd6038383e9d259990c38cc61975f6f;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4d4b4f1be5a8a3122325d98e11767efb91d95b4cc0c0ebccaafce797d3767a83d6ffb781376d597ca8e10491249b2898c9903e733a9bb12826360ea8b17d645ff4352263554f9ddf81028c6f68c2aa964325c59a519092e0c5d0c8040eb1fc96a053;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h283a1ab05707ba2179427db7e419be25e41c26e7ee1a57156c708451eb74cdcd8db395e0ff35de1b6e783403ef0ecb2b5c3f3173b7974e975d17c2f520187388b3a77836e14db27d1b4c253bc610f4c0b825cb3f893f96343ed2ab0be4843e28d92d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8de7ad1fccbd1fa7c10d5b696ca44025121d8238c7974808b299f7650d249d1fa2a0c730d11152a350673844a4ee33c18ad5c698099b08fdccbb78ce5e330b2c99e82fdc98b957544a16c4a68b6f2d5c3a28de0d7644a90d6fff99c8d8f29e00b357;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h388ed6465f3266a70023fb2f962475842bf4c0d2749b377fcc78713b7c78ab11986b0b3cfb0dc47099ff5110c6eaf140f2d315cff7e60f1fc6c5bfc44b6cf80eb31f396d926dfd6043e2e7c100e8ed8020e81d5e0397ab872b968b8d120c81488593;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h943ef949b70681e5f6ef6f821c99494e5bfcdcd2eff2990aaed6919b50d8680aea151fd38e27b573db43d5bb2dcc5b48effc118a4a7ad3bb762a857c632c900fdd647894c056941e77bedf4f56e8c6ee0f364c5b42706520dae877c4b85c6c939206;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf8ec216066d18e2dfe7b29118dc474930bd7e8bdd56787c565146eeab30c267f26cc4fe834676e7320ad68782c2de7e5c23bd6b7795acb5fca3e4deed2856d44268e5b97819a77894b8cd59c3e26d370ae97621b463f7d867bc83cae6dbe2013c84a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6aefc39e16645a9a40717235ba00fbd06948461809bceae877a50d864808c8d648d40a6d09e7e8e28aa5749d148a3f459d485f1e836eb8a8be19b9bbf9a745db223d8bee8bc1fd3163c4f7be95d8fd927ca2d5fa69071a10f3b328ad323f07794597;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6995a8dd12dbe0a3a82b1846e58798ae2079757e0f104d134e2bf8f688952b3100a44784f0c5d5d66e6c15ff643865d10200dafc47cea3b01134deb8c640f96f6f5142abdcd7e1376b604ec86d6b06876906ed14cd336f22ad943b41dba3061bc113;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbc3e35cc98efcabb9afe250dcc650490c9aeb60a5f145f170ac6929cf0242ed0f3c363ad5d711f837f60624a8c42c31c158548638da46b8f7d3112e4a2100bc42ab0b883889aef524a32a8b77112e132aaa3ddb1584f4854c6629df914099392f1d7;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1b5711429cb8b168b75149dd08bb70d669421ae44fd7155accea38bed090df8b1e5b56bd3245507a160023844b9d5bc5f63e16e623be22abf14af02235cf2c9bc638c1c781630856a5df2f14c6512d108b8477f3cf7599bfc3ff0cbe43fcbf3ef0b1;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf5f7e5e942a603a2eda3379dcbdbac789da2711e5b08b6b08e8f9ee87a30a9e782eaff3c96c75dd62355ef5c4836729b5119c42806063628b3a0e5ec6a7da0048559b30a061a8f8e830e9649636c60630eedf4ece84a892668e8e780379d760c3d7a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h569a5826f0b504fe970238c95626c7efb63b1d73ae25d3dd66ad352002d69d015e998ccbc4a34c26dc7d918dab14ebac0e56922f8c8b1e136f9451cce2bbb1b0c813432fc237339e8a2120f02e5072a130eac95767c7c32270c9fd20ce38e7dd1779;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbd2f767d397b2f95322bb4c98aa0f47b0dde794dc7ca7ef5ab5680ed22b0639c6a79852395e05d87920a0b98ea79f945de4b54bdc7cba008968929084e1b488585d65750aeaf88459bee5ef9b1bf211774d1a533a4210a50e1fc742018dfe878ab87;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7092288b9f6219a1b2ecf9c593b20323ccd8af7312152bd5a85513a02fce43132f37819285e1bb758af17ca2fdf056c473d9fd47142569269f3ae6e01565c0b7b25a922fd84164ca4a672241ff31ce7bec0252685d60072ca2e06c40f2b96482ed94;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4f4b2f79373501c2b92a83c30fefd01dacee5033ecd6982f049133ed3a4d95a508185557ad42a9f5d79f751bbe07ad3f42c22943f23b65dafeefa6897941ad68b6132c2d0e66159db40ebdf85a8cbe5f3d7c1bb9680b912b07e3d41edc42adf542d9;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd71eeb843d5ead43a2d2f0e0a745afd18714daa05f3ea4ac8c743f24260e568b047364b0f23a1621941d6797fa463e719462ce697636a14c3d0cf0c763ad02c3022db07062212cba03132f8344a83dbd46836a0f33c551973d897eb7f3893e507473;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc36d4121af9637523ba2b799ae4bc4388adead0e89778483d7b4438466cc60cfc9d5cc988bce4a0b69ab3438bac4c4a03c04b06520ff87545c703c0b852760afb2df1b9155acc6fb687b70235c0b1b889aabaa0fb6be0e83f7466b32cbbc901ad82d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1fce5c33b4f8bf62caaa5daa0d541afaa65d23fea219080ca72c02f14fc467b6f5545281c09b51a09e1feba135bd44e69a8017244430e7b58fa704feb0e4f11c9a905e7e07a2b1a628648e1b717d7c0c57fab6dcfbb6c19bd68df40abc3db583a86a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf12267ff5e3e4034884e2e88c732947210de34ef8b7411cde8497de1e07c26dd4913a45d075ec885758f846a5c0967e37a1db49aa511963c99ce2d59120924521401ec86bf27eb316a40edf706cb939c2f25a0502e6413b011d5938749df131e3c69;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he5ba92f1d027745c8bb99ea223f02f7c453a456b228220fc29c6cc95687eab8cf2955eea48f95e05a17e189321310c54cad7f5be842c2945efa77dc2caf9d0b5c579190913a4ed4c32081eb18dcd1d6d63e4e7ae08ce6478806e8bee238e76da336b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hac518a3bfc368eb666dcd1b85d1e8998ce37172f99c8c4f1715a9a621625f0efa0934aa4f37e3948ef5d49647a1bb68e14f55ba6e2dbeabf92f1cee1c0904c7ee75db40a450984bbb6b6f99503791b98005395751045c321476a8a2a726cc28c797a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb15c294fd5bbab450fa6ca5808475872f4f93103b9605a1f93c2338177ab74b39b0b108c889e5de37ada97d13e15d42291c3b51a4a0136dca93680ec90bf52b517272cf7df1969f3343ba423c9b8f582e7c7869d25681e56c17cdfae578c812e93c1;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7fde53553b08d98f27d5f0592e9d26884d4610efc2865bcb11379f603c4dcf95308a3bf4d3bae7e3494fc096dffe3de12fdbb47e162f3dad800624f7f39df1221e937f6d15b136bbd0a09d6fee006d3a62cd79674859cd3f289f42c6c012a6ee2be;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h62c27c927a68469406732983375e16a8bdc089287bd82b41d103288596c1bbf513652a73d508197232dfbe1fe5896dd062eca336a75b8f52e378a2a87262b66c3ef346f0acca07bd711cb2ed50e3e7d26d337baf4dc7368be152e4237f1e4d3da455;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6b72570c8cce60a3b89eda1824f0ab04bbfcd5ecf53d57ebb73415f8b92377312c0d464f8bac39421193ada0a085b39c1d005d4a337469869747e1af8cb9dc437afe524be3a14390b122f003014a58ba3959fcc055861f01424cc572aaf4f68d1b42;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hde035e62fec8cf5ae1978b0c3c917eae778981b9ec6c8a3e0cc81b3422fc98465c4f6b5055f9151e680a508c54798c70e8a137e019ba9afc04f13337ddd25b22b24397340658aa8d663fa1d4d88ef933799aaaeab99d1d022f800f5b821169db2afa;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8c2c8797d4e3aa597414507a687951d36dee7b4c5c17bfea331a0faaa4014a0b702141be226749e3374db92186fdf9c90dd81e1ec1942cd03542a57eec58739fa84bc10ec12d5dfa25e94ede844f979770038eb1582de98c45cf14d06aebe73b3846;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h97f62cbe24d5f7441dcb8032ca33f69b0f4d46d73c3f31a8bb5f90672df174276d1697e4f228fc5cfdbf7f5eb610cf856ed7a1c2c6cdee7dbbe5c2ca91c3409250aac3e37f8aab682295371f21a78781eff31f2c0b238fcf3abc6c981360ce39a7eb;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h506ab425b15e418b0badd17652303dc5f2c471f1b0dbcd4c60e5327a1fa961457e1f53d093b183d67a3b47b661db8173d7c662ec3788e5ee072f7fe256d711143f4bfa622231dbf39950583a7c8dc7cce4915d15c30a682554e18b8b262520da7f84;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc1a4c206793139d08e9f9b571da2fe38d81e9f2755f4b921d1136e0590339b03edebd44f661afd13a3bbdeade22cc97774d07fb12801b062912862a0957a6840e32214f24ba0be543cd8351b53998f59aa755e29cde8289ce6da3147cacb7b771c38;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h125cbff8c7efd63a3101700f17601bc0cd2486256a295ce60d47576230ee3bc436c42a951de0cdc2e7149a69ba0a52c98bd651ae3a1a3b4d73a69e59013fe04c5e3c217b08189ea05738ac86644a43e955ba0a0b2cd6798dff6770a5a28e17cc4360;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfd9f5c6021fe5d61a5b601b379ddd0e8704682dced2f299ba7b87589f1693e0540088e44582a6307ff38a1e004d3cbcd1c7eb974d84c98809a89eb2364790d7550cbd7bd9c3441bd4e56851724eeac669e609edcca008be19f8b991df97bbe24a422;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2ceccd6f2d06ba56358221be963252c88c493f63803820eb693d0e87b2a9c4f1c34fca9613304842894d03dc8dc615ced1e30d57d966fce6d1fd85efd1098a8dc909e5594d9ca2c6b502a9c6d64671f2753be4637628b7bd87ac04ba4a6e75f6a0ae;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9f8ab67dc3e9789d2bd4e95d33ee75d6fb42660a8401f95982708bf9f25256d16eb0b423c1dcae09c96254959f12f3038645d15a125aaa202398a85cbbaa4c68b3bed3e2428f9d7a19ebe7354e23927edf1f962c831f65e93f6ea7288d392539dd91;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h38f7932e7956d3e5b0354d409e8b9de8dbbd16b76809c077e755887a8e64aef509c8ba7cf1731bd252c866059ffb8eb2008936dad55794a9e700b0583e676f105dba99b56a9b1fa7ac6b8805f99a9157f09f9a20056a1aee8306f020a4094d6d09dd;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h532283170f944834d36ec5b1e36ec97ff8d460fc37fcef76d37c998d22e80f995467ec15738aab6b633259cbff25779b0997d9c228d190ec3fe2af4589ccbb29fb92315f7fd9c3098c894c31504ec4cb0eefff89ab5a5e92ef472e391acf217d174e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc3aa6bd5e8745c8458530d0cad7d4d3315b07110f6194daccd1eedbe089dcff16d2c29b0d0b74596106d235da145244e7a729948492dbd24f15af0f9b7aed195230a1c611fd7b3cf1d770ec3ed3c4d430a9ac37545cd2da36e296f4c10ffb3cf3da5;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7ed16f650c7a0acaaefebcad1cf2c8d5fe3fb74a8fceb5e17069181e86fb85e514d6d520038ee61a36134a1d03b6242cde3c0c70b8f61c364a3a7c26b0ff33a0f5865a59791d7306eac3b508f82494b2a2ca7e7310ded416387f567b1a24162d3aad;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4a74a1020aede3146449961edb26a74beb2638e605966e03f95902ca8f6c0e8c375235ff7708258ba088ab81e5aa03a1ce1e560461e254da2731d1d91c40338156e2ee9bc86bf5487d5f83d5e33e8131f2f2c151fcc7028b7253008b6b4cd6827d2b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7a00157a5af716e66d4547abe714a620546a970fadb03a74f42cc42dfed32477086e0d83a0ea2f4af9d11923caa5c4067145313098d227629f2e5b941a8c8ab715ecf0ec672d09492d5c1a0b5b2fd499f39c82b2df2631971b738a4252100c701f7e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h760273a2fd3305562a114a9c522d5905ad796c924dd45e4c25b2f4622ec30e87107e5eccd031526063c7d4d8f1fabfc4b5f0735fd2a723bcc4526b69e5f3d9f81159505ddea87c7e70053bebf16f48349ec0628f1ace9458c28b03681e53de30fe;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h428844e6dde51457d57f8563e6a82f1c7369f50360c628d952d765e6e3198e0e06c76b6844e0c9418e4c77f41371e5fbb837bb145ec9505990dce5879819f07d820e1a9649fcac8f448232022252322bc089f602916688e00ab18edec03615bd2c2b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf170a25dd9b7b6cecfd14baa35535099d908272fada84a69e80a35c230a1077476a53248250ff06c1cca48627e7d371b8e143641d99abea09111121fe18755b4e8ae0fca9fdbb765946fa639e34d9f54482424fe5e314428a87ce5b45261f75d5b60;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha3ccd42451896d6e8e11343a44e03efc7f2123c19a43ad940c87811a966f9e281ba698e757bcba4f0e598c3bc3057e38e5365d19c241ea0b19b66db6842841b680d7a7a1b2caa21d5bfc83c59452fbafd60c14ebd26540f2b17da651bd652e555f44;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'haaf37b69fce9ddabafe6adb5af6ebf5a3d130d951b4e2b7304f88a7e9b2c8bf19a98898b07958b8efc2f202cfe365c3d1d95a678a7277e1bc8960f9009c525d3389cb779ae7a3e8aafe14508ede2e0e8ed545ecc0596d0c05564b11cca2cd05dbcc0;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfb24721b10e7878fee7d794b5d2587344ee80729bb26e70bcfb21a763dfdc97510da2cdd6d247cca5c91d8ab8b8d0a0336711bd685c0391c230a246a3861d2d7662089d3d3d6de67d53ee718225267b013fb6e661f113064c883c8b86bee76ca0815;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h677c70074f6252bc8db7ecdea979308d8bf963126b3da694741839ac7c7a5b0b572e9116925fe804470c8d22d33bc5a0d66e587d0bc84b3f57a5b5d861c6e274d41c863b326e2618d29b160279c12eb08e30eaab83b48bf88253191a110d508fc838;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc705c73292ec24963b6d2c5d5c975b280ca6f28a5526c731ad9eba1629261970bd32c758121b1aa9165e0d05d124849706e5a1c69f565398bb725a4c847f3dcb1f8817e69c23f469cd4982e5ff0b21d9d4ab43f0d0715dbe68a2332875aae43a107;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha4d381b9a04debae264304e945ce9776390cce014283f986440cd44226d8f80582bd5e155c17791bd5dc481a9a947c514e0a79a47911c22d8ce9a928cfb902a5c3a01faa2f89f2f48c0d3eafb15161a14ed2d8aa74673559ff66c6b7a4c04ae80a4d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2f9a041250c16cc75c72498c262190241d2aeaa6c15a2560f5078f45d198ed8d2246181ec81130f42e8e8a7bba91ca15436df582d474cd7a0be311084fde70a135fdbadcdd83758ff72c332ed27f38d878cc527dcd714f0f3a18d170cff870df6d9;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h597d69fbac3f34b7b2802cbec7f3053c1faaf4a07983cd6010aa1406eb9c40bab493e85b53d7267184c3b4bf8fbf02253859d20816afdd519313522820464b6d657f15ca54806d6f13dc9266031de0806c34d7f278cac04dd34bcb7726149a9e5270;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4decb4032b0a6ed8c01694dcd7a7a251e089ddfe465078fff880f1d3c2cbe849334d36d93add1846f0093bee43281380cfc9e5a5db937d4627f2baca6a59720329024fbc3f980ac5ae8d31f018a213d277bad878c74b5f7f5781397292b0404a37d1;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2033f463a7344ec4eb0e840fb1124379805b0d0c98d3ec669f704302e1fb8125215413847617e25c3411559b787fdcbf7bf8424d0801efb2b45caf783f2e414092e11b9d8ee808103934caed53e2ee0e75cb035ae6bcd04522a4232ede2d1ea0dac6;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h567df3cce69e9f8f8dbdbb88725f3fc923466b0c5607c9924aa393cb012412ec6cc867925c5254472bf932af7b343f4607e3c10d66e387fa8ca1911fa20d5bd326b021cdb66c948509fd4126f5d97de0fd66885252b1e3d45db4b282283ce1b09048;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6ad3d20da8068023aa5f73d489f22f3ee62c4837c76015ba54690bf6b0fef33bd020b88ffd7d3a505219370dba7376d94702adbe792d6bec03c73bb1409396994e885013b63c9128847aa6b9a3612ae15085cab8fc1626d999a6e37e840030187a88;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he494a2a90219f4ebc75f4a6f0f2c9022a59d393f608cddc823b88ae69f0ce90282f6a3d220ddfc39307b73af27e4d7356173ef2edc34cc0501545c0ea60aef64f20c588afbc7f6915dedb59798e3542f2967a9d1df7b905f3fb8a154411dab270d3e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hee9fad2d07924d538a11f9ef30d29622136499e2c91b95beb4dd18d088da551dcb116325abb2781c14009531e5421d221c63384acaad7363030b2174eb88aed0a5b8079d6709c3d687d0b02b0d6df5460e4823d07c8036ed876026eb1749752be3c7;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h33d66741591e062d7904cc0ee6a646a380bfd27fb0962008765ca5041f11c360c9326be57542e9c6e0b283b25ef7c2b1218f8a0217bb2ca9c10ff4d64469d019235553c89de242dc76998d9b2b73c4d3c7eb222f0b482208ed9a5fe1978ab653aa2;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h645ccc1592a1ccc00a2263d9ca0d33d3bb12008911b6d208f0fc04f2bf4f11540a2454a0acc27a37f6f8f52638bfeb20a45690a7a7358f3a95848f532a865a3db25202e30fe6faa3593c6dd743f0c08bcea1ac62d6167800b219ff01daf50ea6094b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9ee2f07ecf345421f36f84fde075397278b3664b0871714d6f2bbba608bcc683e6ff83bb7ca9929a94b6a98e0585743df6a0cfb5d3ea99124873a41f04de73f70a02403e9be857cb64534949adbe5a7cbc88fd366fcdc0cbc6a6ba1b183a04d786ab;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h13cb19cf8976edcb4a57743961cc2426830216f466a6155a2f55b358388c475c955025fb56907b4ef13367aa2099e8eaf6ab294de0d9fc31ed3a891e44f2a563f29ee8d5321cc5b5044680f7e18796e6298634078c9c799bf3aef8ae39986b3823bb;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha6f8d5984118881ad75c628e3dbce7aad52f9842f5bcf13c990fbf20b7ab2c32200409a6ced44b55de19d059ef6bed4fa0360dce9f89179f94ae7c0ca9bc6cfde2a1f37db4da927c77c69ac3175fc71942e879342c77c76493b63b1f249dfd8e1e0;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h131bde59b16ff02b46eff93933ef544b3c3936b79b80b916726ffd4051565a181090cea55d3d535d72726f7f157d4fb4458fe1ae77f97efcebd2ce26956b5054d9042e6ef67973af982d4fd08e2f65bda7b3adab297013cbc8cf0051a31e9d7bb75;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9e05abd5364938cb4ac1bb8aab39d3b51013f6f9f86b76f45f9792c182105bb95dd4f3729c68a833d5d3653827a1c37820a47ea0191d331a8dca0a7db95f81f124287d27d22be8cbe3a6403992044cf8f9eb88b1c1b532eba97ed5f930020926aac6;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h23e6da3142f53e69015a00543dc4d6b49cad8bee5ca66f38e9ec143526535771b613b06f2c1feb7a792d19144787d6e98fe4eb19d8a23de1a6245f6d028a9537ccfacddaa00813276ca445485d86765688b2aec8b1948c50e20bb8c8c870f026e9b6;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h79510ee28eea401fe96756f534754a9e36e05798ecf888b99773e91c20d641bb7947f3639c4dd2f5e4ee990d3c4dee93a30725ffad8d648c35271445f8fe6653d2cd390c5a605c5619ea0e48e1d54cc08802524c2e4bea2eedb8ddc1384c4a056162;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3afe1719982c2aa76be4be07b49acce1db24b6f54aefc5a7029d4189af24e7e44e6ba593939add52342b23d76eac665dde62d19becbfc71e366f9e2cbc08e144aa7d80c4895e62619a4056714b6a8ddddf2b38fe7db598b75a1ed8adc1f81ae5b79e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h12f6dbf47d1dd771e1e3b16bf3c4391abc87185a8bf55263a4da955fc35c2cb868fb3b3b49e0fe2ee0065812ac9efc01910ad270edcd1525540ef228c849e83aa20481a6389c8170e3d7691c24c23453f4c826790d0ca0ced5ab67caac0686328ca2;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h455df6a4a962062a11f0c3b109ffabc76ae65c04b61081ab24a5f29698121808a7fb87989cc6eeec7b74cc9beeded3d6bb1f6da915d66c700fa91bdc71787ede23fbfae51697a85ec99d49f6fd3d9c28a9d6e18249395cc3ca6a748b4027c011e8af;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf1aaf77351ec83da97a283169e50ade0e099a5c69126ae8e2c736dbb2b08e1b3c898fe71865a74860bc30dd700fdc29841e9b6c7ad2e46589a4da3297d9621a1d65c7c69f88961f940455da60b675b477657a8b8befcf4c08b7cf60260022b9603ba;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8d7722a78cc5f7b8ce87bd05e46e9b06f32236c5e2d6686cccd81c0d84c789d5b685c21ddaba5115a45a82a88affc20b15f9e12bb1b18a5a597979df2534049f820a9885f4aa5786f335ccd024b92e60e9f93d9c2f91a20c74dc1fdfcada1fff5a58;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h24bc8585575cf1369a867ab93a56646dc7e4a58d60fc9dac6d25be6f915c3f4458a9f473382db095418feb7947fa90adad8838cc1dbe418dba2dcb2f46dcf914fd66d74143e95fabe518485f9ada73cd3caea1ce1daa6ca5df26b6924f266e525a7b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h345946d5a629fa519ad614aa11c3cbeeddf3db6893344fc31855d02fd9a9fefe8ca0e7981f4798724791257a2d0e32e9d88c1235d06651a3c72124c6c16f3c6b292ba2479321730a2f1590f95380e14c3643600dc811e99359be45c19bc49213a24e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7620da103266f4d607cfbe3d8998738fdaa1308082ba96a9f09be0bb772ed870b5288dbabe64ea32d529499ffa2f6980804a80f44d4bdf9a1cea6fe348bffbebada1006f07d14e0aefeda385c6f96c30ecae027842d2682e2256fc42a910d9da1efe;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hefd9ee0b4b6f4f098f097606816d70001b11e37335f95e3ce6ba232bb7ba3afd5e287ed77e04d87b85afb3a2a62df9e89f2c6fd440cf6574f8782df6d97afbe33cb743ea396db985852ae47b60f5d2194fc5ab606ba8bfcc8cc25053c67ce934d099;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h459a3817a2340ed5d3cdd09cf0af863d04569c18ae4ce927e4bc44f6f20dcfdbf662f6f3c76a87b13252b564560f72cfccc7a5af23d754716cbf630701e8338ae638397c7b3ed583cc0834b7419c30bbd1cda691aad8c1b31531852dcb5563d26b42;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3ca1d976926bee23b223ab0e80ab10f66224177059f67d2ffeb31214f7856faa6168aa36a790ef4f4600df9ec2173d6f4ca0730979694b27e5901a4dd5dff2af6a7ae7604ceb6a739ee94bedf804c5145f25bfc386dc9e71198cde7e624b8b114fa0;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h931838eee1497097808cf722ee31b7cd4da67026e786b9c6e7d89a6662db9bcfbba22202d78013fcec9de31991771bf2aad3faae250b7e04f8444d3aa6e4cd2e011a8b4a2dc5012e4c38daf38dd650e62b6026bd429e6178febe3d1aac55fa61eb47;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he3196c3b2f7dd92506bc6874c1ad0e9e3bbaa61a5865d2d8bc7ddd499d2a678dc91c6982a3f4412bbc7f5918e9076765b311f82d5b2f7b3a18a555d34c7bedac860ed3fb23b14b2b454fc76c07d933f710046cb9331bddbb7d3f3633236c467691db;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hcec8e017f7eb9033d3183d080c5253dd4fa5754774ef493e858fdd4150d80b2493eeebd18e41baad0ddcf5d8e1722d1f83fc37b3f2d95e7523777edac951f1f6d8f110ea74ba651fb245ba65a20033ef29eadb29c476119ce3f92f9fad2be474efef;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'haf0b89b126b20cc20acbadce144cf662f7c27e0b55ff63942c7f744ad5a42c48291f4e5433a97c59902ba5b1c32f4305151df468a35f052e806225b05168bc2b68ff757489a46aaf5217ef1f40857f9fcfd68bed8f57260391189773a6abfc9edd13;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb9cd2609e47770c36f6584b17fc3f03d2b7c5bf251cbb8c5ef72a963d7211f1e6a147e5a71eb70ba22f7a4b2253623a04cf2e2291b8ad6b8dee5137250254bb98ceefb3dedd8a33247b40bc41296d55b6c6e1174f7e47f5390fa20adb9b22c89108;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'haed0daab0f16e51f259e71a0b04a39228940c109e72eac6f8fd5fde59f97656e3b3e4aae6ab8cee9002c34a8aa662874f149ae98a1bd6c2d3e8f76f27b65de56b097fc510799ccdb177ec74e61e161a17737e69d06458a8d16dce4373cc0024f9568;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd8e334523e27cfc78d2359189114473c49c8480beab4c910260da975829e8d464c119542d89b3e38ff8bb8c0e704e37ea1b3749b30a2e7f30aa1c47e02da4819602b32fdebf1d24c54a980990fb44b930d0d4a676dba32ec71a7e405c308bb79544;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfd105e2006f3db985e66b174d8eeb44b0e6065b7c3efe60d2c0a86b92ae5fc1b7ca9e5644d4b828f19309b8ca3b6ca31176ad916bd20dbb543ca34366b41474915c3b283264d3b3e61a60ac7cb8cad6bffe9a66a7cb21c3ee633a779f6b52bb73776;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6b6645a98351502c44ca678fcfd61bbc32b9be09eb4cd1d5a36a65e96b6686f88e979927c1fea9e1f1d5f2d75c7f27bcc596fbe286e98fe863863b9f27bcdbc930959c028f8d918159b0fe4e123ada30925aef8a2f9c93c03f8f1ba5c0318fa3f06b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h68bf1823d7717f3727269e29883499324601e7896c4a35ba77c4bea15c49454491948dce65f25682fe7290e5dfcfb7fdbe09009d0618d2bb12b9d3c2542b8f60e4e60279ff1e0b3fe525db19d838f9d50dc8c23dd0445abe85e84be3a4fc1e6fccd0;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h74c4f7143383cc9dbaee91783988eacd31caaba174b83b36aebc5d2d9039e71a2bbe70bc658ada75c2e9c0d0cb2a031f66fa04f0ec40f81c84f6a2f2c72750ebac6459175db7a8b28cefcea4dd1d8f0e0992931271c6f387ce01005c0146233452b0;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hcc7a4405eedb12cc8582266f528228c49f963336dd40c7f448ad8b80f06b636a1dd982287d10e2c3e67e1fde795e198842f95f71c554d705003501b788aec004e40573afbb4476450fe74f6ae807ebf65de34e5f7e8d66e1be2e2a4c4e798443c8e1;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9e0fe5b1dfbfc4dd13d3841c6bee6a26b273cad7aa4c8ddf1c6946e5928d0a45bcc107367057b089488c82f1bfe0b79eb28e1eebbb25a0cf3764187bd3b2721d5ddb842972f02365cc8318536e1c48d428d251d2e8976c408ab8b00fa94d69dd1d13;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he8354f63fdcbd37cba418f49368bf7dd75ef342dfbfaae2b623256be18e6d56fcfee49be0b7c3008e85505ed9c6daf2efad76c9b2fabba55b9c3e7d33195728484070781daf6b65ab3408d5236ffceaa230148e1b92781b06dbcf622bb85cc9d9193;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd91b3e61f13927cf6dd45f3ee67475531b8092bc1a58e2f8fe7b483b8f522df61e7ae1f85ac3c3f77abac13a41e216311c1a44233a95eadc9438bd6e4066a5256482ed151564b2ff002d6887f80b026ffb5efeea65e4cccdb00de39fe66fd3f950bd;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h29ccc9b541478034b9bca554030afae321b36ec224562d7932963ce68d3c09061807c89b2b9abe0eb4972c9a2804049bd94ad2d75b944fd1b89301eb1286101e700ace8054a565b060f0da48ce566b27b8fbf550bc1015a81baf71f0ad92e311adf;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2dd1e674d1beea8cd8ef325fbbe96e6209bd9d4a81df0a2894ede8dabdb00ec78cb9ce559a63182f3fcdf2b4bd7660c2a316e2311e3797f613b79d0d745cdb53a5b80cfb3699ced5b091fbaed0f296e4d4449fcc2fe35df656c213d3ceaca56a8c97;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8ed5fbd4d9c883401a933469cd3dcf9a2d1d27a5cb1320aae37b8d6f56e83de515a417582d0cdd6ba57d0182ef4f38888de1d92db6d22f35ae477d61c67083f024ca15874c2f6b7463ca07c74cb3d57587f51a60c5c5835f8c62ea518f38863733f2;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6723a5ee1f88604c84d1c829a4a5c2d6aa4aa21cbff5e6e7713c9e31386e1833d5b9720f5c00eda95c77ff511eae7cce1b6976d9122cbe4ae63d22d78caa0e0604fac5762d709aa31439c2f8b8adc60a464cb0b61dd1313475ade746a1556e532d69;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5052ab430404c1b7e7ccedeadddfebf8a62d1049b81c762b477fd7a15ebe64b6051227ecf48f2c3bdd9491172fe223159601b451a27b937332db071b255d0324641c62ab365b28d6e59ce3e9da819807f3351a56cf3ccad423e90d0771c9a065deb6;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h51cccac2b32f6928c86fe5d8889747b6919865e853beecbb65cd6ed65722362939ed0106f0af0f1aa988ba8042623dd56c92de5dfc82513e79b05eb578b174e8bc59514f9832e89ec8b6d6e015ebf28b988054c33aae3d0987fab620a1ae6ff100a1;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h93f563159b963723fa7e01f7281ef09457dc9cba7e906e4eddb071c0c1cca9a2f90dae7e72b709698296ac42be9e0f3b09e5a4eb4e2e74665b5091d6b73defa24123a36f0663a3a9c5d1ab10eac87173bd2e00565465a53b59664f13350813280685;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf137a8ab632041b1b18d76afc7130566144b5c6a92ae2d381f4d3ee89570ac64fe9669477ae2c44ce8111735313390be752e98afd84fdc2d5ef873bdec9ea02076dff835e829b265abb24b65742732d2789f8a0bfee1b77c60ee446fc3b588315d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7c80af764ac819892249b9f067dd3fb8467dbb67cdd73a7f4d3d4bc3dd833cce13254c932d700b2d30bcb1094d00e7052be1861ce618999c419a7cc8f148e32272ccb405d0488f6ce659e4e55ad6c90a84e7bc4376bf23fc5d2c8f67e59c917ae7a0;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hff705824ffa3dbb3bb6e058850d89727fc2869d45c36e1b33ff604bb983e7080ab23fe7a181746675900d787eba334493ae2acc934af7680bb36d34e2c453b4cf91058171ec3a98180d02b17a8e79176a201ac33f2bd2910f4e536ce3c407249241;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6dd616cb3e31d5bbd8a2209b3b775afcf84c002a64299b18387540b34028d9a73ddce31ef41e53a469952074f0c2372c015912caadb16ebe212371156487d96748adaa789661bd40a7ebb6660f63ab888b8b6bbd2f91095907a4c43dd51c18787af5;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5988faf0a8c19432cdea9f21a4eba0653ca09e9ed5509c187f3c870fc5f128919dbe8bdfd2e2daa5a25441f504441a43aa2f95e4184d0aa256c122cfd6bbf03ab31c214512e6ce14b099ffbe3aa075c647be9710f51364e0bef712afe2faf017fcb8;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h605c656315d25712fca53526e6e067ed14ebe1e47c5e6bccc2b1aeea077d59d5c0688a47c9da0992f775b817abd8f2cf5719716c21b35b0c7317d1babc6abcd5b541c3bd9b81635ab3a97443c2475fbaa96bc552e2b61867abd5c5d4ce9a056921a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h94b56cbf89f12a8ee911610050119dc7e527372d4fa80a0dc7cd218f41d1e60684f95ba8b52f4aede59eeb56ecbb2e2cd81d8f761595265cf949777a264b218c1124207143e414f530fa61a1bb1c9a6353a561985ccc98eeada017e04e222e39c75a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hcebc925d4d46be015e172defec4a8f8c33d3b3ce67701eed0dc73ce0d45cfdff5b7e436109b9b158801b5676bcfaee99751ed2a6d8ea2bb20b11b52158969f965e2ed22f8700552aecb2c21f5050a2dcb3435f40f475618126050bbff35a6a18e06c;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6fad09e2aa599ede4d37721f99539953ddfed7fc7e96162bc8b9db9019769698d428e3e519a2afcfa49366250707a5e46794a230efde3ba37f98bb895f6bd1741d8221d79bb7b361513d8b74ac7b4f118b9fe43712a14fa974cd085a71d8f5338e28;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h79b5f9e3e2020f2a00727b0f0cde052bfed689b03c528a66de2d6901ff06f95fb9bbd3e11817947bc5b2b9eea25ef8c0589dd10d946133924e55163d5630c764b8145a3191b1e542c3b9ad6de89ee06e12157053018074eb6985189d45b30c96929e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha7f15495aa8c6fb39136d3e8ee65b856d6a9d2f30e4df776e45982b3e88e0b4bb2075ea565e98c2ee19ce15d1b21725543bd9c51a7a16809ea2c8f69f9bd3115ad5abde03ba0d042645785e89d0b5f0df97c8402055bf717601f8b3a017793f9f701;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7ec919a0d40ad26c9bfc398caaec1fb45d40644a0b7764012a7ac1b9a4011beb7e034cb0c76909be20c5fb65d21ca65ba28a91b518322d04c6bc4304d3b5beadab3eae4f3712d662abf5490e7a1dc310ddff51317468570ba1a1190c161ad9f7353c;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hae6f77fcfe1f700332fc98c5db0ef873748312d2208eca568566c1be7c6ba4fa75d1b6ee9cc9172ed68119a868ce9a8a756434399e514296cf3b8651db1da16ae441091c4dddc128e0562e9d9dd8a7220ce2f1028939e351d6d82c5c1daa9c2656f7;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'haee5f5c9a71dd6437b39a569fdbe29e897771efe629f83d4ef1d11f7a15e6875659918c6d1b8fd4fb9c95401d9a90ee68ac3e7ece2cf0703adb812af2cc02afc5bad24c4f141dfc05f74a645934df589c173625dd7397e38df6ba31319fe7ad06b89;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h66534648f6736cf8a7e0b63aafdaae426f4a0835382c97b2b3e24c25fc18365fc760629bcb7979eccee8e26acf363ffe0ab9672d2e244d8d8b4a9a21e31a28b2e69f1edde81181bf633b775c61f7dae02a7b4187767ca940d296445f3942ce73fec7;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb35e1b8e91f6b8e9a0895d776b316c6dd6c37b0f4a1dcb32d176da41096c52705ed84a8fb2df288e440eed1cbe666e0d909e14f0a467f7ea9b2752fd6c06959746beb7060ce3917c150e7b372000ec8d777867c62f9dfe7f513d75c27393f97ed64a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h35e585d6866b690c092a3e6ad71f0a10ecb68ac20d0eab7413177dbaf7ea93634e9e742c1cb7b9105de81d1daf9f70b239535f0dd2d5f9ecda9d97588cc73b429d76727b93323274db433825a4bf023fc1107e9956bf93eaec1bc1156530227451b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h195b3cff1eacd11664f8af51a1b79dbabb8f0f46871d5efbf2c655bd36e4e99c906c96009108ae3e7218fc0c982c449e9737f283f5c97054b313714b5622ddb83e8181fbb7f2929388da1c71acb6e6b6f34e0992b274f59fb55f5aaa01dab86de04a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hba69e80a38e4ec49ff689d7443b2960406404e7ec93d45ee5e5fcce334a9aec3c5a18bd17caf3d1f1b42fccab8920d28611d8be98c9a9c6296a3a15bc616f4c7a6e67e0911bf158146e5f464368c008d7e72f8099c03af0a39fced35301cde7825aa;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h446fed026dfe3d216551b4103027889801af6e326fd4221f7fd841454503952d8a3e00ad2e9d07cceaedbe21b7de9bbec3df2d74e2d8fbc597bd7a597aca9724f98ea23374c879ed06009b981a101a6a0e70e32e9e05229569a87a813298274ae129;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he155cb52e41142bf468a535a841641382551e7d5d4cb7e6d35d2458aebd6e293e46a9262a8bcdf657c9e6bfbab1dfacc0e3af35b25889801e1d6c69c60c14df7bca52e574aded88ff7e2377048a7e384b5654c8bc14161c12db87550da2896a527ca;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h655ce473076118870357f2fa05c55b3af10e1b63a66590e6376ca4a912e8c6618417cf3e72edbcf3b06f10a7286aacd289fd8192486f3abf6065521df4365febe37a21443f75aad33d86b38a22db98e6003a93ace49384ca8b3e4e614dfc6f7bcfe9;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hcde6c615172da5da79a052ad99d6d2e3859f2a46704344433540a68856028b5fdc4eac95d8cb40285562c61fe1f4642e4111ab810735f0180ed599ed69657726c16bf5db0bdea8e425508dcf9263cd2c706dfa8fde3e65cde415a6ceefae01450cb7;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1cde00bdfbcc146a9c132691cfb533f418682a16418110a72a35f8d70b859d99a67a50388af97d21813b0ec963fb339ec76a4c37400fc588df19b149a38d3de65290ea31909ceede9152da5eb8ebd377a50633f7acbca623c80ffee59bf58a308690;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h900b7153952727698c15b37db05019bfd71c070da8f056ed382abade92e18a29acf0bec9b8efe387a85471b58b18fab915e46f3dad8baa7505cb67d2f350598539576bc763306dd751fb9f067ba2ecdcadc0ba971d3fcf4b2bec94b67b93bee84ebc;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he4009f61118d5794e630de6b3a61df4c1b0e563565570369cf6cff410c73be066a1f4331288e3113b6ee4e5e1b8e47e4e9b7d51bbcfa0cbda97cabf751ad96ca82bbdcc724032b2c28d33b4510dde5092b25292d552e9c7c9deb4ea7bac5d8c4b67d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7083d238ec68c7573906c4ae153d107e77cf72c1d59661001e437743e20e2b53cd6c277969e4da2e927483740af3d1a022571a406bac4e70e4f947f472fe99935af34f2569fed62f893678f39c4f67bd13ceb4a87ebead2a55737bee66ee5590cf13;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd3fa65edd3223cb993e374be2bb66d5d7a27fd9c1a1e4b6ee5571455e092599b892f840a62529b0de77cfc2ccb164b27cea330659e64a46475cbde56542bcb88e432824c6a97e6c6bc04141517da035c6f9df8f69f472c3e99474af6650cf23325a7;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3bcbf875492150565e74309ad344a4bb53569dece005d12d17e57e2902a952449b221e3af07a35332da041e0a104d37d547b2c28a2a3335ed3ffe9380283d596d78905807c3dc611b7627ef3be4e78707e24361a4baa32a004574a3d252e70965b77;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h66895a06b9bc33139ee50c25f00c79546adad368e305a4e6cf14bac64c6c30c39c80992bb9883ac3f754e9bf1a637accced5e2252a6be810f569cc14c68b29ec203e206fccb302dd626469ecae0ddcc036c87fff9597e4545f3b94d8471470c77417;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4d2dd69647d15bcb0d6aa272ee0390f0d2957ea9b89aca821da7ad8642c7777e4ea42c0fc9558e67c898ce5137dd21f29b0415bd9f59326c193f0ced03be83fbc722f7fc43ad42bb88c2e818feaa3a1c9482d6087cac2eda7b53c88a7513fcf90304;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5831d8ce01258531c6af31d629b6739455f06804d358bb888e6b72e59efc2783a79025edad3040818f69ba8d8da16ccf57c6e2949a51d3ecbfca53a83da6fbf339c415ee92336a5a828e5bef6a1cfd7bdd03bab0fb5f5414fb88c92bf4de4c807e65;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hab1d2be48ddbfd958599feab812b4491b076222dc4b410b4d072b80b6ce4c0a041a433836362c4e49e6c85407738046ff9f2ac76c0a5a3399a62e9d3c4d098f01091634463991f083bd83b1354331918028e4d5ce9c0c9c695298726daf144e97552;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h487ab518ca8cc4cd6ec9fe90039d6550cbc66610d4bbf65321a48f3013fae953801eec9a1e3e3493a48b9eea1acaaf1bcb5636b6810dac6bbac2c1a7e699e687aa17a72e822c6b7cfdeb199a0dda9f0fab7d900b3baf3525bc9a2dfaaf1bea86aaab;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7e9f2b064ad9a3cb581816cf7d072cafba1d9bfb3c43c5950bd347be3532287883d7c6f541eb454e1ed2bcb772dd1176ca1a21b6a89b2235ef85e70d24449a0f077275f3d83967326e91441c4b0a6383ce6ee22404d6b11663a11fdfdad56fa58631;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1802163ca9aa8de3758b2498d9212f0cfbff1abada3c02f4856f12a4cea8fb89a909ed7fd277571cc8f103faf2d9ab745159006ca67faa8d59122fff6168dc0e288a4e0a2b368d61631d013cceba33e06e4d13d16899ed5a34ad07e551711b0a3ea9;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hab05b64bb2a3bcdf3461efa99caeb3809182b484149af20b23a1deb74f46cebbff86c2ebc468b6f69a44ee00cc4a0ae0f33d93d40c09a0add2d70d9682ce043294bd324692790622a504cbed545c01e34448caf7bde8df4732879744013e8603f4c7;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf8640e6f391314fe763d48cb70a836c45e90f06b54998e55589ed139384c99c36d2b4c48d1cf8e7de6b2508fa85804786c32163663a473c12782dc9aeb3612625129daa33c8c513d7261d4c01e1b330456b1ba120400dcc7a77f11d2145a1fb0f2c7;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5585fe236a97f7a22598f78f2bb30b95fccb9b811fc24190b497e3a14aad32a7fa3be8c8d43fccfd9ffa157da9cd6a9e94801e89a20ddbaa9255b8db720c67746ef89613b32ed659b7f1913b46964615a5e04198171f9ac03d8b6bcb2bf9193e2c0;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb5a6c83b32da3768b5639c7b26fe932d8cfb6ab56c06758487fc532934142a8a42a2a134c54e50e97d02d0ccb11455f30b3a5baf84faeb410f4bfdf06f32065bdc088e82e023501c74d92dbdbeda12a8f27e4260c3b01f9fd893a6cdaf368f3606b4;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hef61d2b0fcbdea6f6dfca955bd1c3533b04044ad36360e483d09cff03e95e6a13c1d6dd676c09b2b9bb489803ca4f401acd10f5ffb5db32001b8841663876d4d42b6128eeec6b648330f6e72e08347775301c67c790790fc1638185e2e0ebe4de4c4;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h94e21f8022980c1760944cbd5f963f91486a2d42b494f234d18b1d305a0982e793d72cafea03170b3d9359c484f3e2cf4348e6aa57de47a084acae853457eb323f30ef0044a0077cdd41c3b231c1c9a6a258de48b9a3028d99ca786c8e5067501174;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4da5c052db6960ded2a9f9178f8e0009f3ef91f05947cd2cd3bda48bb3fda638e5f7649851e92935900bc8fb6f1edcd9c9250eba2b8093774ef0d1ea60d22d1579b85802bf660d37adda58e87700c4eb688b0473ed6090d33aeaa982cd9d1685bdda;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf86d3105d1931969c3cc6f44e0dfcdfb8d4f710b880672dd7e769b17266d15b5771abf3467e2a906e1e2f2d3d84348cd32c01da4b0c719caf904ffb8509491d5f36c7f4604f2e75e38628553054b8e6c3c85d57785487b7f512f0e264d531ea3bd58;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9b65ad5ad821bce730b93e0b3a09fe8e73925d647519fc3348feae3daa441cd7462d34c919c06340de96f0ee9b70571faeb452c1079a8da38156385bdbd03bd9a5b9631ed838f30b0a9938c65144ce8cc5646e957c401e09373eae963afd3e1351a2;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf687cbca306114fe99daea67fa0f14a68adf6582d8afcd54f525a63c826e792d1073c4bce6eda04bc0dc3dafdd8b26ce6aa5219147413a3482fa4080f03bbf0606c74cb2a28a2c9c01db64f2a65788342a06c8720d24dc0ad6f181721bbc1a4ab8bf;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h49ab64d1c0c1ded490f2eda2d1b5fc4fed9b605d28b9b83e4bbf1aaf8154648e3ce115500c171eb81d5c5e1ae9ad29cf14cebd76512809c4b20d5e19c973c7d2a8197cda59b9eaba4989a796b37b0a9ca6620d2e3b86291be8d0ab2a2d68f5711a46;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9a5a0e52a579af37a5fff1145e3e4a22f947c580f23a92f6a484dda75a34a8fb5e520c6386adaa27f61442ab1a0bc42d869d561f569285f33c5002df2270b918c346526c355b08089a49071bdab6c9e48dbd2f49275586e68b5635a3a7c167748a56;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3eb1b22cde1c7e4f62e8cf206e6c346856cf7195672856190bbb3992bbbbadb89514d60f570f87b6945a1d197ec81b3a48696f22450279b7f5e2ae37596854657ecc79a0ea2783dd8442fd0b21e5fac697e3beea1e147e8a0378ea73c0543f62e608;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h611dce29c839b2c201a319d7bfa161f54034d9fd41368f2df52931590785e20c61454e1ffb96574453a854ae14cca0076c2e9b11cd1cfe675be7095737c1e4db51b0d8aa5fdd34f0178f837141580316237048a392c224dc86d7c900dc796347e748;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he053d829df67e6d85efed61afa63920a762b96ef0a9fed7713c00cd557d5476d286723d23f8438a91b42c4ab5daa821ab0e3569e856d76016580e2a7c24913da38b6c309b1e32095180e086a36f7d6bc8d85bb858c8ac5f99acde1a018fac695a444;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5a0a66f9f29db8b09cbce1d85008ea70ff0768197ac6acde0b916ee44c02cb338191096c99c65878d1c3257de7562200ecfcabc0436ae28b48c39306dc94a3e78c53a42907436791e4efd63b1dd3897a88fbe4a1c624acaf956f0897680b910143bc;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3c02c52d95f64e922d5e0ea1ce6daf78b6a2c688b0c66e2f27a23ba416e82e82b93ed620fd66b6e128f0d9632ef1c033602ad46a114d3ede47c6b095a3ffb87a31f44c5e9970a0af10fc7c8d01b0e84f5f4f51fc7b8ba89869d7ba48b3de505b8a76;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb0171d6823adccc5fb38b3311539229a2bcc2aae7e2de232764405b212d628b2ae1f253d574aaf023a9135f65e31b274e08b26e555eca042a1ab02f79639bd012e516a44896eb1a5a56bb0a61e3a4ab203caf5d76fd33abf40279dd5523a58505077;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h768173818516124f90f55e51732f2e88118d8809afbc62f2a1b9d85159e0fe1aea6bc8234c247460c8a13dd0d017e5cdeef89d81fc50ec963ef6869e1bb268a53bbd36dfbe895c72cc971bfb844de861fef804e4eca4771e10986567a39c11f0ce76;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7324e86cbf6cb12d7211fbc4ed50d35219d8594cea35cc79df0c31bfc496b21e8ecb37786513e1ca21780a1ec0421e89ae6f9ab3074ce3f22b28f06096e9b078889dcce63e1ee16c38077b5dc4fca61bb77cd9c03321791cbdbecd6bc4ebec7b542c;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha21de7a05732675352cba503c6ec54a02bf8595cf6ea6f9c4d5a90bb8d4f8f2a9d9e3dbee8649afa698a0a73f95f80cc17821bbe56a0ab0a346659602d6a309d3d31eec0aff9cf5548f873480689ffcc41d95103498caf71105161ccdf8f3a8490ce;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h929a4fb26ab6fca40e5c663efe34b75803d86e029c03c9f5e9aef09be933f342a1417ea029adecac85a50867e767de69e9e2c58a04aa1a399301ab2d4578599ffe977d0390ddeb7b4e89836a7d5b674ca7937b715f7a84cf62ef1a05216bbb70b98;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he3a70a923b0dcf757f9e6aaf6a4c31ee3e19fe5f5d21af74cd6a35aec55effb8f1634654871b5a8388276caa77d63fc80bc40fcf8eed1d00a91e5f3c72e5b07bc690169f44f3a875fedc7425aef55d8371c5d56614e27f1fa30b4b07351611723f6b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha8c2412c644390eb901394a2216cf5a045255aa8bb28330af4ce5696eca6336e8d98611e6bc0fe58610eb1d4fa972f77977ac454f532890e2198f79355fbbfe392bae9ef754acac1c3119805ede018d6aac36ab27ea934877769b35a84ab5b732461;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hca2da58e68725933d7cf6999825090516f06a35c9c8d3771e6bdfb8e9dca13831b527fdc0c1b07ecf555e512c8ecc4543dbde7d6ca37882dd81623608413641563af964b00737502c3306cfda21c600aba62b4fa0b4d505d27bf7a5ea840736a6f95;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h146d763716c33e305993856b4c11817fc00f2cba49b4c19faf270a423b09a7eef7c191394dfd70d20f12024cc22d185eca07709fb15501b6954063c82117d5d027100691de8f23a378e22a202add01f44e6c58cf07b0642f06b81cbf0fa8a5de3519;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h86b4368b9a111ff867b3323378b221b05157bf75f161bc54a8f26b3fdfcac1f5661efdedacf7a37e0a545c87f51de2008ee3e9fa4ce7fd8310e8dc31ab0d500bcfc9b3686285c2c89f1e827ccb89582ec77a197da67de1eac5840ab5ff4e61534ec5;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2a054e67b9701cd586b8751bbc6b460035141fcd1138677f41a1f5403899f369f84da407f94249b1ef87559113757a58073e44b8b1ab60f191db1b8fcd70e5e970b157a3f1b3abab08bb07eb064ef3fd72c588985476017f3b5ef81d3e03b04b07a0;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4cbbec7ec5cb0a3f5f4d22b372f780d73a6c95b8595ee74d322aa6f20a5d75a78a7ae751ef7df8bfdcab16b2ff9bb86b2f01e708eae6f1cc211e03064c1f1dff29509f217280ec6a6c9147a81be375910a381833a292cbe465841b76f22cbc2fd4f8;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc3f1382ae4ce00669c2e2271ffa4eeaeb5111336d4ec74e87963dfb1fe12756dea705970a423e08b836c4122aaed46b3cc0f23bf202087253a9f73b119869b1acfbd76d6ddebcb3297fcb2d56c10e65aaf574a0b432321d92639425c13a6361ae0b4;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4aa670632e610c77620e55127becaea6d1c56baead3127065f46d9fdeb19fe57dc5feea87a16266eaea3e14345d04da740d5ed9d1a43ff5826f7b3a94728c1e5e6146a1f49e6e601aa611502e245967a477e114e5a04faf21cc085eb6e9308915a57;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc5db712b1468177074029a2224946b78badd338c99fa4f68c5531a28f55c6e7e084173a7f6f3e24a957d89716bc031842ff2012357476033218e414d404b939cd419576decaa386340a1e0e5f52fcce6e73454c28ec5f1912e54235929f898d92aa5;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf72e741ecb2e08575657bf4dd377477c4c10532665fb7a1f9f657e874dedabae839e02692d4c94c421f9dbc31b78050c3abbef5e8390b9e9040304455781ab886a468770e829e3d425874b9c3dfa1b09fc2884fba79235c7c5a111bc01d8a155585f;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h41f4f14ff06b4c7c6a59d27ab8170fe43ccbbd9719d6bd8b0280a1022e36a2321bf2b930530a926808b036e5335ddd044cdf3f989d994fa8af074a4e00965f6ba187cf1924727ed54bed4c3923aa141ddd9f185812f49168262fbfaeab92c28fbf56;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd1ca3999cacef3d0ffb23977baf46a2d09623bed4167a7e1be7800bb5aa91b7988aa68943242f69eb979c6c7a8da0480a7c7b55a54c5f17e93aa9120e46b500c349a785ca0b7e327edf5c9eba3ba7af21f326be4868aa0e34e3e0081f2b0b2a5ee0a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1a8b282200c6d55e2989efb64f59e124299d49fe21f6485d9b4cd8c827953f504f03b64d99b23cd49ceaa87dca331eb5d1289901e98da2f484b5a577e64712e372a3e9e4c96597286c836041305ddc0a06a1b25e2a473f414f3060e8207a1b58671;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h23d33e0748b28cdbda6d6288cb6e5f19669967b34ec4ca0beec1515c0e7f1370998cecc52d64fc1e7dc7fd17d186e9c74bbd015aa81d8ccf48995d5f1ba7cd0cb021a12b39f651515f9e265b225391e70ba95b31f95902aeda0ca077558ed1ed1629;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha0b93a2d83eca4ed88b2b4f839fa9e07b2a0a88678445fd6d0d3976d531ad23232b18109208472dc8c6ba05815dee0261a41f1b7670be4aa1306656563278a1bfbd9b3239bcb3087d9a2a21046db84241c5051c144e938a1b8a9a25dae595c365ada;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7bb5a7c69402747d22dbcc93e91e5b99e3e338db041c71b8ad0de0671f5ac1625d356274f8f7f3cdc6b55a11aa17452eab3f91a3eab3d5f6f672877d23d1cf87deeb504a6efd0fe743f7d6bd08d11033b906b8a953af89f12aee940591dcd060d47d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc9e5b13ed18d91a7ff4c45191df1aa46f52763d20da00ee13da0eb3671caadc1af15234c2a76ff43742f26eee3c7d83d54e7cbec730f0c1372caea5266f386be20daa9378b26bc0e79bab0b6265ef28f5b0f2721e548b4ac1c6cecd894b14758bf92;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6739e3247f7daefe5697fe0c18da218e95ca94eb4706ca652153b5293f48fb1053129ae820a08f8d092acd6ce0bf5499da122ed7830e9d7dabed344ec7820a4939a9cffa8daf4e8b2ee8b5e22a40f9cbb4643acbd771f003d8e561019d253db7cd66;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha5c27ac6371152c6cb5154ac8f4349fac4e2df9eedd42ced7de872c3d239fad34a5db4a04d80e9b62cbea9278e2ba003afab076f955e63b9f4c95dbf9e246e8ca38a8bc2fd519757aa5d7b12051640e158dfea46dc45f29c72eeea416670685ec627;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2e89fc02968defa94f434bfc44b9bac12975cfb43ae92ce4a708c1e3f6a90ae40a90d490836b3bce1ca2d82fb3107af8e04e0e3443a2c59dd00d45155f890fa4bebc30946252d999dccd681372c408a7600b4de59ec9ad86df3277cc43874ae40845;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc81cdb4e341dacef1b1048810bfc16ac4233b6ee8ce01ed66abd2ab24a636e67c786e70dc6f657a766d81cc5b04b098fb9087cf3745dee97af5c1594cff32bea2fab3da7237509ba1ca1e97ac44f7577a84aa629479f2b7cec30bea895c400a2912d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd067f4df3979ee8891bac0fa7d7517a05cb305311d3d7c27279fd9f94901fcee2848939a17d668039842e7955fb22bcb66cdc18f4524a562c8849f44533b07d2005506c938e3816e7cadb44eff104b4c03a95fee4f95a99556ccbe76656f29564f8a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbfd4f9bc06bbf58216bc171ee38946c3a3310a209f0f5c5e1ba0e2c07dfe5c3658d0678819a2cb16db886cab6165b6c000619a76257058e36a5469d36dda7d78a4dddf882f1ec07060198a44916c156951c60f06d78b9b9dacd81fd2d7744aa45be4;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1efa075250da6b775a505c6ad0046144fdfd0dcc48afc6c8bedcdf6d995d0da54890370636bf16508d22a2dfebc4afeb9b89953e5540ee066716ec1710e8d0dce90a0133497218b54f02fe0351a1622f6038f54d6754aec8604ac60cf73b7897bbcb;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf188e468f113619569b6ceccceac6390d54ff0b6a7c2dc7a36edf3bddda41705f6b402224f95f129897ef2f0825a543c9cb6e0f8a274e3a0e79e8e47bd52f7e9a20fff862b369478c4960e4b20f50d5959ffc0c790102a72163949a9f1313ac9a58e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd9020baa087b9967f9b6c408af5344bed16eb65881ca5e5a08a2560ce03252ce040caeb016b134dd19c9fcaacf50c988872b9e322f9c5690ded5f369b395061d836d6982db877f8a5f78e1477e633ba95e3b1a8d2618296c58027029402c1b0c32d9;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd57f52f5983ae4dfe7b769151af1957c0012a2127b761db7af9638fbee859ba6be5bdecacc8b4c7bbf6c952710b27da505c0cf29721378aa4767f039adbd90819776f48903d7c4874d28408df6069a18501aa1d53af03a49e8b52e16eff468adeafc;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf3a6c2fee470e0f1dcb4ae257f95c97bd57378a653053dfec256dea1c65ac7fe816389454b2e62b090ab920c515ddd60de8947664d44a02946ffc04864445c25300d2eb7da6a7075b3592390c4d82aab2b84a1acb1c197307673a03d902087cc0a89;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hea2cd143c9a7160c5e031397bd5de335618497f1115218214a422a79f70e4213e34f4e759cd441c78e90b22bb4f0d9d619e4c051794be9dcc6b37aeb4a1cb30f0b67ef284032961b0aa6228ff53167ce4c55d68a3c107a480e8ea6fa8a5267631a9;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1ab149e1bf877d706b20bf449b681dc3ab25d30804ecd91e47b55cd9ffb7007e5021ba528c7f2bdf2a086ca56f0b904b36ba04f4647fbe1b958ee9790df779c5709933d687aa955c120e52932c140256717a8490ec3d1bda778ed433436769fe673f;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h790929fa0749641f6f1de2088ece40465201f4d6052bf49035bd2cf1d5b5cc32f913870ed4adfd1e90a6b54d9b295da8183233afb14c445f5a1b0542711b3e9847203fc926f1704f55f3c13a2062833972bbc4a7a9ad8bde204c04dc7604dd7b4e8d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h265c0a191cccd0c4c74e2e3fd6b0878a3d262b9709ff0af5e974ecd24b66ba3e1c02af1cf117ce099f88b0dee74bf86542efe2b490419014827aa72375e34c5b990c5161914b9abc7153df8bf487cc903909ba693ec5533b02c14df2b77aed4fbe86;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h771c9056d66bc73fd62b81e4a5e890575191bab1d926d2617d8171b6b72cda11ecccb6086cb3a525df6c9e3690d10541631a78e32b7325af52978d3d533a98986bf07782ecce2ebcc5e3febb9644849b57bd1a6fea2f090a79e2715e6bb566ace6eb;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdb1c3ef670e4591f7673ccc100cdc6526a8874ad94976bd3bafcc09fce9a6cf0c1b2687ee0c430266e79291530733adca859a1ba2631eb6e15b43605902b33738d1c530e976d69f976bb91a272703192d1858c76091a2e09311cb2974b8f168ab76b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'haa5221468ddd99c80aad9ec4310983cefaf82328c10eb1be18784c94f8a385a24a2a5f580b03040cabd28725b956e2eadef6a95e009e7e64b1cf3fc6191530f37f966853bf2e88154f46e216918d87f36ec76328c88f593f96cee2f55477dee72d18;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7b0e1c232bcd0928daeb0e440cc0abdc3675d00f29eb1f376fbd82fc35bcd3a200c29b97ebdc6c968d750a41619b35d8a6aa4e7d9b01c7f5bf075b41d2639a3b098ec9542d8d4bf45f8279351c0883b5afbcd412428b671a583f2e9d44f455077144;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h581dd8cff6651dc584ee7967ae95e27f1a29051d9ec4b8ee4d09ee89729e31765030018e11120ac147a9242ebec10d0cfab138d0255eebdf5ab160e3792d4cc49b05d3d888bae6ba5cd0b79e0799ec6d318dd4ae4ecef8e26ccf560bc15d37dd626f;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h146fafe221f051027e6ba978b62ad22fbaf4684cf51e620235c3b716691395027a48cc4ca770a67e643f3aae7599f40f43794b229a8994f083d335fd47ab21e1a8826bdd28f75cf21422dc8dd1752889af5600eaaae3124478fc9665e60192c8c5a8;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h43885a969090cdb4e83b925af75bbe3357821c2d8be032fc4820b275d39ad8f6ef5fbe74af9f1dc1567bb203365ea19131ef7adb87cd72979757107613da09521627b7f5cbc71cd5798db8bb41d20d1751b28ed6f3556a08a50576dcaac11c6af3bd;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc4d3b7ab865bfe5bc33b14155ddd3cca774cae0ff3fc12da91d912109e74380da3dbd96a434e3284b97ddc4651e55806c8757c1fc2af7146dccbc243c32cf0f5e21f7877df05549a8fb81ddb56d06bbc075ec797c4f8fed61e428e9d55280be445a2;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hda57eb0f1d9a13eeb7459ab2b603a32e92d68ce6366899db183778cfd56cd6bbd56b86b4d35991b4dd09cb8ccef72a4b60f9b70b259df24f8f961401ada7e545d38c0ef5fd51dd997da75beee4152c867426d2eee9512d5e0f24bcb65bd829957c58;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdb4d6bc2e3a5a384b255477e81470758b9535f4dadbc66a4a5862162513d0451af41d7c6550a10f025991db2ec1a440e5ba4312e63fc4a63156542cffa8edfd5c2d1582eb97520fa9075dc4f30bf08af11a2dc7c10ee45149cee5d5d15c6e2947a35;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf470fa93d71fc03455870b3a64f5d3e90155144f15f0481670a69abf2328f7e5f7a84aadae40c30f38bb31ddf5199a9534822531b1f1f41d01b2d10e39abc7c517f0aca8f9e833e2b0b4b7bf257f4f3592cafdcf5bbaff3eb41b7ddccba6f4726cd3;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbb2522d7f6f8617b365812a9f91d8ebff22def68275d9081dc68177d12301812a80647963b628d63ee0004c0ea6f85a635309bcc90a2c23bbdb21c06d9697c5cdb3ce1562095deb576dbd0d29f54e51e167ac8295d12d44914a680bbe708a86e37bf;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfb90f7f96e7c588fdcf0525530aaea6cf8904f9a0ac4732daa22f7e6c71914530313ab22f9eb91b12cdb1a916a3859a7b87115f1d4600539afc2875d8726d71ca457d8e4dc4e2d1b7114deef839125ae50668706ee41477b7b4e6e357bcb25823810;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4ffd9c583a6a85664f86edcb7c4824ca862abf64422779b80523910120407426991cbba2b8bd8a5a5a684f66915acda0df45bc6156faa5293630960befe84da2771ddc8dfe1d708e61eda5ed5a345b749c98b7aa3c344279d54b7cdf496b25b85046;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha2ce1fee0b262527bb11d90bb78dfbc3bc588bbdde1fb26912fc56807fb1abf1fc9ee663384b9ac0319893740fd7f8c802cbb5dac54ad48ec3399fb380b27a2a6f31f018bc2c1783a6379553bab1c80a76c5db1ffaadd6bd5a4a5c58f33c3aa46f84;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf6ccbc9c1c2bcb5c68fe58dd527541b93ee639d4bf9fbba19abaac9198c021e719c58a6a432de2409fb990140aee8e7977612047f1ce4b349c4ce311a854e615999861d6b2518c32e618ebe7821b061994180601ba13ad917af300dc732fdbb74b70;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfc791c234b33c95d86b3225bcad4692fd4d585107bef9a574e432ab2971b41fbc9c45d970778a40e4bd79f992008eb321dfa0dca5ba92138d37474e3b2de2c69f1b7581c4859f1d50d601596e7bed82e15210b9f95af83774bbfc388f344d33033b3;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h44cf63e01d16261206f9b062a24daab2cc6c5044b26f950128045db9749bab2e1e7fee0e375368b5d765edc43a8f642c52bce2fe91df710dcf0a9af607083b0726cfdbd4d11c7ba2efdce558aaa5334dfba6dfa101051e85e58945ae0f7ff05810e0;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc44aca3b95f4105f2eabf5d1508fb3feafdf3ac6402d00ea5eec8965f72b0de4ada6686f789c81396cbda8e5a5cb489d07c5553e781db2fa5d1779d536b26bf0328fa4feb33dfe56e7dec7f3a1ed3faeb612601e2f94f133def6c511a2a6ad3ff3f2;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd51a0737e5ffca3aa67f37feb051d1d2c781a6d21bf6dd287d7f4ef41a4763a7229ba120e9111e2f17ad3cecfa054b46a8c234acee309c80b150567af34d1abdf085bb3da6954dbf5e0a2941897c6ec2c5c285fd7e6a0613ce921127a75639382af6;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb8916ea209ebaf67830b62f2d20b73e8497e148089bbec8246a05bf1e54f75099794e493f33a6c22972f5b6849e1117e901c00ca35d06620ceee6f04dd70db448d406febef6f955f67cad3f6f7f25f65f1e56d97d292c885a23c9cfaf2095fd0b278;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5a41906027bc4ad5b1042d4b2d0f1899b195ea4bdd1c9d35bbcdc1906ca1a0effaa9d12d86545657fb2d37f8c2526de84aa4543a0cbc97b654cd2fd42b3c364f1f077a48fd48e27d0486fe58de6f0e2710a9cfbf2f8cb695ed9e4db115a1377c9ab8;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdb6b73a2ab0b7450c506a1e4f6d6bb2fafb9ed19da8bea09304ce8b22957a273dd8ed7873252856cfbc1da4305e50ea49b4aa2fbd4e3706d67c19455a1fe98c8a0b14b2263b42f1407bc3b0ba8e3454efc27dfa3f9865d202c0140fa84d4e7f9c1ca;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h469c94ead593a4d00381f206cc88bcdcab241014b0fce960e5679fcd9f1e511a45f9effef4fbae06085a687cd2e95ec4263e9e04b7f7d0efb0d5b61658ca1dd6e1c5379c0a1f6af409849d2e13914ad23b3a001133d86ed15de2705ae25a85cb303a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbc746f88c7c453f72ec1b552aa891ee47d8f7c1275a9bab2c1b6d2ffc760eaafb56c790b0189926593b88ad89bfc91d2090fbeb29425b61203b2b5accfaea6d107b97dc695111dab4712329ca6868effbde58a19b6b88a63b7e368a433f3157cd113;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha63cb08786e33f5f445f52643404190a50fec937a94d5f3db647d095750bb945b22648d797e71e793c12500de196ac64eb95bd58388e48e61dd919433687ec929872ddd91137e967b3aaeb7fa896db746a90d36ca0a922546ffe5003b07821d5db8f;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he57ab5a348ddada8a0caa20465615c66b16652ede35ccc4c8daa52b2599bcfbe8f9e2f2e8a5402fab2d7436c6b5656b910a842c21e7f395b4b13d17e74c3361d371390a86b724cbc92c40fc984a86e6ba086710e896fa659bbd0c00cd31dd6ed63df;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h606b08f5dcf3bc97a79e9eb57ac950094445e1594bcd4c2332df7922ffb906fa5d65497146423ad6333fbb8f5417fdc7cd3ef9c4ed12170bf0652b94c717285454a08f4baee4d7ad15d8a37eebb15be3d54b8f32360454717ec11abb951f7d47712f;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc90e06a487065ffd0ffb5086d8cf3c8b221714fb5ea57524830aaab59846a99d9eb7e192a0c84ca5801688236e0c9c99ab564c238f8b915d37446f3be07c2c13437108890f984b07bcb181a81987a5835dc23020eac4acbaa7d327973b2a265f1435;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdeba82823190e31f180093ceb3603a6d10fda39195941791eb9724e52b77c1d36285aa885f4d97d35b0aed8400f5d7e903201f5fe4c64020c73a12f1764859b7f7ce58f2506fd4e3f59949637a403e9505aa971adee100bdae35fc2378fbab9b63;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h93df0b937b538865c2a2c728bf4b9c76733dc6db042d2c4eef820a65b193bc14eaf946490db990edeed38bc6c2a681c61bcd3b246f5d1fa77f0333916431fd38a80a54e7f874ce316eaa2b6e349735edc2c70687cd6d5c54db35bb83c1faf5e0bcb3;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2bb8e433a4a9cc7ea0ba09153ffeadd815220acc7018e2fdeba6b71cf9a1517f339cd392a3b07ab91de6c7f58a050b5f40dba8f104d5b509483a99e4708bedd591e98a5318e0b676ffa5677abf5d89d7cfbe7a4fc4ab11f91e3e4866994dd1e02094;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hcd2b368bbb679302550f70726a2a945e5388f1b488a11299a1e22c1bd93acaed49fa02ddd06e131c3b981535beec1938d47ced5d583a3962a2b41246b5cb94a8b0fc3c97f4e3ca223a0198b23b63c049d3c269f899b32a46f8b5141dd2006ca90e9b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1e5cb77e77f5b3cd141ea9949373264e198fb2916c5a5af6d40e60fbe8e5e5426ff449a0dda7d37dede293df8d593dffc5229e9b11d5c957088fc0b3be2cad83dab190681c71efc3ba8e89b700a438c80985ac2a3ec922f8be32c9861a66f55ef29d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdb08237e58fe1aa9d94fff4f2d6a99a6eaecc3f1b94652f54a5ce5e4a81e08456ea7d7e9ebe2934665780f57b9675b607225dc1d52a5cbe85b5103c2437916258b00f055cb0c4f0ad44c298bc49a5b4b1fe0c9a24efa186486a43d235a002951ba2c;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha234007dd510460b65b9bebbeec1fb4348f98238729609a262531e41b6806b94330884246d9383b77cd45815bc425cc4f3342e235edab44a216dbd97862636c8988abb05d2d9b11acbed30ad2c5f33ee56b8362a74e571b660190b1e943bc1cc5e7e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha85e159165a44a46aebb411007642bc087142044a9c0108879f817fadfdac9ac5a825c6d339509c430274f195bdd464790f93ffaa3e07578038f784ec72a3c68aaaf69f1a80147683181b8d5847c21f53cf867796264ae6f10f29b91ea38d759e306;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h747b56341440be8128b10d831a90b928bc88151641e473c2ce1fb8a5d0c3518bf035fd77a6fa0ef0c10bf991f5e590dab41da2aa054ebe0a1a4eda810ddb1467c65e319928b4aff0cbf1bd9c3cbd04f2647d361d09c5a037229015179ff0cf2fc1df;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7f3657b951b3a3d257b25fec8cf91b6a7b4ce24f441d8b7c71efd7cc04532e83b8387a5a9b8f613248b6970b405b2e5f0d287f25f18b84bfcd70a580cdbbc55b93ef1a7b630bed43f6af3daf98b9f7f87250c02f3815ee0877adfa02e50d49acbafb;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h33f012ca3cd4d3ca4ba0cbd82eecce0e162e7f5a799391c3fef03c9b883e4de42a2a4fe4a8530e2dea926f2c6271f7ec0811c6afc8a03ed365658bd89f7059a4c781abd1707b08ca408c20e53b6382ea30d9d3c34747fda15381a97684a0bfd3cfd1;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7b9ad7fbc2662316682bcc62353b9bd0b9d58b9975c9a4952a928996f785ea481bca1a5dcd4ca1eb54b7db456fb7f57897423c8fb46381afcfac59f27380084ae5f02608acab5645758eec0460fc7e6a9a91b45f742bea86be01ae670bd6a0a9884b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h63f0123a4d3b1972e6d59cda2066b6af245c69d8266c7aef7c998bbb0bd1f0d912609434dc0e030da63d7a14b2094dd9b81695dc3c142756cd3675a2e9f79fb218426a5c19cd9999f106004d65671ee12429bf72db8a4ca85d70ad96bc8e1d1f9382;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h78482c126b74e5fb72454657250b6eea14e139e88e360c0f307a6a6d45ed9d774388efdb31ff0624220bc3cbd753e88f8156f5a3f45b200daca43983dbdba5528556f373187fc18805064165e3d45eb9cb12ea9c12928eea65ba070add854647c8ec;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1edadfe60a1028839c209faca279066298a0c2662c860fd105a607b4ff7d575fa3aa14fec53b9d912f4f246e8d383a53ce81d14c05e2e8d7206529dc3b8a5135497d9b1f2ee7220bb4f9d74fd6b86e0be37f9c27f086956158e91ca7a1fdf1f66ebe;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf0f665c10f55c810c7b475b504e2602aff1ecd81d61dcbe4c4e83a86bf14c5352f63232a9da2abd983c463c0e2fdd150a4202f019741327536141b52773e86538a509f2150f5acb4a4141f8b0208383b08227ded09b4d98939f5c74307e351142ecc;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbfc507d049679ffc945eb072bfb71e811a7ad6809c14168cf5b92b397d556ef2da609b9d8ccc038fd9682fb8016683bac823223782ade365b20ea9bd5164f0a445041bd02efbbf5aadeb507c69475c12eca8e650cdf7b860f7975cc73633249ad8c4;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6f51783da90444a32488df5688517ef722085558044991e40c00ba8663aa8645973ba655a087a30b82dd7d188c7260a6ca4bf2f59e3c2f63fc24fe8c354b402cfae4949cc831858301f54de04719a592f4afa982fadda7e9d7a56522c76071bc8713;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h446937ffe6092eb1ee7bf9ee5bd43eeb120fd6d61a8c5e1d0916ed86d3c5d25b27e5aef08ad57f68764233749d82328326234af63d59037bc1db2c156f060be594c4cafac54aa66b5e0bc044bc8ffc7454ee6936580003940f97abb7014b475c5ee3;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h77bf683d592115ea53a9f8e0996a29d6a6aa09078cfad1f0b60223f83f9c88ea1807e08ff258f603fb74cace12b6be0c283f9907bc0dc564eea51c66499e65e01b292beb67618be6cf71ed65c0965d20f6fd2731758c3a6fd8597880c6fcda785d7a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3249e4f5f9e0dd393a3781cf8729fddea745e11a84f209f09250f179e3b8f1ec2598a316a218011af8b7a79093a9739fe7daf96bb93c6d06eb530a5647407f045317ca1f51c06b8d149ab6fa19b217f7b1555cd74b26201ca99061eeb76f1b2763ac;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7fc26be66689fd4c744c4e51f9c1eb8e7bd59ce26195714120d876cdb5bd2c7211acfc538f4e4deafd8322298e516ebdfb4d87c2f51e19f6c6111cb49e7310b0be938e7fb4910a70a0178ed3879148d6e527342f4731f4a32577f3c430610c384550;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5a311b3b5ad3d8bb47badfbe9807cd6de99407da41a2b7ec5a780268de16558bb0ae83dcc2a9423c894f77a11e9bf83be54bb9ab1c2b71a11d478ee66c0f7fc198ecbe3c827d57d09eb33935b36b39373823e6d769c208fe94fdc56694be0ace8509;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hcf8dfbee0993872161a74376d4b62564daac450a293e188f819137616764e05e753e94420e385c9f7ebf87e4f8fa98f6593d4cfdfb1b30e662b57fdb68e228990bed6fa159282874f7b145f22b677106e454d70ed367f2d71bec2a3fa92bf675b78f;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'heed437170a994314816804b85a6b811bb8f697dd3e0eb74987b399166dc120162d29c9f770da01d00b20732db4f7a36b9f722faaecfddb36a2488e9778625c5e7a9ce3839f714d55e280c081884f641083c4aab2dbf55572c1150ecbace0e926f5f;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h873c76e13c3339cc4b8632b92f760d555749fe06b15b924c12c71b7023f132cb56069ae8e3ad22f76633d940a9a2203c2bc66da71f43cd9c9fe7b5db11c8e9e7e7724721cc9595abbfb119810955728e6e83907f08a71626565b10277df68ee9376;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h42c3e501f31d2dfdbfabf45e79e844694bb75355ff227090a01fa5c9ede9a1aa4ffde0fb3d979f40d6085bba72d26af407d4bc17892dc6153e9b880d29f79211bc44bc84712f3bfaa0fba251b8b9d44a3994c2ace6073cf09ba3f79b7461777237ac;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd307ce235b8042d5ef819ac06c04e24af81f178aa2d70957a497e70b0f50bd731965d4ed3332bc2e652282c7d2d69a7820f4e8ac184f152ca00123814da207b703feba7d1fa9ea3d7e7020345847dff9b339bb9f1eb5d5c36add55d282c120c765ac;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h59f83d36391e0fe166e66e3a8113bd7498e6e9a779a2d78bc4e3085468b3dda195bd01900d3dd1c3132e1b08ea7288048d33c685ab4d858ab93274076cb09f73b74507b554bb8fd4d39c1382392a8528d8ce1a6a8c7b2e48f4820d939e0f01f06ec7;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h25d0829e36c1904aa1614dd6410467683898a0e1855088df28eb7565d385dc393a693400c88a8ec232a5fe94a940ece407abb41963702ccb6bcc954b019d47c3fa0e55c373cd57bf4575feff449bcfeca75b4f8ad7a54bb98b88d00b97446a252d9a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9d89d8d211731788b3c3b08fb6c7560c8e03a508099d9587a8143990be407286edbb8759c588d2e5a517d0776baf4f56c2b5da4eaa9187d7065685126e2ba137494f27a7d126dcb1562e22975868021733c18ed5504528c4678d1ba252c64fb09c50;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd427b519353586f8cbff69e2ee41fcc116b0d85879dc2becd4e1101e52fd61f8f0f43d97705bfe8960860d835fb3e6901ee9f789dcb27697e3aa4c59e2b3c1affa564012b38d91a4e3983e860a1a9d51900df982bdd72b840851210e9cdcbaa4afab;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he040be6219c233cb74d6627ad3b5308957d3870fe05c490145ae018a247a3deb3f5104a401187914888801480b2589e4ed1d6c4b17a0d5cc1e81c9098cca55fcc0bbc13c63acf783d3990c323e92a7c57c940f65cd0ab9d8cc4d1e29cda07d7b4612;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdcd28137193f322ba0055381447756450a82b770a2a333f99527b32eb5b1d8cd01f52df755ef0670429e1d1668d9726e4cfdaadb568fd6d42b44411d29a042b75f640cefd08f6d576c2bced1bd6d0d73cdecc4b82a1ce1595878ac7a733cf62e84cb;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h268e1d5a2866a6a37e3b0ccf7bd53f89798f2dbebe68759776d7f6ac4954b911c12e61a666b80a09001d80db5effe16f99792827c2de9ad0b1708d953dc830607f3564208ff8752254aadc4a28361d3d4be6633b56222b9d88f5768cb8b0be839037;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'haac44845d002eecc20247cebb7ef8f6c586204a181837050852babbc276c30b0867d417d9c3c91c644dcde1a25410e2e22c410f72ed49fa38486959467a9eebcecf7acac54a4152ee3fa80a682e6d252400416a9c660704e3038b4e7bff93c6f1264;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9b0bc558c0c8c25633c1fd758e4261a7f35a96359d428c299e07002eaa9f44e0ccc603144548a4604fc059962822c70190177551b2cb448c1665c4c1fb3538d74db34e07b1b9b6114083336ec315d80d445a863936ce16f739169e09eef1fc8ab6e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he85cb07a864550ec63bdad618ab76536f7f65c38303ba5640c293bd35c10c3033357310df1b69ae52f8f9dd6ab880e740d8bf5f87fc71b2b2c0a74047caf22c6aeddbf6c58a443aa116627ed1aa4298cbea0306c23cda30e1e9c8ba3f85b8dee77ed;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbef7ad3c6d579416aedc8c6e6cbc27ad401feda1d2d0b77000e2b98da197a7f366eaa0059f525db2726486f19b87fb63ba7a8b176630669ba4db5e79751806dec53409f5e9c1e99f6f8b9dbc96a8a85fe87189bfe9191114a610a2ee0abf602f2b37;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb77fc27dfa05d4d39184342bebfa580eaa0a6e5a47c6ad761c5c9e0574f3331565a10a401d20f8f538d5e2c4bc3fc789a41a76869e7484f4dd880d88a8a079025f543a85cb162ce6dc0f9b6e8ec9158ff64ee137536df02f8639baa9225b5a726e04;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hccc6190a05088c2ca0856f8017d7807db2e89d619a4517fa6b68a239ea4a9cf9e1607cf16ae980da5bd0c4a281f89b6971cf626bc65849cb73b5b319c2ecd2d84d98cc6b9dc46a48073564a093ad1032fdc59e061d7dddc1d5e7ee4c76304b7876dd;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc0ee6cef39a7a92b241053782ccc6bb5b8a0a9839091efe370f8f0148c0b79e7b70f7a393d9fea1783512c4ff556bfd0927443bb4a8d620929d948beb6775d975b2511ee5627003932ba63ea36cd50d76321a2c2a86d4565bf180dd8a2ed095b18b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1637214e7d43fe6a817a78c5b0f817d1e73fa31aad9435ebb3dea476e8f65bb40e7d1af25df493ce1065d5f4fb157ae7f579cb57eed157d03b2a103d8ccf9b82653f09a9e7cd9a56495c0eef3ac69302fee41fb098cc68b4c67bef3d45753ae6c636;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8a7995091a5bedb93bea1a38803a7b089cd1754d963dfcf872abed1a81f94f831236af85b96302ac2586cb5f4813e27f9e0c48e414c953c36b56f1c98655dae15dbe67f04eaa4278f851aed931a71b48779c044f76ade099934cdb99e4d1b0e38681;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb9f710b17c1fede075945a70552143020d545c69d670974798904d8c70288c333a4043cc9c760a65f1d6d4bfa61c28328a047484e5e77e4131dc2d4134cfc0cd9fbf3938431a64dbbea542c96079d97c22d052a3720b44b0acbaa232689cc11f9603;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9b5086b0cdce587c4b10a6f05d54fe00207d7b8e01c619143db50c3444817c63d36dfd2d850a70f533f31287505e83d2adfa4963845ba719d669ba0f99ba1cff0b32e292d50e2ead5cbf6a90946237ef6649b5269562d11b40e0372930fc2c0294bd;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4912f3917f915c4a777f474c0594df291b207d12e4e302114fb42a8b1d572be838ae37645f30f36716f6d1df9fe04110326cd7e2667f9a61fc74eb6881b39e3e4f9a8cd72efb991cad6a7201d54c4156eb05debefc86f56124ccde97d0fe531d3743;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h26a5a418da94fef1b1f190ffab5aae07c5b06ac012b2bcab9cf47b1c38dce4dda1f8af8ef38cb149f6e3ae036e4594bceb447608f6655aa5d295cce1c3f6ee528327d21ce4f902fb0877c99a939626267b079ef9a4d7d62bae865b5db606c9a8f4a9;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3f13c2f81271fe3c64a57bbbdd01204d3f00d0f2fa9bd411097eb59843906a93ba4d642ca3f8a5de100bfedb53e15ff75e2c2ba24da7e333ffc1afb63cbdf7c6d5413129f6e41db9e18dd1c89a1cadb8a99e2fb105710c330fd27ad88181af888c0f;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4b37275c29645b62a97c56035b27a9f92fe0d2e04f2db50b5d08ba9574b2766ccca0567cfc13f519eabd4abf3fe7bb0ebd3a4625b30dc5b0ee44ac29f168aa404a68d2a5eb97522a5a6885f5fd8de19aec14cb03a0500166b4a8833572894cc7381d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6d9977561dd327797ee4787f6ab9becfcae15c766ad713c22a252cd45f76b690e303a52ec96c8e6f3bf566158e266dfb1f4435332f6803e88338b4292a2b79c0d2d9964aac406aaeb238c0934556cd3423b381b3f84ba361530762aa1931a4c31605;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h50471bd6c62c98c97b970f4e4cd0130e11b061ed53f0ee32a70cc9f2cb06ee468a4f149f3ec2d67cd3bc15ec200fe75c2a206804fa564f4b794c5b80e37b833b0e8358fd53edbc034b2f214d85059d9a8a7df33c27fbd29b5d83cf7eaed32b7d1d1b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfe9f8252997bc1e1e60d6a184e6d501cb8021fe4a3745e847da3e2232c3554c59f9f75a03d35be2cf11dd526ad00a2cbd51f6448035a4b9105f2eb41a5f9ce7b8f5a299323d1366b3cd9c6382d2f32c9d3b35e3bcbc233757a2d9afcb6ade3de1214;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc17207662eb2f357392339c61d1741f6a8c7af86709efec04b806ac89a670435e35c300b4e655102b938c660d8e054cb6acfba06942022f8a59839fe8b814cccaab90bad2cc8d7ebffd1e5cdab2b05e0fefcf0a6c4092eb3337e4fd0f3dd71b142c4;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h306d7dff4319a344855d6436570a6c27f05db1bd0a86118f95572f004575d7a6aa2c5b2284cf74199496c3e87c9a9f38939f310eca987d77d13e652f590987b38fd65f0b9c411f78859bfe21fad2b56568c1e96b0cdd823ab1e9cce6dd4341a559ff;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h413a0548e4d5841d52c6bb3302235d1acc9d9e435808857cee0a2d3685ed62eac756c39fa26fd46512c585e139bfcaf92046bc7b911ed67137ff8422a272c225ac707bf241528e0b466bd9ced9f2352e31877b668e09f4dffbeff92f8c736d761a2c;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hac23de4e6153781410c1c227b68cdc86f2a7b8f59fbbc44cc4930289506d19b209ff03ed231212e6e273936c606bea32b3f28741c73121c27ef75af1ed276d3a4d7ef65ffaaa9ef4690fc1ab32e92b7c83bd8c6c698734a082d956521b37ca9d4c4f;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2b13e00cf0c07f6a1052b04aa704c598320df8e863140af693a2cf259ca13a11d91b6acdeb925a62e0d7b540666351e26775c06a78a4d30e056c8be75eee42def69b88032ec8f58a25c6b26bace6a0bb8f31a9a28a04ccfe740892d1810e3461b150;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd97398eacdc3493adf37e0df0d7fc602637a19c1440d310d2c55eaa1759d542efeee00e8149653387540151c21a24273a03d897b54edc1e042c134f6d05a1736f9416a5f81b880a029fd40ef1ae06eff8e8fbe4e1a43441005533fee316073704e60;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h45f96d97fde647e078d1d13d3ef5f7144e36fdfc808494340cc45ba1faa2cf230407d79212c96c62771e79be77bb7094f4ec94366cec16983f8d348729073a4e90f4bb3463089292e4f826ceed8494b36062128889dc3848a4db1f2b166619dffda9;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7c0f117ff3d6febbdb258d4d24555a8c9ebf292004798af180a6022231425d5b9c51b0df206e3d8a2593a127ceb222e3acf175926fe733f6dc16f646fe362badc0870f8c449dfa742ef6878675ccb6b5e2e1ad62e81786cb2c233f09c2555c7a858;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4d2f9bcf7c609cc89123607f7c77f69f787bd68ddd5bf2c8cc68bc47626b0037b1338ecf6df8ccfb72745b8664f006a236919ecc8a8a3c7fa98724d84925205b112b3bfc53d4f68e39d01ebb99e5fa2c5acb2ed54ba138cad8eb8d0638024c08d36e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h120373e36dc0924237a8dca7dae194748ed22a06b6491680a011cb37d4b5cc88461a84c9c670272f9750bd23563c41817c59f1e6dca8e3662f00cb1ae2835fa6ba832f216b92647f0d9999375ea870f7199bce73b2639b2544dbd756027becf945d8;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdc66e7875e126560734dc3f8fc27e04f8c1f96f896a803ec3eeffdc449edbcd5d188df647a12d00f044b682c1f077e54a10597f552884756482e87f163ccc8c73a371b512d90b8f0d48844a0307bc84d1c65b0dee584f886e8d959ca6a8ab0a15997;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h46cbe4383e0554f19c306b176ea00827a254a0e6769dd12324365f023a67e50dd45565810be937a369f92a3d01ae8386c44cd47c9065ed6c2b153c094e6ff1a6bf4ff8a6cb0254ea0d3160e8cbf0110d00717daf158169a12e91714e523144f8bd3d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd38e4777e04033eeeddaa864709b35b6417c3ed2b332b24cb5cf8dd1cab3b72974f2fd2a296ef0e093be7a26c255ab69dbed46815c46b3e634ef2cbeb475d117993232ca696af0743ece7df60d9c7d9097c28523216663dd4977f9bb17178af48d03;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h84d5fb9da7286648ae9f5fc266cac5cbe116fc4086b69e3afb391778d9df5bfd94c0dd49873ebadc5d10b6f2d53b2ccfb1d451813e483491069f54ffd3c62e58e47e5ea00a7061dd9155367b3d59c8fec8b282da8edaf8702496cd9cd5598092267;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfba94fcd67aa6187540f9f813baed316eef022047afbb85cc13814e82ace127b7a4769b31c32c3dbee7e6e4f7953adc78d6bbc5a998694c5da70a5d96adcde930f15d6d3a1e79c6e3ec3b95f54ceb6074db153f00dd94a470ebe708f939c003fc04f;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5652406322c7e01c60ff8500fd2b1a7f20f7084533aab34164830d11849f9c7da692f0d0c38f01a133a31b22ae394fac8ec076137ccf4d4adb6a4a71aafda80e0cf26758ebf0b9c22e2656f2698ea082bece9dec9697cf2027cc5b3631c6d2d0668b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h87cb9ccff6b5d36198fd224d5a1ee77b33a24fc3ebd3272d89a1e22373ae4c0dd9071c5b12ac6b7eba946e5fd8c67da3435f56c473823e0028095973af4b656544cd5df37cf4ed66528dfc930ef9b5a19fc96f14734a9142ec89ac0f0923eaeb77b7;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h27a464768dbb28118a0c35419ab84227b33fba8e81f8e2292a63e4b685683ef529be1bef974e4f935a5c0ca294b07360708af9114429eb702a5c44c0d459dcabae4fa0c1f2a33631d78800cfc283087d24dc8ddaeef0e8b6e1145411b594bed0b51e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha4fbdf6928974c6a95beeb0788b30e7b04d8fcbd96e400bc483017f3f9ed5e23c5fdf14849270e917a05df56a5a7ed914138303650722595c75d29a7ef22d57bbcdba0ccc1bd0fce6704709608a782f12c4610d6da219b3641ae7abf3d0fc6cd8e75;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h46781a3e47e795e8d74c9ce77cffe66fcc48ea980abfc4018f6dec5ea13716184e85ea10929e1ddc5896bf17ba0368a76166ba7e660709bd3f873005fa82593defc2b55895f5b21f13f16fbb73d54baf8a279d1639573c739c8dfcb590dccb7315e2;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3870d9b76affe0879c7a4e906a5d1d49d0a48ec353ff0f1f7e1074e31b276b812a447cfa642003300c3c30017e969c73f0322d4ba6ad6bf972b1201cd3429c080d48e2a187d7adb721d5603dc3a35af02ae7fb411dab5772b9ddbacd1ca7b9535ea7;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8cf16a9da4b24d1f02e1da2e85ae404054445892c29305f87d088e40596ae8060401f8c87d881e29c13e10a909b3e1fd52439d592405363758d97f099a9021afdc0d720d9c7e120fda7d03585c29a32873481f4f1c4d1a15019b74e20b4155662a3f;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he7d30c330742a42b4884113637fffc1b338f0e462b06202a7e71a62f0168ddd12fa927d265cd55f932218f4e3ed8d885042caaa4bc19ba27719750c4ce3c2c3a9da18aa6ac4fa53d9711dbe69f50a95273cf98b237e9e8ae9ea6778ec5d50e09678d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h99175b5eba21497374d66333f80209253619b620905a8e4f3ade69d7d1fe25e5ad2345781d279c38a7164fcfc9f9f793fafccfaefd371c2b977d41e24f20cdd5b2c48e4fc5f2cb36ea38786ed635765fc09b76aeb92b45cc28e15f3800682148e552;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'haccacf94ac39ec8114c4221ac1dc1fa16ee8fd0d3de0e6b8e962cfc8364b824e9e9544187faf4f69121ebe0d9dfd6d50fbf5c449319625e0d581b0660edcc48c3652201f47574b08260ecfbb1497a9085525e77bf9af75be665240cbf2ad1438c7e5;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h305fefb46664688853292bf74aad14756bb65ee8e7d1d58c2ff6cdf7f5ce77f8230f3cf5b715899025bc52b0800e5193a8706450987755e3168c468540342c09bcd754c862ff2526fba934735a35616f7c363e4a13dde39a313a916373bd7d03d6b7;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf0c8fc942fcb0705e4147df321607d5b0fa39be05173fc3d451f96e6448d319ed3135979bdfd2a3bc20e7f2fdd14aa14dca61570788966fa9a58022c1a72b969b77b4e2802538d7008af22fce591c484c07af4bd6d468e8543754839cabb644ae188;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h564e5aa5d06d0356b3213c01beba430842f385f02b031e907e18e7a79739e77098bda86342e6ce2b8fef1994f466d0195570b489ef1a1ed144a69b3e3978268dc1c9d16eea3142eab0e6d2c25fd2e102d8e52490ed52bca89e1eeaff2cd1d131ea24;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h492cb443a795db8cd11646ecb7c027ca169e114d9fb7ef84ef5c7309fc1a785a0a282a625f727ae8b4463ba4156cb42043ab06f775227dadd28d8986f703e513a3d5d7b5ee4138d52848454c077b0de3e589d1223e564f7199fc7df26dca86808d77;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb6091db84ddc4381a18fdf55042aa6dda6acebf3703995b2aedb2ec1e17b68fe441e967a628a45e53910ceb653bb0cd30539c04b8b2ab38c0551c29ce2bb9d7e7446d249a9c467bf408b477ba8f4d1af8b2ecf1bee357286bcde7ade74e6719d424c;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7f86f87eb464cb3742f7b35f949587ae10af7833e11712748106d5fc8a0f3f3acb116bb742b7119dffd833385b9e1d18a4b4c25a2d3ef1ae72fcfaec48456876c7420253b2387f713d459f4326f463736f7dc56cf2bf617be2ee60dbf119bf979ff1;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hcc1447b7682beeb8e8a5efb9a371de1ebf62623b97f613f4b999fa66df422590518039b87326cc284de3c4de75de825b620ef8ff6d68d9ec5cc0a56f99dc6d06905ad19e547a1c1caf92c5a755494ae4a50ba7e85d34cbb356754bc044cfeaf5820a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6f9ddb10038eaaf72a3ff2d060901e9917e4e0819cadb2f5f4a3aef2d173fb22f78747e7dc27e13fcf5f49d928597617bfba88fcb836a521cd0e8dfc2159f41b28a0f850841689b256b5e50fa92420089224991d017a93dbb3d894fbfd4bef78f86f;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd31427615d9c683fbd4fb0775ed62286d0cf2da0ac92990cfc42ecacbad0ec186115f919895528572e22f1707ba0ea050e2305fb70e361151c48236003b7b10e6aeb45908187de18bfec757eadb87fffb9b987e4af4a2d752853ccb6d431bcbe6700;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h75f8e1df077b4c6f44ba6a1c9e0bb9dfdc63f76a40b343a33c1dbf8cb383b476cbf9dfc711b01d568ac42e0772ceb43cc4dac4a6787baabccc9edac3399331c39447a52f850de770f6ba7235841afe45a84b87d6c38001bbb9bccad745f2a9be2d6e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h801b28c8e4fc2856ab7eea345b23406df0bc4b38178da8f0dc6180fe124e7d4b96151075cb2c7036b8e749ff2bbd0a2bd47fcf63f17f1efa2531e54517945e53ce4312ac84aac2c525f3b621faa80bb15a33a42168017676fc0bad1d3d98f4253027;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2c5cfd8f4a122da1a2834648b60ccd20ad415a2121efbcfc8c480e797dabfff488765f27adc38209083ae6b183b47e92e987ec0306836581348826a737d341610c3589438ff666e2616333fa824bb61f26129efc3ad52443e1fd90a76322a0f49168;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf7634bb290ac6ade5c68b3d41d3f6ea53508f4a1c85da406ffcd17fe52decc0b654401e7e195f85a6f6afac282d2d2dc1a0087727cdee57b15c9bfce1d80e06bb03d8dc03cfcf395d2866567a6e79e28e760360c362bf0692b2b219b8e3d4e7134e7;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h755ae6a79e83ef270cde3fba37f46ad175031f307bd4d5c9b2797c5e113518a4359246829ebd4219b539907e4ee167d981c27a6b5fdeffd4ff2d9c9b5b037a0c843cdebb3109b67c325a7ba1eec28b819d9117cc90b0f1a5b49a8f67b94f43cf700;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h48c5564ad1603657b3ec7459849dc6a5be635fb403978f6a081f0c9b54bcd6ce99aed0e1ec723617ef688fc896860d50cd6f99814e68dfe2270bb6cd2dda0d6150527e3e1590a5b5baac6fb1243fa2c4b7e3fae518e7f389e6ba8f1eb24c60ef5227;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf404fcb8ae06ae88818683e0eaa517697100fb32b8a8c70bd6ed8ddc8280c2df15df0e44779bcf811b8bff4ceff3736889f6fbf0fc3b960cd058127d4a328efc248172619635f5906045e1ae5c12abaea32c84fd3be93b31e53a341f929ed2c3bfc0;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2d0b12f2c1472a576d478d6068f2347bd772a9642ff5abd565416836e4521866b781787442d18a24a6c58c4c3ccfe45dcf9a04d962dbdc5b402f3ae7d83800933801ee53fd60f2d73b323ad35a54f5dd0930c40068a1f6bee6adabdbecf09966d4ef;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4e6daf81e00cf687aa21c4fc3cb6b98f63e6dd1dac16f7a9aba834c13eab46c3b52718e627f42356a075fca2e8f62c0cd70939c4f4b4d74684e5295606b1ee0c3164d4f76ee381d281500cfa38b52a611c5aaa795720833bdfe83d1432a22f98b5f6;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9d4fe197d95d676aa9f93673a931eb04e916428b38127b9b8878264647ccf9a9d9f52a1ae2eb94dd8ef7b55634b335d91f837915a960f6db2e2ac6cd91e9a4ebe0f69c9b77bbee1c507b83606a8c724450b1564d7f4207589314ef4fd4c074f519a2;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h399362a2015e12c443548d1528abfe5072b56d3ad6aa72aafe84c286e9fd9b8096a1e402a3ea613136dae12318b87032320d8d4530d4c141495bdf71954399dc4f72cd2882a843d6e39ca732d02c92b4f9c9108947dd3e5f3955bdf8ae6732cff41d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3b0057e2d7716db69d931c2d51398f02698eebc515ac4bd83e1a3dc260489e8788b30dda25ccf7eff4836f9d5acf89ff6136e91ed9defa8db108c34db766f25aa42fe9130d05bb1c194820a4b590efa5408c045786e265b690246de49033431dbed0;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h58bea2ef92d84155893a6b30d151492216c2340cbca8c7616ea36551c2a7cf59cbe595f5d9e2aa19b030189b636c640f8e48810e13cb5a29a4aee38ab075d21f7883e3452b0ea3e53e0cdccd5b1a93d51e14fa6d31a56f429be0f84374a8ed852d98;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfed6ef51cb2307c1ab1de0562b779dbaf3999f064892764d849183a229bfebd84a130e50a01db9884a117736ad28a96451da3fb16014dd4aaab4ab3a3e4cb73354b48316e33d673df0393a6a5f8fa29420546e3a865525b94ead55686eca6459d470;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h81938e70673f5d63e380e0a8960451322c2ff9c34a17c93fbfbfdc2eb5d8156c678ade783d234b3d60a552ea18b0298f1b9042fb87d4e4d6b0615ba6e398b9479cf010a4e3e9405b2f7eba7307f4b0a6762f179b8ee126d34ce87e17835ebc822079;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h60b2a81c170aad5dff56e5843b6d93dbebadc1ba8107780bd18a3b08a713a27f42aa39eb1a9ae66e93bfb90a3f99bf32428d35d8986ca9c244be081f590c9246c959f85065416837d65a951b80149129e3e5c1e342ecbf1a1f18131bafb429864395;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha91a4135105a6b5cf02d0ea51250900558f9492a171d5a4d203890b2d5de0846f4e8dedb0e432739de56e4b7a28134f547647724462f3ef2f7fab378f5140c6115ab52ba41eb4f96a7b245c5cbaf29d5df45783bd9ab04e469b7dd15d283625e39de;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h25505486aa6a7595bcd0cef547c909bf58ca55e3d3f4b1e8bcd5b3cfe8140d3de5339257860dd1e709d1bc9f44ba3c283c3a1d9c54b80296e45641ec1e5e84e946961e77ae0819936e98dbc84cc819fbda73440ff495f8c9f1ef0e282393532c3ffc;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hefc4f5502fa1db206e3086bc5fd29cdde83d865026c94d60f613bb385ac7d5f2732b83e222007323e522db6c5cb411aa2b362fcecaf7155b877409785b1e4446b5152a9f92e774f45ec2de130bfc4e1e553f0e1fefdb7fde3c5c257384e829c22885;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6586eb8f2451723d2a2a846a1751d7c3a65995946ed78a3eb52126b0b3a596809cb2751187ba91f2334c946dcc06bcc23880e54d28667589d1266951c1c77a5eb7753daa53d338d2e20b0fa58581f61beb1d6a82b9074808bf4d8b87c51750216411;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf25607f18db11ff5d4f91bc34a1d7521a05f53921aeeb79082803877443c827d63037c37fea8ce5084d26bc77380b5724dab1e27c2986ef2c2142757ed23ed2ee22cc335bfc2789d7e121d3ff7bcf96302604862b8fb19e7d5dc806734eea3107f81;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9d15cc257036bfafc55234e194992801422251eea30d0cadc7199a63a685548d191a2d2498a1a7c6616aa569e653df54668ada7b2472318aa11dd84b0f7561076cc5614a28b7bc2733c3d138fecdc43395597382a423791684ed239569cb28ed546c;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3feaf581fc7090ba03f4e0522e1b0e122e4cf75a91fa65efbe1f8b492f7dcee73940902dd4fd474c1818ee3b7c92f26ade5307cdc9336be7df56bc47347692c3b899567a4f3c8a368b3d9f85a69824a55bb2eb70c5ea0b105a7ca753fa4e3d162fa8;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7a17c36476b30b074317b6d250ff53552530c53a70944ed1d65b0f24bf7a244902bd4840ed6571ed917eb3e4395a698911380f8bec11fc9f86dc2fe683e9bd918b918a5d3451282f6d2f28a00e03f123c364c3b383fd50de773e9d390488ef47fc36;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h882f6d969c0350ffed0954ebb9ec016a4bcbf898b17e2af74f48e990b61cfa5d9566f0ad2c99c5ffd74b10aacac95cd6e8d88bf34c1d72f027439edc54da77a4d205b4dcdeb787056cf12d7520016038c0b1982307696bcbb3f1f8db7b91faa59773;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h20cbf23282aa933c7de882ce256fe52203cd6340a2236dd7bb164bbaed25446ce542d68bc917b19c2f4282431647bc8465b794b2318b5261bfe4eefdc939bcb4189a266e6781a51647b39c7f12d259d8b11192e0e2cacd6733d139cdb54f6fc7b2f3;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd93cbac240adb37feb729110277f58347989052926ce7548f0851146a01ebc8e9d87931e905280663706d76218e965cb0cb15f9dc6148b7087bcb9512b3d4ab4543bed04aa11bd90cb2ddf0cb1a9dcf1f7933656ab6e6f3c816a6852171d9c989f8f;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h683ee7b033d1a1e38f11451fc92e024105888428d56669bf462dbc120671a600e81d09eafc01477217fc2e0d7c1c03a69fddaaaae62ac54cd91360d4e784c1f26246db7563f0f8fa5ccda9be6dca54d218500b4b9b981c49721dc66f5dbe2f46741;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h60d6ed664ac3a5d8042ca688c547f0edf64c3543fc133a6379583a2c6b08b601bbce32ecd330262e8184b3af73c0cbb50d81e7e168236e4578d8ecee1cf78183912ec37edc9c5b911c5c8de52b0fdc39c472d961f041f8d9258455712f6b18392ac;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc8d01322d0457ae27033e1c8c7a83288d5e314ee5dff717935d38672930c5826b6e140a80ff9b0fe61a70539ae15bcff4e45dd1ce0fc9c47acd8a7258e3a1b872672721cfef75efb9dd13360a312b7623e79fde9777bf7ece7f002d3c420c24b6e94;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h89cdb85e0c62e25f48c5559bb1cdc13026e654dcdaed58c31f6a230e9e7812c85bf7dc8fbf61ee9cffe1b4032282b2070ee65d5d930657031a8712c52e335ebeb414085ca974dd99ef0369974181b1c21a608d08719a0eccd5cba668dbd35763fb62;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb6ae4d9d2530be6e89a9f75fe089c777ea44be3bd787306e3d763d9fa2a989d02b60ed4d599a8796f44ecb374f086b4b5087e8eff142bc25990a694a87974744db0d1f9ea7de0d99da2339d185fddf460ed30374876ed9cfb3f0a2b5538f996d83ea;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hcced3ffb3e5790001986ea9f590e456b1e2c3b6ae51b432f53ac0a5fc1570abdedf71726064d717add5e89276d961187ae901881e761e682a66fda1e3b571675a153ef7c340a301a2cf14f94025d2c5e576d3403770700edd883560bfff8faa12823;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2b9c6ec6eadda6c0a3a3e20015bba1fa6ec994f87c50988fa40cb0ba0b1a041e327c6b1ca72c39a899520ffcab701d328212253cd68288cbfdd4aa1fafc23cddfe018eb88cd2b1bf9a2be977887b4651cc3c8a1cc59dd3bc183f38085e150943533a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha1fddc33f0c26dcf851ccfe33141d2ac932e8cd3cb88b00d5f9d0a67bfb3fc3e63dcf6171e1dfcfe87161cf7cb5890b5a179a545aa4409704ea0d1d9cf95605120ae494b9cfa74e01df6b902a4a4fa2164ece12ba1b9498c8d94444a04bdafbbf71d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5ba7c1a7129f964aeb3028ba6c3fdd2ebc057beddd7f13ac40eb47d134b71ad96f83b578440fdc78f150c30ecfe481752abfd9e37cd6cae12ea2c605cc9aad1a446f2db6256239606bc8e537ad7f643eb09cc4d9571c3f2cee74dbbc9077a71ac323;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8b2e3c1708311ba852bd81a1014e48321b742032059be0dc7389ad69223c8c3a893613488c804048fe62e4cd6ad1e759441a94c898e8f8a399f752d8c1a5ec87b6306cc200dcfb07c7eb4157f86ee742153acbff3f2a29d687100e4518894ab3c2f0;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6b83a19edfcfb4b6c296e648c86047afe3975f62e2babfb6a13d39d3cb15e32bd3398b56e27fceaf10e28b34b21cf55789c96506be69cd85b1193937aea86b057a0926f358f2bc876dad536d771c8de6c410f7b61739f07d9e420f4979fcf91d6918;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h39d808d9ae506ee8965d1a95dc11e752fea8d9686680d7bbcfde99fada2c98bb59e770644efabd28e478bd71d6c28f8b419f5544cbf6e0f8c9c35000b8efe8a804d0c3485a37636e936854fdc1a841d0365f6c0155f815de7e6e9de57f32d9f8a793;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he1d108e4c45c081c62d65079e519365aab79b06e58ae61e5edba198f6bfd1a54ee98d15364b56713179bff2e95bfa8863992f828c39d4453bf6c54933eed7fd89da592c2423eaaa59dc5cc245bfde907c149f07473388479078d30b6e11bf1cc5c44;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd087f140eeab2e5aee68ff6f79f89dc28ac69377e8ef27a6008b6cafc183521bc45b6680effe402bfd36e8ea3b28ee286fd9dc3f04ead14f6a3dfacdf3a842f0d0d88bd7404f3a51fc508a1e9a7a5c4c26146dd5866bdea4399c698b70ad2009390b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9e6d00689ec38f953d0e37661c758bee8aea1d192ed01441480ccbdbf116676618dcf0bbed9c60da63200c771ae6cd0b978804e74797be30d4043c2e0c0a73601b828d996a3ded667ce0e624f693bbcc4a3dc596bb66bf6feb708fee0373cc429f17;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9346447a35450d1d076041ca1b420b5906c8f8a8f3f07b9f25bb9ed266e82e53d96afe02e9ec668923ac2d46069ebce1fcda2b0d5116a66281780d1c69ea03bd7745b7347886e98fafaa9aaa2e7b46f08725914d155e7fa2ed49cff038ae236035fe;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h40e80ff3ccbcfaa305cafec92c3d73606a4bc271e67b96aeca92a90c15ae3e9976b05f098eaa8e1dcdbc46070cdee1838ee28281df059760356e05edd89d4868371f2690654268d6ac183e9b0d3ed63e38101ad643711c1ddd0ca81aad5301eef424;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6066f55205950a144c9128c14bca25afc027e90e7b25a6316bb86510fab265e9a671d8699cd117fce46303c6e1fa9bbe71c40f0b4626f0c5c10057e79619ca90d0c709c642c5b7ea1ba17fb01f7f929af258ab5c1e43eb67420e823e3d198a420855;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3b127a8601993f8d5a7e3f2b0290a2b9b73c95838354ae015e201522059fcae45d8a4f19c03f9e3a00341afb92ff4fa448ba95669b074082988f103cad6814639890bba5e43ef56c8b594790e5c6f2b0d0c3b25bed4ee28846c90612b83eb5041c39;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbd141ce747d8d7628c54b712cc64b7fb6f42a9d7b1bc252c2d2997b535a5f426d72aac0d6151a61971cf353757700a5dd9d422e7855527f803ee04a6a20aafd5485fa5254110136b8f5e5b86dfd4ca4515429390fb449992d103fc011f08f1a500c5;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h644c4fdead933dc7eb7771ee8dfe59d56d096295ead35544a52a856adc13c636e610882131da3da765868290993fef5009108c21e75aa16a493b6f4e5e8d086ea3d32e0b1959d1d3e92d8f2353ca8830625949116bf9ae07a63f93caefd1b1c25f63;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2bda219d90bd1a34119bdce56f6c72f9ddfcc5526206ed03a0d5513348d5c241dca6f9844f8e1d55bff4e7585ae26f623ac178489203790c7e57cbc53746596685fec8c26d12356be82fc50bbf5b1695098e73968239ea20e83c1d067843721bf1ae;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h76adc6f65937b312ac8626bf317bc249e83ed35e15209a0258e5d2961eac0932c1d050761777074a5a6a8e26f3cc6b1f40184c8386937acf94688d433a7ac2dc8c6125dc93a9b89da70d70541e4649f33c63b349f7ddbe04c004aba71e51b68aa9e0;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf756773b55c74affc3dc525941c54c2afdca3d24c6128626465fb56cf14bdb8ff3bc9ac8a1bc3c795808f225e1ccc0e251104da86138d6cd4cb6b388bb9fd8ff3b941486c25ddeb0b2b773dd62e863748ee6afd30668fa69f98a10d180112a41ff13;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6060cdbaa9cd44cdbe7b8f61d6bed442a22fd1e47c7be0fcafc9f02e9928e91522c4df2611995ed11f181e5de20eb041dba9f70b2a14a77493d173fa950c915a58c11f579e6b520b8acce3855a39a51ab2618059742b661c0c5f9681320e642f6efa;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3e7f31d91bb3451b13b0302b0cee2af947c7f64e85221fbe00d0497e6998aa319983f47dedc11b269fc6037db68a95e228a178f17b5b2df58970b301472477bb2eaace5dedcb19c084edc14c2afdba62bd75213fbd96c61831579f4a7a2fa7dd73fd;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h81f2b4e4f5d2d6f661fd05da8f63734896b5a7e8a5c26c20e718a5c4f95d5a1a998ec533289b91a35b2e39d500eaa71b6d8d3a57d5833b1c67cf23b053f0a95172701df1490b6bf02790301b22ef959e5fb9aba636ecdabe597745b658af2d186c2;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7fbd3546c5d3b6dbd42aa0bf2f35674a192d05f562ec634c89898464301e679d5fb8d04544b3a3f3a6dc2a3bed0bbf57ecc07203528da4e4049ea4fa9e0316a935b94576fa51dcda1f356c044f22f24349b105cbf0ab6e69059d002b13f0f64e77e8;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h200837ed6ac9370e4dd4f756530590af16aa6c46c0651bf49b0d77a54fef204f6bcfa74cda7dcc482bf3137da4d86ef959d947e10a2cf261ff6e448a7dbbd5c5d0be7ee70b38a9ed65556e5c69dd95e3380abaf87ddf8c6a3c88b949b26eedc6f0e0;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5e722d3c238127cc37bdd36f4a20202a7fa415fec42104d42eaadd3e97bb8c886fe82f1f457d5a665bf336913e0bcead9173b95c42454879313d4242b4379375841d31ff325a3d59eaaf7bf03c9312bbb1e8e0bfcc0fca26514cb96be1a9dcab0a9b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h94456d6dbf6cf019212025572ca61d267a80fe68126fe51423a054826c5555e4133f3e46e88dbaa749d74c3011aef0f272a1e9414059cde002cb678f267ba97f691cbb876eef2749b9abdf2d49ed79dcdf56233ada8cf72d7af0eed7faec29adc5c2;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h434b421097d45061bc3166168a822c5bb629d9926b64646c7205dbb8f2bf6fbbac4d239e6b357bfa4ae3a7cca1d81c25a739da93b449b372bb6746c233baacf78aa32df9fab6ecafead06c4e77f5a5ee0acdbd18e85ae7e71debb5ef788bef3b9dc0;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he3ea4243e7d15d178064d011594216f110c62895dc653c1db93cbeb57995fad09e5c9c8f073c22916a0e87052894e12ee9b571c93f9303bc11caf3a09ad673b5ca4b95963a0a8abb26f42e8536f59a00e03442abe4d1c6ba36ad6561a66b381c49d9;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h648cf2eaf26542afe61d12e55d6d15480355fbd88a0ceaf02f3ea70112e15a0c73155c2a11e627df4bd29df3ad873b84de6ed502e2063be11320809a3a62ac012d43782b96c60f85c6b3ca82957b62548dc10b686f3beaf90f61eac7068660fcdd40;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc89610925e77b145d6182aa1044058f96feb4bface60efcdf1f26f2cf6cd742d999aabe155595bae882fc6cc1b5e2be2bb3bedee0c18417a6865c109b1f15e203e833f38b7f55fc9bb86045770a03ad8613ad94f2c730e975bbe8637c0f7adc06f52;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h95cce97f6d145fd48b365d028a067671a6a6944cabdeafb2a88e817b374bb0965039cbfd4955297f66b6851212b015debf7f0713a019e054f5b8e68bdb8a5dd010aacfb9e3c2734c2145f211f24832b25c9be4001dbdc94439e30ff6a07d57927639;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h59964d83af57f347f4ef73d77fb79cfb55992267ec10109c68233e7e641364a899282c24f6a788c05471531e96cf70ee479f204cd3a383de9f0e58dd1511ecc257453b9f4561c513770ee3b724d89c9958c5a63a89aaf33ceae298ccf82ce0611ae8;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb1fcc30a065e92aec8e48311a44d06c4345afa5984991e346d61c9333de94c878d35861c5933a0982ac91fd5d87dc7201a3843380406a58abf4cf190cc0853676a6f4de7360c03aacc91d3750f0488583d57dbd333e05db4bab822c129bd62a1d1ad;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd98d8fbe132c6e5d8ca5dbc428e47efe1b799c2546662d425113a75576fe305c56852a62d67489e9c13bab0c8c363390b9562f2e8a2640737517705ee7197bdd7f671aad2557a1e043c4f2eb6c11563515d14687e20422ec4f35256aaf80e73fc839;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h500b5a8690fd9ee4c5f086c52bb3f8761a9182f1dd4137cff7fa0a310f5f407e18115d908983f2542b4b2cef8bad270d8b3ba5f1a673554336f6bcbefe1dc6cc7f9b9d193bacd8e27663138b3641b1a70747c847410c0592ad1168f5cd56565f56f4;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc2d39e50e3240037bd9720045fe0153ec5486fcef57d5c98d76c23bf438a4149d7f8ad1f0a304d081dfea4d610f20cfc8b45ecc9cb946be63cab6beb8a68cb0a0b4fe1c991989d104b149b932d72f6d2fa47a52b3bfa6e0906c9b0603fb7030fe3db;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfb275c8cbb7b98be28f4d7774e67fa8e561b74394babb7b650878cf348b6b08b0589bb304465defb34f076e1ef0eaa56dd58d2d7ef0e87b0046b3404c15e2010daa0b1a2998ba346123d8a5727b31d59aa4b4b40b9cb4867e1f2ec9660467c2c45ac;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h36ee39ceecd4a9dd1d02b54a18c63037de794fbe9d47894ed978b47d349c111082b4e1234ba9658c432dcb8a720bdd5374946b0780d7025da68e1af972f82010732bea946429e18f9fa3b73192be0ab51b1741b1b9300f108e0b52782b0a90b518f6;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7b662cee3d7f4b6ec22a4ba37c32681de677d8c949527cc4b31f648d05f349f8db63eccefded9f34e1dbe0c782f5b5015910fe9f1453061c50bab564525ebfb708e8ca455d923e9e38780d1fbd1b338dcd3357f622ca5f8bf108976e2f12f61d07d1;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h28dce748ae877436459e9a12ce0d717f8933654c1e484acabd3c2d19037e9529bbe6ee143a60baa57769251b118edbfc18c69995fe3ebeeae219ec987396b214200bace84f77086575eb6fae0599d297f409b26184d7cc1280d3311e33003a856d4;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he724d09f50eff9588f4c993b51f02c25df81e4b3562a19a0d94df39aebab61226234797c40e19ae9232e70603553b085bc63c39dfee9f578e0eb65d911eae6f3a623e9b4268bf86be9606fee43b34f292ef9a28564fad4d3c284993ac60cad9a04e7;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf1fceb51103f02884539883f274778ea938853b93f079fb3a2682e5983570d617b82c2c4d744632b337ed30ace5222eae23f736c997786dd9aae4cc7514439d71d2e038ce10e4cb11d0ca6a9f681c7812a821faa269de32f9f0333b5c6d7639602b5;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc20b87df2b8334890090494674d8d9db82752fefa85fd2b3141b216b50029467f306d7b56d635a1ba4de9655f9f17750328b972156f97619e7ebcb6a3ea82872f8575fd725b0f0cf89a6841466efe740140010672e03ebc5832825b36acd3c6c1b5d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h244630eec65463739e096f29c1e1b148194cd6e02f8814670ce0360a8f281e266c43c0e99cd565b0211861b0f6852724d5d62d22e3a137d25c544382e8585b7bc7be4bce96e699f70672e0f3bbd821b224af37748e25e166e312940cc23aa5be9a0a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h919ce93fe0893f97a2b0cbfb08df41f79d27f722515b469fa06a3e2872e710c15b36c0f1fde1295a4435ee018e6c962cfd1696ae0e45d48c30970b298701aa9574d6fee2a2941de19af30db369566e22811a712dd39d9d54f578b6433e88ef7df466;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8043c82d0132d931e67b2adfefcf6b9c409b2727e8fc0871b163061de7a606eba6e370f3f17b08f18f24491828bbae624cde760b08619eaa773a41450dafeeb1c25f66e5d6798a7bb4a4988356d234c8f52456ef203d2f52137be82e60c7c5bfc2b8;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h357f99b65da85765cbaccd5bfd0d6a5b14f9f15901f1bb46cac79d8e13edb0035e51a12c87eb2709db317e4b778d499d3324c1a661aa271b6999d30fd3ab94d65db1c5af463bbefe66e57643c1b772a5eb1c87ddb78f9cbab958a71b2eab13685a6f;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd5e3c84cb299ff3df8ea0191bce1df388d9c393aa920e59f1670b918629ae64d82d5090348ef20d8b196c2035a2d2c04d92da1812dd2b440c5daa15179f304b202ac7554860cd055184c6de4e3a7c2b87ba432dbea6b7f5d9f68b536b46b21d174c4;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hcfc021833edbf056ce347e4349d55217806d13e41105295ced7031c23489fa5ab1763478179c25d70c103ba591a39d3ca8d931fd595b2b23703615d90c5baeb5e9d36b03a62a8390c28bd51bd6dda2f4d0a155851446af090fcb69f6b2ef478c9512;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h52e68431fa9c9183a262b34aa617446837093119d268ee15fe49da33c0e7d03b90ff4f2b0065dd80a39184311a56f346b03535961a6db24e893a1874bce2607dfff70a190276fa125f7220a730a78e4e86cfc28c34d3f3b22396afdf7a5460c05003;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h497a16126a235fe91ac1f50e715ddf357f50a52a2e61eaa46225338603b08d621321e551d0dd50d0cdaca03e431ce68d166c5420087b287ef34a97d2d2efd9a7ee354b58b52b43ce1324e3820ded46d3de12c32146606839a035d75f840b5fae388b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2b422cb9fca8343804159873db77a5e9c9c36078bfa0855f61f7d598ac7797e3fd1a5856cfe8449d93054dc13d529e7f781c701a77d135ebb09b82ca853c1dcfc06d6ce396243d2a47dd51b34892518786f9bba9773b4014f8219b2c9eed997b930;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd477e9bbeee272778d46b87ecf506c4f00b06cbd5ddb51b9fdecdde3a2cb3897723c681a80840a45a57202d2fc1fb3c4cc88bfe08d13e027ca8f7dfe401738bb92acefa0ddbf5d4673299e416295ea8d46d50f589477a7ddd4cab8b6b2227bb16fd5;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h318824e067d38ef8552b13a3694cf159d54769c86132a40b96afd04d3ffa49c4a92e834e0699d479a96d5f263bd275b03b9e7890c318fc92f4886d21c8bc029c25700932ac010903790ee442ac278d4012c7f159eaaae889d25a430382816366c81f;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8b5bf1028671e752e8eaec9d005c3c77934548288891b82ca43d70bc74649fde9845b56ddb47c5527e17c5da4b5bc818592c2a04bb639f2e7ea591bac18c140adf291c67245733ed7bf39798cc748b08c233be7063bde56b283c37f23d73a6952dfd;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3174574ae98f23a4ae7fde54f164d79dd58139f61c2dd7e7d8066776a53ea641d4698da94739de58e383919200cbc8fd6381ac5718cf690ad0569c5eae0c9821e96f1a5202d0c14525e344ad6980fa81da1119773fb3fd6cce74b23aeb0870e4d008;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7654a46fcc27ff0325bdde6e314e95cfac473d58f9baa8633c65176b612cea80a1638c6370b47e532d8da0efa7035167ec5fce7545252fbc890f81b0b8ab33ff7236a7ef49381d6093e3f1fceb250f2c0b601c01fb4075c6c0a922ade941a1da4ed5;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h82ffa46b0c324005fb8efd8016fe83c238e6fece6f4fbf6e2fd5703a0f3bfc11cf314bc795997034b06df4e68544d0afc1da7eb55a2c432feee0d247146f7e148a45d4f1949a57e8fb0d9e604d89c6b805c10974963b17a9cd403aea0e5163308c16;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7993b9753327f3744df7504f3344f4e5dd3b5316d06191a9ccfdd7605cffacfb17d57334b611fff7874d4f1e65dbe089c07eaca572bfddfc6918618cccec01a1968a2be29258fb306829705222ac66eb204ad312e75409039c0b80d676535b9e191e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hcaa8f306101340e06a50bd37ede6fb01865e44991c6bdeade74ad489c47b3cb0319d378fcf7607a27f3b941cc7eb634226c560548f67ff952f1a8619f7ea71dc379f797d20dc2317f159a41a10529a28bedf8356a00eb1214a14662f496ef0262562;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4f7addcc4b197f3799c345060553aeae88042374a15bb7df68887ecaba8e3a6f96240f8e065b341e65e99354caca5267b6c034dc316f8ee876c46f0862c5359d9d9384766683968317ff99315097b37de4dd4906058f73c8372b28acadca830c1635;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1d350cf689a6def884764fdccf38c0477db7a5bddb1aecf8873376cf813c9fb67d309bc8c3858ea7a9949a6c5a82c7dbc1ec60a6210059839cdcbe27e73e5258131c76930b180dde881a18fd1d12a0876b0255fe0d7bae624d42482e7710026c82aa;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6bc8804d4cd7ba7f50dc2fccba88477fb3e7fec7de43800cf633a2bb4ae433679a72e09a6bcf949ac771155184ffe4438bf31585f28953858a726fea56e3a33a47302b3db0de2339288c64caa41cc77a7ee756e99deb885255f69b389de29235df9f;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h660fdd22e287b2240f6da278d3a246d4d8fe81ab4d367fea14e23b42f0fbab4c82892c8215947a4a1c1b7b114f5518bf0ce72de5051a4cb524eb70407b30df10f2e89d07c8e7780c7e9e9a68d990f2801f13ed219c1d34e5f8c43d78410033fe6ae4;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h63df0929618c81800de602071ab82111a07348b9e64fd3728e26af26c3a2e498de03b69ff6518357863069e8c40af0f462921dccfa7ea13ae50226e48a066f749565c450b873da23844e1709f029538398a48dfc703bbe56481c1b72cf5ec1e8087;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd3e67b4b6e93c13cbf7b1b51d25d46122b55e8c8be15b1487fdce7405aaeea9f6ac8c5a50eff2d5570bee8b27ad15c2bcb85d7b5d23121417e690e7707b0d2db4098e5c9c4a633b1ce32da38a33a9d86684c630ddcf0b24454556df5a789d6529ad3;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h831a80c17802d683bbe13600191c6cc7aa2de1ec1e14a2a1050c3a80b2b9faad5da41664299bc46ec44df840f23fcec9421f00f236cf0f5170aa67df40400c726df0b35e888d0ae3be1ce6effb380275cae0d44d8ab11518b1a0d65e12dae6183f24;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h830c4faf2be86bf2f57c224efaea0a5ad46c2892e0bae04b79eb75377542863d36122b151f55e769a21b1dae0302d1e5ea035e427ef824c73fa9778c871339c4a55d77a07a07c0d6d45ce3ffd920c47dcc11d911421de3528506d36bc7fb043898a2;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h59b6a69bdd181b5d7778aa7ec6e50798f48f08199fee0f739c10182ca84fcd312d302cce247a821e4ad1c57965b68176f499279cb7c58b9e691150bc9e6fc893b4c30d986fffed0896a00ed488133ec2921fe70f9f1a19eaf2b924826004e6f227c6;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h53865f5f700541f758de41e2ed3d0cd47bdf39e61d3b02eb651cc05164033c5acdbf9fe7a760228a5b9086e66422189860bc6fc313266be639bf1f80b991159f1f88ec16523404bff620762633dc8b63e31a1546677c9314a0d0532b442fa5863306;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc7140c02a1df31c1c8732f3778d49654408f7d33a6d77eaba496f71f5012731e174f7f1db0f72f652aa80430f2b5f5f163f0a88f8e21e89770ee07c771ccf95602e94eb9e7dd8462976db860279297782f12e9730ec9a3039a518f30889cd487503e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h27d431c5a6d54e81844650db29133943a5afaa00b55dc2badd899f6c34a690ed69bf374864e8d0e16ed1fcb735d1102c590ee56676461ef774545a1031fdca0b00078effa9d37049fab47d89cf539e419ccb01cf235f9d98f21a52a6107541cff8c9;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1aa722e3fe0abb0b6d3f83b4c2f3d3f4d3043dea98812ddc5729b3ac419078dbfd8a2d8a8260b6a1a6528bc8ce655be70005f497bc018036d8ba0288e90c37799a8c37fa759809df5b668cbae374309468906335141c2b8edd5b55e1e4a23a830dd0;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h738d72820d396a7a126026e32638a0ae612ffae3d2d73c93c19cbcc6d8998f854681193352e0b323454fbb86acc18aca58bf132a0ed6642429f3701daaacd373dfd68bc3affcab73216cc35033fa63743862bb11ac41339abd604e5655d5c2b18f48;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf8d8ac6197d2ffbc88bd2a9e0f138a68c5d10bc669e91f98d370a69a2caf44e5232defca9173c250171bc78a954017900f37cdf3fe66681a1edd4f846c99884d20d7a0c508618a47388221e0fa2fe3342887a79b5b59ad6c0aac415a9243ff3239f2;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'heda5291479f56c020fcae8cc26ac752519a140e63561e874f13f382d9bec156382a424f9fd36022266014a1754ae6f49a3ed8cdb29701854ba42b674a62cfac21e6a9bf8a55435e623129167ff272bb7e44329829e84ff14d31ccb9782472d05332a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h19ff83d15f10a9231403d05e855956ae8b7290eb47c8d345cf7aaef442b5c7836565319f2a27871ff6a4bb73146d9fd2d2b43ad2609c48fe6001be9a5dec5d69ec3dc67dac860dd047f297e36f661b8da8fddc0d6974e547dea0730fc76eec07d009;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h22340abacdf0cea56dd0fbd649fa2a81111eb29682c1c71c54527c53811f263503e39fd2c3d849e18ead9d3e6cfba608205b88c3e0a20b6b00ba35b05e2e8a56ef0d2728aa6f83a4e7f2ba9fb9652a476e51efd98d58db8596d3d25e0d907a91d099;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb2cf265928c9cae133f16f09a8d6fd62cc5510da2f957007a83f6aad43ebd1d60aeb4be75515054144bc57bee0ce98e77cca2303f8b67a6d692fd1e95dd8a229b6fbd6142492697011574db386df7db58d1442b21021dc22cbac95e4a288aac9d47f;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3506cad72f2c4034db833a0a7c0a0d1c68dfdf38965ffc97499d3f55375f8608f291975e37b4735ed56034254d047b7a266d82c2559241b759bad6f4441da6a6bd13a4b13ed7b9b7040126c7cf2dafeebb8df5e441c3bac76496511a7ae74f68cc9d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h94fb3a633442aa7777b7ed5f8deadb619e037b2549bba4d75a109ed8eade386da73e71c3185dbe9f918a781b99d4422f587cd06d14723da615f573929b9ec706d458d99b7feda2898deb4a8d3fc1ebf06787ff5e823ae506d34fde1208cbbd2da8d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdb8b404a12303e9de0d707eca1e1af77067da3a40e8315be08e8ffe67981a2425ce19044b69ab9efabb5f84921e838449367be601610317f3ca52a39ed10c3d5549ec4e28f93ea4bc055b4f1b7f6f6c4885a9c142c7dc9f5231e2f35471b125bf9a6;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h90518d4d18661ccf66649b43c0cd35609b88d8a8ca79fefdae949cabae454de0d42432633ffdf90717656f1b28a7e1aa4b4ffb80fb4976e3dbef0e8d02d3eeebf4e530c5e4bed10bd4ea4751dc0e80bff78ae5074f0084a65567e94e9005eb2df09d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8fb9fe6045039b78be8fa352c21f1f9ca0b3a9dbbcf8b9d4875fa31a81ae2084d12378996371ec35571023fc84bcadcdc5eb58b470f35c1a81917c8f6e07808a87d577f11f6023cc8a246676bc830b01c48814838d2bc1811f72ebd4f54bf2a0f3d9;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h34c619537081474941dec5c87ed886bc906a9357b3dac865d2c2643405d689037cc58e3b47964584fe9a72273a830f23010fb9ae2805012ab0630d9e03a433e54d74bafd002f10cc4c6bbb3537ca5e75ad4996368caae88fcfb58844dbf66d85e8ab;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2030aa41feeaba72ac0084d8fc8630407b4092fd9135910a5b1e1a5644f8eb51da8d44c1224f58c7f3e84a3520c0a77ff3d1a8881cbc2b4b2b58157724b20eef0d2f7fe4dd79f3d9d20ea5f3499e5b5f3496fa8b452f3bb14eec493006a56d5f0bfd;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1d5de741e108832831030b6a2e27dd22f5ad8a71713efd71ad80328a7a2b5d331708c355e246eb450e507a7877e9e08aea382b671762233216a5388b313b33f79ce20c2f43d29fc6ef1558d7b16df206491b4d2018a389935019170ad431915cd5c4;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h44e4a4da4ccdb737b24ecb156ebc65011757388211d310110805a968bfeba7c6643814e52156849a08adaa1a33312094964f99649657fedfa2cf2dc00ef69386862e85dd1fd619fe7d6b2ddd18694a04da194980b60bc9c021c4aa1b0581f7f09346;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h369d849e9ccd4b1a86f732f2c8daf159f369bff75f15640e92763a9dd02ffa46f05f25e7df5c29f8c22be1ac9252ba92aa6d5ee70d92744259dfd00b7afbf44ae6a756ee1ebd6a24b952be478ce5a0c71571d360d7b9e939ef28a2bb8b6e693ef389;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he043791799eb9200a6de23039e5926e221749e76684d5b82e4e3a88dfe0a2872dae8ccd39928ea0445766699f0eeb3449e8f940b58742e729106f7b3a0269ddccd2995afcbc25e97dbb8bbd0e9bc03b88952136d843d7183eaa9bd0472e92f1afa53;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1a1ac3be064b8ac6f3c6fafdc95b71477f8b5241ed8f6607f0205ae761716be314fa4f8474ca36fd9e719ce85a38a13bab0ec4e555cab7c5e373121c0c6b084cf31aaa1b88c6ff288c390737eafe77c34a4716604d14076d4b77e0cc9daab498775;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6434ff5fe3035645854c9db55f9cfbd6b6ac3a20ce2fa5f2264a9cbd731f060265ca988e96fa5c133a55883933a422e20b4478baa57e544d6e27b193f3f7a313b1ee6a26fa42b3a77443ecaadd94f48b75f0f17f1dd0838977c4ce9d8d4b7ae7e56;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'haa71ab70b350218b3e3f8423f015f637f6f5e83ab2a8f4739b0467757f50f11da8b77ee6fa05bc02be19b82da9213b566bb5270ceb207ddc0ad69ddfa8d3e88365f9b0d50f8f4ef38ffb6042de794c20b84e0e10984b6203de018767c4011e0e2aea;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd98d29a2eaba79c823138cdc31e9445887c89c9a2d2ffbd8c3642097039ae829e56f8128a018e3052f527c891522e6e3a650fca7ea875b9c7c31c2cdc7a5a521fac7a053dc23c645a0bea322314fcbccbeea719a4e56328b2b06ec5326a8c4131734;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdb40d4e3b0e31cf5d714cf9b86c2ed7c9e36e88aabeb3be02fe5bc8490bb88f00dd7b8781bd8dd28278f6393b1299bc402b0043f29b7ec7acef017bc86234a6612bf287e6b6f577e118a0e2f2b7f376e46943767df424318505e2668a83ed324917;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8e3d05edbd31da5177708da324440764a4ef638d18628829855d30704d1f10a0efd5ec740a1980fb2ef4b6c6c0df9b81037f662972ae4690afa6120632ab1b4ea088d1f1d63702c26166bf39c9d21974a9c2480b5d5bab6b87eeb35d3f5706a3c913;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4601003b205fcf5e9a07e2d8e4b14053d97c750be1b011fbc918ab9bc7fadc31eee65074ca059b3b1df9b0c89b0c48319809862068bed4fb4765ded540c7be136d4a3bd2b85ad038e45ca05cd143bc559487dfc6819679567ae835e16344ef7fbfd7;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf71e3189c5972b906342c4d96a1872d56e0b377bd1acfe7cea259c0693aac1aa8283d9e8b2c36dd967bbf0db9c17b6f578e9a5909e42be3e0ecdbb9731ddd5e83b7e8b3e8b24f45f2098e7c7ce0a40af6f3aa06081edc94be5a29fdbd0771dc33e0b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4bf234bb3788697e1b55995225dbcf47d803f2307a21f2a6eea6465a153f9bfac62b4f8e0b4392aba8990ce9b20e9f2679f82d8a919703842337864adf540a385528dd9319e2695137d214b6d7520194d799f459e7b312daa55f3e0940a7d0fa1cda;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbc387c5f90c3ee2c332c01c6839d17969c2c6b9e38f7f564149c5b7e4e66568da21c8c39832d0685dedebae6b781f911fb6de53c3fd0494bc97a3a9f8e7b3940628661575f6477ccc6ce261c95bd45bab69dfba6b6389cbc8af907f1332d7eb448c3;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9bddd3a8ee7e63ab6bcc0f96aa45e48b815041402d5e9155c3fea0fbcd80919a39d4b96dbfa51d7cf2347f0f26a16ed0db6f6b27c8ce323d9785f1accb1401240ca1a46080d7d46a4677a562c6112f75f3e4d5ab4e00080eaf18ac687ba15e2d6d48;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8dfedd91029952e5b0f820643c9749fdf5a95d1d54c130a07eedf152baf5ab2d4eb1993d8051ba39b22c2bc6826e901ccd74b5365162c57f69fd401d3ad933d2013eb8dfb0af3f0b223ca534527a87d93cfd73b6ff258775aa355d8034bfd7b0f515;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h596b056390e83604eeaa0536684b4ff781c3d7594db4e707ea7f97f4f069ae7b03821675ef8d350ca78d2a76d22f95853633cfdc49487f53025736ddd670ea7a384bb1dd8ee6bbfccdc81f634c2c2ca5406d757136b3d1f7ea182f2732373ed773fb;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf92f9e3252248c3013b665d89e1b359facae535c45ea26729193c7cce266aacf2473a0d5fcd0fe4a946c879dcba6bfc9f2009020b889d44d107bb0ac9e2c3f2b51055b9ce04f08657cd34fccc8859fbe2e9412f621154f40d10bf034c0bf814c91c1;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1f425b6463d46c9a9b444f896c60e37738c72e46b4c53e7bb1838ba4ffa69c31896a83fdef07e03272d167663a24da0f27770a0ce53f15800fa9f942c4e867583348d372ac6f44801476c88d5afbcb6319bf2fcd20406d6158c7e268ae91bceb86f4;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd7c18f388f747c1034e7a480efd45ab0070c34ff5c807f38a4126b11b6e63d407b8ca0d3c2c4b0dbb5b5368d6b5de12563c2ace42185471dc7b27d301169d028b4166a444bbef4f2dc809453a4780fb5b76bd6a026d5f6ff046a813d108e5bce1314;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hea74674221ae65945b87bb8c775d00731e179d68cfafc8b81da58c8ec9e5744d1b8a0ef76e2509891d0e8e7e38aaaf838cddc779ed055ab74145d95db44433d8226793912f5a25ab917fb3099fccd123ec1217aadf119a40912f794029f541822cb0;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h36cc728fdf4a13603300c5ae856ab415d260a7c77c6e736a6c34b2fb06e92a6c0f58e1b0e198d99774fc46bc59ac3eda43f3766549aa703cd345322d6ea8d0445b68922dfe51ddc18add65182220d4f337287ed977d8454379e6f6f3742212aa0ac6;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbcdbeac49557be08fb1363e944f1ae4e1da15151ba4df3f66c647f5437be319d1772bee5a70197216151e3f4c4cf21dc845d4d38f4a84983f445efd196a6183f917147f52eb2e6381684779e01a5e110011163f3c6d6a05310b32cb741eb16bf0608;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb8ebdd42bf0758df16c1b481b2ef544a1a5b75d244b656f28faa75949dce4d1059b4da2bcc6433d8e3c4837ca891374a0c65a7c2d59cd276b8e815f8d080d0c133adafd037c87e5d92b854674e6e0ca8486e123290b0b992988a6d8e3d89caf8ec3b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h25402d65c55fae5cf6a60acf3130721675f92d8991d2316261d221ff91a77e36d86b6f46c8124872d01c98a6d13d01e35a99932caa7750c770976c989fe0f8f17548a35ea1d5318ba9b33e8832065b05c124534481c007261a99dc0de037f530d8cf;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf83c1f64b35e2bfd1fd797e55e71fc5c3f03cc0c6f1291e9ce06c068cb4a08df3a9364332e33b236126b2b78cece2adc71401ed225e2a385d76f716e53932db1f65d18cbb70a404d31f0babeeb02fb0d47ad4bd3f52ecd4c33467363aa8a954e128e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he537719bd42e88e21dd407e6aa6db2e6820b8d566ce966f1fa647700480a232f0455c04c3e9b2f9dd2bbe250ed887de0675985cf46fc2081365a957f485fb571ab7c9cb0d33e33cc654575b5f38479e22efc80683314cf21b7e81ac98b380793a0dd;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3fee76f9b6f1ba5aea44c6eb8485e83b370046d0641fd180aaded66ed441c8ebfa62afc1d8aad2fb2e2290076e6409987b209681435d3c85cee295f17aabdb84c84d1c480fc12f92e4fe2733d499a2018587f5bce7d0b49d13a455de193ebdab0fa9;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h31820de24faf8f4c8eaac91c2f92b86eaee6cfa2256f275819e5fb5bb825d1f218b9ed04ec1d07e92fe6c28ed1ef98eaeb0591ff5724c6e7ff248ec0e4e0db2ad32bd33cdc9f4f5b2fb6cca25e6148ff3a7f3a7f95ac70a11751ca6627df222aedd4;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1e1691a4a6dbb65908c1e3e6ca1e79671a33938166de76648500cd782d6aa01c8dffc8f15aa97e9a2cf8d960af53c8299a87fad3c0bd2563002f20447cfe60767a6e877d4a3a10c4770131b6c5a1e9d931a3546153c745cd2f33c89c3f757eee5c63;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3801653d1685c477fc8389ac1c032a9fab31a52810d831bfda5f87b8569c27ab9afc2651f14ace51f87b16207a3c991a260795fa34289b77b080ddc78eecadc040a059bd97e8180a1084fc31aa5c71bd1b64908cfea4e1eefc13134044d7761abf38;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h177215dc0ed1e937050ed422ee84361a066e8fb5e24be490812469986887cd6bb532c51c0c944f960a3ba9362e60c4e83382e482b388f18486607946342024fc372195064d6656f4073d96824467a08b729b38f28855f54772f1b16b19e02b0e6421;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'head3d14b6b90d90f68634ee507c39c5c9c7e3da685e2facf63e9e3c83cd0d080c27b58e9dc41ca04515a05a02852e4b8e233fcf6cbca9b548046c92c0dcedfb99e356d0571bdfca6ea2bee176812c32ce3c07fa1120e6f6683da819ebd9224368ccc;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h96b97d055561d604c58595215c19b3acd3844d19718a96d85fc3f63de4a16acfbcdee08ec3a5101d5996d94b9f5aba6c529fd4a72010119aae85f46dad06bd033ca4e526a86caee4c08059c0271f3fca6b3ef703f91b8c3ed18d09edf7a4b14e32fe;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha7d6ae4a209b911bff4e1b1a09b066751f5b32b46644eb1c47067fdcdcfbdb7004ae147244a1061577ade9f940b2852a6c88b24528f032fbca5e7592e8a06ba6f6c01ab0f5ab4f38fbc7a4dfb2dfb7610e859ac96604dfbf39a661f272cd2ba0b523;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hcab4f86309a5ed4eeb96350eb70f1f02eebf548e4d6b13ac63f81e765a36956202b9284cacf5fa5fcf31c3c52c89d0a2af12602191f58b7c7ddc0f736ba6c48cf1ad870014f1a4050e25e8d205552dd65ea79433511a4e06ddf075a0a04fee547e8f;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6632568e92f7293b5e3732e74f38f1516875b5d9721d4c60cc6c555214fb1e3bb69cddecea93ccbcc9e7f891c7a8b13326c46d7bda22a09521c1be97beed2ba07f654c6c3f1ebd1337992dd6a5f550a7c323bc79ba4b34166339a155fd4711188bc7;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h57660df19a55e2627a014fd23cf0ff571d09a9656becf71e428c9a0c3b4f1a10769a3d8e66460a4e2abe47ccd46d0cf2279a31d793a533e34cc8657038705d04030ba48728794fd6507fd35d0bfecf7fd2a5c4b4b27611d124ae6621379e0242f45c;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfe07916fa0f17ceca65c3ba8dc27deea81a3bb0af7fa2739785120ccfc88b44803d5fd5f191d786e30648e6cdf7fdac74f4dff862decb60f79e8b92fa6662d3c2bc6bfed0ee250deef8a6312cbaa51a56c87f414d124da4888d1dba1ca4bdd621e97;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h626385971fc1e5a2f4306b3db60547891ea21226e668faafc1651bee527d172bac2bfd224a2bd092ba3e8e9b642fd80f58dc2f5110f84ea4258b5c2dbefbbcf30ea2e526e7137752bce14bc50a8e607b4dcd7f9a0d60ac270b49f3606e7d93ca5616;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1b66ab7d4babca41f1621f1a9615f2042f48b4f5b5bdef0ccb61587371a491cdab1ebb96ad957ff3baf4d2be0ddb7e577f790e1e84daae2a8936a6f205810bc7e5e3e45120d5579ba084b4ff56a7387e821a6860bb41be3ff9aebe57647920c7d782;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he6467faee572657030e6db47ca3b743ec7e780e236fd7b429b9c13d82b3800c1b91deb476e3cbf04ad838ff76ef7f9e65a6355ae28b683537808d45267136b1693d2df6b1fc4dc0c711611d4737d7accaadccfc38be5ad84cf90195f395c99cd9ac4;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he411a0275989eda9701a942d3eab6c9c0fa3ee1710f9c363a5f2e8c91d27ce7af3fe99262420e480ed2d53db26d33f67467a4f959392c5e7ba33105a5785654a13d58c8389a7ce6e971ba1fa41033b9598535327cb11ef118818e51a1f7559c429ed;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5490a70005ab85f9df744b1af357424ec93164583b3d250d1228fe8f60ed4c8d9146632863c547f8bb06b75cee99931257ac4a900c711dace6bccebded8b550074cce4400867b32809fdec1e26beeca7b910a5f9c237e618fb49ebe084b5ce6b76c4;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hcc448b52632b7a81467a00b46b799be0611c314ac5d3790d0843155dc5ea4674bd62c419c486e83ce8a5ea8eca13163014e0fd0963acbbc89c418840483f6d2984511de471d388f9008dc72ede31d6f99accd0570b9db07d1cc7ce5d5f04d632284;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h596dd61f0e7ace495505f65767e7513e76268119b7e0e230bc9e3c122124f70c420801aeb37bf2cca5ad161407130d0bdd5418b24c8c84257f871610076690b899e10015f0f27000bb824c4c0cc1a2d326ee3651d2aec62f77b36dd665849ce22dd3;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9a39bfd2b8b1cb21057ab43261f883c5588b3ff540bb0233d6464bc4f5afd8babce3f507f1265e0fcabb1bd15a5d45fc576ff7de1f5108bdce0cd01887269cb3f28066ed60c299927b34cb8edb5ddb6c7b39c234bc028eed5b2b7ed11e6825ee70ee;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5b7aae510006264c51dc0b41efd5ef8a16c72f378d445971d0fd3351a35fe4c6a37eae95af48653629d42994c279ad9778518b2727247e5281b6db3c1b049f75c0a7eb5c6cf7f9adba3975c28a24c8049449d4c6dd65f2b774056a0113759fc5f41d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h92048c73f13abccbe2a6ad30922e9c2c9180409e5dae9a4c7deb28bca1ca480a7a7887d768057d85365191a7614e864c7499491f4ffb4d413dd8aeeec8835d8b722efd1b1bfc16418283b0031965055edb421f1c7bd8e8bf0c5ba64a28e2ce74bd2a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3b1a5abcf03c900c2342761aea6cd6ce8605f599e6af3004beb04a5a3241131f2f01a88206ad9f3293674b71408204244d07ec2c60db9bb3baa51bf2bd5263decff104f8dc32a01afa27ad28d3f45c405557d8b08686814677ea51f21a6d034ca836;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5ee47403fdb7bb07fb409bb5b07b67ea45aa31a663da1b28948de0aa413162f1ea3e2051a7db12996482448d88ff5b2fc8a9debee8bcddccd7e3ca43a7c342baba8bea275897f4e6f88787d44baf533ae122764b5a291f8782fb9221a6fdb95206b3;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9bdf0f78e0ad178f89cab52bce49e66a42444d3ae7ac6d27c4f0c548325ee49822f14ad9fd3103382641205b4ccf9a57bb17723949ab140b336a4102f7deba033ff7a76ec8a60c106fad754e00534b71b94f66bcb6becef129dea2cfe3539b3baead;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7b088d167a7e45fbf36b347b1bb1ce3a702b9310f846b2357b656e95ac5b79953ba321b5e82bb901290007d263c3d5bf97741ed852754eb983b1fa2ec376022e98d809fb063f30fb4bc3429db4656f7ffcf810579c12161e57d6c901060603d8ee14;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7cf11c2ee0fd397fb06867915dc15efef95437ebf166efe5a56b35f6625fcfef91c08fc2f0563ea55c8a7f86acb2bcfb81ccbcd030413edcf7b74a93a7e18da8fde9902fa09a8499354efa203ab6bd61e1b726ebf6790d57e5f6392b92c5557cab1c;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he0df00183ec5f6966c2fd0f874ebde93ec9338d06283dfb25e6b3a5943d4f61152f41d05edc19323b8b28a5c4a860a5cea5cfbd6f39b89af973087effe1a97e1a6733e4a495476182a290fcfe33ed0325d3e089e69af531033b4e9e11a303640e3dd;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hffb89e8b9d4bf4c88d821e59282c4c2fed2937fae1ac7ca2ce0f37ef5cabc7288836fa58a4cf9a353cf221328b73edc524754b8de4ffaba4faa31eb1ddd8cc530798586bda37203302179c6ec24a541454b63f32120760783282d89423c16b7a8079;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfa472868f01840c90c7c9ba2b88cf04f6b65e06d5444ee8a2dca3e4d8a58df5df2a13e9983ba2202e0ec63aa072a92b2b0d1d234ce565175c6214fdfc9edc6b4685194e3c4a06e0b6be07c141c68914cd9e4d6298ed55d434d8829d53113e98d7e3b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h50cdd3bc5c2b78de5d7ca2950ef918f8c90a496833c3926848149a177d68887c9b0f14e1f2c7a8cc622c9eed07f9d79006b05a8560f7eb20b33f3694b3f88c1101edbbe3aee2b56a8b81c4b6ff506ad341e3c1244a74633c7fa986c16fa87cbb494a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hce169b2a5208a9fdd54970ba1ab9a3e24860166de34937de0b8d6346bc76211e051687104431c61942d63709b849fe96a7d6866ea2b74e0d0e8f022b7a0de1ca69621a4dbb0efb345d8a84ff9f658bb32c03474e6b9b5f54be598d21eaa71d4b730;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h153997fe359d462471481234fe93a230afe931150c29bbb85d33e1ebefdecbc87e4fb01f566ea239f29f68fe9661d1f6f2f6fda2295f581816e9ce2b27dc2724bc3c4449c31b9a9b3a29097bc07a2602ee604f9385a08cf9fd82adea9288ddb24b54;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h29a7e227463263d55d6aad7752727507c4482a0d43c5495fbe8f41661c719268c6151a9834023ce189cb66e52c943f4d74a5007b565a4c0fa840575b812ac7333d508968cf1b0afea9940335f43ee74859bff5f7c9872bf53e2d9d3bd085346ed1da;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h41d9e15c4292dee559c66f036c15a0cf1b12b33328faf72cf46298fde2dc21d42cf9123153d6a79379c42a3207a296dbaa89e9c6fc043a4c6af814770aa0a11fb5037344c2870e94017edbb50aa57f111bd0f175492e59de709dd98e58ce86500f24;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2be38c4a873b5cdd0428f02ba23afd252f64f57f34cbe1bda82826b35932d7cca07b1cf0f7526ccd609eadcd3ae280603e683b0e99b0c6a0803de82f46ba31054af30e502686135a58d16e114240e8a2774754531a226b822bf610e6d80098bd73f9;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb49fa2f7da4a1b527afbac7d9b08d828330be853c1f460955d8c9825920445acec20d0394519856a9bd84b6db31a68627c45e3af705dbd3a26cb73ee1a9cda07604152a07d5715782e3cf90f50490df9e8f40cfcf7c5d6368914a7562157ada4ba06;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha949f95222f5e9e60e33d8cae8ec101050a1922b000ab97a8a89172e690a9b2ed6a11c4cfc1c665aa858ab4639e447a4727663c8d24e376bf43b615cf936d2204d7722d8834e2f3e5b97f0b95bbeddbb0393f267665bed00b8a0bb36c51babab1be9;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc319ea695a51ae15b7d9662bae14e254422a5c781d9ff637862855d5c810005211ce1e3a226a78a14d8dc8197dba8eef51bb2a4f634fbad527a4d67de9700d9e61c6cfa9c19fa0f540e46e5ee411ba0f84525cb6fe3b5d64cbc096baf84bae37993;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hec64a5690e61521c54947dda4ab42b468b1779e5170f04f0f6635e094d38b9d07dbbc45600efbbfd95d37907137c30c8e26273f5269e66e7dd96f1ed2d65a5cf360b6487e14cda51a1668579ef19ccfc714597271fda76738269b65d3d47f2392700;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9ef2bac9390d8b4f680d6a245766bab626b059a77b855a4199038c7b9b2378ab39922d28418b8ef430dc7f2afd0a41efe73bdb68a1273343da9f084aac2756fd08505609d1bf7ded8eb06ccfb99f295437ddcbcea03563b288749cf076f226564b1f;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbf41f30a8e55d8efe5ab07cc2a7373970c7d56185ed3fb38e6abc4dd6624c4e77e47edcb808a6864e75a75de72366ac0c1ffe668347b51d07034a8da50359a43b651ead66065f26fec914ea4c1faeb313618d09196be81ec14c48373e06c3bd18629;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3dc0dfa1a71f4f65d8de0ca06ce6cd537a4e2027160a099007011fd477915ff0650edea97d36c30a01c0999c6aeb9dbfb76e691b75cc0cd58d9a31020b40b075efd44719dfd6271a7ddf275bb4c54f525e519d2920c4b03a4db51f52ea854d8d234f;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'heb18a4eae5d5549a28d6746ae30e28df626cad8c21f034a26cbe876e334d527c896605bce4ef482575002789df7484dd3d0605f7b865f6fe6f9edb4ac0e22dd7a8182ec6abbff6306727b2f191313001e703f4b2f9d8697c057354d62e4cb5e0f6b0;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h45a55ef520f73676dd21e030369162b064913d26d0774d4987bae3ec530a7576ae4a4e5d188b9b84e025a3a3cdee326a1ce2138a53e4b0d1b653b18cb45fedb8899ef76881d747e24eee9fc63eff993d77609555e7bd9652351004e14ec37a28051c;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h56d602e3e4406d4dd1f8425f8c1d15a80676938e11082687d6b1eef76c0b212b50797a51e3d5acd9698d213bdea7cdfa1e2c568ebc0c0e8f34e476787fddfa89bd8b0ae66ba53039e15defe0e36c9a11387fb4d69f9cb527b1068cd2903eed01cd5a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h291c8c220dee9fa63155794d94c7238e428d628750eaf586d47428271cc33f233a076123a23a20a2ee21079de60a8eec653f1ece1281af527fa6bb34de2fee257b72bf7c91d8cddf1a3c06f38cfcf5b66f0b0b4fd6a4e87d8c770d558149a2748fc4;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf541e2a7c0ac21c15d1c972819881aabfea919657a9ac3a0bb9f8fddc808a797a24b6b555cb21ba9947ed3dfb7fb70f15e52ef52d5cc60e0be124f3edf093ab5cdec9287af29560dd27809602d66e00344463b7e7bfb67feb2ca8662008b5c7baf13;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbf4fe29b2f001f01474de6eb9eeaaeb00e05b8553c3993f5fbdbff520e3ff5568d7d5dde7a399dba6e8fcbec610d2cabfe5daa3b4c1e29f4c5e9de9cf7d133bdf7dd9f6e8069bf1cc6bb7cf706b9ada64323d97a1441ebf5dd4b66d65160b91572;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h40d391d607e048c35f76b8dca90fff02548aacf4a67936145d8729bb286f55d91cef2df5f05926e239473f94804cf54520628e8877239f7db2bf51ba1524c8950a72be2174a8eeb6445e57d9fd4d9a715757ea0223ce017cb8962e2ecabff8603d87;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he0ce4ee4710760e68c3ad928092810c36426079d7e582c4fe317cac3427a4762c3f4ddd9199f39a036aa8d12c1c1105e21ce32fc37d0a219a9bb86c13a1724f5263dbcc8437373436c13b9dc11c0296e91bbde84092ff3c5df9c2fabf5addc3a8124;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'haf408f3c750d76faac927e66d52f605a1686acf226ebdd595e06beec0bc18fcc6f27ca5965a294f4a5019651e8466852b9c5eb64b34423d3e8f559d10fd041a336ec9fcce721b570e01b933e5310b65b06a03f92bf447fb40103d9ddb2ff0b00b262;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf8f8b302be5921fb32275c877989f8e6c100fb8ac84dba8b10f2d588050f274b2e907f25e5c6560cfad34f062177f488cdca0da6e124e9c41562548ae20be840158b479299508a627e9757ec20b7efab3e2b82385f09a415acc322a40c65f884ec76;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7acf96cd3782acce8f5925bc88f017c473bf9195ce9d4264732ba65ce0df431d687287f50947335f1e3106b83aa1c4e5be10dbc2f2c57ebddb8e361ab7b6bc129f9b0de8cd525b26735c3eb3986282cc27a88287fea0e6cfd93619c4fdc98261540e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfa98ecc68cb248e699b6032e47cf5f4ca9eaff09f14da5315172b625235277fb2afe6fd6f071b45aaf36be9be3e9e04bbaad2e5c393e6eebece8e7b1a3fc7bffc2b1da7940547db04073216f60aee9ca92b9759021ba61bebebed29eec6a3c7d4e1f;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he3a68acfccff79e19efc12aa4cf10cedc9a91b369cbcade21c851f20805a2d559f1ef7a87cc7309a383a529685cede6a8dc951e67458b2f4a031313b1ffe1884b76cc2f973b4da0c14267551fbf48671a006299552f057d5e5d6b99a10e7ed42a712;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc0c4d6a96e0add65ded10bb253b002aae432adafaf981c2c32da9c5a20c8f64be8dc177b0745e7f66013c380cdc80f1438ecbb2ba5c7e43fd6a5c1daae14a31712ebb00e93544f6d3584acc857b3b8e40d1b9d742b75a1a72ba1bde43f5eb8e08e50;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h62117d993be890e2c540b8d2e258fc563e05b6d4cb0bf904c38dbb028564cf02209f7069f2e05ed7fd99af732659521a0cfe6fc67c3f30f4d1c0000d9e3eb5aa64e0d587f06f6837a121a9ac5626a30c210e9845f8dd3b1876d9d0da14f038dd24e8;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha5906fd7f2210a85581500afad6a575f8667168cdce35e579abc89dce8766b45879aa87581e84034276b4c902aedf7faf8963e73e8c7baead97bf5c57557989277d86e5a952640af04907ba24dab37139b04711efffd501c797720991f2585eb28eb;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h89db7cc3cd12f460ca1e5aec6736c50f9d32a806596742c996316fd9bc99dd4d461474b9b1c755673d76a66aa31a8079a8a124dc6bda9c754aecca3cad6b9dbe33b89d82c1ba02d38300d542a2ea72ec48ab6e2b545bf76ae96e2dc55e601b5d3da4;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1ff0a8da92bf311adc9fdc52ec977e4db10895f125d2f28942a244e5b2d03ef8c171413ff1b59eb5d1d5d90b570167aba2d3a4f79c8bbd456f3dbc27e91ef2831d243032b5d3cd35281efb5ece1dc413d508bb8723ed9711bb6f659ede1d7fcf914a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1f017738decfde004948dbb4cc34f37dc1acdd6a1064f8bed1638cd60a27c9d97aa965a647d8adf2f60974b6bfc4f0762a855d699934314a20bf39e1238268d8dcaa49695b835ae67adb9429a03717d189a47cfb9538dbde6a675538dfdb7da6570d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha0cee82b7357c220c048f0a8337fb5cf05a05c9b44ac815adf733b030664948aca7d395fafb9ddfb8896d53ba32a3b2ed0e0ca41ec6768a8b5225258f781647dc7638e51b54b0582d90103af6c0da237c2a6e7a3a5b580731b052910d1738256f5d6;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h90af49ebf9419a4ff01d6336d0801afd0864b924b0eebd81d5c118e87c251ab3fd4a1b0f65ea3e62dcc7662e6ab5c79a6a16a3d21c7f61fd53b7d1b362320bd55a29cfe9da0f586aa36ae1174d0310ba4d1d6e09ade41bdf1c9b6c28aa7cce207e55;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb52ffd3d9e584d65fdf91fbf538e3c8410bd098415b62c5b5bbc766c7c4becef488bea3568c3860e05b0e99eeec9052de2f8aacbd02981ec3d35edb4440c8646bc6fe33d87dc5a748f063c12372cbb14b2938ab58488119ff207e7266fb134fb7af9;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h62790d81c005f9d82ae33e476ecb5901de15797d729ce3dc55d0c1bc56003d2cc4d98d892cfcdf9df82c188a349ba36681e9b25a78724e98f0e3398b666c502557048264d359e6ebda6dc1e20a3e95cdc15ab4ef4380fcee330476fa5fa02784019e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he18ca3054ddf5902459e290be3d4c6f51a2eddbd83ef42ddae6998382b94a240154dc31b49db9528f5f162c7a50c5182a0dab718471c44e207451fdc4fa043a7accbe3658d7f1526ee12ae51f57b56928b1e3e5aab2c9d4cb72cb636cf574a739ce2;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h25d9b0c671af5dfc5f0336af26a3a5bf11b987cbdd51c6ddcf7760d2c7226faa20893d9ed43bbf9c2179799806f2daa6ac0246f77544c6179539a832cae7ff0b5f890cc595d42a5ae66dc011ff0f926f033a7ac2143a04584dd24697e4c73de7200e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2678be63781eed1187cca6561abbf3dedbcac6cd9ef6e124889ae8e776419a682ebcbc30a8b997b35ab7364bf81c039d0e90afe5fd0469659620318c38475d766dd51a16c1fc951dbfbddb8464a104b9a1b7bada4239dda09260cc23ef799e68846d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h405db71ff21461b2421d3fe8670d043fb4690ff40e09fcbabace3f9a3cc5a506ffe1182e46ad60bb262dad8a1b953bab95382bb2388a999cd058e71d3d5ca95b427902e9872b8d8efef4c7bda2f13b985047d39261805c911f89bb6355a5f82d890;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he53e97b5ec7deecba4161cc066ca71b61c7a42fbe76046baed9b4f0c62b534465c175a1f3eeee961ec5d32012624ce86725772758f100d3a530d6344fc8f7ec5ae45c7d4ee74006719dafe6d9bd1681f4084615d258e08206d4f5f83c2786cd29f79;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hab61c9cab23ea9873fa1684317a49574f627a3a3e9ad303ee47d1a69cbbe61d150ec8efc69d6384d5ceb64361b36e4da6dbf23084a3bca92cb11163ba2e331a571b7ede0a92e2d4095a0c03b55e423e5282c2129ae8ce0003cf768a495cbea2b8f3;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h672cb40a443bd1eaf8a651cb6522abf2d5af64746929d0068ad98a08852628129417c51ffa95fdc1e5a403d63aeb346d9b58fcb194a6e937f3bb1c4316704af366b2915ead097445c27584a2aff92eaf3d3b3d60d38297de27d142542c1ce9e160ce;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6726408268fcc4e349048f96fdbee1c1d929abc76610059bb982d420c89bf6939df203c12f76cd7bb4217ad2fb2f1ccfbf9250aaf364c9bdfaed4791c7aaefe01762f4274673c1c7955a3eb43258b613d1a3fa6caf79e5e48dab263ea06cf441b3b7;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9afef84710abe8d469650d11f7d9ba21fb6bc3f5244a055a7aefa308573212f73a7d0ae61e93d6de39503cca414cfb60fbf0f9b8c92c0f9d77764801d9927ad2206d0a1a8bec67571d96da986c6625a91794e1341624ee6c7ee85b09a922966b330b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc0838356f4195393fcbf081005ab73099611fdecd54feafe2787b850fa9a2fa45e1acc4fb4cb4dfdbc7f23da4c5c353fa0969a12d83f82e8e6ec70b7002272dac19728e5bf5f7053983860862716580fbcea9900ec15936a0bc67a3597c85ea49728;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8f37227bdf29851f33b32599bb435a2bfc368195a48c586aa33dc4dbc8e67103ad64b43a7b2b85311e657b50a3defd8f51dda3e083a0aea8bb16758e42d483008c4836ce6c5ebbf295a58ca2341073b59867691792f0a5b051a1343920f61443934b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h215f40f65e977e2f6b2fcc8159f13784ef867a989e3065b2fdcfa9cebf22bb3502d3cec3f496c7ad24a58fbf98417a03b15d8a578932c229edad9dd240a74bd7b11c299a69d2d423f1e8d7cff63cf6a0b1964acd5824f3d387a3a877114579ccfd4b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5229fdd1e6d5e7243938ac7ba89c1e9033c0c4b288b82c7eafb288f2970f9fc702ef8d8baa8f88ec0ebfc5affc906e0502e22ead1d6b81fb138c2e8a778ca385c307bac4bab808f85558df664dd03db1d3c64e9d39fbf2438699b8df3bcdf1f047c8;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h370478a580add168ca4933665b81cb92212ba36da8c47adf8c4ea9bcc379de76f7048a4ae3e9e311edcd508a70dace6be14401b20d7e8f68c18ca44184acc84cc1107bbbf655a7635e455d0a381c85f595a74fa98d4cfefbe8b28472a8c297ef3a72;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4136f535fb7c3e45ab7a1f43de3de3b791f169cdc2bbcb8a4264712d619012ccded01f471a6618b7c212e3737ddfbd2a6f110e65d66116bbc33efb9e8b416fdfabb63296b6f43fd3a0b57f05fd65bac6385e38640d376e489557cec2aa50461a64bf;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha3caa7c2589568e35366d433f2b60dcc0499c2e456362385ae8dcb161814ace83f64fda7eacfba0c44c1bf98c3c348ecd9e9e614ec9e4c8fd19907359d063e1045b506ed297dfc13bc8140f1d6240fe68c74514f297d3a28c9a4e83f5952332ec317;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbaae3b54b3a9c417e7bb0ab1027bd0b6d54fd6b890c51fe737e2d8fa792adde3b12b42511157090e6cd72d2faa2db9f9066aa27a3970fc7d442eda1f83f3c7a98bdf104299a8998237405a59a7b0142a0e2753b38ade998d4122fa940f8c8c82bce2;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdd68933b064511b52e48a59c59ff5d7ceebf86ce7988f3e61f61bd55d7acd2cfb3dd21c214d541d545dabfc6e6c3fb11e6275eee13c88df123854b7cb0cd74b00e57adf1be238ec01b713bbb6d34f862239c84fbdd144c4342d31169898c9958f58;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h957a25e625f8b481571348dab66f5d7faed43b57eb303a3c07ef2563a3d793529749be59f18c05aa95afe33f04c3a30747df2ab96552f0ddf465b0108896fc959b298810e7b46f46b1b330c7cd1fb263ce53ef6d604619f2a6b8fd4f45c12bd52eb;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he551301ad64f02f4d63014400fd95840ca357edbff5006f63d6b6ecbf47ee805210f56b4a9952a3cefd61d3bed7a43a030e74e450b57eed6b43d968c6436669899de44814d108934aa0d2da6352034015f2c0ee1c332901e0d4926a57dd8e1aa75d9;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd7123a250b73c6f867cd12fd11028dc6fd9301a372a07c7914bf760497ddf4b0183af48437382e0d565c4bbf863a720bbe5cf2208d364a7b017eb9d9f972aa575730ae0dd7e9624bfbc71eb660e77710f42c456c5b3b0dc1fa7e4e8081ea124236e8;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7fe7296510da82ade4c0e54924b089d646e5e14acfe1393a418a01767765d58a47e88171658fa1449bbf495bfafd4a5733c3d747c0e8b0fcb9ae2cff0001bb992be677dcfc427c130e93da5ea8a4e1682a8de6d9af48a8c0fae5aad739646326fbcc;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9fb9f88e424aa18729f5e82e439b255d8505a57ac025d06809aebff234dfc366784fb3d0b830be002e7c3bd749e6f37f02d762662dbbdb7b285c963fbce03bf0943b8595ce4f6077ada7dd2f59eff16856804c59edf5546e8e28dc787c17a7474396;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf1ea22ed0fe87b2c0af754827df9df8c23bec13e0fa5d45b54c767f71ac97db68e382ac8a1030f902182df6c457e685a13602ca81e6f939198e5973b4f58530de597a63fa8df154f04db5c99342e1d058ce6c09caf76fd57cad3e05e4c1eea739b05;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h819ea45b6c09724076b8c2d56d6a3df80c3ef7828bb784349f1e714342840c1810460a0b5d0a4aef30747229465e1d25cc6366dd684b67c382377e7fe1aa7974202d8f7bc1cb46976621809b76fe2db0be923de3317ec8a0482e29dedeef57ba4b03;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbac299f6f640e287659fa00e758aa8919756effc2a0a4f3690831e087302cc999cb24cb975074c19c2b5800d19227ee6bdeabcaf8b092e894c175c4693d12cb0d9721de5c70f4733308310c991118ca9cb465735112aca910bc3819b477e4ecf1b9b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hef074cba683929205a1ca1e972ccfa1fc9b79f749605c883004b5dce84fe9ea24f1f4dc43e9ae0e1e35dd5264dd73c19d77450f6a0c8b551441e45bb43d6b78775aeb1cd460972f8583ba45107392ef205686f06c495dfc09654f3ef4c7318f1c174;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3cee516a263a3da502511aecff3e926cb35240ca6745f0d56491d6c6a158a87878e9e3fdcd619e7cc6c24d1b9b62248a6107c068de087455e19e8d96409d4ecef58921e493150091c76f7854a4f54bf3c8322ffd001ffacff7e384250572fb44ed35;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc93015ac19ec4b518b0b8818c82a0f0ff4029d9bfbdb3143556db582817be4b6aa22be6c4b02c3b69c835d7ffa2562d8f812c9c063313d62a5d7bbb86813d455027239f6662803033521f06c7176aeda4e5415701545d27c4c99222e1e2a700928a9;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h284982faad65c6d92dacf3c724f9a03979ddc56f5ac225867b2106238b31ec23edda10a55b753a2357d20a23492dfaf238ce51a208a4ff5f450a706725e62efcf193ee46d27d3f2a4ef5a8f557ca6be3cdd00b6372b1c5bd8cd37cb1d3b4df946e42;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h34696b078fce15e536bc93729b2255a0d5ba26ecb6ccd94a4a632c36564993d1070284baea18c2398c79c69b3c10ac4b7bb5a025deaa64a72da1614168239e49afe9e1f5d6f685cedc62517330b8f96ea1ab42e297fab3b450489a9b8fcd7e2055bb;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h637be12293673379710e2a3e76a2e30c22366c0103e4d37af245cc2345bfffae6722578ff2d4fcfb96b763b6aebd4aa11e8409befd2823b4777b7ef3b5fdd37f7b21ab95b07abfde1068732b62596e695cf3299006ea5ec7d6e67f1305807855f8e3;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he599cb82e6baa4ecda4326207fbb878fccf266429d33e4b3c5fe48f988b2480aac9a114b88381e4ea81cc18ba468a441484ac3075ff63697e1eba2c1d7fd019807605797698614f38dd832df8bb26d643021968c32328dd3248c1d519e49ee23287f;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2f11eda7bf9efee895e1728fb075d2bc7bfbda36471b72404eabd106d0bff44f1f8055b211ea94fe7aedb00dff0ba25e07a44254b100ad83a910ed0d1751e300e5dc25f27398c157e445c473953f73c8aec5c9cfb4ce448ebab22db131076345137f;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h946b051536bc5c7d6857f846763beade017bd64bf9c1912629d2878b10004de8d29c2f7a28f43f14a1ea067e3663977214ed807213035ac49d554eb5cf24c9dcb4807c2f39a0de7558ab70a6a25b4cfbc8c84ec725b5479c7cb70dccf4cb53a1c2a1;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb00084c0cdd348b3c70528a3c6b59231fdc2fd46746464078f2593278585ea2dc3197eca2e9f3877e3c3c20d508b0ca77951e34a8ac8dcb1658046d7f8a35aa6d7b32fdbedd07d6df2e68049382a1d708027f9b4941039f8e126f2594ef43ef340c6;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb8e58fa705f38bb26bcbd0ee6b137c2fc2b9fdc82f82c439b9146cd822b64363101b5941d889a634691a9ed41e6be06463e6aea4b07b3a680e21f3a919eda6cea33a5e2a8fbadf903591a4d0536eaee77c41035dab4961f6cce9a13e6b713aef5288;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h931418c6a69711d499a955f2827de54ee496c0e1d9f51f27401087136fe0dd6adf79833a3b1d57e4f6a0b51b686bf161e904f63165edad0976c164f3dfb1663f00f1ca787c406581c88a764a66bc000f692eca09637814b14e5786b29971bfbb20ac;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h904a33e11233e44f8a41f2529edc83edc59a5ed6d2213c56edf327973ee21b75fc35e01593d37db76d2f1431c1e6e7fc89e74de0c96da4964544fc1e6eacbea32c2a851d964a477c6dd30db8315087d6618646a7ed0c1d534773f5b5891b19bae35e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hba8bfc1d9e5b1f74dd76b129f8f89dc9e2e859487089531f6bb70ff8472b77a1520f6dd43c8ca0e26d32d7404c6d09b60bda22a649c7382c5187073638fe8abf6d460965365bcdef8177491a2602456d73e0a61bb099be212aebc292c6370007e472;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hafd6e1293aec9f08cb87f23e5cf4ca0d28af7fd935ba86706e6d97527b6885d036a53601a4e3a8b006d2552f425b22c26dd6f4261413c4b65fb353fadfb9b1c712b3d2e08c8e56b0c1879ceb77cc2ffc1991a31615c0b5acd4c8aab06317b6699af4;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'heef54ac4594da75b6aaa698ee813003933fb5b8330334502388cd41d34e7f0153845612cdd259b6eba694d625426187b369732742a187da767577808384cec1ba6bbd461688ea3b4f8b0c15a52aa47c27640143894e18f4272b3af5801ceee201a33;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb693389d57dd4ca6220814bae78a30d9ad6c3383e4c8f1bc9279acc40092083c5ba52f32d24197d90d6b39fb4c51ce09b565d23ec1796d94be25fe351df70ba51e8f137f5e99002f6e6506169ecbf259a74dcb3b1ccc9f0e10e0a4c96b890cc8fdc8;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9e20a9fd90a488ad6f9a90c7d1c693e5dfacbeca92e5aa0e9ab10c60227912dc2d9407f6cc5b6b963f43f099e3b64ab8f2107bcc7c30a0a1b8fa66506161ccd53a26dcb4201b54d4f99c5ad3fa8a6e2cd969967196f697f8e64b93f8a4b4e4fd900d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he4435aa015ea2dc1b2577bfb062a2878d104ce245f363af8c082b559cd6778acb26c695d0875ef0c1aabb9de8cb48eb740c144d7de02e7844dd86e45faeafc1c824bb683ba7f5d97c575e67bdb90689924cbe82f3448890ab346aeb78c468747a6c6;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb372a5e9d527aa89c1c3b1540a5c68b18eff7e1131c3467db70db575d4ea00d8e56469cd97fa2066b32a7f56928d2dccdb7dfa0075545404ea624a8cb6c8ccaced1d3e78d2e3ed8fda4445882bcd6fd93e74bb9abb6eeb0c540b337182eb32d9c648;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1a8ae31d215e04fb4374c32d1f5f3e984e14173502fb2677e9987366c2f45633aa55b2515b8310b49bb946dc681dbd65f4ce99b762e93a88661c2a9b2cafb9c1a9a598c18233636d08f2adcc9ee45c6bda2264e3cd73a9e591b1b10ff872a38bd4ff;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf7de0682a2b29cde7e2577dd372d5c1cea66078d4716480db9793526f497f77b0dbc5550634d9d7e82098972b3b3b0ce996af2daf865479868ca73b032b33013397933c1c6c43ec98854465d37ac4ab2382a81ce89940d2a7d841f6878997820f085;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbd7dbeed76430a15cfca33187465f38d23df52675e48a87aa5d01c6f284d89eef2ffa7efa4546500c77ad3fadef2496002b1e0f2b3bda642dc25ad9d699be6a20622cee8a87546a5dbd3beb83248b06323b00db1c6112ae2a88234633ede5a369ba2;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha6f8f9a948ad7de0d9643be76bf81a2b9b78185f75362f567846288bb6e0adbab6490afb576400c84261c00e500a6b7dd93115c76d275acecde38468cc4984ed6d34b8d3759fcd52736e1c150c3ae5bfbeceb7c30d3704af876ca13b42730d36bcbe;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd4282d7b81f697bc581ef71e61c2a3e128da87a4f3f143e878a0b7bfb54f00bdd0769fd9ba275a86fd3682c936ac556826d943368c2f9c0a5dc103c1a1e661011f36045cc3345df454ce787f994d0ed8ebf78d83ba8d467ccf338eb27ba56de3e81b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5e15bde9422f9b70ef9db016fb5c36c515f25beb02b27f54b0322bb1b60e2dcd2980cf0599e0d64e7550e527b74e88849c1b44755704604e22f9e7d2bd285788cc21dbb86e01599cd811249eb901bf1a87535e359c159d92b6ad9c3ead8f97ad4a3c;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h262df23322e2e328c882227d35bc99aecbd92b6c585c685a1ec9864a53e477312699555e1d0b1af791f37be8c25987e4291ada1277565a7fd8e7351a95228b5ead2bace64d6812998cf9063fa3b923b2f22075b464253ad3e3866a57cee74cab3c57;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hcc3c3b00ee7adb9515bbc79eaf5c7d26fae14650133ebae77cab1370e53869508e6180aa54da88263d325a16536fa349acbf5995da4e61c634e2b90604502584fd6ddd2eb24f7705f4107959267bdcc2a3e5b9594e72cfc5be309e3f5b5ebb6a1bac;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdd3278894eaf9f5cfc774aff6f338e9f648b8d01bba6a882d1125a2910dc4a0fa97fa236480948b4f5397c13d7db0b3913afe11716d5e74f4596f93231c69e40f75770fe22d29cf24da0a3973284854fd45a102ee7dd117f555878e9cac797ea773d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1761c25b582118242b31dd4f15533e521c1d645ec9f69ff893d45e01ac8cdf8b1fafd48e89721550a1598cb61fa3c940a1b4a1d051cf7127b8f080c8248b5a0395afcb53b59640054d4fd14f8abbbfd844b9e768762995cec9ffbfe374809e081b68;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc000b87ca954b78a7ad96de0d747e386dd4b770db627aca125d86582225230e41067662cbe8e0befc21894d23f52cc50adc787cc92494d09a8fa527b8657c7947527e3de0019826e7f08800f7f59b3c5be47c882abf7747f1c3d41b6a7fecb0d4360;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf06ffccc8c14c5c524e87942390aaa86c9ed371e0fc85eeee39d12e4d4e493bcc02db2ccb88775cd0533b8c07b03d7fe2cde2bd28c9b71d18c4467500b8748389d13de6f3ec91dea65a6f56181d0166cdc8315d3723ba81fe87b1385e877a404db04;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h17f9490a2fb6090b4b0a54c7a0e60c330c6f4d99b2dbb81fae2bd9280f23d56fea5d04f25c9b9175efb1a870bd4f97f5ac6de14ad017eb4d7d388f06a242c830a207edacfdad78897a38633d30deb7a32e548c78b60cd8c586319e968a4a088b31aa;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbb72771cfd72378c312451be02bcdd27b7a1cf453e89294ce3809b9c423a1cb0a1920e438d96af54018d83c061a494cdce69cdbda9985d6663ccbe7f6fa6b2daf5aa55c0f1dbd1256e4e20896d9abc0df29d9bf7e60b038454ddfcc1eaa67717183f;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hacf3398a0a887e6f1291dfcac49c0109d1279247cc2b16aa396a518344c07219a839d12fe74e3e4b935d026424a7348cb4a9028f053801003b8c78ac4ad28f525d8f6c666de6321147673f598f8c5c43e2111585e3ab7a3ec4792e38e0a01c5aeabb;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hff3d8ad6e08419e7c13e7c2ae9af173631e4b07b59418cca47a6e541a846167ab31e06363489ddd96c42c76a3f20323d3ac8d07cfa6f6c44bf9cf0f289cd163db01d07e6aaa6fa00329e902824a38eb2528fd261886e944ae078fdf69f5932fcd81b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h66abdb14d7c698d78b58c4a6757d13ec26f41ee2ca25bc9e2e97c966934d16afef3f4d26eb5412bc0ffdf9d63b4af0297426e3ef94564883cd3b7aee4e735c9256b04430a44d6aa4f8ddd31d1c80828b5246b2e4b9840cf182de6311eabab73036bc;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h985e6f5eab330534f049d59a2af2abc6ede52c0a37d289960f4a931215318763cd5caf004e631cdb21053407f72e354352d3ca76caeecfc5fa97fe40f406f1c59e106a188595d80cadad8174fb5302ae2195505c4a2d42ee5e39765c7f1f1c53215e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha9193eecb133b6428382c0bce8b0e577de543a1689dd2d7c67205bda1ec64af79278c5976e6d0cda9c926824d96f48f940f27bf6c79d99f2b355063c347dfc5cd32f822f9f28f060c98d41676c3ed54a0f7b12f93d5a95b433bfe970e520de5c2af8;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h623da05552699a98e4c728fffaab903cd5e6882e9aabd0643fa85d9a1fd9291087f3d62c638ad9fe499ac5b9d4ee6564a981d86a2ba6a8308e6af16e052f02a92df466cc73c4f4cbe50b8923bf8f8f55ea15c10e491cd3e9a47ce835fdd183ec5e5;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h374db072d2e5b7ec490bf69e0555f9cc3bd7eba0068e196561915cf65cb75f1a7590b2aae1b6157b47cf2fca4583a6b4bde8555daafb4c9612259b051ccb302086dec3a14fcbb88febffc3c7601753f0e0a28469085b0758446d7d9878f14f669eca;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h89c27ac6b0d584bc07b2446be11719985b80eb45daae3e8ab45d4999c6e3a155e7eef20551b902af9c1181d94b1b24a7bfccb354fc212bc5194567ab1d66629f7afdfa15599c21dbe7d1bc3c33f3bb9f76a584d177bee4f03af5c00a4fbd2b8351fa;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdb79a9271f3c7e9b09546547b86d1f080535445ae623f6fa1af1b38814635c408c04965d300335682bf480c86c2ba16c2f5bcad825842ef0c2575ef40adf9aed4c83867eacad36f374bae40a9c3cb02cc53770214f3f8e926894f6690b9e94b19f72;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3921544607f0f7f11fc8c8005780595efaddceab2adcc3352a0d035c508116c40215c30150b668eeca1522958487a7d214d5d6cd3934189229649c95ebdc57efeffcb2473659a8bc3a0dceb9d8095bef5958bfc9f053f903b5300bdba8d9f1f6ddd5;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h933cc4bd99391de35a072abf069a65346540a904f3affae07c48d5630dca8f6ac7912a9519ba52b517402789241d6a7a87be6121641bd7d20ebbc9b937ba28d4deb8683b770113d3d264d790cc8c5c0856d777ad5171a36e8d4476fb81912f60ed45;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5574309cc429d5915224cfb18cf6ee4fdc20a2ed3bb6686e3a66e1a3d844ea5e048acfab10ba28289d63721a2493d9e2629532f12db983fdb97d641182fbea96371194900de4fe67b998d8ec8dbbe2d775c10ff54a7b4dbaf155a89a1b138a842a2;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3f0d67de3b94b780c5db0ab6c6766d6719ad7a69088e9720844ad67f5bdc4f70e2137e9e501166441da974b63e9430761cb579f470d2f172c0fadaf04cd1f91c4a03ab297773fc1ab9e9ad74ae60a13832ea74dea798bf6cadef0a26cce4b7138ee9;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he17d1caf8d23ca88b9999ed28dd95d8886e8cfc65374248002c05d1592382748b12f47691b276f963df69c5abada4e01a944826114d42365d9b4defa612f3e034e96b661e8c57dc299444652465f843ca8fb89be85c090be7532bb06d56bd927237c;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h712363497dc8950ab2745309e3dcd47529ba958a0658f22b3a1951a6e636163ef655f6507b6adc7eb845339d2515659d9327f93bfb42ede76dfcf0f74b565e823195fe77466298ad63aa9cfd51ee8ce8f6d7c63661316ad3e630b98a7ffc7af80cd5;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd879067f274dc6d3d22b3109fa884bc8ce3735d7a85d56f656a2297b67bcb201d2ce346bd4214393fa5a35645c550f74f33afb7538f274f3db7e07ecdd3e1e0f7b477edbc22d66178882e5981531f1ee9f733384a72af1774735dcd37802da29a38d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd3c958dfca3c780774541562359cca7065163594768182d29eae7537562dbf98b2d48c2b873c6f8c180fd7b1e887c4d828ea59fde86c9c82eaf3e093c656b21c810ceb648e6074da89ece0a21b1efa2a1eaa0758867deefb92060860b8568d04dedc;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h414b45f398411892a9db3812e003ec0092586f0f310d280c4fc35b889558cbaed907cf85059495c7623dc8f76022087a64c761e6787160be34ad97267e5d47920fa8e2b748d2f635b04a7a2613fcf280a895114d6099554c2330c0b6f04434a31065;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hff083865002a2794b9888a2773b97dce80296ede06fb82302e4162718de56eb5f9d108105c9713b68926c63616965d31cf5447154a81cbcf19410fb8705f36b3c0226877513ffbdb545ba1286897f21a5b56b9d7f0515dd9f9dd88fa0854dbf7f738;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hef1b56ad182cf6341ac4a84b60d50e099812a40ca439d27a741442df9750965e54b42b8e4b040bffdf6ea4ff0f646003601bfb1a09d700ee1b56430ef2ad7f677a65162d7010bb6780623f1cb9bb836636702bd92019ebf8da5917ae1283a382579d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8af0d8157067a86921d9c47254470b494d87f26b002b7ea796a287dbf8ea811f627150a82646b1aab2c26251885b54a1ea80f0fdcfc64965d2269e58237d7b76bb277d35af9105dc12e59581e3acf94d6190c1725c1983f929df2b4c3d2148c921b4;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb1532eec1ba39ca4f1d53a15a6f2099800f3efc4febf1c05647ac3ca81b167575697c298c5321851009db131d60a1031ea6672fdf9862b8ed69eeeccf16ba21f3679468555508c01f2fcb1b7c3ddc2a2613ede74099a33ca2565b951d4b19438a44d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfe27ba69d849f11e081ba3fe9dcf25543027dc43eda5664df1a7817c87616fc58edb385a13c96fd2817ad38b5853dc96fbd732c046855d5d2a7d2c2d25c5f015f83dc7e402f26b7f1d3eaa92262bdfa12f79329f2b96b2447352b94a4fd7c563c6cb;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbf0c72bf99435fb5a85b6d02cf5a5cbe6a0416e623b5b590ee3464ce5a0a9eff5a38a8af05de9bf271c5ed171a0611e0331386776b67bbc7018c03cc70bb8ce993432ce1e1236e9c1f84fa08506a0a714e6ac1a9a94557de9f727aac9ba2175d4917;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9bb3b8ee216e4ed896c4526c5d42b17fbff56da7bbf2d69803bae9a3ee1f5578dc6a71d8811ed038c0e8ae9800546f8811bbdacd96c16343cfc77811f07611046e8c89687c6307c68671ee0732035556f5fcd64d346f6b3fb12bfd035cb0ff36fd95;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4043eb8b037481e9cff6359dcd6941dfc46a64a0cf5d3cc1e3e6e5ab73dd1190066513ed8dfc6b03b819c316937aac55019942979f2e298013b841b3c15737c1b4a6c0ef74d514f2aa32c00daf52e14f4d34a31ffe9e4371de34f3f37f046c879ebd;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc6be832883aae29b28a6aed7d4cb2f03bc5ddecf85c1a8b191964ba4178675eed04d4685322fb0bb196d5993523f69f190fb1a4c11c13bd4c8000bd5d924ebfa3fee61f82ab5bdfae4ad1ebeb5962cefc48f5e5d9c522bab91843c2a9f7b036b1d4d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3236d839af8c3ad6d9f5d8aee3289f376debe087305d825c92d9c65d204875236631091192b5079aaeb25b666bde290e34bef6e51dce9604d71d2a2b1014b1926c6eb2e9394b6f76af402a69a3736719ab02df1f634e6c39a3b74c701b4c88474317;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf541d00cff39a4834dcf3e24f678cc25dd26178d1cd2059413dc9d53679686233c8f1522f05f4fda0720d48d61e94e8c3da48795e752366ec9ca0cc093bd70aa6480b229e37006e2f23afa5bf898192abb099e973c41469900ca438053d4ba9134b7;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'heb49417e2cebecb10e14e5436ff7a919aa6cbff799308d7c478cd6b44319cc5f0cb717126777b94be435ff6d717e93db589d6195d49094c22ce3bec21145822510a91890f2eaefdba0f1f9445b622e6cc81dafeda81b233ab24d44a63c9b3df0ef8a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1606db9627d28d703a74cac9a72352c92a7753a2d1c21337578620aaecd9bd50d5e0c0abe9e7a478a5e704f99c040d290132b6fe49b308d839b3d2646b7a1bf1da081daba9d1b2123ccca44bc68a31b12a148757c0cda25d5bd41c66306f425b9b2b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdeaa6c4e03849082eecfe1122536994cf26f3d8f94b637c8b46c8da099287bd726686d82d1f3a334bec2e50aedd6ee422dea607a8a23b88b80069131a5ff1e51da7dad1834bb6f3e3aa141a5d27a6d244ca390bd095f885e887bc21c7544ad452ad9;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6e6b6627149ebcafbe1f0ac4b0b3d0b415b9e4f12a5ffbe69c9cf849c13e7daa8d692704cda7928e734eb7e7a91e4e100c8b8b799e242baf713d117da70319848c1125eed3661b6cab90aa815d8372c5c27088be3bf19ee9b7f0c3639a0d9fb002cf;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h83af683fdcef8ed8516dc057f229cf8b0f3c44a15ccb84e6c4842058af95d42d3306734ba5fc4afdd8665320a4d647faf0dd536db2b80c41cacb1ff1d2f93df4d93f8eea7b86a956f35561899da28d855c4465507ebf2bfb67dc6c1fcc57732b37ff;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hcb88fd04c7ff38ff5159d67443712f300dbdf4dac871742a7d5e43f5dfaa20366436556adea10a69d0598904fcf69c8216d05973aec631ab712551ef2861def0af31c581ed115c8322a309febbe7c96736f695d1180aeb79c97963985bb9ae340692;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h32623be1f6a2dca6dbf60c83713cb9204bda981a9d43a0ce93c3ec3d9da87a9d7484796afa04fd6a72496344121db537bdc10237d8d80bd544308aef95ffd66793832e7bdfdcfa71eb73cd4038fd253f63f8a709e17a86b40db5e2aed9adb4087910;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4058aa36f2cf64074c8ddb1cfce1012e2119e5342f9aa943bc594208328a525f5b4ea2f2843a9569cd74feaf49d25c383a95200192b67d79afd232bc486e1704fbf4be7edc997e3d73b1a6c88e54c97be2a3f7360cc0a093950564a3b62e9c446e8d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5102c8617100de811a1393e7b03d0e16610304300b6399230c513bc532a16e41a632a1ffaf6a6b5704d71c5d41e1260f2c4a78245f68658e6ca9ee9f156842f73062e2a14f5bb6a16cf7ef40a105d0da9cff762ed9af5380687eb8b73a35aec7d55c;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1ac4e4dac4753ba3ba51f091fe916eff51be72c16714d33839070a05ca2ee58694ee2b840de86bedca96513157665040f43cfc752fef6b9a60f3807d7ea3d995c1aaf2fa5e22eb86b5c466bd73dfcb37a6cb130757048ec4851d88b93bb19cc9aa2d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h63a4030a632d4345aa7eb87a9488e10f40a3a128d54a75802b6365a9f99b3ab97b6e4d7b6d419027c86e7a8d502de5845e0ecf5bfd1d2cb3226e90517ae987adc4d225220661446ae16238f93cc221323f2a919507d7014674e6b206a858ab6cd7d4;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3c73d8ab315adcdf8347d37bacd86571f4df496ebe9e4e9dfeb37cb484bdee0188e333ee6156632687df0bf672ab3669beca70abd6a9d5af0cbda673e420f720fa99c304b220bfc458ffa478b7fd4efb7c8bbf3ac3012c105753d7dcf4faa2732168;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha721e18e26a46043ef131962293533275822f9a7d15724e27eeaf47110c2fff7d3558e0b792fa969562ffcf84c633956196dd320531173f43a0749143b04d38dab93fee4a3162f2dfb100044cab854fe8b4c0f13465faf573a3eddb3847178b2e100;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6c30229332cb26f60a3d270d912cecc2b3636e905fc3cc7e3e1325acff13c5af89744726e47514fa599a7086776008640aba2ed05bf218c69fb90d8f564b18b6416360b923b935441526b8c8e0f00e9f56271b2e194cbbb15cd3e577173eeabbf46e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6419a8ca3b4d5651e6fb14eda9e4c324f0f9deb2d52b9baab91bd3f74181baafe7e60b8f0b4fa85157a65f30e03a0f40067a6c13f22b85cf75fb3bda2c5be87c05004fc8bb8348416870687bebd455efbbcda7f840a2b3a18f39d93709852e9438a9;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7e15dc705111d5f9fb8a3a14c841d6f6e7b1bda0b954b8fec78f19da041779248e82617b4d2d067302a294f3705b1523bb4870e422578e8ab67610379ccf732c34402733f2641e0d5ca6a723ca887e24b95abf870c058246bdda62a671fe2b9b949b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd66eef2ee92886c6445409adf2daf145f310ee6021ecb74379104e5073861920ce7a6f463105143c0c72eb57fe9eda174b8a98d838772ee0c2548c27b8836fb5fadd0d7d378942c28e7e3818131a325f7d8efee89a9173bf06c077a33b6a9e56b5a5;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he1feac1082f6133794d79bae20404f189f3217def6b3650459cef9a497636520ecfb6a0d390943a569c87f0ddf4caaec2b6c908c0afa061b340343b443b40ea6aaa5b2adc3040928e92e86a51ee673d19e19a9de04738e2a267672f75b59a7387f93;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8add5af0ad569307274d60211f9b73f1ddc8abadbb3bb79c424fe7b54fa2e70fb10797af8c259c5aadffd0ffe100d210857ecf12fbaa2510aa3b23504d11496985ea8e05b6c35bb68a5a6a4170e395a152fd1938f9c59a45b46f10ee959913fb0590;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc9fef4fcc402ccb1fc40dbe6db76e6432a13e2c6771364f4e50b28d1e12313ebb31a9a8a5ce798fddd30ccedc1f7de09539d18c3012d345bcd1ce7eee2b7c6e9d08beeaec7499f3a2014537fe612e16f24b2124a0082690cf4f4780d763c98758e0a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8b2902ec4488cc574a36bceeac8326fdb36db6b192c9eb52686387c941f43cebb9385ba56c7440a4c4e927bfe550617b3430e5b0cac01b71f43abd64f964a93447e813390f33f7d0421274a0f99559e5a206743041a0772b2efcd0eb8d2d8534e851;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbe6c8c5129dc80f679f1fd3bc322f0ea65666ed565ada8ab7f44602a6d4460e36db045abcc54943ad630aa152d4dadec9601ca40cd6768ed07f14eecd0750b671364566d385ac6138672fb90dc7c5e109b37b69bd15fc9d633188b24481f0ec449bf;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6665ea9507fd4c1766529b43e6b20c637f86b742a9bc82ccf7a3f3b7857433608081e8b3b798ff27282b230653278332b2d3473dca4028e8607d86a3dd1a4bec616313c9a6d61910dc8d76a8d075485ca27a2a91dc4f892ac4dafb0348d0711aa7ae;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf65a83deb68988f722a7bec607dda351be4741f1556cae4a8e28d4d91727ae8cd16fc3cbc8a3df73f4451fc19fa43dcceb805c7cad535320119bc3e36baea76adaf469237210394a26984d06290b99520d7a2d2830df8142bd8ec905bcf92655a120;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha910626bd507f8f549fb7514677758ec12e0e4130cef2030457654858fde672b36174fadd5157e865a55ab9a5026d618ff045a810ad6f5d7b72308df4134d756c1e931a4f819495f3ca21c8fb038e981c70e1c15c6a0e73f1d00453e096a903fa962;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h30d4e616cc3633d21e477162652f708c7f6e599a857f1194b2ad6044ce2c5e4dd014c34789cd21634e12c5f373d87b65d3ea7281002d8e746a39bc884873ea116dc99e41893325c2206a45f5462e1195320c58573764af3b3efa11f082d436d519bd;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h20a42af633a3c19903d82626174821236b4233c88b1c89c0512bb9d4e684a32f3d3b907afa0c01f59c13dd6e7766ede6869655bebee8ca59e3360ccdf439657f02e70de4d72fe802df5670024a15e368d66638b975fb0a3c8be4600e36d614a195c3;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h23053633cd41d43f00b9463c4ffd889f25862833a4fb984710dd45503fe4ec797aedd23c82014e41805abfd52243069db524b2a0c7ce132c7f3ca8db611282cdb4c7d51c78a6dd8427f1c8431f6fb2047a4b0b4203d3e2db8b74981f089352bca6b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc66ce309a7684aea8f7af735db8816290eb7bfb216cb4996cc791307491a243bff883cc4e90029bbce7c781ee6cba5d86b62715f0e649f7890bbacb7cb15a31e7b7c0c0c0427ab6d17ff60bcd2f5189933652fa45315a3bd702e0e87508aa250360b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h73cd322e96bf71efce01760dbc00e86327a8cf8190b2cd7939b524227ac70b90b9a140f127e74893ffb67f856df243c06a52bad39d7424d0f9526ead2ccd473c0c8ec54f8779bb905f8f7eabc30a058bd1ebb65e0f5cee48de0fde363818e8c9a99b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he3cb7c341d58b6071ff462f18651bac0bb3d7d74d6ee9da59b177b1097157b7a2a2ccb3cd7d62bec13ae3c3a2196651731b1b5375acfc520ed1f9a9c0cdd0ba0c5d5156a3236c565a7a226376e592a00664d753bf20384710205ee6ad06278d98227;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h550659e78cd62d87da4d9003a84b79e050fb26471819696e4e7f173a77a7edb0896a05280628bff5398b042dd64561e9ef3ba9db81d49e4f67d9d087278dc1361316ab549d01975d61169d78c5f49c36ab85db78f707820d1e3e7f2356548033dc1b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h12e47c294a2ad8e6b03f76072f8fe71bc8f60d1c5f4f01ccc49ac5a3f008a3db41de6c7bc06462fdbb64082eac28850669b99a27dd8097d5faf09eeda31be67fe277f2365d9a14965ae602a6d2358ecd262b2f38bfc54d6ec4be86908ef316255ecb;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb6b1d2a542c13ad78540c42f3bfe640756fcd33037204a24183a5304ed9b71362b2914fbb654dded375eb5010916ae06d30ad3ce6095570bbc621928c8ade5c1ce52d0475e521d7ce9e6f9f98712eab5b184ac4d039f56be4d1f5fd68851c1d1981;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7be010a22b6d1b42bf61c2cfc2c17ffac429261b665feb3d6b2abc1bc06c555c7589832718134cb2bfe90ee93aeaaa8e0ff73dbecfbb99121770384168b4c54b3f7436755e6ba227c9cf29b1d8cf8945cab933466e0644d2a3d144b375a00acd125e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha3d793a13a9d997c063e6c1c3ba34bf6bcdba8c254c9a4eb88bf7c8a1b38b462fed74df5d426518522a56207b660c66ab139786af0563419abb73e52f59842cbc2f9f285182a07503403aace7d1dca882693c5e8e6039aabe914d067509606c93a72;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he1e4fb1b781e53883d1b5d2f8b206afae881aadb1e666e7b04f6e75b0e007b3dd99788fea7bac77f559978d19fd798f1b3094813659b02cf3cd637365b43001bf2b9d64db0304cb1e05bd08151a096de4718f76a07894182c267e9e5374e43f37954;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h54653dcebca34c90383bc0f70c800fea6fae1879df28f218395b073e4eb43ad00320ac44b8b8407637dc3bcb0891362f5568c8ddb70bc49c1586a1098d8f7536e0ee99d080662ee96f4f9b8fd1d90602860b17f2683ca28c8a52926b9fbbe72677df;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf924526db870217e9b13f601955104787b91ab16164d605270825fb70c1fb5ff8472651b0bcb3bff15f413b7fd4819999e08558df615b5cfadc7f73ea34f0b487c3df376035056f5c66df9e3bced45f249159c5b9fd07573fde040f62b3e163d49db;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h47743538c482c118898559f8fd81cba61c01fef547dd47523ca6ab5d653bcacba78932d2f4a9f3fc5b939cd6bb84496cf774fcda6d974d58aff086ef27eb6389ca63624374aed968ee419d90fcbb76da4b858b4048f4b1d5a74a193be6d4a399913d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb9b84c8ef044553a27c2acc9fa69d323290a5a90669c11353bdd307717f303108993d3fd96a8eb892c0df790213a837276cae5c8c471d9fa04b86f96957d46122e63bac96d340fe5c52daeca6d97341e7abcd6d8dcd0f217d69bc2711013b64a50be;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd15bc87c0ff38096e43e2edc60716a3bcb7ee84b84f529ba09d17e969ea51f57d9497fe75622824d8e7018ef0235326958492cb23290d738325af13c9aa214379e952d89c1f7cfc283e440b1377d6e63aa1bdd3f5dfc79f106c0ac5b66f9bf5d66dc;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h385cc4060135f6acffe63bce614ae270e6555454608c718c4298fad53f5e2a4794161fd875ff266f52278ac6babc92615b2ba428133040dd95ae390ea45ed90a22b02e539e0a8cbb8776afadadfe54e481dcae02a363b7e78fe7f8cd60f55e6c23f3;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2fc794f9b208d0e6c7749f6b6aa5e750275d66e33bfc0ed3e6d88c41ac08e676af507acac9e0a9ce8951ece156567fa2b8f98a06e7e1f406e5461b9caa87a8e8f486329bf9a7d6ee2955a82f6812f82388adab1ca98e9002af68b8a7cd7f6f371f51;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9ca0f19760801ecc11f7e616edddb799de2e8280d723079cc71dac1a14cb8141f585765432b90b8808ec509520972afba6628c8374f6218312298d527f71d0facbbee4e84b4c632198e1b21a522ca31b55307dce2c5d12372b89e50ef317cfb42bef;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h55b97eaf5b4993558a25991b1a5fd9d3f18997b1eef5a4c199a1fca84318130f8d2b524ab5c3c581e50ae33934d0979c5bb0f07420febae4a1f81fbf481792fb9365ef483067e893bb2d812d2e5cc46fc7e14f7b748cd68b8acaab4f0fab7fea58ff;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9c87945f3c12174efbc15158347f44e501a90bac0701b604ba7cc295ed561904d929a151464e056b43a79e9f52895c94d11b168f6f2e9998c91b461624442159021e0ffbd20d5d9f4f202dc614409c8357cac89f4ea51d8415c731a97932f650871b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hccb136a485bad30f7b3742109abb41f686bcf9db1683776db6f19e46fe8dd7c716afc9db520403386eb97bf21b3a28d3df11ce7dc98a26f2e713896bf7fac66756870eafc9d68f81535160002883d833fc3abc35b44064b40823f9b636965a934a5b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h29ec5c949244736526fc8cee5c7e09fc29276052724b06ad627d06b6419b5dfb82c069fa7a5605a6f4192262eedbf247d8af9f930d8991fec10f9f0336f88477f357526dc5130ecc9c9baacbd84ac414fcdb2605870f4916122d0e4b64677be1145c;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9dee2840bd8e4698d583fd1488f068efe877973d4978a7f2da678106ba1bbf09e9e1caba9391512f99dc0417a7ec86778f57a499366afe74b1cf8c15c58a75da81bdfb9457723e4df294639831499568b035b5a1d0908a56475de08f7bfce5212fc2;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb82b9c542ded51957288a16d8fd745a8196df068491c2539d078c462fbe0a261937664ad4b4cd40edad6e352eeb99ed25101b1a13b9da2ea1426ddb3800672511e7cfe06f74747e41537e48758e15a6e14f0312aee0a24ca22688c9b98f696b833cd;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h422a196158344f5932d4f63e8ada5a3c12f619074a98fa02a05956b7bd04625b1674c07445b3bc2ff632128a9e029cf407f126376a8298864789271da9ea38a1e5ec455944516306c1e7e1db71b75c5f8df20d7a44a71136f38afdccaf791d60b0d3;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbdc1ea454328e9751a94bfd15fa9fb3ea45e91e66200ad2945d14f15c99f69f118c5fdf3ab8caf95174e3f1f07b4dd5e1fe43eb554e13d30b0e78b374b8cb200aa357d8224aaac55f8a9c989f5801fbe71a9a80c87c7bcf3873ee2a2fb40631d9c60;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h49c0ac844b92f01ea0f817b33a09e920c1355ee383d48a8beb8593ddd0a38f68d0b2f4191863415a31f3cd9fc64bede479739c3e2eb71a2878c0052f526c5eadb74fd4eb87ec6f841999eedb89c7544d92659e83347a45b9d5f6a884446fa03abe30;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5a4fc4207e7824526a4ec5d74d225f8f67893df950219b9ca84af1c98e247359c96a49ac7f83c1da69c238960609bd3b9a15615c387c83073267e21bef54587ee08483ef37e1e3ffcd9d13676d64e90ef1734cea957480aee74bf4a9b0f04ed0d7a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd61a233f69328dc402a75d65c8338f1fa9b527f2c8d3e477b160d6f6761bcd114ee71496fa4111a56cd7a2d4b7fe312a3f6521fa512b223ec17653003ab62565eea27148a304a04b02a8daaa80eca0b0cf5465a33ef7458b1a3db39e0eb0cd88e1f9;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h70b14767597382c302bb333a04df800cf03a42c7603711feb779cf4064dbeabe114a8b04d10324ac806803865747aa2be2a33cca22f0bceedd96a11d29b8068f2430beaf8e752811e5cfb633cfbd7c5123102a5fbcc3231c447307d33e44331fb126;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hecf1c503c07b7ee482eebfc26e007f57438dd6655b7963b70bfb48c9e5b1df5535395209d2cb79724c713cfdfcef38cef2ab4ac77811640741649135569bebb1e60573fadddd60e561244a4578887ad91ce49054ea1e1e860302b44cd202fe42cbb0;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5b0b9d3e340df6ab8841c4dd5145319669366ae495c5acbf57405a6af384abef63e1ec63e3d99d234847ade206ae7582f8179575c3777df4984657d15bc10710a4c286204846bdb791eab4b1cdf21392b841de9df5b949c1c1f705d0d39cebdb0e2c;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hacd75d441c3437dbde90e10bb541a6b955ef60efcb9e6c9a1926bd3d46d63c87d29dc29156a022fe96a018eadbcfed472c82bb5a16ca5ac0077ee34682302f454c0598f8b33983616f6c18d82f51e1a22dc9e82a2ba0648bc55e2e77a3239d6eea36;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5969d39813f333cdd97bed68e53a3577a52b781069958fde5f52fd47dab9779d0750848b4d7169327ed79543ef0f4edfe3906085c97d1a55040a6c69be4a9e17e55ec970fb313c1c0cef95bc1b7887f9d58ddfe0da94ef9fcf701e7819cca7cd9c2;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1c68b5cacfe92650f68fdeb5bdff67694339a45136a0c5af822c8d499e4bfb38818158bf2e4b6666baf0e13cc9d7342e8201cc37f6c05c470678205f303227ad7bb84d5dae731d75d2b744c3b3d385f5dd24774a865429015943ad549f0a89345b84;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3e98373c194af53dd8e6f4c1b294f0d3c91ab79d9c083ab9bf5e86560a9ceae1ba3ab2781a7f3fda672b25ca3ef144f047f603c76e816f832b25da2864fa147a0826e5528c5fc9f970842d41f9ffa6df03847c95736431655c5af337a5efee22b26e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4d749fb289d29aa22d50853f8ea5661ace76741c67d2ae89c66d419e9c24ea3c8d83bc9868df72885669695990571b145a05549b489f34f39c480b0f1f001f58563afc925cba20c637b856422a53a6dcd1b7f9b736d7d605197300d05a3fadb3c285;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h730e42b99446bca94adc204c6d804fe914b25b0884f8a5121fcd3b330fad7de60f03d6a4e101eb0747aae301538bb579bc4cfd91e0d5a1064ef38dbdb3669b15e4ecf9f83b065cf9867deac7e0581b642affe5286554b9ca372dee1379e8367c34fe;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc95e4b3cff4e6e7a4889eba4f12ccaa4a904c1138362b48fdd6ab2ed7a2ddb4b97734f8c3e6845ff198a3d60648e7e65ce1b7891b54e3b783944489140b4f2f138d352961c009d83e0517c96e9c730b8eb967562b6ddc77ff9b639ccd5420947f658;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5f3fc47fc643380305301c03ff2097a08467db0f8b0c9825841d96167fa43aba655c45166d6c6267f107224b079a3c2d4d19c3d6cc89b5f30dbc0374ca6229d62bbd233869f0bfc84eadf81a28110de8a3439aaab3ea8ec869e86c21775332593a8c;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h173b879b62736b27953cc736a6a64b169a61c25e0be11dc2bc8c0c884d8ce3935e18b1cbee206e71640454fcbb7df54635fadf80c00f928bd050797ff162a0d8fa4a441af137fea5bdddf6743f0cf6497df42d6c1bf34cdfd5629670c63c3d2eeba1;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6adda0e6d265abc5a6034fddf94dec367a81eeee4d6571fe2ccbb10e980bce76f6223d882ff1450e593a24c47e73035c032cd62cf001f346f4ea95969ee863fa7a90927d0f42ca130335647fc2bccdba896b80eef31b6c64701281921fb6d510baf6;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hed3915055a389d0e6aca94214b176e4de4c40e794dcf05c73e142bdb9c62d3c9d6d24712ab901e8d127103dbf94a32cbf9bb85fe8614fd14e17a4b829b6b29cc5da0b501f3df31aa2840f2cbdf48d20ac9f4800b04a2a7a1aee4063ed1974de1622e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5bd0a5d234176b5237e031359adc39f695507460eefcc5ad5c89208ea8cf4a28a5f83ee2c465ee9afb7ec64954a61910b109363bd378113fcc37de585c345bd2835ba18c82e6b5028a09cf54cb3022eae4b4c5e7f2dd963cd94a1c48575c58d4ebf8;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h940933dcd9b2f6b1120544142f1c1ee167fdd6539a96b75f0cf9568704b2764a2561552195185aeefd8b192d08f0e243ad0836aa6a67b9da1777363dad41da7f46471e90b2f74014b8a01f7c75563fa29ba0337b48866db91a3cba3daddcc3a66d59;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7f07562b9bcb09aeae5b13b9c36e931cbe8ef58d6b85e234f8fe133ad4f1dd78ad4285e0a171ed0ca1b0660a66fab92b00b4369fb928ab3a23cfbd73e2df68e285d5e46c5501233bab7ab34af795484feb16d8a90b8a7716f4278445a355eb709599;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd3f11e0129066377e162b0612d5ffe68b8cab0324bd1df5e2ce14e15382b764feb6e7ddc4ad37b3d7138613270c822c5886e70633f7e4749b7e6b41986fdf2e0f1d174aa73d1a7b8eade7845643b3eddf3349d476341777d821f0527e8e06e98ab22;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdf54c14c9103fec9e41bdac066848fb71e979068239daef77ca7c8e347b471cd6c5ff214165930869c8a898942e6ed4a649ffd4f7aafbde020cf1d776c995f6a87b530adc55c54c1ebb76f465a40f7667898f26b4d9dbc454b557e98eded71e73faa;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1c094ac0555441b9f67518e4a23965d182cef56357d05d4d49fe7cae1e4c0d3999cfd9039876176370819321957c7688058db2a7022f676f72e6dbed2890a57c08d8ea747d2c4319ce123e227195162199278f53855934883c02c7a0d732fe20aa2a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf58e996308638847aa330121845c4eae44d6e94bf0179c81000275b4d8da4b4d6009ab21cc87d977fb5b965085be6f1924c8a751170d3a9a4b8ed01f028091789823a6b60b86dcfc704b9830ba47f787f8b0843b5e1f235772c4ae222dd738d173a5;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he1a26f41fefbd6a9ff72b5ec00a0b9319d4c2dad53cd0c8757a8bb5ba5b9e65c18adf1cc862faa2fcf58bb4857ea56aecdf5f923f2fb5a34bf8a464ed0be281a1707aa551bd2c0ed88c6d2dc66d1aed53948c348832a34c822695c1b425686a3b8b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha69144324c576776a5b690f5453c537342159fee9f909ff3a517bab262cd800782c505993e643f2ed65399980a7b5a75fe24d998865c3b7c1b75a16bfaa035d2fe867432af804ea755d46b3c00f17c9e47cf12563a2aee76c019b14f5d08b62cf9e3;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h68012c93a28c9a6fed0d372a428af885d9304bbc67fe1cf7ec149756dc1d77fa80415b040f55abb9c6b8db694fe9235cb83a2539110508ba21e09325fb784e82f0f938fcabf15ed18187cc09f85e09489490d1d48ec3b4633329c3520f9096e1ca02;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3dce96f7ae6d6099458fbc8f8d487ba2167a3383c5c3a768cf8fcab3da0cac35d351ce7fd991c260f5c0a5f1032cc3936db09bbaae01842d15021177f17a5e2ecd6b53ef417fbd3417e2a82295b738f2a0b52acfa9fd57b7143ec1e4ba3bdfd81d05;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5b17578036391aeb4cae0e4218c3d7d5ec8477249ea057d846adcfa80c1afd9a288f27d999d41b0de94378769e89bf2abb45d2c5cc98e0fc346266e079cf631173cc43e582df8e29ad3c660ca6776fd016dd86f635d4ada2888790de2a7709afd0ae;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h10b63b0c81b733f9c99e9edd825ec91e6b2a24d73c106abd6f47d19eccdb1591e3dfb4fbe0075506a89614f8f7487abc1bfd46870591d09e8dc761c235d31e0b5b84d2162618218b5de323e30a15a5fbf9a556de97dbc5f9654be76e16e831d2a9ad;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6f3758e5cd64c54a5d22b4959dac1f0641f5ce3a17d4ea0ffc73260c89634bcc9cd6289aabe7a4f21ed5b28ed49fdb33ba53615ca5d59c9358b724d05fcffbf7449194d242ededf5249fb895222e37aaabddc6bb5fa881ce2230b93bbba81d8dedc8;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6222b8fafc37242173da0f7881cbc6604b28601097130dc62613827677846e4528d692ffce004bb9655364d6395e9637d445a57a4c4ba6426fa99a7bb522fbe203b2e13861e7349079eb5c26d51efa79ce394eb697e2e335a77a131482107b49ca9e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha2a7373dca7b20b65d4e1db35a52dfa8b8185587d8e794e314e30431be673fffe76a712cc985e6d42fd07174e177674f71976fa66ea13ed2d24b779cdc4f735ebe964d7e3c7a327e68456f1546262a78101b1bf7c603b943aff5f1069eaf46a982b4;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1ff9ccd8655a1026b04d0f9fa8bcc589b64f4edfb2f1c2305e1a4d35abfb4730299c778542eca6f756d4411d6f2181f2c8242a1bfbef9517535084171f5cb4c1343d793cbcb782d25f1aa1346fe15c79cb865bafdbc6023ec6bb79351bafb2c8a866;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9d2ca16af0a6270c58ff790e60d766b187c66c4230853991a347b2676062bd90af188b0c4197ebbc63a5f36083d9f45f7179cc4e1bff42b4cac85d8966c5d68e93a3e974d76df042689565e9690898c6e0e7c77df88912847e8841687585b060258d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h744e06cfade74717ebfd974ef3869dbbe8d13cd16b74524565e7d71415d3ebe65d97ba545e32968d78ee3d75ffa92224142f80ad43bc09571559cbe3a1d4034bae84967ae085c2beb8468ceead4359cad28e8143d23f2fe7194d99c7f052a4977af3;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h32d79331937825ad9be53e9be11c05a443c6aa34da43d714af31f6378e095d198542a50b30a59b657d8f1e5e59ce80f8de8a1e4e4661a544a5f6116eb26e031f5d24d34c8b18bbf43022b769741ff71817820341e76cb2b2055004b03cf90c7fba6b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he528d41a262c2123cd804b50853fcc35b16a654376fb77699b22d7b6519f5c720d85b7a7ceb388427f7f7ebf60af46cbc481334ffe3587727b8128d6718d49b014e3e264b087c65d2e6bc0e85dcb780ad4907f4868eab744aabb33dd38fecbdd2975;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7135d404c9d5df38378374e3befdfca196f6ba60feba0b0f499426a6c1e60d35ad5b3434c7e522171b235371b2c3d0a8467b154b25f4133d596a5032bde66bf81f21949d129889ccfc922c95d1a7aaa454641962792be21cabc4a5316ef5c3cc6a3b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbf38d584424c2e635d08abc0cc81f54c7ffc1c3691d8693de34910f69cf8bcc9f089fa049208471c50d5d43d2917e616296d9fb16e7c6cbcdde3ef802a1258961deed68670cc0ea63315413c19732c22921d0e07ab3f814cdd9fb2363702ce5114a8;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hff6527f6c78ac03df1a5d86fbfb82211d1e11b8b79d7d42ada4d890fc4caa4b98c0e95c67fd883acc5516f86ac71129344fcdd56f7b9f3936ecfb1bf24e005383bb0beb8fa50c7c0e340cba804df793990e51aabe483dc848078401d8202b694d489;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h98977c400928d6414115f35e2306805404bbb357bb675231ef6c9bc61fcb8bfe26e43239fbcf573c9803d7074af273ee9f3c20a410317fe24c0e705aadb11719ffd7779699760eed07bce4c44a4cd2694d5981fe2ab9b07a5f32b13c341eaefbf129;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1dcfa6ba482f6a8e3a58f9659debda0a721ec0374c7fb820879595b2619c3e97eb5d89f2ce25ec58070dc4bbd7aee2b5aaaf929940688a80e274b428650da5d0f16c94c63916474fa8bf2b785e113d7a37ae172ca37bbde9db357f4c7c6cfae06574;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h339d75b0fc6fa3215596dc107f677fb30f158ff6c186f671a3d0187c2d584422eef5d8aed96d6e5e406e038f112a537b623a8c3634504e1ac1cdc9fde8bcb644cb578d0508e5e11fd130dc5659604456275c64491eb2613e2b9911b4084b93c78ff5;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h723f48494c49aa73a6c1e1e6626b7270f78b1a8d5d484a6b713ea1ba20d9e2ca65a00d07687c9cb02d82490d25f31b6660e5aca34735e246e86e9e530257187fd96de361632ddd925f80b8226486d7fcd7c68cf40c95cdf413e5eab733d1606727bf;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc71b3c5ca587322bf3043292f4e19fb3ebef239a565cfb32d8c8907498ce5be294b2407e4c227550d268a60229e4bc93469c4c3db181162462264dc5f7693e3ee291abc58f2d999d4d97cba0aec0ede6317df7732f936d461676438a41c7ec00386c;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdeded916d46ddb09d659f62b740b4593a96b59f7c993a75e106db58be4260b521292d17de6e7b1d523777ec485818b166ea2989aaf8f8f01f4256da265be7b2bc24fe8a90dc0e52d223ec84f8552551b0793365dba07c3705d9d0fa741ee36fcc864;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h95397719c08d4608278a5dae3439dec7fb9ecd5642acc3a3535c09702fd398c1fdb9436934614f5f8be4061eb458f8b2db0a8adb42f6706a85f5467ca62e80a352981c4f6b12f4b9c1a263caaa9df57bab5f3bf83b25232987a2478e9ae9d69ee109;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4f7a53f426dbfce181458b46c78319412eb06656cb6e4dae0ffe6b45ea3fa7bd0e1689510a396b6e18cff4127f419ab0514458923494faec8fef61b72d3439394f49947963c03d3bd82f91364d7f721f1319948d99fc9fdb8c8e53d53d3e7cc75da3;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h62b34714a61b4b0c9874eaf477d84e7453adf4326542dc6db15f5ae9176a0c5fae74ced8622297b2448f4bc898fef3d3460c5e2117ee8f01dcd0044ffa17bc66e9b70d95a653ea567ae29ce41e2ab310533506312cb8d977128e6a58de2427ab724d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h880f9614c485589241320d111a4aba79fac16da4196653b930bd313b01600a9f6ab9060b386f6b0e041e1e6759c907a13b06470ad0752d589f5e2a93f7383785e5e3c2182b4679a26c787d5d8cca399680173b7de85774c68a2097ee3b280a95be0a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha166cf2795d45646991bac483749b3ee73589cf27648b678144dbb99da8b3fdf3faf38ab82a84dcb3b4689fa9485b362fb1d772539de2f4260288ea69c41a7657fb64b055a32b71660abe5d1e8b19bc6e276009542fdc2c804dcd2407709ab12b6bd;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd51706b29af7954d2c23cb889b3bd033fc35aa21734b06c830f394689bef5f867ee987e5ac595ed05c64221b0b3a9230522707ec4b85089149521cb056e02fdd1de67af18bc298817d380a006baa3571ba47bc6d21f69a753903dfe5cb08a73db852;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hebcfcf74c70740ad55baf3aeaecf900fc8ab4e6420b757d0969d85904c02c4c19e4c22ebf56b50385af9f9bf60abfbfe3fe51b9f0b6bad2cc3ccc76a4a19c57381bbecfc9cf47e4fc0dd4659598056c69c0f20a45bb190c2e777d2fefac0cce3d863;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb4808ccd933938f8519291ec0af88987636635842a7b95ec36cd6254200000e95f5c87f509b15f6206c8b6de8587426bd5a735359661b814ebbf1526ee7b0131a046deb60e11fdb255caf439cdaf20ee43b280904ea05530b68691cb73bd7f93c14c;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc72e446ae2c261bb1ae1a071d72e57e95237e8a875900f99791e31303b0566991401d308124aff732e941f08937b2f4b341891020d269dfb60b71339069608d94339a615a5885b00f12213d28cbf001001e7d636720a8c58766c5adc90540710a55;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he94a7cd070c037f6e804d4884d77c671b8adf41e6f58df1831bcc80659f90450d4fb371c87d0df17bf47e54cbd58035b4992944cbb84699045d8f45e12911cbe2aa4c95d4d19b7c439beb3ebb86b2ae620800367b86c7a5c96bfaf8802596cf9be79;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb6ed1e0eae040290d6061b23f2fc3b669b6b773eb9bc24ccc6746161e6abbb2f02f701393ca0e8cc0e3998b59374564cbe80fefe9e6f5e2dd46cc5a2b2a775ee870aa4ee3e6e340ee98d3a12dec94125b746d9ec868f57a6f60e315564f3ae55973a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h57ff1c993861ba0b75a55c1a37d1a210ed48365082a873bc8820e84af48cde16d941fdfa5c29f7c787b07b5691f7a431a57bb1fc3cab349504c778a1528b7718f46cbd3e4c8ef3e8b1aac1d608a440fcff5bce72648dd31d3970926d9313baf2458d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7f8a6fb66ddfa60186994982bf2b3ddc971a0e832bef16deb05548635e3c63d35f9091642d9a81848cffcfd875ae24ead42db2a0584407d38a005196c6c72cb1c155b2f4a67a66acd004de962734e69d25a630eaa2b2e6ee39a0ea8c5efcc593e0c2;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'haa5a342550f3db002bf9f119deb5fdbb4988987a875e25ceecacc6547291d40ee3aa4f274c5f71f11e22fcdf914aba505f988ce9519dc73792c450857d425bb92b2d7628f06fa5af0c08bdbcf857152e638276a1e135ce0fb8cbf4bae78b0730df62;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h564aa109364644e9fc54111cdfd6d487938e38d001e3daf588a1d7bd33c05dfcf553ecfc473783f03ff490c323b3d4f85d79d85a3a8147f45f65703725dc35090fbfb939cce80e21d5713a0077805e7cbfb075876c84bb01ec734933065899183b62;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb89ef9e152916773f0362722825a6f379aa5a378fb306422973c8eb2f04620818684b2a89e28647c394d3758cd87f0897f9f1cb0707fd84139ef1c2c07a41e824bf9ba4d89b3119cbb72b35de39073b3b45ef664754f753d01bb65b11e780e04bbe3;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7e922d183063b0d12b6533a76a062e0c7d8b5af795894f169ca20aea4365c599b0095bcb2f89ad9e9f6a61da6ff7818e8fcefca1323b166826efb76524a4a3c6b8fda5badb705e0d5c1f0ade08e800894c88feceb8620d907ae5e69bc92fcc8ac49b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5ff6a09f315a97f510915a43fd2879e690f966e7bd17512d7e1619674ca53221ba118c7fc537183cb64be0e267664ec23c52ccbf06a85be4b1fc84afd222c135668bf8c7595bfdb7b45ba289476c48ad9b8276e15e62db1ca321a4875766e7f9823a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hea9efa3436d11bd4aa665f8b1f2873e49947e24055acf8c445cf1bb78afa48802ef23b849fe4da04af8b0b805bb9705507dddc62638a9b4e6fa737334a53dd46f4529a3efc21195437a02e0834903e35a0aba39b6371dd872509673b406bf6bdc66a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hebde2154cc43be63ceee3e3e2379a5db333ca11dfc62c400d762bba2e0f8f8468f58877ecec026d06f7f91fe7f0e0b0d9d43b2af75f02ce89501763953749dde81f095e3f3c9042a764674e7b7846d6dda7318e6caa1268b2b33d444026df61aafa0;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb4193185eb920fcde1d6eb39a92321afd01a04fc207f682663783869ebbfc4d832201e987b9ddcc02c4814031c3b5e2d85a27834f4aa39a60d7d5604ffb6107ac258a885688efb6fe712583f8777f5c5392466907757fd7eb8ee7f4dc886b1e14fde;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3e4bbd43735554adb12556a859f735d278b537f9d77e0818f13328fd711b04b43ec2f6f5b4107167b99a03411748a718c2f8bcfa4d54b0b495d6f22cd120077bfc1599164a08f89115daf3919a15f0861b3240570c40f87e6a6830e69415c911fdc0;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h33afa60f56ac390c702731244f09b934d0204180ed72cd1a37abc9dc8e3220d86b6d1e425bc09ad6b6665387b8dec2ecab43b5c561a1135d21230b1bc5e5e3cc03831d71b29b903e1558ba6517e58062924e3c632e5637f71c27f1ac036a31e348a2;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h814166b0a07b968248013ec34e9a92e92981a29a9d8e20e254333c6f29a4997ea91827175025749e0db1c6b5e815d2bb72a35f8bd444594bd7eff63fa268b2bdc76a64e2598208228074fe6493f3cb41ad6431df1d19974250c5ac4e4963c5e93655;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9ddc380253add9e921b42dc65a71022c8051c01fbdce62b09275e730e606ceb76f9e9de48f09fcd953a50dbfb90e33f81355f4f8931e4ea04afa47e25d40b9c694a05180bcf365e7efa3e55155e7b79f48666e90215ba7570a03ae2c3a279b4126c3;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7db37b9d713977261e9b151140ecfe6f5ca55d39a86254c57c62240cfa79f370844797f7441072fa588ec084618209e8df107064ef6066848270de7811828d1d983fe78fcd07fd31894e1370445a7a66dc718a10f537f28caad7ec1e10db22f8e462;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3338bf9c7333ca60f130839f974c6cd507da879c8360c5ba78e0ac1a5aa178ade1b60df7ab3fa47f8b4fc4ac01ab39c4505f1a0ef2a1840c32240661cf72157b2779d0b9dbf774f03c711b2f09bd3c894e7bef5b2add5950bb3ed92a692880136214;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6d2dabdbf907727948c35d8c26ff2f8f9e526e7612b6584bfa34408095dde9036e352beb8ed92545ae68792af422894698acc3af71465cde088e1f829db14c7af74bbe07f38a6ecf00fc4acbe50e8ca8797f6f7329d51a17d74759380d9787def4e3;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3f4b4de20df3a3190f4cf7f32ce4af211ba7444bc321ae430bbffd024eda7bdbc595548a80bd4ab321940fff5c0eff6975eb49f8600a1664527fa3044605f97e5262c9077b50afa1fb6c54898c48907d88a1a14440a742f704b8d524e05b5aa3f87f;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h553e31e7479edcde034ab0e4de7a76ee2521dd43142bc6e9c1ebfe0f09bd213297fcad9fc9dac717603e73b48dd5698fdcacc53226083e816b97388424a771a51e0ed09761470853169242df8e433aa51fcafe7eea5403b60d90e08e8c6493ae4e26;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd2bc56053ceb460f23745c009d2b3f6aaa0b820b256f71ac88ff581cddc5fc97b8c86e5c54de65477a7f72f8c6161307eff812c41ae82a20addea3005f2b152e042fd12179a4903659977557cd1d06c2f91667e444c015f3aed08bc588dc78539c94;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he7aab0eeabce0197bcb263f690c58a74d1354a597062e9155ecf64eb94ac480de0a8f192970772c7c5fe5581ea82f1883cecc798b0ee6e129aefec358ee03e220a78fe524da267121b5f3c4460818ac0decafce82510f7ab713dcf1f8ca0e5cbee71;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h84769217b0978512d213311d5792d213d6a195aa2a4567ffa537d3db6afed4ca66f3c4fa38074161e838bd59e6cdfca73e75675efd12f072391eeb7eff0abb797517dc39d929150227b6ffc54ed90083c33b88ee5cc129e51fb3db5ea62126874b68;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5cde786bef4f374a9684edfbdb38a4e4102ca499535ed1ac96d164ee6b1804d6469831dc7651360fce41d7996c90d37ce3300bcb664ef0e99338f59a68adca8a2575462c8e5e073162def5da474bad873db1b2f84065133e4ddd5a3e8556756a15eb;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd5db0b130af094978a23844282c7717e7592415e52dfc939a048240e07948e18f60b19d43d7da24866b18562d5cf5dbf551246cf32639a26d96050446c28f722d19a41dc7873a0248aaf6ac003d84191f1d4b378c93b61b1f85e06954409ec13cb8f;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9b5bbcda02f85bdbe67a0f451f0866a92a1dd93719bcb2e04194ecc024f4561c03fb0eb29a6251c47ffd1bb850369efcdea35cf3f62a29cce0bddcef046ad788451dc441ee5d75f6ef31e7d57ff249f07558ad2701078a76620d2ce9ee44e9d7704f;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h74a8cd32ce8b98de89f9d20197c130bdf7f4e2b2dea8b442b511dc304ee3a85b5f5034f9d77077addf943e18cfd79f65da5d0e9cc050af23ff6e48f9eeb90b0a7001e15ee054d55ebfdc416e751c39169e8af3f0439e9467cf4a9948709dcabf552c;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5ae991ea9628a1c8b4ed044b1557b1c7996d28d4c728afc3ef86dc7d6ea50557bc72c5ad89e315796bc5b5470d35897e373c6e87337de2c845ec0ec69f074aca855e18287d9e16e77e71fe3b3791e2844c8d06999e22bb586dba86bf5b18b7fcd7c0;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc42689f113b8984b95555f70109ee8c551e668471d4ab8119c256200f571e971e7b291475f46687c41badb7bfc6a148c7aafa7b2a86605cca129f11a02eed5ab99e49ca9c8cc8f6cc8826e7864244565f70b681f6118ab55ce64424efd1ee0378470;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he622b0563943a03a7486d2a942c649ae3d02beffe0bdb68215401abaf17758ee44a78fdc1d501e704af68e9556a3b269b4c8a403614623c34ca05f1d66ef523d495f26c2b1d1c577604b0f15f20aa7fbf2c8af956f923c72f7c27a5cb8c7679e4ce3;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6ee4739f4dd815e4f5382f30d01643819857209e1d747baa1c5ab24316dc6a0910e13ce3a49a87c63dce3bba161bb175ce907476a6b5e7c8d4986387fa9d69aee44b789c5347aca4951344197a20b4aeead419beb02fb99ed07277f70d1cca38b402;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1988299ec247ce8cddd10eadfa28f50ddd7b7222ec4b55f1cfc73b4c7ce3e417b0402bc273d1456f66804ad76eeb26fbe298008d258f918a0577e7af115f57f659a8bc54a1126b59dcfce07e49aa5ac9eb1f47ba57f78a5f5db3ddd7b5551ada2227;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he2cfb37dca297b41dc14de0c310646eaa6aebb111a2a782d9e6155df2c94fb98680d3587f67805165129704db7d21c88632d4171688f125658df4ef115ff0e203578b9601297417134a4bec9e4317faa6710da5bb9ab23f2a069ff7a8cb388ac53bd;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5d86ad23f01d8b980af95fba69dc50b64b453e3e06497edcf3d388f94673e703a1c0ab7be5e6acdb2aa705468fbff20f0629d40c60070f1c2884c01a9021c745992e4b0c2d38ccc3a7c6c65da070a5bfac764bfba3ac6dff11c9e5e03e05d3c3db7;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf80ba7c1cff2ac49819705c2c9379c839b56aa8217ac8bd4a031cc981eb2d5e07e353f29d52bdb188f0e1f425547f01a71106571b928de33cfa1eebe3670c724ba1aaff24ff5e88ade5d06c9fccde811a0f30b827b416dc2f6f64bcbe02b055fdff6;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd23541070368b139185c69fbc4de5539091c961e57d797333e7b0fe22420c5b36adf12876a56db2b2592af4dbd0a8bdf87b3ec0d5e0e3884048fbc7862fa0aca51b4460af912ed94572b12d55327d9f3cde46d6c8d3bcd2ed77aac03f01053e95923;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8177e1b407875141b4a13e30ae8b064f355729c95db31300923c37025862fbdfd5ff20d3bed75658a77062c5e89d72bced8fcaa802f6518a25466c19e5f3c78e14dd89ab95d715ffe28d447add83c8de57407a0ce946a8790f9ad92da3dcdcc6918b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hef58be4a96f333f2d485e18181649c67bf58db443bd8eb6ac0b2cd42bc3cc903cab889fa986e16c5de6197c469b1980e3e61e6fd1b8e6758c858a7208a59c26f8362a9fc9bd9600a3ed3f9d57eab9a367b11778f6b99794c05e401ce17c9ee4046f0;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h265f24c6234f7ba51e192972a2938fd28a78a2fc639975744d7bf8b88399ce305316082ba126593df263aaa0967c9a0022ac6cf20bfcd2b92316e66b278ddedadc04f1d6387e58ab599b8a42b487b30b41f3173c750cab6749b0c73be73184118261;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h69c1de6f557ebd8a85cd22e1c7f72c1a36a07e1b0636d7820b6a3e704e959c7c1ef0620071fa16b84573b912183d797f8880471bcf9df9aac9499722ab63b220c904b0efec390908acd97d5525c6b4d3933627ea66809b3c620050b63b4fa9305b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb4f7e35415745ce90a4778025976f4a2c2dde107b177e8c3cf384f7246ba29b67e5f6e204c09daf565a6b622f663fea6fed19e3370377db646aa82601828d9043142bf77719ed1e61ff187660b32c9e611a28ab1c097104a2d4a43951c4141e00f4a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc8fdd636111c3c437948521cb92c062b645804a520227e4888fe0933c6ad215c03b8163145de3cd7c07f1cafcbd0caae0a3915a67abdcca05c9de5b8b2e8bc30de647d552c4b8da36fbe30de627a451c71461a53d0609a8cd9be71b0fc1e774d1a5a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h529d522d4ef1aeafa1bacae7e6fb2cc344cb3b2ef0b919a1bdfb688c10b61f1c8e68833d9bdefb0ad1b171ea95d6b456098f5ac45876e6c3dd6637fec1f39ea9a20dee68bb89eb38dddf4ef534a1881bbe6d2744bb0bf8db7d48e1abae63100dcb26;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc20e26113ea0079f651788a0c515ffe4032cb0db6131c0656e46ea2842d0cc9dd610d23718e5a24eeb34ad360fef6905e078720aeaa9b8c4d2ce9f17d45570ab641df7cccecd10b646b141e22749f129c6f38903177202cab155685abeec3ae6d0ed;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h30f02e44e5dec417be9f40056eeb703abb4d6318f80cb9ca1772e3b71319a5f7e086a0c2741240890a5fb1f5cc277b37bc647b89f6af138d72aaca812e8491cf5090cd7ce1704f4a52af13d098f5d380606a1e68777fc7833f4f7a354e2406a15ed5;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4c839eda14e4f847f888987552bcadf54bee30264ae42be38165b749498d5828e8d3db99b62181567e0f33ce55c4b40cecd05bbdd9148373aa2e786b6fe87ed8efb4dd081896d15a86ba49dc55dbb979c50ecb7bd491a819f8026e2f87ef3abc0c5b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha5c4268a454cd976c3773173262e165642bb63de84a7ce037dd58074229cce445301a8c899887f505069dc34d7de95b1b9601cdbd0f9f6cd7514959ddb7756fa06b0c86e3259fc239aae705bbfba7ff921609ef8e04abd4cbe7c67829f262c246046;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h859bbee943ec502a5a6b338242b2719afecaa73308344dc50d27eabcd67bc02a9a8a8842bd75e2e738ee76094aeff7dc4c13fc242591b0d1d72021c11fc433a58c9097a91dc4174d2293a340ec5a1965ea8c7bfbec5198bffe03d29e4f50597731e6;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he2ffb8dced8c9efe76b2654711074b3636787df8a98c7fed9b56b32ac8329d59ff4942cdb6a0fcc4d09ed42f7dd2c9b21a99f5703fb8058d6da98132ecfa7ae7e90367d9ba97ceef290df888d9b4a05e6538abe07c595ea73feda93271fc9316f3aa;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb49e35c383818ac1b6a5939216bc29171f1050d65bff932b611e4b601482a37dffdfc8771ec8a0b93ac7626a72855b05fd0eb7d3d1674e7a3ba95aefd5f7a63abb72cc0c430a67c96d01e377326a6303dbcb5e74ce0ea6991b946524a9d73a53e0eb;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5aa180e8f26a872f3cf226e1a2445e170c72ba7b2b84d00697c4237de6f85ac2b9855c537daf70d10978244c63c6323b81bb35cb195cbdbf2d92f7d84bbe80ce3f13e89e7144f407571528a7942a9f7b5280417b347acd17affcfc00cbe003c64e71;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h16a78bbd4eb1c5bcaf8835d4ab7a5ba6077558df7f49262111dc144e650fc5c3fb8968b88df622b60b84ba78580b8890c8f40a2ac82be1ca5ee490a64500d9a54524fa7fd1bfaffcc6985bbc53cf3d4a29a5ee353ca0978f18edbe04f9c1c710f575;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h566519fa3e621f41ce5350af2a1b6d9f0c77dc62fe979faf8be2a091928665e267d96a65a2b1f088779cd636ad673cec94b3ec812c489d7204b43c9109479198b1cf59199cbb9d8d41eb9d2c82f9e8a842c74cbd366226b09f8ba1d11c727ad9d10d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h13d56f6ec0b071e9a04d3808d266c2f6d624ae08aa2d030721e9c424887001de4e1ea70eab26b4287ef8e668e398e229a0c3faf6cc1581216ba0e3e38d9780900afaf9ab6686c28b8451baa3b7ec6eb9746285612acfaa6c1b685d18ed40f02ff4a4;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7c752f819442caccfc5ee5a735a631aaab0172aa35ad48ada154e89b827d697539ca3e2a9c3aa9fe2ce872e05570f1e0aa6f1bb2688692d2d6e282725dce2532aeb332689daeeb3262e043a5ebf294a43cc568b7daf51972d85d3c1be132b5f64b8e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h855ec728604676f9bc680d14c93f0c1d9bee7597227e887cb9149f5f136c543407723956b34edf642fb228a2f3b1f52c5b2c61666d07f8ab167e0d972e91a2fad08558b3cba7f2fc1490bb6d55f4a4b3829c351753de817516e4b09f89f49098767d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hcbc5550ff176ec0b1c7703717655dcfdc8379d31cee912a6710e87f9ec0e5a3887cd01fda2a33096f2bd771ae23a2a55069db9e82bfa6fc972f0b75cad99c4e171cc31d367155d69ace3af55e910a9d07960ebb0547a880c8934453780a917e94b04;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4e1b251d55377987cea4f7760830686b4b4110252a762aade54ae45f6ed4ffc9bca4e51970242f4ddf8ebde84709e261cfd39cef4c500592b15e45ef199097db3bce446a4e5f4a8b9cce93b632cd77926ec231df7818b929b422cbfb3f5c4a3f9d28;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h59c86c8f78283cdc6f11352a5da870f7e7d7c2e9a94b878362c5fb70fc1988efeda35182fed648c721de4ab95e62ae6deed38699d361338fa1253cffa211b38f6841d718f6bbdf72f49c69b490d1b601cf94f433a307d858d5ece5c25d564e90f3f;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7bf76e5ad0676f4887b6a889a08e3932a24390137abfa2a68621a69883a3d75ba9ea83b92a4c4e67f0ce5cb79afc3c7c48a2f8e044d52dfded721d4cbf2b1a65e63f3570109dbfd51f2c97b7a5eb9b43ee3878f3b2cdab5baf0f1151b7e4ca15d9b1;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h48f6ab0b98d53b25224c076ea665ce7b00a4d4559ee65fa8776ad47c5af199484b283b58616dd7ae6f56c7957e358a03b8ba6c15b428c3c9051b28f20aaf5d08def70c00b399d5d9f6d51aa376ff38194a0838f20e5f1d215a0e6f1687c68e1ee6bd;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h90549f5eaeaf428bd11ab3e7ef32a3e6a7c9249a995a67382e25875fac5d30d07d4849f79a24a409e7591f0270b0d01cb200a8addc0a503add02c276383059dc6fdba130e3775dfa681c08560e3d0c1313fa8cb5ec25a1d396efbb967c885faa14d7;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6bae32add9565852511244d1587fa40b28fa2b58b3990cdb8c671fe5ecffc52f54ba041aff6b9b3893c3545dcbc7bdf6e2bbc874da8b9d3d2b2811ecea9fbe448aa85a383daf0000dcc3fabf8527d132b4774ff3e92aa0d926ddbe8699e28e07522d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfa30d8a0d1cc17820e2282e1a8cb29bcced469c7541ba832765c23148230dc61e052903b2b9bbfe2bc2c345d4b439fbcf7508e5f949392270f01e7394737a99f1e56361d2fd2e0a8c0bac73f50fab6ac56edb3352fc001f9d962fc4f73fadede3af4;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf84212279cec2a3178015887b61e52556cb26c802caf99aaf493cc3f6a9b0f72db2578da900c052d5d0f4e44fed1caf4927ea16168b67d01689cf0d9e257bce1c5c25a6a8100485df6b064736bdf5ed5d11877da19c2cb77e9007175bc5f5d4e3b2;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1564ba783442382e7a30e92196cacde6fe1840137e662719555ec7f697e39572677cc9879a43f444cbeec8b9c71092710794bc794f4dd75ea9c5cb8966d8df55941029343a7493b2b55f6adab43b44d6635fd2131e9915d73d50e777be38ae88bd87;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7e2e20f2c19a65bb285bdceb3614e6cecf78d1c1b48c8daa8b9b2b426fe3ad4af06f01e9e8cf47ff29e1f82bf70cc81f97a813b7347f0c21cd079138ded973edf347e422563194150b0a80e350150eb5d74d900d910ab1881a1096b7935b2658759e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hceeeb5419eeb8580a7668d9a5a15d7c79c32a24561ec8457e6a16257efefb43340951171fa700e0c0478427aa03a55da9921a3aaab8f036a59877fc365852aba0b99feb727520305a0157d8570c15158dc04f2ebc2121b70b19619844999aaedd2f4;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h76781761c1fa91ab42e64b55fbee5047367776b3d5b71bd32f8246bd6b79c15ed2b5c6e69f00befcfe421f414045fda2c72298fcd96bc5126bbe5781cd4997ab649867d812ea55f0600564bbcaf01a6c2fd820fbdd9a69bf62da719765e6c7297e3e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf14c75f79a1dcd21d8fc8a79d7c07d2eed03e25837bdc3c50d4db833d1e00ec90f9a5b1f45f2a695b11c7f0b18424f5f705f40226194b1dac3dbbad6cdc0b0e1d568a660ddee568cec78e2ac18ef3bcf47a0fbcb75a379f21fe6c5a874048e83d25d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h25a712ee4963b026c2c97aa9c1a281577d9a9de8cf3ddbe7ce32407e0b56fe324c02cb684d394849d21fc436590feb9a0ed68781e8399f6a0a6cc56d904a43cc222fa2e4390b70e81b01380b8071d98badd7a3b2582e4a44ef89e41b8c76f893ffd7;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1f37dd88c6ebe6df6f44bc6298ac066a8779bfb6856e438718330d993c9097c490f6f975a07b6486498649e3b1f18a2349b6e7f3cae12515071106423c1ab419835094ef887f00e7e348c5225736a15fe0fa1ea24c6e6811c2cbacddfdf39f4a6067;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h49c02aed87eae9f3555d2dcf0b9a1949e9713163ff0f0a269bad228f558b1e8bfac32f7a4786c88bef392fe5232de2f491425a7d1a3b979928ce26edb5080f22301ba7f7add91b5ef6ad44a65e40b17ed8281b5f3f192df87d99d5cfd206b025c85f;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7a543f338a43f8b24fd59cc7a6900d1a9c9d073fc6dae49a2ffa3bfdcd4022308fabe98734ef21c0acb5d207faf040c8a20c6a5f9be694119b6791c5d3441adfef885848a31ccba6c63c258155a7e2bb07295807a845f2d21a56d64b67d63e2f9237;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'heae6c9024e9f051249b616ce9416c2a7e496dd84057004cd36dab1340927c5228b064098d91f1404fb2b7cc7ff049eb680750614c58d17da9d3bab1c9118c0c32a606b2b85f5334c7c751e24fef30ce1385468ecca26e3e1957d0d764dd2fdcd830;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd4b355408bedbccc1c5328ee8915eff46557aa45fd7175f43bf2752a39822a97d4bdc3dad9687f3962c2d1cf9e69a0613daef809687c92b236f574f8215b5b356981f549f056c0c5a04f8ed0fafba334f11caf35381ba0497a60accd91a98680a9a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'haacce418bc05e62b22283fb855dfafb53355e32bff7ec22c1206610dc8f55d1743173a67f3424b68f626cb596bf02609a64909aae6087ba000829992de97af300202254d5172729ef245bef563ff0761499ca0efab92cc2b5b76b26d7b9a5f03386d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h933e30167e121bb99735adef1f0ae56d2e363abdec0223c3f5a3638d3ee735f9459b41b63d03f2ab5ae913e933153a87c17fcf0733b375491723e5a772feb8e87ec8b777be439684d00b47918c75f6017d835fcfecd17b874cd72382fb371732de40;
        #1
        $finish();
    end
endmodule
