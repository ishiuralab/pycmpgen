module testbench();
    reg [0:0] src0;
    reg [1:0] src1;
    reg [2:0] src2;
    reg [3:0] src3;
    reg [4:0] src4;
    reg [5:0] src5;
    reg [6:0] src6;
    reg [7:0] src7;
    reg [8:0] src8;
    reg [9:0] src9;
    reg [10:0] src10;
    reg [11:0] src11;
    reg [12:0] src12;
    reg [13:0] src13;
    reg [14:0] src14;
    reg [15:0] src15;
    reg [16:0] src16;
    reg [17:0] src17;
    reg [18:0] src18;
    reg [19:0] src19;
    reg [20:0] src20;
    reg [21:0] src21;
    reg [22:0] src22;
    reg [23:0] src23;
    reg [24:0] src24;
    reg [25:0] src25;
    reg [24:0] src26;
    reg [23:0] src27;
    reg [22:0] src28;
    reg [21:0] src29;
    reg [20:0] src30;
    reg [19:0] src31;
    reg [18:0] src32;
    reg [17:0] src33;
    reg [16:0] src34;
    reg [15:0] src35;
    reg [14:0] src36;
    reg [13:0] src37;
    reg [12:0] src38;
    reg [11:0] src39;
    reg [10:0] src40;
    reg [9:0] src41;
    reg [8:0] src42;
    reg [7:0] src43;
    reg [6:0] src44;
    reg [5:0] src45;
    reg [4:0] src46;
    reg [3:0] src47;
    reg [2:0] src48;
    reg [1:0] src49;
    reg [0:0] src50;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [0:0] dst26;
    wire [0:0] dst27;
    wire [0:0] dst28;
    wire [0:0] dst29;
    wire [0:0] dst30;
    wire [0:0] dst31;
    wire [0:0] dst32;
    wire [0:0] dst33;
    wire [0:0] dst34;
    wire [0:0] dst35;
    wire [0:0] dst36;
    wire [0:0] dst37;
    wire [0:0] dst38;
    wire [0:0] dst39;
    wire [0:0] dst40;
    wire [0:0] dst41;
    wire [0:0] dst42;
    wire [0:0] dst43;
    wire [0:0] dst44;
    wire [0:0] dst45;
    wire [0:0] dst46;
    wire [0:0] dst47;
    wire [0:0] dst48;
    wire [0:0] dst49;
    wire [0:0] dst50;
    wire [0:0] dst51;
    wire [0:0] dst52;
    wire [51:0] srcsum;
    wire [51:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .src31(src31),
        .src32(src32),
        .src33(src33),
        .src34(src34),
        .src35(src35),
        .src36(src36),
        .src37(src37),
        .src38(src38),
        .src39(src39),
        .src40(src40),
        .src41(src41),
        .src42(src42),
        .src43(src43),
        .src44(src44),
        .src45(src45),
        .src46(src46),
        .src47(src47),
        .src48(src48),
        .src49(src49),
        .src50(src50),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25),
        .dst26(dst26),
        .dst27(dst27),
        .dst28(dst28),
        .dst29(dst29),
        .dst30(dst30),
        .dst31(dst31),
        .dst32(dst32),
        .dst33(dst33),
        .dst34(dst34),
        .dst35(dst35),
        .dst36(dst36),
        .dst37(dst37),
        .dst38(dst38),
        .dst39(dst39),
        .dst40(dst40),
        .dst41(dst41),
        .dst42(dst42),
        .dst43(dst43),
        .dst44(dst44),
        .dst45(dst45),
        .dst46(dst46),
        .dst47(dst47),
        .dst48(dst48),
        .dst49(dst49),
        .dst50(dst50),
        .dst51(dst51),
        .dst52(dst52));
    assign srcsum = ((src0[0])<<0) + ((src1[0] + src1[1])<<1) + ((src2[0] + src2[1] + src2[2])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15] + src18[16] + src18[17] + src18[18])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13] + src19[14] + src19[15] + src19[16] + src19[17] + src19[18] + src19[19])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6] + src20[7] + src20[8] + src20[9] + src20[10] + src20[11] + src20[12] + src20[13] + src20[14] + src20[15] + src20[16] + src20[17] + src20[18] + src20[19] + src20[20])<<20) + ((src21[0] + src21[1] + src21[2] + src21[3] + src21[4] + src21[5] + src21[6] + src21[7] + src21[8] + src21[9] + src21[10] + src21[11] + src21[12] + src21[13] + src21[14] + src21[15] + src21[16] + src21[17] + src21[18] + src21[19] + src21[20] + src21[21])<<21) + ((src22[0] + src22[1] + src22[2] + src22[3] + src22[4] + src22[5] + src22[6] + src22[7] + src22[8] + src22[9] + src22[10] + src22[11] + src22[12] + src22[13] + src22[14] + src22[15] + src22[16] + src22[17] + src22[18] + src22[19] + src22[20] + src22[21] + src22[22])<<22) + ((src23[0] + src23[1] + src23[2] + src23[3] + src23[4] + src23[5] + src23[6] + src23[7] + src23[8] + src23[9] + src23[10] + src23[11] + src23[12] + src23[13] + src23[14] + src23[15] + src23[16] + src23[17] + src23[18] + src23[19] + src23[20] + src23[21] + src23[22] + src23[23])<<23) + ((src24[0] + src24[1] + src24[2] + src24[3] + src24[4] + src24[5] + src24[6] + src24[7] + src24[8] + src24[9] + src24[10] + src24[11] + src24[12] + src24[13] + src24[14] + src24[15] + src24[16] + src24[17] + src24[18] + src24[19] + src24[20] + src24[21] + src24[22] + src24[23] + src24[24])<<24) + ((src25[0] + src25[1] + src25[2] + src25[3] + src25[4] + src25[5] + src25[6] + src25[7] + src25[8] + src25[9] + src25[10] + src25[11] + src25[12] + src25[13] + src25[14] + src25[15] + src25[16] + src25[17] + src25[18] + src25[19] + src25[20] + src25[21] + src25[22] + src25[23] + src25[24] + src25[25])<<25) + ((src26[0] + src26[1] + src26[2] + src26[3] + src26[4] + src26[5] + src26[6] + src26[7] + src26[8] + src26[9] + src26[10] + src26[11] + src26[12] + src26[13] + src26[14] + src26[15] + src26[16] + src26[17] + src26[18] + src26[19] + src26[20] + src26[21] + src26[22] + src26[23] + src26[24])<<26) + ((src27[0] + src27[1] + src27[2] + src27[3] + src27[4] + src27[5] + src27[6] + src27[7] + src27[8] + src27[9] + src27[10] + src27[11] + src27[12] + src27[13] + src27[14] + src27[15] + src27[16] + src27[17] + src27[18] + src27[19] + src27[20] + src27[21] + src27[22] + src27[23])<<27) + ((src28[0] + src28[1] + src28[2] + src28[3] + src28[4] + src28[5] + src28[6] + src28[7] + src28[8] + src28[9] + src28[10] + src28[11] + src28[12] + src28[13] + src28[14] + src28[15] + src28[16] + src28[17] + src28[18] + src28[19] + src28[20] + src28[21] + src28[22])<<28) + ((src29[0] + src29[1] + src29[2] + src29[3] + src29[4] + src29[5] + src29[6] + src29[7] + src29[8] + src29[9] + src29[10] + src29[11] + src29[12] + src29[13] + src29[14] + src29[15] + src29[16] + src29[17] + src29[18] + src29[19] + src29[20] + src29[21])<<29) + ((src30[0] + src30[1] + src30[2] + src30[3] + src30[4] + src30[5] + src30[6] + src30[7] + src30[8] + src30[9] + src30[10] + src30[11] + src30[12] + src30[13] + src30[14] + src30[15] + src30[16] + src30[17] + src30[18] + src30[19] + src30[20])<<30) + ((src31[0] + src31[1] + src31[2] + src31[3] + src31[4] + src31[5] + src31[6] + src31[7] + src31[8] + src31[9] + src31[10] + src31[11] + src31[12] + src31[13] + src31[14] + src31[15] + src31[16] + src31[17] + src31[18] + src31[19])<<31) + ((src32[0] + src32[1] + src32[2] + src32[3] + src32[4] + src32[5] + src32[6] + src32[7] + src32[8] + src32[9] + src32[10] + src32[11] + src32[12] + src32[13] + src32[14] + src32[15] + src32[16] + src32[17] + src32[18])<<32) + ((src33[0] + src33[1] + src33[2] + src33[3] + src33[4] + src33[5] + src33[6] + src33[7] + src33[8] + src33[9] + src33[10] + src33[11] + src33[12] + src33[13] + src33[14] + src33[15] + src33[16] + src33[17])<<33) + ((src34[0] + src34[1] + src34[2] + src34[3] + src34[4] + src34[5] + src34[6] + src34[7] + src34[8] + src34[9] + src34[10] + src34[11] + src34[12] + src34[13] + src34[14] + src34[15] + src34[16])<<34) + ((src35[0] + src35[1] + src35[2] + src35[3] + src35[4] + src35[5] + src35[6] + src35[7] + src35[8] + src35[9] + src35[10] + src35[11] + src35[12] + src35[13] + src35[14] + src35[15])<<35) + ((src36[0] + src36[1] + src36[2] + src36[3] + src36[4] + src36[5] + src36[6] + src36[7] + src36[8] + src36[9] + src36[10] + src36[11] + src36[12] + src36[13] + src36[14])<<36) + ((src37[0] + src37[1] + src37[2] + src37[3] + src37[4] + src37[5] + src37[6] + src37[7] + src37[8] + src37[9] + src37[10] + src37[11] + src37[12] + src37[13])<<37) + ((src38[0] + src38[1] + src38[2] + src38[3] + src38[4] + src38[5] + src38[6] + src38[7] + src38[8] + src38[9] + src38[10] + src38[11] + src38[12])<<38) + ((src39[0] + src39[1] + src39[2] + src39[3] + src39[4] + src39[5] + src39[6] + src39[7] + src39[8] + src39[9] + src39[10] + src39[11])<<39) + ((src40[0] + src40[1] + src40[2] + src40[3] + src40[4] + src40[5] + src40[6] + src40[7] + src40[8] + src40[9] + src40[10])<<40) + ((src41[0] + src41[1] + src41[2] + src41[3] + src41[4] + src41[5] + src41[6] + src41[7] + src41[8] + src41[9])<<41) + ((src42[0] + src42[1] + src42[2] + src42[3] + src42[4] + src42[5] + src42[6] + src42[7] + src42[8])<<42) + ((src43[0] + src43[1] + src43[2] + src43[3] + src43[4] + src43[5] + src43[6] + src43[7])<<43) + ((src44[0] + src44[1] + src44[2] + src44[3] + src44[4] + src44[5] + src44[6])<<44) + ((src45[0] + src45[1] + src45[2] + src45[3] + src45[4] + src45[5])<<45) + ((src46[0] + src46[1] + src46[2] + src46[3] + src46[4])<<46) + ((src47[0] + src47[1] + src47[2] + src47[3])<<47) + ((src48[0] + src48[1] + src48[2])<<48) + ((src49[0] + src49[1])<<49) + ((src50[0])<<50);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25) + ((dst26[0])<<26) + ((dst27[0])<<27) + ((dst28[0])<<28) + ((dst29[0])<<29) + ((dst30[0])<<30) + ((dst31[0])<<31) + ((dst32[0])<<32) + ((dst33[0])<<33) + ((dst34[0])<<34) + ((dst35[0])<<35) + ((dst36[0])<<36) + ((dst37[0])<<37) + ((dst38[0])<<38) + ((dst39[0])<<39) + ((dst40[0])<<40) + ((dst41[0])<<41) + ((dst42[0])<<42) + ((dst43[0])<<43) + ((dst44[0])<<44) + ((dst45[0])<<45) + ((dst46[0])<<46) + ((dst47[0])<<47) + ((dst48[0])<<48) + ((dst49[0])<<49) + ((dst50[0])<<50) + ((dst51[0])<<51) + ((dst52[0])<<52);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h0;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8570196967ec62e536e9c96611dce2c0f8977e173aa3f4ebc3935fe28077f5b5a092c68120a6007ad72de20ec3e1e6e63d69577e307b5d5677d5741972590d692c0216f832cc0cc89535e31c75dc4e5acd21c4321;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h54f9d77011066a31702e43c80be06fb2c2d09df1ebcc95ecf010637ed662f7ea6d6cb8d7ce420333e8e82039ba0e2e634a51b420a3e72d6a2e45710e954fca2b31c65b1c5219e8963ed704634df48c316ca0a1e15;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc90fddd0d4994f0b1359cf10ec4c7939fa561b0250fea9488cd600b5183db661fd8132b36eb686e278b29b4787ab3e0b41b93ce46eb494e11489900a1c2a9163a075c116cc97190c2b6e18b89e0ba3f5a9bed09f1;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfe6d806820ed638d70d90e08d977cf617ec0a4e73ac63d6f05f65b306ff5a08d252e04cc5ae4c31f9d012eae5c862a6c33f699b9b2662cb390ccd3975942f7e61a653c2412bb4c672c7ca7e4bb88960271647de13;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6b65620763be53f3fefa76099d1569a5b0ea1e52a82857378ecdccf8ccf3b88438cbdb08fb15ce404386d9fe1de72d7857b9d01de6994d5757d48f0becea1de4c360bdf715c827c548084d8a9885f66b2b5c64220;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2fe46ecc779de589e360c7cd3f01a7a37417c7abc7c2f92c79b34215b07cdf356b84f2cb17dc198c6c50ab66a843f675f153257ed36d31d8408a344a20c79fe7c51b02aab4657e7cef4b3530061c16926e6882c60;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfb87c0f1cedf454e2b91f9a08e11d5df1bb04a4d168b289803923ac13c3a568dc6609921f81a3f6020025f9000da26ba7a326d2790392398516e25b2b7855284f338fa6cc9f11ac1f5f55a6453b1728c377ec5695;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5ca108115a23d899ef4b59335d57ed85e291e3748351b41a97f664eb92b8bbcf432739b92548ba563cc3e3b32626f50db9bb7a7be6d67de12007db8aa8f1840cbf23abd893a695ce569b5d5023ce337f696afbf81;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'heaf10b87500e5670898dc0cae1c2e6bdc4fa456ca1c4dc65db01a270dbb4792008d4d35dc217465eb1045c0c28d999149c11f38d26472386f768765a2ae6d86544e699357d115b294460d0d6278febf733bce6d3a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h59f51d6d10d92a631f9e40c182d8a70a1d97ec79ecd0f7ea718f6b4a5410b71afbf2a5d6de0653fcef20901ad21b7544726c133a69ed53c924ea4ddc4f175cb5b3c997b7589ab2be1900ebbfd800c40135f7b7cb6;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf03ed2f65a5ed99a9b53cc7e9578579a27fc55846a59d1d03bdae11a1028f775721b3bf6bc564b96c021f855bd713d46b00b05797e7245cda891c05f52970aa43aad4a976ec303b5e55321c9bb04a3768830939d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h96ee94e5209351dc2c376a616b9ebb41370a87c994fd54a964e4d62be3791b51e47023fc080521289c2cdb36494b9cffe2d8a4041920fe546ad5ae3f53ccefeacbf887e4bc71dacc897195640208dc52157c71556;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha889c7b3290897398dce5ed9942fc3981b864ff35a5045365cabd463fd468f310cc33484788f45c6e5ce53ddd076c96f077d82f60de11b0e07c847d0ae7009c99ad9f326fdb55451a7d03a85a402ce899cb44efb4;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc7918f19758c389c76142de2aa2185568631ae04bb12fc0ee75bca1f2255e810567367104f0d645fa9189f202f59ec19b8ae71376089324bd62a214066bad60b8be67f44a13ac5acd4479345c9b3328070f3a8ca4;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc2f9c5efbca4824b67fb24dc2a183c933e5a1fbe7b1e5c186516b8c6ea5c4af43d5546d66d51340af2da6615a5cafa082e7cd5ef629d25213b67f48669f84e4d32285f8e8e3d0a21970f1f0edcadb1145181b7fae;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4da29b8153ce4d6d03208ee69c5a01a366cb614da88c9011b7bc7b9b47ddbf715349ff34a5a4004b4c2c86a260bfebde8244f7aea609c5ac7b9c8c81fb31187e890d1f723a5a8a96a997ad51180a46695f65fff28;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h43760983b401a22cc731d6fc976607e8d12f8a2eb520dafd6f468559d91ac0e89e45e2b7144f8dec8e96587f0a4d3bb5bb6cfdce61f1987974c49dda6a4af59df66953f1b187f7025d13179633b7006c6824ad675;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7e0952cdd16922ac87177411a92e358cbd08842495f91ec642d02d509738c9ee84141f3b4c37d5b3a9ef64067bda5df2e20e57c5c2b3f8d720cd0656aaa0d9cc73b2c6bc04c273a20f35a20fbd256d5ffed3108af;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1ad609134c73d8d47885c8cbb4e9cecf38521bb4b34628f7bf69be0e1f8f978392bf871dbe43efedd4febf328f43cdf8e80a78977a55c1fd8fa92e4d36b04db0253ae6b154a63b3308083f2f7a87d37f23b911c17;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h69457a2d836175de2bd1e8b5a65832694655c83ad14660539b15d2bd1cba102f12dc24be5b04819af24ca569692d36742649e5c8ec94f7bfbb7d407d33c12e1e11bf7137b67070bc89f271488905ce10e360c894f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6a49067b691802111b5f3a9890d9b1da9c2de490a5b0878f93ab8b458b4b99418c9ed6ba7af6595f15575897e31064588be295a39602aa4d7362a4133bd0be83b73bb6b1516c55f0bc1d64a84aaee1f5f8e21cb60;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h140511345bcd59916de5cafc7a5ced26d411010ed3ff82ac30f6ce09696576842fcf4d39deb18a31a477e7c9271e4bc9cc614426cff9c7033263a1f0307aeb45429032879ebb51f76bbacdddc628e0b3d201b742a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h19edfb00f6c8d1ee5d6e9e253bce83d57aa0db3fbb0cea1e28906786419a2118844bbb0271ac4f1150a4ee5d26c4363a1283806e6239f90dc774937c1c3fb54475f1f4aa4579e760e779f6b86f1bbde44a4c6272e;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h15284ee90919a3b3d2602b22f492b6e0ee5f15f14aa213b624ba2373992559272cc675adb895533bcd081f101189c761f241518f3e3cc08d26d3f98ac10d861437c7dab1fc4912681ea8720d52ea5bf52e5614be5;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha340e8ff7c7a1bed761f3eb59a665f82cec4d62bf4a15d5c3407c28c01a8ad2fec87cec3e24190a1fcd11036708522e9373b92f45afc61a1739e4fc0631d38e21db69b965b85e9b0651f4dd6b8f5126364aae76e5;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd57747609876088a0bfe556af89e5afc30d66069a8e814ed1a9ceb6504c1d9bba9b12c3638cb3a2b19597bae9b3810c4e619a118c30646fd489a9c652070d96fdfac37e90aa3de4e9348b32062979edb1f9a2953d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc140add955d3090bbecb89fdb0c94c53a43041fe244bf0332bf52964a9a7b679d7a06adeb5b6c5295b70df32a302f5f33d152ce76ff74aa7f8132b4b4ba3164a53cebe1ce02c9f402c9c8e51b1f611c72e3c4c3f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he3d2756829979bdcb58766172a7c9f4b33a54863419263eabc6b43cd2b15d0c7f672636f6cb4f25bc9030d1f11ca470d2b2456a3dd8bc821df8478ce9925180e1f9cb5085e6a8d5a0587d1fdcde200f2774f921ad;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha93eb63b3cc056365155c9fd4dcba235fd3030f0f753d0dc97872112b14e300fc206be54a7cf2fb76768c8d90197c67569a578653f526f92aae8287e7d08a423e9d6a89d1558d130d9e8f1633d2216f72210ba478;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h91b12cb2005981931a7a7ffab05cdec538dcde0f62bb509b36837e7d26421a101bcefe4b133640f2deca2ce393ca0ce5935b1d3995dcb4aead24f8386c8d312ce9e9810ecf18d1b01427540188ef92f9e0b713163;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h72b24be47d11b7c38e75077bac2244d64d32c53ed3c51710d18bca342ce7800377f714beaad195a19aba03cfa92aa5dc4198a068865ece94b2bd7a4e337ca98c0a0c993b9f9a7a4f99c6563cad866e0c773692248;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2bb1385de671a3c9512eb25845aa6a5b54306fad78b3d34168e511ecbc0d16508b727d8607e30eb6d598069a7b3968d0e5fdb8dedfacd9dd8f5d9719216cf919d064484cc33bd370c5209d3bff06782cb88906aac;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h846b87d6fdea02abbf3645a446ddd18dfacf0964e88a0e87adab4eb53ef2b8b1eb387e186f36079109e015de34c131e3d3a2b53bc5a831cb59f5f3c0098194b75837c8ef576ee4692815f8d2066bd668017f6791e;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb7eb9159936341a9f83420202fd23582c7ca6c479c84beaea84d280174449273776a189cd1f49657a2a354bae2bfc6c996a31e0aa01575d76101dc82dcfd63353f05028ca39f136f81dccf1f856648ae25619d859;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h73dbec52f02b47b577816a19fca542b68dc6ea74b3fbee3ad80dc2d5a94e1f7a756052044a9c70f78fa3f9ca839af7c1b9d8a54ac9d2e88a5ce12de042a3da25c795190b67a0035cd3a1ff675dbdead7fb8f72339;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4f58161314764d813a4bd67bd0c39b223d448475303cdac15f9a2240fe58414832d185aeddf69e1c13bee1a0ac531ed84deea9032e2c76a15dcf80b13ea485bde769549b92bc2a90550b79eb21c28644f47dfabf7;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h999d7815bdbc9eabd61755868bef60a475c412e3529c37774f47d075a100886e4f6781f179ef586de648f8098c40cd90767a3a07a44ec0c8fa2aaab0f4f74f86ecd70946e914b3d9973e02c2735f0f4b41bedf671;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h452b95da52a2a0cf6d6ce679eba7a0a25e2364968a88d0110f7450181ca82ba75cd8ac7ae3fab912b1e6201d4d349e3523bb46be7259fe71f0690cd71f5dc00eeb8b34852a6318e4f66446052a787eaee9e57c8fb;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd36a547b70ada620920598474138b2e868299548b56334bb8663df5667c1685823a2ab9b2efc905f8e45e436bbc33a7d90169d895f3361847dea7e9dfc5bc926bb19391299f1295c427931e530334cb0254307fd7;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h568d4e4d9933d800b8113b0537a2356410c7282244daa441ca8b8f84b006b257b3011386d81e9489e6ec1abf30ce184556de5a5cd78eec73841fa895702a9394c960a9f46a0357dbf57f356e01596be22b1b46b7b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h80c0bc72cadf086b48720d58de16259b0a55dbefd04b451eceed0fe3dcd346ac3cda5debd550f90594bba4e050cca6e4d71d4a71b0f6a17754ff13dad20b7a9723341fd7a7a0d6a6eca408193c318cca8100f8847;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hddd5b22718d72c0978be5b769dabbee4b039b5a2cff9462316ca4547bb2ec76ac3b462da412ed3e916c057c38a926e4c16f1b3c372e8e6b97b872ebcefb45cb7f7c95068435024de59c28ce7648bb95b25a806d71;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hdf3b5e5d0b8c8b6b11e9f40f32c4fc9344d984848dd82fffac92d39d36a3e93c34b00df7490884d1397198ba65b7cc811c3e323e9fbd7b95ea3d1360355fb88c05977303f1ce9bf834bff7237aab8ea7ecc6ba64a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h37b8be337969f56ad7ff6e5eb1df6275aa2a985b7b44cc85e0fcd0eb4b5f3031a4a2277533752cd45a93ca59a4f752d11cd0585b14ae01e420f7939c214b30612c9e6d6f844ce88638cb77b3edebc3d5f0dcec30e;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7951a68d524635794660e4252690cdcda6d85844a60a9c8a876f2fc88985504f8f7ee9b9dcd2a745d830d4bdbfc46c3c15b669bc22f71bdd6e3ade36d99b50b0412959def036782692d9d47d242919e91b7a1cf63;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc73fa919f4fc32a16538677ee8fdc8604833b8e62fb825929f1b1ead7370284615a18f296d0a83063a8b25913695ee58ce305e9d5d11f51331e175d51d06238b18348722fb505079cdec9e803a0f5c839a881710c;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h32759d66fb710442ce378d1161c101b93366d0b438cb73cfc01ce6dbd115d6f662a9966fa7a6dfdfb9ea3806a6cc6e653cf44548b50e679a907a428237ab0e6368940e3c6772c21eac6363bb02e11da7be6965bf4;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h40e427896174769744666bfe6da4e2139822cc2fe568e4b11d53171a8b8a0817fbc0551c44638b4794f91fffdc7dd95a90775d66cf12facfbade90c2138e2c6b289f03f3f49d4cc244776c42f38524df87668be91;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2586dad936ab2f0faa47f81bc5f7b02b8b5f7390ddf44916a89e139658660e09a0119ed9f5887ce87bae00123747e7d224e9b6f64281c5b736b31a2c36c58c67db264ce835e654a16932d38c19303283485f8168a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5e8865a69158e23157d7c688141c361018189e825e06f1e5bb02e16d3857a19cf5b70a2633a24d59b671609ce9381571a31f2089fb8ff65f9623797a1ae1ffd4485b3919dc86d186333f02d7e9f0602a474c24c87;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd35fe9af3c3c9357d9fedeec388c5683667fae237e879cc0e911c93c19692d610c608cd18faf609a818fc2e887879346392d3032880ffb8b678e4bddd507357499caf7e84c8aff6b63bfda84723bc5aa1a6a8db8a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h304800208b68c538d1af6e426b834fa7dae102605757aa9bb297ecbd2f89bf3653530ed5e4fc29462257c040acf2ee8bc69c4ba169659cf150262c52550c303da318c814971f30e55106ac3f1c3b9991e01e9cdf8;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbdc0c918dae3513c4b1e261066f22b7bfe1ea4f6a7aece1a5d09fbc58916d59be4c7d64fa9b111131643f189eacc50ba51b2cddf0db797a6262b54ee599400ae365a0d3f7c7c5edd66c88c9ecb1e04521f6794676;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7e155283eeaa1c924bf06b40d9f0274c1965fde2f7be2324bceebb142952c586d1d9d1b4c7d32e257f42c4ed6fbe5275336ab0cc07a78b156b186958e0e048a573afb4e0ccbe8697d41421d1db927d0d05ab13f77;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h50c7076dad45cb62e546e0cb263f6b596c0eb047243aec5c54ab1205f912cad88678844129c95c5ff1cc01b76c86bd732c85463717c67c8292d422bc9ead5b8701f11259d561f43387b9e1c7dee0be9b5d2203dd2;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he6ef936f5214d24120bef09827253941e3b4971323ba02781334e1a574858cbf2b9c8925135326016d225775ccafb0f17a3ea57cf405375283146cf622931863025f97f0b73c69f53fdf58f3b0f81b252aa2957d6;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h293ddd1a968d28908fbadc843d0399c134809a57d780d2de580b1841685948d14de9c1948e7515e80c49cc0b32246e9ddf90ddc6fdeddd63c0492a50037c2537f0b4deb2a6dcc1aa989c5c383ccbb094a985fecdd;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h82d1406fd0a4dba5458b31dbffc2ca2993ca87312ae76ff66d61d2d153474624495231c9aa2c885837537b0672587ef787248b82b1f52cbda78756540f5de8fa43516481a9ffdf9875bc0614efadc6a8f72b544b5;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfe247ac81b2497870fec6245c271d4dcdb4cf47ba7a12f1ab62a5744c2284df78003c350c75b973ca3f06e66ea42ee72b4ebaa112b19797a856e888de3cbbb2fc53bfea77626947f43a2ac8adf81be4254e583912;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h91144d9259e88b37396bd9444fc995f6652331592d22f0ae494e5126b16b6fc97b7267368cb46b0541ce64704a710ddabdf3a7b4ae34aa3b30005c1fe6ab1d20d2b68645257293b9f03a1e7e90410462a5b0416fa;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc8da4dc9d585a3fd6210b251050f49205963664119b79052b91ecd46953ad59e4e33da4a2656a7b6c31d96fa9ea3caaf92217c9605ac8716b7f0c089de321f04e2fe3013fe5567557e32c0553898437643def7875;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5d3441b929d759f5ccc1a19603af01b68aae0e9f5ca4219eb2be2a3c7c4e6724184467ad863b7ecd58836c00a28244d1b53b50abffa816a10ff589b29fa8aad8b72b667f7804addb9d3844dccc430cf16e2b5d188;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h47135820e0f07d5f48766be416bdc1fe63df64fa3e4fb40232384053bbc6233ca44d277fd2c71a3d9ba265d5ffaa2871add62cfe71b511938ecdd1df80a3c4ab6a1b33244e0d274632e20a1334a38a7ee48cf1da8;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h27cda59aa1d3133c9f1c469a4e849567519ac4483bfd49aedf4919490f7549e18afdeb3146a06abdafde94a24ecdcbb6971f5a2ff92f0440e2dc4a83d1421c3fa1dc01b0b6472976bac6678e3664f9825a7d9633b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hea77862b3df4b7253998e66a82cf0e27887fb5b802fe7596f8088d72fa12888a0f94c375908df267f86d06a7f90dd7cd604290db4d8dee5106a3bbc201988119dbf41503a0abd069a3afe5b15ed93ce587b62dd04;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3b96f590a8d499856f5336c3dbafb7e1835bcfb42dece5cf28351edf0d05a14942b0143b2a54ba835acc57c75ee483c6d2c51e197c4bed965cee791ef6c6e86c870e33ae62150226d7fd2b193b7e9d9f4e574806f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4eda899eaaee76ab60d9bc7519acfbf2078f773ea31809ed2a27f1379061253e5e78a07d38e4ea6114221e86262c78674c7557453b1ecca6217e7be3b89cf0fefc34f86af146040e43e4956f8e70f901877569f47;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb4cf69fa1ce7ff53f2584159df3c846b6be88c2e300c3371b9f3d8c12e46706b5a19d340bb8d014ad459cba6bf0cefef784030ca2b0832a3e17a214f5c43927edcbf0b8bdef8ce476b6ea4a7b2d30228700053b44;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h886e7dad9ab427be2d3dc5a883d95b83b23f504056592e0861e5d466c8797bc0ecffa615eebab9504f9c460bc6fb23cf9ca5912537f4600f7bc2249aeb6044b56e3f76322612292eaf9de5d9b325d5c13c8e18f38;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h391b0ec7096135858597bc4103ddeb742dde29f1eab5bff0e630abdc300a0a37378a2502d87cdcce27721cebaa82bc40ca2c932247b66d63e5225f30924b6ef73e7d1018745fa74c3b3a100b43020b48c03f1c71e;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc717c50bc05ae04d42847181085af387088cadfaa5ff9036bcdcbbf3477d7dd6f3ee653886dba02ca26b5a63acc62d29fe73f3ae0477d5b6a2ab2bbe29d52f65b3fa2f4fa9284f5889334cb6967d682b0465cb61a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5cb0bd84de1f8de49e3c5f486b2936abc3fed341541ba0fb7524109dd3f528d4b4ad3c3b569116fe413b19bcc7d392becbf80747cf0dacd44893ca8289dc042790f412ea8ac2899ca2d9d438a6322cc3622e89ddf;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h28f0bed895df902b0e4685651843f7881852e7b5e235434b1ca36e78e5bd772beb5c7b454367e71d595a320ef4ce51e85552b459f3b634d9000bf6e2ae29b3f5be3e9e41467e73ddca362721b9c9962afc8c1c719;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4138697d3bf3693cfd97aae0a11c84a94bf77df26622dd665143012503e4a07ce330f737e959442f966d328e6fb03b7f8ee9b825f1e5426edf05170ac907d5032781d58db897b2cb03829d52e1bce03bf7d56f3f2;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he10d39aa78212e340e35d2fb56b0cb296d729740f9417f4749cb7b7d78f6a6f7b95eafe3f32b9b55ad7f899613d4ec40b965228bc827217cf41c1be5c5fcdaa819959699b2ec98c4cd229b4dcff7820f59f75d6c3;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf8871eef803e0cba9bd0e5d3b482f25684c1c923ea20ad6f972236cbd6ed076c62082d2294fb543735bd2a91801d437995a35dbdef6f9dc371dfaf6ce7cf0f909f889624b667ce65bdb6443f163455d010be419ac;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2f1685b916f6d388337aced005d4f852d0147a24d93be7831005a11dd21633f0095157915fe48d0e702ab1000aefa25da1273ba7535a9619ba82775086b644d7b42ea87f4ba876816c4718a820d1f4bdb58131cc6;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he854a825e4b6a7c89f481a8b882a5144830965422ebb1d38b99acd7c691741477d640f7ae7dfb5733519616c1edc21b7f05ddfa758078fa79b217350ea996f350f0b084331ed34bf69acfc08bb531d3ad6f76a2f3;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h58920a9568c68f374e58092cb7fbbc618110abfdba3eb1e82c0fd11a3d9583ad92fbc0ede6d87c7ac43f03d07fd273bba259fccd7caed8d33a82a0879ebdef6466cf9bf592bb472c686f6e2669207ee13b25a0901;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7d71ad23afe49b64242a7b21724baa15ef98c8702def5ffdb015802917ac105e6466d6dea12d112358c42eb5c49e8458a5cf210c03cdf209dbe72d7fb8c738e4583a6d1ea86241f29dbe2faed3bed1babe9a761a4;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd200ec807d99bb4173a3de93332000f744ce7f14796e76b644a76834fa78224f269bb481be23e32687a029905701c14c5aff2351eb534f4a2384a4566a16e4488158faa72c1c056a155323d62bf61cacc8040e279;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h47ecdb0ce0a65c7db282438857148c2ec2f15d253e5abc28ea7c50301c075b7e2f234266a7c3c55476859d5ff6eb0265a6bd514bb0801e4d21f7186b067b9d34417515587024ed808c3df5d2eb27d619b3f533a6a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he39be573618f0cf23dccb51f41121f1d3bba5790c32d28ad15146538a72518d48d99c04ecd547dfacd2e5dee45eb9692fd1b436f6b63cb5efef898e11980d952f94206f0bb1d75dffbd5a15cca6518cba6591b309;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha0bf12ba11df9779efcf3d63604dd87fa056f02ca70899683bb66635c5c8310f654774be64e7923d0fdd0c93ba98682f57a9d7777c8774e228c8568cb9cda7c099e8515df34f2905807dbce36bedc9742136b1672;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbb4633ead771a9d872db55a2c22eccbd08a2c52e638260b5a1bfc5a17a6c488bd15ea4ffeb6e5358f319dbfe68d9573b42d5464d8cd6f66974f170c567ca6e38c7f6f1c4aba09f7d4959823147b1fb98b2d13890b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h17a5f46bd773060ed53dfac01ab93dc8eee33cfffc16863cd37bf6456941512f810048ff30fa20ac461674b28d7acb10873e280ea36fdc8f272ebb7248ba0273a31244ece56f67ea7cb0d352e64a4f144904861fa;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h790f77fae353b50491a044e29184c172cdf326f0d892e1b02e7a81b46b7603b0499b787186c8a3d5bdca2ff237b0d39180b8ab73921727a75fd24dc63f4db7f7a37a33568129179ac5a1d30d85bd7c0a10dfecf68;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'heeced21b01e7d9e0404bb7440bc3643e549ddefec8ff90cc81b52f92e67952970bdfdeb7154538e7b570e72696d2586d8d524b42734e64d9d5838bbf0dd7250b4ecc2bd301f70c85af02021de3fd19794619cc441;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hde86c4834f104c89d8206ad2cb17e76acfd3a679039c9a90f6ae22db0429e3b1b36d0291c2d62330841e0a81b5d18331a49cf9beb104497afb25ac61fc693da8c4bd21fe1d44e38874e0b0de4c1e0f033185b36a3;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7656ea9799b4d4b80689581948caf89ca6e2d168f94081f7a88deee0e198646e77a917157f1db7cc0c8d880dec02847a3f2ee1d18cd63ce8449cc0d243269563fe1c8715e69ae8105e7473b232b5bb3555fede7af;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h586237c4cd6eff30d9282750ad28a946cb37fcaca2096065e080ea283c09a8f60b9f575f5d362e02b2b54ba643430ad3c6a2a240f5732fd87d6a7c4ddacd44b27d6b350180859092070b83649ed41f1e9fb3aa93e;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc6a03157ccd91f63b650f80c39345fdd7c05d1dd6162ab48cbeb5c015b089a3789a3bf6ae880cabb9501c1a3bccef373cbb9d505b54d92d3f8a86b651dbfb64ef2371b15c9dccbab912c3c4e2549618c30483114a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9bc37057dd1f69f1236c7496dff3c2df923d38b571c9f417d179b3a333ea96d9499a802d34ac15bde43ce71eec4d041e43cf11612906f4ddc0aec91d479da2c358e56869a525625c1547d1eed821e376ac86685c9;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9bffec1a789e5d3015ab8b6ab5014372b33d61c5e07248a17e71e444f0daa313c61e5c7412b02526adf7db3390875ccd5006a6785100c1ca42c9ebe0d6ff7ac1dafe00984b7c5dbd9e504e182f7b268f13f7225d2;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbf5b7963d5376c2dc9829bc5548cd0828fd5fc6de8f1d2d84020e92891dfc776fde0503843e85b7e052eceeb11339c4c172ce3fe9cf7bb10ea034a1da93f14f69b3e824082f84b9c6e3c30f6030d925c2b501ea8b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7de077a61cce44afa74ae143f4b9b17ec11e3d46ba2b437e495dd6645987cd174da0d5e371cf94e6fab9c5df0b705431539e27f6fefcb80d8e75c8a4c103e60db2f7fd5a4cdfad67ad89d07570a17ce5d99deaa43;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h98152d7a331b7ec2ef373febda7484037b4296c66fdc1b39d4c66851a44106ca00a0b214d7ab8cb34dad6b4116a7bad1e36273b87be8807c0a4b21dde395ba80c78ddba36e55499b0d55a67b4e2c1698a38f61efc;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9e8ed100ae220647897cb0a6c2712c4d97a9d33507d6a2d84df9e65028f1ebb25aed1c39bb4ffdf5b868a60f3153b6bb7b584151247fff76e65fa31568d29b9c6fd3d59f276bfcd7c230d35ba291f29c256c8ca3d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h75082553ce86dad1fc22325087e4f34698e84223be599e0a0c1041f1067c457ebade78c2cc7591066f58c1b8552855dfa997f70888663371c864310be858d06a2637bba50ef7f3cfca481274422494b4bb21ff163;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha7f92c9d117eb9d72b00e8b5dea9f5fae81a5f9290fc828e39c7867725b8606019920aea44e7a83a38c26bfd2d1cff011c6bd52016fa7e537a7106dff6af8e50d2db0333b70ce69e5391352499fa8e64eea0bad3b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7f3fc0b0b315964d0deda8da72eec56da2a2ad82b7a5e2819d265150b165ce9ad040f8d2f061488cd5a59febffd0dbcd9f7c21565f03679bc15ab7bf7bb9c64655fe7a089369ba33fb91a4b62588399d27d352447;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h92affea11a8133f0596fd911ba72625711670edddb6dc028ef7521ce4baf931336442f4bee08b0a6aa1305ba3d43d1c86200b8d08a4d48b2e2524e3a9195ba8cabf7a3bafd8f6f1e86ad2c8a2feebfe550dc5a554;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2500c4ba21b94091005f1249aeda22fbfba73810329b05636d2853b0c2b52b77383ebfd1f04e07ceb104fcd3051c758542fe17b990322c6eaf761a90be0308aded04118c94a1bb3161f793d12573b8f1e3bf15e3d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5874ef4f895c0d031918d2e39af78c08b43a5c24d45fd6c1236c9e503d0c3ea96c220ae1d06ba5ac3671ff3b73f90c4ffe4d76c86c48cd66514b0d03754b861393d5b7c7bd8fbc2e90d556fb49057ce42ff1cda12;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4ae6bdd3c4737ff2784dbbdd933df4a4a01a9e79f7af18e75416f281f997b80ec4825a379e1993ffd0e80c2c1ff713a479322685ad6fd431526bb8fee791c88f6f497e787ec9fb2c0e9b2f70451020c4a42bcd3b9;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2f3eb059e8810d82e594007cb3e732b6ebbba58b27e6d9bbd0e5b49810939b218f1bfd416836e68a8293e417bfd20bb7902bca0862e25d687afe9ec1282c79431aace242337d6e341c386232d98dfe7b5673b2dba;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5b4e4d14e122853dc5b8d0ea204e99fd25144a817b605cdae34d1644bd77bbec1104081ee07bfb703c53b579406b5972efa69ed6bbb32f8631c5209c8fdce99d552aa4288200354951f3ac2403ad672eb635be266;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6fef89cacf7bace5cefb0f493685a3c37e2711d7dca307291de1870be5a2bcc1df56eba2684a0061ebec77087d00dca25854db20a486a9bd7bb088bd8a18c4617505d9842f1fb6e676fa21271bb42405577861853;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7524a611c346be3fb784240c3cf62301b1323cc92a5127af4c3b580299ff2282ef2c1dc38d60844f3e89414172c579f8bb6af48ed58251b9a1b6c8f6e4af5ae620984ee5ed33317069dfd2f5cdbc682e8a047b085;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4f67d89a05c2b81c768b4c4d3971a3dcf9728429c65203f7c52c3cdbce68d6b53c0f1a92a985239b4f299efba651c4c0bba2c801491c1acd76108b7ec202d070719fc1272b4ca5681b78d23b612ca2368cefc350c;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he6b5cf1a2ce9fe97ceb5c02f106e49ef29556d978afd75e1c213fe03f3ea1d3afa38d8cb79fba9339da740ca59da0ab8569042227735e1eea6428fb4a06ef0a6085c0b81031c292e92975230d8fb83d837fb51d64;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he1e05303b116f7e80e3b6a646f8ab75438344dd9e61533a1bb592a4786740d4ad8ce91f5f9c1d554c92fa718d0430918864dc7f39e1bc6be1f5f6e9e8b6f9e5472fa9196db17c84d25ac5bd81ba4b7290ce0df387;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5a03e858b5cd636a80e74ad14a91ffdb33f9c56b88c292f0eaad54f6a6a9dbf846e5ed442575e29902ff659bc9067e4098142139833e6fef07835668f44f1983bb9ee8d068b66e703e2dbc24c177b2d27edfe8aca;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb6a9fe3bd5428349d4d38c8a02be7aa7506012fcbe898c29d0de220f7bb778f99146aa8ceea39461c379cb4afcc7671ffadc56511000a9242431f6ba5601b886028164f2b82081fc521cf955564f2bb08cf45ff11;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5b173d5b700959fbaf6a94dc4acdf24d0d60cc4c70d4c45a8d97c9bfe55638519d8b5105947ce8d836d9a81c9410f668c4392e0859dbd6573f3259bf1e52cffd70832ae758286d0578e143990add8bf9355b7c813;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h56c61acd1567af1fe2ada704813db580efe9c45134f84b060e3d57abddd5b436c2c0737148e7b1e783f403b083d8f8e70c380cba10e7d82b0bc046111ec6dc0d99ec95da6210a5c714a568d4c2d0923d547b12d06;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1086c5de3699c32f7e92fabac32328969bef60f2d1056203e688641fe117e8daee816a9bf624ef331d79c441cbf985fe30bc75f212bc36a947d7b52ef658e3e4fedd394b49456fdc4e64a261617570b6a254d8be6;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h76e9de0392301236a8c7e2089dbf78ad858b8c08d3208a784c5329d7a133fb3444399773b8e485f3880c4abc5378557e8302cfa38c8fc7f05c75bb58eb397a16ab3cfb6a225109d63c1072cb3c2dbad8b9e0968ac;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha97c24e551c2302c3a6939cc79a1714f33fc4ce2cf2a78d643bf0893828a53fdb3e54a1953ecf9ab6a6170fbcadd8684e2b484e55b42566ee0915074cfa99f68cd4a3680ffd305122845d9be2029cd660cd2d5a87;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h710c18977e2057bbda9af4665392a3a7f786247ce9d892272066d62b0a0bf6a7ff8a18abd56572610ccca06959576ba60659af017ff29e053a369178336ff5a068b67af0ddb39d97fe6323ec39238781a26b87494;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hea5bf998a590dd14d5753f08a3ba4f52ff1249a04288db1ff97348d92e1d86ccb4b9b27d1d176afb3391797a5c45db09afbaf049cdd01a8994d47915e5bfa1062cac9c401a2ce64a15d502f254f399cd37fedb98a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h47cf8170efa56ae6b50d2df2adbabf2c8253269ae53daed9dba9370e53dfd1c7b02d737ec1e257c8d0241e3b23bb521dd028ee066bd8dfdbfbf337d288c174e299040719169aaa59ce906a4592679909e8dfc84e7;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2558bb287f47fd662c618c1676a55d3f20bfbe5d8d856e0b523f3b481893c6eb0cdbd8c93c97d77946ce572cecf09b7f2fa4e88a9bce5b1abe1c58a9fee459074f5a5f8b22d2ca457b2a2258e9643fbb43a2d6f41;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h45a0e30c0e915783816e7a01693837be8ad0aca3809b12f3e42f8339673d5342903df0ca30ae1d4f7c35b626539ee8e94751f53800a35964cad78f58f38a467a15919c7ed6ba0b5f363d15fe87a31e15e31423cf;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1400af1eacbca11f526c9e97e71dfab402d69ce2ea78d13ed266c05a388ea33251f0cc3c79303356ffe9f51b23cfe302bb0a1021110a456251d7e9f0ef734d5b3c23188f13238eb1394584d52fb2f3a518382e950;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he46f6a92e35eb3ece38018f9a8678cfa3d76f64036e20e501cc37d0b5bc17f213393f5effc676f5149938b907d9abf5d0071d843130f57945f7999a2c9e5c02041e032c5005fd52a99de2b96bee4f9147d3339ebf;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h52b704d3357ead400245fe8da06323b4386661758da7e696a352886b652f97622f6f3812376922332cdfde2ea4b0a0bc9b63a3ddd08c3a681965648735032d0f623244edba8b8b0f9bb7878f3bcd877456c46e11e;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he36586f4c65e1e64409d996de623ea84b704fd836ac431d098b7a2c6351689274ca3bc4bf909bf494ef008b137ca707f971f265a9bf3354c40c86dd44fde03ca83be5bac2ea156bd394d1326011c4caf5be1313d0;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h850c7376e87d1ecec3d4e989b78fe0f5eacc0ab6408bfb6f69443f6687d4768029cc2a7db87dc5ac440757d89e348477cde7861bc8203051ee5f13438fed7f7778ac9cccba467a3bed6fe547ec88cfe385965e52;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd8526af4e39a41239cf1c9317f80616ee7ddd4388f5e5ecbc3211c1c9b1132ea8319f0ab7ffce5c36dbe5d77738280e8e2c61bdba92494e7c45e5e64f4227645862617cf7ce30f8e54ea025eada1f8cd8d6683d9a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9e421ebbde733a0c7c2c6c796b40cd7819208e2e4de75ce57984df2ffd3a7bf36980d95b5b3a8ec8407534b2bf5b93e3d0af017d1c6320c6dddb8f931159939efe4d36fa16e294333057c1c3ad667c062964ba3a1;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb9adf4124d9d9397bd097f624558ff202e256319acbc7a6866710ba76a50b9f665d08f5372054511dba774bd1a036bc6056340a287d35d26846773360fa41ae14a727ddc32bbe345e0db9d35e89abcfeb7a6be1cf;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf6286355f756e3ccdca5d43187cb92f44490b86527f60ee3390fe6be77decaa214943f875b8c243d7037a6991cb14715da62ce1af91334f3b33db6449bf2d2b6cf331a7bbbf3c8c55ceea202b86d429812368e8ec;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h864fcd92be0302ae0bed911eb727010da875391c033c67df55f4c6b7d2b2f11149a3439c66675c14ddf86d6973a33962544a9bfea432b286d75dd26c3a4f40cf856f538d955c496726ca5c3f5392fb4a830b69550;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd307354caeeb4b4ad214e28fd6ded08b814c9531930a640c30f23c588dedabfb0b5cf664597e3d6ff67ccb6ef9a8b6ad6c6f5c1be3d5c6a927a873328fb09f2eb8ca7e70dc956fdf88969dd009d9c497f96720517;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf0722c5eef00303591edd160f06539a9409c09450dd72eaf0a93e1f5965eaceb56997d528c5cd17d4c27938fb7a5815e316e389e4875fc19269125061e35356932f9e78c893859f27551de36302c9e91353eaa672;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6a823c680d265bb6bd1693a8f68709075593d56b590d9e8031edca98b3bf49a9e0c92452aad5897486fd30f95a86a25fbd7a2d5b2c050d31728a4c81708447098b807c5a5f7a83b75f370b78ff54365f1dcd19e70;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h57a4d5ae0ae87ebc69bab9edc1a6ed7279a86e603af3c9491112c878b342dcf319201924a2480dffafe0723b9ce9016a50a084dcd52a10485056528a0e939494d26bca0217490063c7b2edee2520c6ef17a4dfde2;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf4304d310d0cfbf96824e466c8a195bab607422e18dab2647524bf97d4a8bcf6c45b8cba66c820dded118dc7d55de1f107689affaf98ab3075625a03db819041872e8cc1225cb8f06e1ef0856062a6386c9e27be;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha288ca2b2f8b43be4375449f956bd10b8405f5d5e60fab138bf6f4d8b1e742a19fc221170b3be08513e368e6c41509d8024ca8d86cd8ae498344a1fc316744f7921f02df5cb1dfa4bc593517efc5748258babe476;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2d879245a691e869a7f9c9dd61e6e94c9b96b6c8b67025e0cc90611265e4147d4de55b1ed3142dde406ab41a915883d65d210dab37fc2534ddeaa2ddb9b0e3576007d7a9eee84b6af5be3d55b04ecce606318b96c;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbe11d52d7df33d3a515ab8c08cee66e9ab4901f43f00859b4c3762095353db14d979f196e86c4519155a0401abfa5474df6ce90a758e11709a3854117338fe22759860ebbc314535fdc0dc418c4a2fc70a4800b10;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9ed72de156d7033682b8338f0400c2d557e7b096016b34ef3a71f6404541195ac6b7b6a01ef881eb87957e776005eda6fca602f04b63d05dc2af58c08d61d95a1cdae771d71b01b9cb1d24acaafdb2c60652ee465;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb48eb9d9cfcdd1f79db3074fba394070a056daa04d5a6dcc4e9afe6a0af869249aece437fcce2d73a065614bea09cea24b44a4d6bee395e508aab03cd6c97878ac64bfa11cf1e537b71df08601cdb4dfa1ae77158;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf1c2aa3c40ce26d614c4d1e7e39e9a05c784ce30b9110e5386c1e76e3210a6adb067ed824762b166d2192a0e7b53d27376a5dc6efd3d06c2f8f9980e716da95575f33112504f058a82fc0ba0c623d314b0297d2f2;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb6a2da341cb9cc71095003b35154afc704407f090cb945ff13ff8d355b71da52cc936f31d673e1bcfbe996ac81b26648551eaa6fa08f44d2f410e48e29f8784f5a16bf6126c8f3f0ed5f6409bf0fb157a4e7a2ad6;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8edbed6f8909f36d99949b6e368e4725d74e4334a1008ea4f15e5749499edc39c36b203a23bd7c174ac823124d4ca582d012bef339d18de68f3ad1a3f8809998190be93275b76ae015f493cb398ef2d1ea2e6c9e9;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4b04adf6d94dabfdb090e69ed926aeab48d4a0fe6666e0331af4986991ae54520f614821b74520b04142d777ead5ebb4c1c657395d7205f59b0eaaff46ae38e139a0eb55ca61c34f471e0e0b608a6bf9e12220a20;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7bccc26b3f7f2b3baa2eb3ca5281268af3f54a9e60e80873110094d20a561b2744d716bcfc78b4dea4b2401c9664b47a7d49521525ac42671dbad20123a6cf9a8bf7570df8f65f4314f0f238c946a788e8a0da19e;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h69b39d47596a50784298905d1cc673a6dd5a181ce23287c9c9c8a962b0f635e88d8c472322648a2cfc3f1fcfa35c8d019fc9b0a350cda82f2a095b2ed224a8baa309c5a875b0aef31046e01d93e490c2888efbb53;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h10a9138fd2984f58ac8be37b12977bd2270933e049b56b1c0272f3267e4a8cc8c5dbec57c1477b980c4158c6d1b075424a6f2dd0b969977711e0ad374f125079a6b6c6615b8da2cadb871ee45ac814ce7a5dcd929;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hddfc8a27ff36177996ebba00cfae2cf00d6f86238324473f3283c565292d00fc733c74d6e735d1b8920a21754e33bcf93d964eb7bac4219aaf3d0c51da22dcc98c44a80d7963107fdfd0d073aa4ad556481c2c0f3;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h90373e1ce36146c6ec9efcefd30be66ea587660a5889539f322b6a008defc7c10c5656cc9d9412242c091e81188f56a7ea786b687eced26945e9431b8ca44885d459a43af8d0ff1bc6011c3e9c130cfeedf9ff53a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb205b4d8c885c73413eb78766f90d17d74953646d20f36c1da9fae8c46b936a2b2fc513afa109704907d73080ccd4b58e5bc4dd8d315d38834eafc89457e5e8d20ecb36f6e9952e7ddffe07218d449f6c2ce6a32b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha22e6ae8855a6151c950b1f6761fa4a66ebd215fdaf058131c58ca14ab54520fb580338a006776124b116511cce031d10a77a9201b9f64f3ed9ef749d9922dfc9307bf3533119a3ccb0f3546b5fe03f1f8b0c045a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'haf5e1a9d9e465391195779b9a479001cfa163d1f13592d6eb166af9aad392ef5a8e2feefd3e668e1480a97e188db02d2e07771ea7b4fb17fada8f81afd520915c45804dbbaea7fcd0c4c8f84d9c03abff1e6b39;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha5ddb69e956d7925472289098063cdd89daa16d61ea5599dc5543638489909ea791adb7deefcf8d59584bf3e0a6a6e9bc7a72597a79b30066aed23ee3836992ae058c2c2924adb6ed8a332531f9c6db27dd86a980;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbca5d65c303c6561a7636c47aa9879c645a01cbeb2e81b5ddcd58dae8d650b1a8beba5f942af46ccc8cbf33f8482411ed71980020b9bb0b082dfd9c5952df2a14be2145c063ae5e5e497a610c03f13be2879186a4;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hda6a76bfa1a4a6faaa95e3f4526842aa351f77c1847ebf7dc4ec96d140636d6c96a2234ce5d9dba8a8d4e9fb3ff03a75ecece09b38828ac73f596750c4eb8d1cb9c6f558f379b237e6a764f14feb8807133c62b7d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd4e3967f2da11558fa53b5b19c3f8728e6f19e6e0f8c27fe8e546dacc131ea0a78d4fcf4a8084502ffe050ab06868ff3a7ca351f001693918610b59390d915341d55587a75c6ac695e3516cc642d8f71c114d92a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3031267342e2922f41e45ef1924ec7c35abb4bf1f1738e15741d27c3b53cefba371bf2ae93e2e00775426cd685f5476037d93fda0248aab664d2372c067941edbf8b4e21633c33bb93935bcebf61fe61f122d0de;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc642749fe7245dc976066d29412ead7693a271b903eb3cfe67112e78b4b5390f93d69996ce6e4987e24bab764e335b3a5901c1a66e2d5945c624f00f46eec3c792b617d4f308130b800383cea66e8fd6d9deb9562;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb870b56b53ce5337360c0531b6b2b0548861f1f571c7e3175fd6ae89ec9a24d5f4addcf453f040ee5cb188ec3736da0792f456e1a72511101948de6254b7258547c57bec7bd56735245a41acb4fa22db7614bad9d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc9de23884d61d0bd9726e13be0749d375bb903a4e73fa05038575b2f6ffd4cfcea17ba010e4160c9dad479894ef110bfc231f65b45fc32c98b6ce3d5126979c5b8ec7cdebe0f5744db66f71b4b8face4c5d6eb8a7;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h923aa563a07125b8cadc02f3d7972388fcabbebef384a704dae4c9067b3ea2fd1a48b0f7960bda8010e74217103f47d12272001311eb89f4679119e03b4582efdb8cac1584805e6a6fda6ab062b870ac0d66f3ed4;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfde136b8d6ec62fc1e84829721fc6671561d0340709a121466e11bf99839201625516b0a610de3d9f6561ee661e053a64c95ef8cb76604938e0950feff567be4a49e562926bd9e6783008492dec7aff518d6dbfd8;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4dec4ae7afde3a16a0d8916b59314073f7a0970463ca4d3f00589414647e89a2da90e04647bce15e1033c6705f6566191ff04199d5fbca0b2cf5bafbbdebd3d0bbe2f6e735b66b3d4e98a17638333f99dfb51fe1;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6f0ad041cd338adc585a5f812237960debb43e077d6523542a783f1694c0f0bb7e9ccd051fac38a75aedb68545a87de6c47141c57cfcd2fb0e3e4e2e3b1b8367989ef5a94488bbd5dc9ba3862b592395d29f618f8;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h269a9b4906162b218730a4bdf2caae299441c58e14b635f8f3d8adbf390f7c7238e67f67b86f6288b7c7dc3608b77b487664969bcf414919b5c756255cf69ba784ff47f4d05c78946721641e7fe701bed38546bea;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb2cd5741fe8e923046cc13974932b56d37e3bcc159aad9d445f8949ab63dbc36cd6b72d71e773b91b98ff52dd81aef65a75e143af4bf044490b452df71026b7f2ca04504a6ad11dfcd3720be26576cc08fafa1eb0;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h42f288c1ffe73e4092b0dfaac5253c7fa5aee6195c422a8c672abea0257009acad2769b87113b0f630c1666cdd0926b048aa29739f3739d02e6cfabe05764ec26c09f779790dde4f1a04852b7a28c25261286b36b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h51fd86d1ec20b67d59bcf62d45214121b0a80bddf6cc1d715209d93dae7873ad51f89865049bbe152ea73424bc2ea58cf667f1df34c6100051b4abde8d782c82f45f1f35a9d55218a56cbb255cea150a9bfaacadb;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h330af8a9f140572867d70368d5b724c6c36e074b7eaddd991027df63e24bd996899c71decff91ff313afecd7dbb94279ce82f93e94696a46d6ad465a6e102545865d18eef807c9a47574c888baf8a531138c56322;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h32ba6af27aa6472892d9765357ead4bedc7a2dd87cb3654fb2e9620855eb47935458ff49025f8e3e47ec9b5722c745f31b1b3abd0f1448dfeb761c293a24c3242454bdec723b14fdeb8af2eb61f2dac38dd4e05ff;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4a0208f3646c29a3314f1579d492909cb835c5a59a9c8bb192779189367ef9ced1acd5e358fe4b423ce653fc8c51908bf337d3c39395e25e7a65610d15b733720ea0598bd0f19f9fc17b9f4f17243bf9f359109e0;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h239f86b75e8cd86c62445b033a5a8038b61252814c0096b9b9e9be4872f090e59506e00715c34711afe4e0ff75880a679f95386a75c573e25908a6eb95ae2c7fa0bb0982163698cedeced6dd15153c73e59c59ec4;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hdec903b340250bdb1555ba19b6f5224282306c9586ddea8e77753ffaf9ff7f18d5faa786e42581b8bc93baf3e5c8b325bcf3696b4e48b147ecc5cc8354c86b3202ee25b392744174f4345ddbf15b9f97ee6138d77;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6e578b749508a98571acedab3c295ac1a0b4e0437510404b3807a13245dc06ee1eeb525548c041ee0184576bdb2e173288eccfa1e999d0fadbf23f7aa0d98a9c5079fbcb9ce2cdf4c304938cfa5a9cd6e7ff3b7ef;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h999cc0f042c49e57d813fce857186698b74e3598f30448b0ae73542dcf0f5edb820f75ac696604a83175219056ed5d7c2e3334aa36ad1b612aaf393848d3bf08453b0bbefa917a0aed6c306538cfe3de252b40a1b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfbbfecaafa03ee2f83c50d1d507a30b0fe2d90babb197785d5c034f7fd4e33391270251242b4e67fee392fe4c2cf7595a19678b2ea3519626315194d294f4c327702b931bc342810c191dad986d1dce962b0109e7;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hcbb28fc4881397de51a318d45ade077425f7bc0e983925ed6e2d1a9e5556bec261c8ce6b23d01aac3dd83f153dd286ab98eb77c88db73e6202f97365902aa4c69e3d1f657a46ee03d4e35e55c093925b319299103;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6ea263b2fd9702e6f3c2ee87fcaf1f5b58f4354895ec6ce2da7d6a9460cd9e13f6c7bae49b03afb7f22c6dcfb98ed84e2150b5aa1db1e268dfa5842a55a39e334d4e557f982d82056b27e57ebdaf2495d53f58409;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6636ccf40b04e43e6e33c3612650796bbb3266b0579b5954910f5471c62ff6ae77dd1b0f0b4118be3f2d4cc45143d7072d3dda7b65921f365cb59583f538fd66840475753874d7a7c226d6bd21c2a7b4ca327462e;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7bde0e8e2158d796e470721d59697e21e490ac8f08968fe13642e065efac5c031030c3bcf2ba1e207b29b2833552f287f02d187061912b5a18f831f0b9dee0e00a409f0ebe45938e70dce03a1e4029e40cbd20844;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd7f88a077a671498790102df15cea1660c8738b4f50a0d877ea10bcb1a53a5c9eb95465a83ff57695ad376c5f5b10990eb2ad32893d273ea50d5bbafbbd872657ca67ad3ad2ee04f3542fb735ae446eb37b0f2bb6;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6b8827797caa0790518afa714219614ba834055602c67ff82911fe3251aa6b613043a03b82cf613c7b12bbd7c86b7bca5490670228c0d0ea91e1b7889f52f6c90937714b2fcade5a038a5ed3279e79e2275818b4f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h23236fc4f70374bb22a057edce9260b5ca57d92d4cc6be9d6e488e7926c8e707e954add7f86cafc1b209c80657ebfbeee150367bdfb0f494c1d53d5ea9f2732f6052433e7d1c995fa59e46fb7d62bb095d2ec7acf;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4aca384d1e8d2bd81bd4e32575773263fbadbfcd7998a5f1d900709326c17ba843761f1914acc8feeb33b3ca8e0f5bd704507352aedf5bd3b4b9a450564efa44199cc9e0c50f03a2d00a049266c95374f3504db31;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3c17a32b96d2f63e8a430475eb156f407330041c4695a83679e768518f3cf6467f97515284a9b562a95f46e3f35cd147c8a270d9cd576cb264fe85872648a40ca0c3125e8ed4799ead5c06aa7e243e771b6b04cae;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2961c4fb09376f94c5e713220479c4356c39c12b95c6d6e3f45ad2f159ebe449ceb12153fdd607f1d5c07cbce2fe5967765e97861b4e9127a8d3deb68b4064f2d79a3ebb807d6f752c65efba199eb68d242dda6d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3993b5c94029a05a7b012bbeee719460cadfa093cbb83d15e4c42de4a65660dd444e3f4a41d62fbadb81c38651e550f5ea244153bb4d30152227a1cf9f7b1d6bf80bdc3261b8bfb24e79008644e7ee6ef8468ad7;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8815eb15999c2f65db03e41d8e3e0f0fdef5b0c7836ccefe8487b103b66b72291f923ebec00b5f07ebc758eaaf7bb5362d974d4fdb534cdc77854ca773fe21862bc1b85999c96813372e2dd3aa01d066c8e8d1d20;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd657ba4195f4037e3c7f6ef580a05587482742febfc91792f2d86fe6269da6614665cde0f093f8fa68908f4660b69a1ed940425bcd770df239f9c496461320f5bad6ccc769f903201516eb4352d03eff8c7ebe612;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf28cdf28fb643f67ef9945ecef9b18e4c5cb131285f9a662072a50ca0a9cd1130d15cb3489db931cbfe0742e8a8a5a9bc9e552f56d148da3bd92c28ee844a964c65ee6649f24142b774537d3961543b1684c0fab3;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hdbb9f2379e32af68ce7481e63c07147fb91216e1a8311a435b21eea89d35c5957d187fa08236f24afde36c3eacbe7e088338638593b939340154cb6c981f767d5c8037cacfc78ea788ebf27b96512a57a43fbd410;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h24eff7433fb090577c5046f9ee10afc5f331e30afbe60cb4a7b5840087dbebc48ddf9676c38803f30f531f486ecbee1d413534cc29de13812a49928eb97d75da0820ea65ae1ee2623304258fd937a9a6af11866cf;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h69f6eca48ea952dd03f30cca94d31402b440a182751f1f584d6a36782a2e776eb71e468bbaeed5743e7440b2c3264e903511e8acca3fe9efdaf4874d35b17eb79d8bb72a19306add4ee1ad01cf4c3977621274df3;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb61f27b1648f04be57918ff68080d5aeebd9fb257dd62bda2f882717b559cc5d5bd4261756b8bc9244e178362feb9b4ec3a75d27f63680ff1c6bedbb15d2ddde04fbb9cacd0540821ebf848621b26f8600cbdcd75;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8ee8164147a2e4d0df0eba60a031e04104222f2f712afb52d28d69c1c1db825b71967d922508774d5c2a9f827f5d8e0a1a807454c27fa01cb4f0d6bc285700c60751ad6d5f76397ea45544e6cbf4862ae9892e332;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf9d56eb6bf6ddc75681af9e1e5e8cf954f29a49a7005ef27dcda77bb339304e08f1cf9833eab19b91ceb4cbd8e8b9d11052ab662a18c8ac7133217caec0ff61a647f7e633c262682f503dabe224f37d0f5d9672e9;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd0a9e90c57be35d4ea5bca4a33094f13be49d5240222de07f65f6c7faabd9740ce128a20eb56d837f855b18bc9fc29962cf8e62f03daf2cd061e07d283682d6367a78d0bb2cae7b4ee5527e8dd13bc7ca9a1b1ed3;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h36df3a28a33488c72648525860651f500663850ade6351fc66cc640719551086b51b98d26c9ef070ab5f09c2838268d18408b25bb9c72e6f5e95984860e4a8c69bbc86462f874f2b6486d62f5a86c05ecc97f8d9f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h48c63f9a32b58cd3cc29fdb9f07ff1612c636bc1c5f4964695b680143af0a92201e9b7039cd3addf172cb297720e34e4d0d87fe68d87d1c54fa6f07889e4e0d956457379244545b716931af0cda15eb472b88229d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h41ab1526acad11b7997c04d7619a2fb6107a78fd2d1443b4ccac1faf64c29526f42297ddc989c71cb3cb245a63f14ee8f6d540ae30a9f86396d6351f5fae73b5c0a47053bd938e2e46dc5a945ec38bc00b5511e37;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3b0a0af65b3180a2f779d98a7fed97220abb6acf7e1d38b81dc86c14138cba874111bd557e878507a72f88e4099f539405d47aec05dbce5e78b90d2608824bd0e6c3c769ee66084b9ba14dfad91e574c7a153c4ff;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9648d41167d29c845f6d3b704cac241a0eaade95f2d46f6079107f671b8940de76eee66c1ee0c6635f57bf052d53e7d9e244f7cb5301dee4a3560ccf6e5ece34c068978ce49a1d11af0f6ea5e14ccb24f358e2389;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'heca752119112dabb5379be25400e6a6bec83942b59eb74aa8b3cdb5faa965389a25bb66a03c0182f441a98803272a7368fef9460b0afed0ad977d10f70f9d0223f42fa632ba766608cad9a4e8a49eeeed7fd2180f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5c9418e65781c3f03229bffb97b23635f159dd5543a3daad63438a2c9f1aaa281604b5d59d80a1d4385fa3d912080bd214f4161e7ca33503b171f4b5346e51574aaf02f0acd686e10d2fe1b8d64d49f6a3e368005;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5d1e99708e696f3589b2ea9a332797c2d70d135e52f0112d59372f1a2ce5be3c5e29de78261a2c42160ff37a92153635afd4ee8af33169ee62ec7051342ba165b66109f38c4e86c60cdb3b48ada6a495cc04b0644;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he7efea9756a52b946ffcd1944bbb082ba76532ffc634ae672fbf4668975eec89609eafbd13669ae269b3f6172a568833e2706003b0b66fceb248af872df8619afe73d838fe9ec00f28852aa7aba0d906164db1580;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2fb9a9a4cd325a45ebf5a51c16d3a493fa554362112dfaba9270d392016b48c90664bbcbcb223a67c24a44c7f1db0f751c5fa9def5e2b46495e97abd4a710c2e136c72d1177cb01481c585e861ee6637464ed25ec;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2ca07a43e880e307d6d6236d9b1204dc28a8706a7f7eae3454444bdc34228837481465c942660805c0309eddac56eebfbcb60c3320c375fc9d9c7f357458670c980ff77c832f542cd6a137d9c7abaaec925107c5b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he017c53418c2b1451838a2c7af37969f80283204ce43d47777f62eec5320ebe6a74f6bf803f725605d005139806e19453a252b42040c2a08270bb2a38e27451fcd4c6b219a57156fe3fbf2216ece470bdd7f037f4;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h11e4621c385db15d91382d15b05d58b3dd91081440179a4789a43b85e19627d6887d5c2e279228fb9a5523dcc4592113f3c73436b97855ab37ab0842b97bef49572b6485879927c30533f9985bd3928ee011aa9;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd9c80821ab19904d6204b0703373b345403b3cb1b7feaa8c7a53df01711f64b04c3ddb24f819569a2dcf8865362ff5b4d70b4512faea8397f9a41cc48eb94f5cc606b9f5ca48f198d90e2c7c2d35dcd746628b459;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hcfd8ec498b7839da6230a4d86cb75ad83e45863f37cefc84d445802d92dafc41a326d39e8d5685b1b468c45bf3e050618c854c6cc9e6951852315b4a2cf62392b3a9ecd707c43f736d2205bdae2d9274e38839e15;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hac5dfc973655f850acf1f1b910c718b509d8ace44be9cda376d26e850727dec97713c91befd87cd235c1f2c48669e31b0b297309464c5ad993acf43572b7d4fe8fbc9b5105b34040ffafb6b308e56eb203a9881ec;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hee150bd5c78b31ac6f6f36372d69ec59b37fa2b1ae9fca68fe6b6a4fd00fa874866e7a0bd1a960ec87aed04d62beb5ff6ab4fc2a03c7acbddff881ba316bf9f581377c46b34115da0d9e48eeebf176764eb905436;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfdf187eb2b45bd17bac15c99991690029b1cc2f41420bbf41953cf045d7c2232e5315791e1923c59ad3f8df54406bbe5adfacd41f4e9dbb19cfec8214de5d074733fb9edba63d3f5589bb2bb5f7d72a5db43d6de6;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc4ffae86797254c0f6761d3b96faa98b96c717fa2cd96ffa298b8c285e72f26f1bba9a43a7d68028ccaeee396e22ab53ccd11ac0f0c5b6b56b22892ccf3c8bcf37716f3c08528e3b3e696c328eaf6b602bba84653;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hdbb5417c69cb92eaa816e81b0934bacf2903a90df7977934bd783129f785b8591adf7bbc70edb317ed3fd919774c5255a03a5de82c29b9bfbd6154ff4534b2d66679bbe84c884dce977cf8e36a8faaf4a3642a34d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h93b611d552d1126874790c22757ec22c48e071f38744b73659a9a8f15684dc4f18083a4b742e3b461a59d332ff32c14ce9c1a2fd0441ebecfa93d9d302f5fe6d8ac88aa601fbd16bbdc37979c9260e3be3c0fd4bf;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3a7b2566559bb326500d2d02178fbeaba9e9243b9959b63ea69ca8a1f565cac1c8039d42b5796839f9f0367d262242211cdac4dfcb82c0df58374e22edb893cc2436a6298d2a6e58d8cee81abeba4427da9aef45d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfed21ac76760b51584bfcdd40f7f9957c2444cce081740ee114518fc7fda05513d5ed76eaa52e9240baf8075eac10d8fa6e0bb5f4b289444860dd512fa12d3a3155c5db0e39015bd0c3673a1ca46a904f5bb1f3cc;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfc3a115505b4812ad859a13dde00fd0eebcfeeec39f92f6be78b7360d47a2da47fe95e115b90eae16c0bd904c5b0deb0b986b884e5abf0fd1c4c6aaf8a620a6d6c3ddc14e59f6b50a4707ebb3f46343d9138fe96;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4225e2bdca4c8613e52d4d0aba2e8bee1b5d2476a4bef00040e83a0a8f76fdabc7b6e0d4d9e7fbc8d432040ba56ee9ed5c7d501d2e9a7b43c6ae0012559208c308e13a27e32bec9c7aa8638d85dde6dff3f4624b5;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf68f61bb533b14477dcb8a23e588dba4c2c61ad6f55fe258385bca2bdb366b8075324392022011ad8c4d168a7bd3b315ec3ffadcb19519008f341fe2a701b72d165db6fd4afea8c28e5a62bc1a899f764168d9628;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2f5a798b860c5e6184b5c13f6a9f41e0a37977aaef693bedac802d2268fa8f155d1d8ea164f347b8e55cfb006b1044b31a53a5700bccb3aa866a43855ee3c220f8197ab825d15043494172dcf6ba4e30f9331832;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h60b9894e998138ab34dbecf00b146cfa18f23116d8b110769a8daff8b7df566e48c820401587e966e13be324659cd4ca9ecbab4d329fd07c7f0b50d1c3477a09073c6d8d1fff82f4b2603102757cf02396c5fa8f9;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf1a95cb84abb626ce39996344440bcdc07fb6c45aed0fe2a3b93660cdebd6b991d31adf4b32985249f1425ec093a27523880eab3b17d4007d2cdd12cb1f1637830246388e077da075ff630d1bfd5e863a7fb90825;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4c12cbd2332147de97dfbc03d4cdd7b2b946a0cca96b82cfd5668b68a7763be92d6dcba3d3ae6f25cfb4a5f9d3b3cec83810853b227b816ae9e4e0375272480c5caf85fb215eef8cf240ad8db5a4d56f844cdd457;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf957a8f6fe747235c7ecb4dcaeff0aa73caaceb9b35b349eb254866d10861149cd801f4bfea97ac551c1fca71a3023f0c73ca226440a33b970fd32b15aca73a6968fff8fb4d856c44ec7bf44eaeab9a5c9e1f985c;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd4434927299df4ef9cbafc24d268aca2369da6f5ad6a9292b8a7337e5e48ac0d7f53788959f3135302c592f1d4b0edb00c20e0882d046ff3a42f5f5b282f28dc711a05eccba20ba9fc665330fbd5411727dae7dff;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha3af6122faeb2a280b8b39586f40a32345021e73b59b598f382d5a193ec3257e602fde0c09721d2787c5bb8259783aac7c95e21c2dac0b3bd6a36a3ca3631465da9fd90fec6b0d9878f2198afc82cf2a0fbee9c26;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd58837236ac2b341502059046997fa9c0c33c63a7a6afcfe0501537939cf9ea7ceb3748481461cb2e97751f9f39ea21628c587a7ce1895c688af4a2ff758b1edf2839d806816513b3155072ebe318d694cd9f4eab;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1ce0d390238a3ca8c4bb0d3a1054268af0f262d49e5fce82b545f879e69a29a79fefe76a6f70523ed91677aee2390b2fcd3569c69e4a03121c3a42c3b3e1cf80c5a746e714d0cb2d9c124efa2c4d368eacb7028ec;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb397e617e07db820768e2b0639b449b0a051ba0837ed0fd67c3e09bc8471ae1d935ade304680265919716e9aada65c342167342175cc588c646b7607b003d3f709f860a6723ef10049b496d2367232534fd544401;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h77ee416fd7bd00990ee09378a68848117c95870382500dc7dde86dc13271e3379f02f89b62805c91c72f38adf3a75ffa6058475614f4112e5313732a5b138040d4bd4418db901d2130e980b0165fe61a5e0416891;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h34a6ccf387fbdb8a68f0dd7e7cef1271b03011926712012aac129879a7a684b8dacf79397657688bb62eabec28d5957c366435800ae506e1633124576472edc74da47b89d377a16afed638cedb187368d92542c2a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd2536821ee0bf492784216874870f7670cbbe75b45ddcf80f23e6ba66ed8bdcf8c9ec93c0fa2899eb2080a721af2ca7ce8d87216e0da8ab051f7242154067d08ed027590e770c4085541143cb1887e1a0c57f32b2;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h44ce8a9aaa8c6aeef0852502c8a49a1937095dc5940f2ab683114aeafe824b50b8bbc9da2d3886397f50944b6e44a3d1d03c9d175fb9235415671676a1480a28d3d8fa0ba56f33c8773bb63cddf2b2028b724b2a6;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h496eaefea13a1cda348a99f6628d42cbf1c77ec0fc2b5fe78fba6ac3210713bfe7ded9d00ad048f25b1e7a6913904e714fd42e2a993eb77902eb66f3918354a1d19e20a2222eba27887849a1acdb230f19f098996;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2be429dbdf16578cc80c6b8db89b00d0ca9afb781ae9f471d348d699efdc4850f4b8a1666a8eff8476e74d7d174343030b0f9e9bb391661ea94fb6909e651947ef4f52f16f13c2175736544caf3bad949448e9235;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2f1e37d61b40f20f144a022e4ed6081fac392301c54c7786ea9d14e2771d44e2a4b2bb5d8506f1a849d60204f721257ef8dc3bcd6346a1aae973135289c3fdc11fddd99ea16bf06098f16313c37c4e483573d01d9;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hde664f6c524e9e548629b8c5bcc5299b9dee87723bee6915ab42be92ea537c080e671ab7a2af84f849c482df830cefe60fb6c5b63754d4eb21fe146e62897ad8eec3d72a209618ee40c29f5b9b5f81619b98c1d08;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8021617333c88740949655f540ff17d68b43cf59f78078acf3f2c70ca58cb75f303df5ae08b338300570217f6848b0dae2b056c4d13d7473e75c58eac1b2a2c6e633904ba31f5ab92c86392e0b74e4aeead0d624c;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8fd34f45c8d75da83433ed59c789b260bc8c63a0c90d7c58ce6b5b2dbe7a5ce3a172db6ef90192c0e41190006e7c326c031d4ec7212ec6becba66f85e277c1f5e1cce0febc4340340206757561b6a33779ada3e61;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd1820c7f5d6a4a3dcb579f9879e219741c30e843bf40edf8d5e422c8f4cec45159ec1a3798360323575d826c7c30f7b70ddfa8283d12e7c205390a0449d586afbba00b2ca604535aeeae58a8b0144ddab951aab33;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5a42803e564e422b92ee2af34e72fbcc855d7a9f104a3fb82989fef21ee8bb4563a0b680a7915193de51b2541a8aa80d9a5194bee9d2521ffc6757311d517834e16aeda43b9fbf6de378470c9d598a345460ce5bd;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbe27fdbdf325d8249b2a2073315f9287578f45aa8bcd69743147c17eb51eb2a4f8b24c8a7109b2ef3bc34317d3ec2e6ae96018ebb75d948a1a4506355c4d1304b6414e6ba220625cfe0abf8d5b651455f52a7b8fa;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h81272ad6b2e6a639545a7922ff237cb3f0930cc9e712f57205fc494f5564f67b8cd1df474476913b56e4543394dc0cf017f3d3c4504c0f426b7ef4eea50566296e4349f66d63e7e8d763c875e9b049f206c85fb9e;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4dbbb43344927f8901df9f524d14bc32aee23d586caaee7db72768636e5c3c86e518297c639e97d13c486c4c886e5169ad43c9863f50fb7f02114ca753a45ef04c699468bdfc0b85889b8f7fcb7385a6df44024cb;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h11ec04877493df8c75e672b7dd27e69ed4b41521edc9ffce0c730d4831d32a2f343a87f727af84bfbbd8b235b30973c3ebe6cd7189a88d5f798c5d9d1faf22a3e0756446f3dc4b208f7a80b7d0ec71f392311a88b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6edbca2e2fe1642829cbe24233c47ef92bdf0361b24d96a1c1278b598c526647e96201aa17f75cb256e12b801772e1d67320d9f80e03c54cd9a71024be359479b1f92bb9fa573de9d8b9d72b602bd51d59b990edb;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h29f1d002dfea0f46a9968f2e0b334c8dd2e0e35e3bc51eb8c352771b397d4cb257f8c6bda806e03f2875dc0aafec8274922ba409278209b658bddcb8a6cff8d7565a36247833c00208f9b89a8515f2f4cfd7a73bc;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc5c8f7fc38fbe69915246f9b11ca148303baea939e4d68d766ce0b5e2f0bb979065a2be486ded5a8061eb01ffd73f513403288850678bf56198610406f0af85800c62283812f651ce7eb7e6387a100954cf055fc7;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hab21eefa17100621b6842224be978e78a6c402dd9940bbad269b5b4a2877d21ec1ed6916194a640a933f8b3fe83a3210ee2440bbcc0743ea544969634818f2595b4d432d57c856c32012b5638a94719bd64f15afd;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hed026e0c1c36459661eed8665bf876db7f182df359cf45498a44a3edb104672b22ae912f5ceda7d3825978594901f4f821450b1cd04cb585f1ab24f529c581887dc2dafc06949870a8b33e547644cefa800365117;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h204017f7278971f99286194d85d9286f8ca334183d1541c30c46bbbbda92ed4f888fda8f38adc8d6c4603f756438c990af3f6f31a7577c950a3b65d66a169c1016e49c195ffc587af6caf4307d3a247da168d32aa;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha710efb3fc8d9e2d594eb7fedda03d684ed807ff0d2d57a0e5fdcf84058ab912aabb56df5a41b1a94d4ab69fb1161cd15e45d970398b109bb25cc3055c4ea58b1dcefa9b52d2aa662e7687cae14a8164a9d8681d1;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'haf79ee7de023329378ef174fa2819e7e02636a63001860f52f7ac9ceaa7ad8971b8d9842e63a725b547106e552e364dbf607d7dda18bf8f8ae95084375f1d8a2c54ef8eb0d2511d76f9cfdf4b5c69ca93c812646c;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4e268919345ae76f126a80239a11ebcac9cfed97308570f6d0139d6c3633397a8856b951ce73dbc93dcc4d71e28f153dafeaaf53f58a89734678f8f35675d26de8f1271b1c199085b71f8615cab977f704357daab;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he1ef04364ad8eb5d1ab1a41fc747d4e053021d466605335963d921e5845de42d62cbc47ee82989ef13c528ecac495369da18cd58b7847c3cc11b28df0baaaec4478623c654aa6e9d2dbae5e69e323f2169a63d09d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha6dbb01664832a122da9f1d228882a85b21a946054886398cf71cdb30203b5227a5c0ab38d8b1e33319a2656132fa15818f0d1abfd20eaa815a653d57d84ee2471df6892eb153ee3bf9b8dd1a9034ea5622f0461;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4b5140637f19cf26a02522bc38e772269f873e6500d72c9a74f3fb48ed38cbf2c9c57fdefaefe8724f03b111191f41b275b13dca903ba8be05e6872dfea5847373674f8fe5be8f821a128644df045dab75eb9f1c5;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hac64a00dd97a4d5e1594a93f91b87286d3967cf5a1b0c470a8c3540ea9f234c63925957b55a1233b3750b84e8a24845cb1b760aad320da774fa0ebd58d63135448600567c206a37634cacd06043a55b8c24cd4847;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hde09a049af946095a8a73bbadf0c38250e12c48b39ad13d9ffa52fd23e7559e968fdcd7ccf874a715d52b09e2cb7b42cd03f205c5f25a8e8d884addb65b68c5d82552e061c1cbf7170059afe0a9e8d62e80dbf270;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5d46fa560c899d5ac7648c32c84976b5642f920dc39c6b865d9566ee86578dd31d8d423fd7c55033d92daeb3ed04157b9d5d91beead31d59ce66a7f8ac6b7ef9fdbf98dd02ac92bb16932d0dc3e5b1b9a07751f43;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h71dc8e25ae6c730d5a18ff207783da77d2042825c6a9af74381de26543d2bfac2fc66d257949eb276d3420bd29f9132a0a7a01dfe77eb2e8b72364f261073db366a3aa850b7bf544760fffeeda03f47a4f25c5085;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h66e38f10510e3db761f86d2accdfa39e88177c7a629dbe4af3272cfc770e2e7a76889314f726c15efc7e3416da47e04ee05bd26f231a48281aa1a16be541b813c650941a775eeefbf16ebdb5fca0ed4c80ba0c164;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h69c23dc05d5674a5a83dc122fe1a0534469648295a19bd190f54d0d464641d4756bcff45bce0392035a377a7dfc6dce7500184d821fcadcbd50e35c899e2a9de2182db66316b829416d200d4d7d7a776a4d49c08;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc93788944b0482aaa4b6555b41930938f537300e0015a4c45662c839add7634f23c110b731863f455e0be2b1c2c1aa8783205a1c94010b262fb6884c59f91668b654b75230177ba6355ec1014eb2e221791237eae;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8d50e06d38426e06318eb83d5a16dc8c6389f9fc08ad18814013aa888338a2861d75a092bcbc79a02bd5797f7c87b12da0fe64ffe5ff7935c88bc9df588c5ca2900acc7704bf0b6912c6f6e1436994fbe306611e5;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hde52d8cdc3c51ef7d7d2663b91759aaf7b9fb85e72c871cfd053ff1dceadd98ef3b2009402caed3c35b5392f1469a666edd6f3bd9c09dd30b775f47031bf1a1fed703163b81c335b7c8ae051aaee701d568e9ba20;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h473bf17758d2aa91b251817c7b1f50f558acc7e9a0ac1775fa9c1667e332a01ef5ec5ee816d9d50eb7852d1715c180f49d9f22ade3404fbae3e06889722f1844b564fc4318957c759d99200c1053ad2166ba184c1;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h97c7f020039bcc1f84c8644fe350c7e9d7b747876a94f068f59c92b8027c5a882647bf9d5889c0b578444d508861cd140a778a6d8a5ab6a3d5e60bb184c6407b615803986901b409341ef60b8aebb853beb429a13;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8d66726c94fd696151b8f423c2398389507ba3561961b8af5e1920baad3883e36b571a9fee3f983cc3d35ec49c4b674fab0d2e14b029300bbd1eb78f8d58c17988a724d1fa54241771d99155a2614980c5bbc2296;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'habe6aafa50a5468b1e2c7c62ad8edf78b7f099d8505d3dfb7954a044943abe4f3004c7c6fb4a43f5a580f35d915ded61b53811a0d0a93e2d98288e20c85c44b74fe024ffbc6ac5ea0f82333d194b97ec1674e51ed;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h850d6138d7ed24c9e5d52a3d93ef1902e5e720620816172742130e3cf24f2daef4966d3f019205a821c36eac72c14e00512f529f3ff88bc5b0a1cba73f4be53f9d9f0fd856cd337fe51cf74b3fcb3e57570101ebb;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9a86b08317c5bca6db6a8c100149fb8d5aed5a752cb9da944865bdb2ba02520ae75c21f63aaf6cbc931b28f6a3d2863f07508ab1ae8ba53fcc70fb89be7f830f09df56175fdb76ceb0ba2c95848ed98b666051983;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha70eb3f13e31d9af7157283fb58e324511663b7d9328f8d0dace548a1da5900efd2b67bb490cfec2918aedf1f0846e29a99e340c4b569889f81541d187b92858376839b1ae7d665aa08af6d62673756b14e4e29;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7edbdbef7d54a3934d658c77113eed4c9152d66aa7a6034630fe740e3d1de6e030652acc2ea02dc7cd43df711bff7d1d925a67866057955d20ebe369dd0b4603788fd40526183f0d01d1efad3363fc830552ad82a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4480507ab428813000ea74032f5b0fc1aaafde0ed54bc9cdd201ff0fe60269547666f808a38241e91c6ae544362da7cb411e57a03ecda41b72fce673463a8807dd4c8f889e1a6adce39dca3861bc8f32da5cbd46a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h88921c62f01db0d174b48c9b3c0e114968c1ce474beac3bd3fe80a7462ccf1f6d99d15a0dbc37b9f9ae898ae38a9b2cd42bcece0306d660b079020e236823117b3bada2a59942dddb93f16f66418056354a031d54;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h47c8ec8a479fd7440dd03370b40f45ca96697a5ec4953f6380b3f47e800010631684b2000311f857a6ddf4eb6fe1177459078baa850048298064f4ae1f1b66a881f7573b4a6844bc7e71d751ca19ff67e35f94d07;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h47fd93f0d96aef6e911bd4f09bde5082af69dc6b8a03d846f39643af9c6c4adc4af4f47f0c347e56e6383fdd3ed0b34de173c53b065e131898d18a291eac2211e5e975c85a6e7a2830059e842f7486b4da4671276;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h409621a47c6e9f903acb37f31695946352a411756256716892659c475678bd7bb8a4a321cf6b1fad3d097c6d0f59b58e494bb95efd74c3f7336c978cf3e9f44ebedb19613055232a200e70b8d138608476823f10f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6da0f1c022988fd091fb863322c607d0cb28f415e86dc8254572b8607d6bfb4135749b79990e11369b5db0deb5d17d3e2d6544415c91c2fbbf5e8a77fcc076768447c42a6c9388747508310d87f59e7b3a773c02d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb185413ecd99abc173166000446568c8a1e36220bba3340084a10a3f0575d41f0fc7fcc10d4a2eee351fe281b78a52454f145d3b2245af6ff6d625c15bcb33272267856f0a6e1f16861dd5c7c5cbd3525a2eb1a38;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha2088bd63f630486b7f1556e7c77d3c74564b3b286b16b2316b1a1f3348dab9a448494c18d3e09938cad8ef732932518f12b067df3f8d27747aded00cb4fe477a18aad7fe22b3db30f509b80019a731ae9421f508;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h152a0c05514aae712bca4f217aa8a0bdf710665c5820b20722e4096353e370fc28f13863e3049187d7f59b50209b8eb0cd876d66333d91400655604eb565574610562ac0eb8803bb9369854ebeb03e3d8cc3c7b35;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha351396ea466c847dca38818a05a89b23c8de2282b2cb053d2e6f05412a63e23086197be27dcfd64b4087ae8e1329cda8ec4b2389dc2077a5b14f431a3fb187de6ed7cd852b8ce13f2246a3ce63cd791f2a70f45;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h61b8da7684f1eb3d167541a6cfd8a062c13c45c94472f5292851f59700e2770ffe2a0a85ff55e107957d740ccf0872587eaaf0ba159c11a231fd828f5720aa372cba629df6d88527c75e450b306e66b2af454bad2;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc302121cd0c3394ab0c36a9ad3bdd70265f40bad4768b6a215d9b0bb8695d235b14cb87855bc762bb4d8011631f1b7ed68f1cdce12c8d773a383339e0414be90049caaba3d18aba36b5347df3d2bafa752be92354;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hda7f597d3d3954bf79e90f40f81e8928065483423b61785dee538adadabc359beef6d2c28efdef75fbcc976e129e06644fca68d38ccc75c38073ebda18eaaa4013dfa33051fb718a73d13fdda42729d50af3d453d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb2e5748d9d266a7453b45b8c8adbc9ad9e7cfd6477c22a20c4a5c9582f54b4448ce0ca2fe4fd980b6d0c7a57791e472797f24da4559ec7a455942033a2773b9dd0d430dcf67dcbb56a2eee1ea20890b23e062c406;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he0e3af8ecabddd5c1a976a71270e081861a39985600b05cb7c35a71cf39271e06d94753c1d1f0a7b0109089630bdc58f19294101817ba96cc6f2b3ce227d8dbf8bc7090b9a0be9e6c4b169a5b3c6abecffa79747a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfdedf6994b4686acca5a222344ef7765e9e08a96733dc78019f5cb7a28127bb5d30b7e1d38fb4312a67753e2b2f15f0f3eb887ae0f7ed1ad51fe0d37a5ec40d682790225b299145c9fd707cb686407d3d6283575a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'haec596e73fc54f7e99a8c919df68ed2f8fe6a80a0126aa7456e55b892ef5c7322aad3897bb00c2e1797fb9c36f4aa4cab97fd4d489f60c49e82f04c03cbc04807a37f1ab82829806199541164b2feabd9ec060ce8;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9cc9d91a06130cbbf2fa6319199f92a43250ccdfe5ce46b4f5a2f6f26f9ae3f795270561e4aa1e8a54d0cccb9d77a373e4eee772ff232ad70e12ff0876e5f890d7111b7aa3136e6bb4884658de57a80630a24886b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he0ec40564430eea552ab43799c14c798f857a991abe009866dd5f3cfe36500ec26f5e5ad3b747aa8bf7b23e3463bf3f1b244c759370f8776b901b34f8534f922db667dbb664f814f2a667ad129939fcdafef143c2;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h72580057c94ff215976f8790086548d73c4da8bd224a3927584a9d0f559e217eccf1a87fb36ce1805f4d300422d72eec082ed27e348c37cc87ebbcc67f193fe48aa893f13ab7545fbd84a4ca02de6ecb679c80754;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hee801ef7d8e9f7fcc063fbf718b7b301dabdaa40491e255dfff11d8f5bdff863aa5a71fdc9ebc230d7922881ffc002cb4503c6205324a535e0b845f5c762c4fc70c7798761fdb7b9198d10657b8299a914aa7f71a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h758dc51ce38ecd09cffe84d59e05746187480388ce50b2a493950d3cd27e1ecec21620b0d81e74ddb0dcd7886a20152bb49e8a6e4722e15cb91a1f7d2e5eadea0e53a7f7d948adff36c464e822569bc64d8bc850d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h159a4eca0d8da3f0c71cd675f2eb39dd86ea1edd6b1dc46ca7d5b54dcc67276102f7ab5b9b02c54a3533dbb4f50405f84449f83a3b9ef6ba4c85df77f911a18896bd496289143e447df4a0fcdccfe2f9d349345cf;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hdf995a343057fb585014f7d670ea9495276368742cb4907a6a0f7910783cdb464ae4eb2b34b4fb117e294a46b91a1f9cb333bb9897c22a92300b441214e1431de69bdaf8f09364325fac1695cac42c9e8f34cf63d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h94b4b2e83eb732db2c4e38f4ebf2094823da948749918fcd3617db36baca361d256119a60f4bff2ef3ca1d559266d553339104e4d4ebd3f36490cb6c4f04adbf9dbf99971b1a01078ee2601b45fe73042e41ec9c5;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h69c33553377b129636f747931c4a9649c552e67941161c20f87d46bacf5ce7b788b75d36adcea5209ea39555d09a0188f49e8082ebc1b5152122ebb21935ccc965eaee3ab8d980109fae0ab8c25fe25deee23d999;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hcd72f34e40e775573428b2217c4aa8c03aab9b5c6107f68847b0f70235b8067522d79cf7c9cb1f44da88664b61549d3ed78ec9a8c75406918ff0b5525bb3cecf3b8f3e3c952b2ba778aa48f1ad35a1efcca6fd94e;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h922b104cbff07ed8a27d0b38b0f2a3a222923d8643277f0772e261062513ef0a2ddfabd4bed72dcb1c01994082d2cfb6c26257f77247ec8ae63ffddb4e669157cf162cc0d36b36769675da5193164dc4513c8feac;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6ce318c183693331c6ad1a3ca1a25e680d7d09be1618c8052ff969cb7bd87ddbf38219645199cb6918aa4c6296d5021cfb478c9939d24190b7fe7d586d35c9513709aa5a9b6a7b774a03c61136f723baca5fa90f5;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hcff20bf4a69fc793d3c2c99fb5a99195207c03bb86e32295cdfdb8390fb2448af5a62d8800e59f4f8da229db7b3905d555a36f83f8db1ece5db246d5bc5327ad562d43d1a8cfbe82931fc5676719c55c300768035;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h301fd6b331aca9646ae5057ddcef7253d836d81f5b565c10739c3e7477ddc60bbdd0bedd64dd45696feb186ff7f4ec2ccdb15ceff9a959283e360ebc86ff4566d6738658417a8518c56abcc7d75afa306d934af98;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h438a7d3fe97cdfaa87079fff955e9c8d9bfc1a75773a4d38cf5200993fef8c16ad4f6396037045d672add9d87d0e3ff2eaf6534bf5163adb2eea2961bf10be73d3347746cff6f6f6317e78da4c06060f48f380276;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h260d6ef3170cb66e11581b06a60d013ae0f6d49d92ead2e10ea5560bf34433634e2408df6750eea3b2a2363305c985ae3fe07be6ffd591cc1d69a4d66333663da6c57109480134d0fbe59b188874be0d909a1b9e2;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc466dbec608e48bff2f8150ce454f84112872f78dd2d0171c2c3cb9336b1a7146bdb9987ccc99e1b712a62696071e5110d1f6c4193994ef47fe81102a9a13d904dc953a69cf498c5cb11fd277a4d702dbea4b3ca6;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h66583df39fd8b68cb28776da0442b167f1d8c8050a58d8125cf3a812926305edc036e9d4e1f58b1841c283a257b745d778c70bab810c6330bd07e61eb5aa4277b067e6d176e1f70995c6fc3dc8011ee4d9e394da8;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h978c71beac72279517c7faa0544e2bcf941ddadac5c1cadcaf7cc5f15788ec993215d2766dbe41f3c7cf0cbe841caf8016d5d971aba628aaa5f5c3e3c59fd6945f00cc6ac131ab259f3c03fe6621d9d55d4c5777d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6872547cb8c8b36c622df4a984bec22472bbfba334d046b8b26b6510270d73b261bf395e5e39539b92b4e5d2257b8b8fcb24d68536ea43946b1d5e96397d28ac98746c67aa7e60bcb706b469457e2612bf633af36;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he7439ef20230f6cbf94523d81c522b546b4364167183fb3eb20d05a0794e1e58ffe47a1c27a1b453bd902736bab6bb9596ae37a0ea52d23abbd4ec5604444fe0f4ccea3accf681304ce413da618658422d8e1e37;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h838ea1a07de8f28116cf3b1858d2017245482129d45abe503d252aa499d9dbe0da610107fe06b2b024ba188c138a2347c7609e0ec7a6d879c2ed71c88f8ac38cdb9c34712eabda9452b290ef3af0c890acc433046;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc8e7263ae683afd5e95266a718411988811b45b1421e93e275ff0aa5387f6cd8ab405bed671a38246be37ec7b01115680a115033c01dc63ffc604917f7ab54f557216331dedaaa58cb849392a5cdb8c82c3e7a764;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbca360eeb84b301aa20ef41967345f2794814d535e798f3f40bfacc154b61d54956745ef53e622e7a0e6219ed5405fb68a2095e8cd5a237e19ed2107cd0add30cf698968b37209cc0c50b16d28b51f74e8b4e77d3;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd42433847ef3a258008b1fec9730fd47fef80805e30b49bd5384b374cc2cec382f7873578a6854c3ee080f2ba0952c039a3a4f4fac55be45469dfacb7ff80464a267f529ad77fe7d4310c6fc258a4710c97eb9e00;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb2cae592355ee50c948cfa568330f578100fa0083cf00c0720736c67b06d8a7d70dea2eafa9b88d7e0dd9ba0c77031a24b7bd22e2a1856ce6cd6384d6b4b255748c0deccd4837f79bb908caf2619fbd8e57a77dcc;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf00368c320c678cc4c797f9f79e4483e575d0b360f48404bd0d5fa16136e60ca039e97d765c4b9b9f5f5abb4ff20b3e61ad76472e8f960e3260d044f5fc61b87131fab7b46a41114268df7cc2ce3b2360ae8edc6e;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf6f54c4f275f31a9e7ccbd981d95ae096106e5fa2bb6764a4e05c9530158a351dc3c7297e5c5f3fadf603280921316c68946a29c92a5d13535390be9f6948330833f5f1ea935f2e2884001cec4f2c86017f123f23;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2b30abd056507e8a9a702c09466ee3a59363f91f35fe1bc849659a5b3d765995e62b62507ac784c675984169db24dcea6247e59aca472b26b3fbbed81f74c351857afa4e05786c21482be2e375d2d422ce42432cc;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4ac62991e5d6207ca5e368442f80187935391b15570935cf73e6e3b98e21790112158d810772012975006a8f681bc1fad4c4d2fce580972b95f8f2d9f1d10b8f73d926bfa595adafbe919fb52bdadbc064eb7d10a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb2eb6c619315a828b909db7448f9fdca77360b9346d15e9ac61fab3c1cc4786039e4aa1fb70ad205925a01553f2f916748bfc4902bbd4e2c99aeb7cbcc42d630f5eac790916153152aee3630154bf1f8c6461cdf8;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd4d96715fc571950b37b392daa874e5a3ca9fc157a3a5cceaca6528e18b1c67a5858e7e5b39dcdd13ac8b915ec8583b4397192c403a2704fa8b33ff7d0bc89727ba6c202889f6999c305400d5f7be7ab2bf19eef0;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h348038b4c4682d827b0302a242e4eca095549d0fe68c7e761133c5e275696ab797d29572a33c213f360e9f14fb49a2619c4a2337955926d6dc92e5f2b0f71dcbf5db262fa0b5df3ed2f5f41e8997ce529b330bd1e;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h96f1b7c45ce6d9b633d74768d07d542a4ef6d8ca11cfe4eed809667c9502f0238458db07a136ecba704556b4d1fd9de0de67a501d7885afae33dd61e135a932dc8017d2c73a25a238143fe1ce1555294d7d9642aa;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h49e75eb0be3936b1732021b1e691403ce3c5766e0a3c743c900f4548e02a28e6b994e0b07adcffd0718c3728601be9222eea2a3da5a0d13605671754cb23dbc5040907db21369488c79ab216a449509e0bb80530;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7df15888acad57d2914431c13335da113a4e87237953c7b0f9609a8f9c5d44326c17a792a11ebd2ed000684e107dfa80aed0e8ac013251ba976cf74d7175cd46cc312b228e21d2f6681bfda8fb742e6078245c877;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hba6be9e96d3470637bb9b36fe58082ae2f1c6a61619e423df98e8c8b5eece745b5f3ac4511cb8fd539aa874ff0b855d145000a4409a6c7c91e74755e2d78e69117a85806ed5ae9e7fe2c6b9e448d8329fc67576fb;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5ed599f2e7f49b0b5d204968d50dc2a44dc7f26acf31708cb84a26c4a4f4f138c5bb6f49b8cb34c57777fc0b657d749e5a6fd284fd8cfc25ec5f0207dcec483f91f998038e2a391edb18cc591e80e27f81b943ba5;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h451a5f4337f9c1c3521928497f92ddf842a9240922d393860262ad97fecd944c68fc98ad20f034b1be77e3da5b5a9c96c051897e6a6d027d945d22371ffe28001e706b23eb4b77996785941b167dbd94a8556e313;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8edc243004ea81fbd48b0bd3f373e96c9b416a411cf707eb1fe1a2b167639593a5d80e82590a5cc2089276e713752af28bab58a1294a22b45a6dad90520b197ffae38c9c0e10e3fead2bc16575e443892249f32a3;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h22e408889e338dd50842485f104551307b373ea40cc0f09aeb05d8dea661825951c0510eae8a17a425e2b6f7d010e5f29bd3a812662cf18c69f6b61c229efa173d557921c78b2ec05e8884bde9c52ef76cac821ea;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h28cab549916e76836a3338d243b7c0867ec9379bc00d35e241a88e4cbbd9233354903c9a0d5859c00b2e2cdd5ca3d3c911af69d65dfc0298f61477fae2d5a39d320986b73859120408884c2a5f12cf9de2389e20b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2dff3e7b49feba1ca611087fd99143e5b29b872506b260e8dce9d430431497d8b6b577b6eb4ad24cfc06dc8f37366893a98d76a9812a6969eba875b956299bb07656111623264ac55e253712b67bb486f7edf4d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h522a34de0ce60f069a5124f0be665d0e9f6851b918a4c8caf4e94eb7c052ab6c533a08688a4e8ee9e7407127e4d30ff084a5f1713dd95b9c435fa1261d8093f8b64e7680f630769b520a6cf95cc8280f51ba77855;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h968299ff6dd73c246fdfeb806014f393b800ffbc43d882cedf0d0bca2af7cfe5fea577803d8b627bb0809d423def57b580154d224ee8d6900d703905d4d2b9460143bda5033936cc897b79c16d6ac25a98d2028f0;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4cfa06f06f3aae86daa89bdad4a70bebae3fe33fc1435bb3eb6ed2d6e1a60544a6742747d69a9ff1a1ed16feef18d521ba6e95a4d0adedce89e7e19ad7c6213c6692e6365caf2dadeb68bd9513703e580f713c38;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h59b689015bb8340bb4d8b5c7030f26fda81e728b8c399ff67341c3c880a7a6904b51b1f8d924648908e7ebf5605ee06333d849234fe05c4434fbd169813f7b5f381e74e49f5945ef6a4532f777e004f8f53d1252f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h535c56c93cb52c7fa15f4f7d8c57674d806103099a6d31349547ff5011916174506a3ccf4bd721855da88628eabaff89b6985fc2859acd488eac11844dff44a07791478f5edf5db6e70cd09986904e5a9b6947adb;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hec6d2300587fd813f7cdef32edd5153c82931417883f4781b67874a5f41f017531edf2935bd1a94de4523a9a4069a8131d51cc9da70aac45e264b575796f3a961abf80195b6b972d4326e83ad76f1dbbe58ee340a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hab8b59c0dd4eca04e7bb1a54c0af5872e12bb9dda00350c7dea4636801481eb5e6cd3b00230c45d57841f17924eb05baf0c4baa062937e7a32274881e8d6f7839813d605bd9afd0c8dafd474d0bc4c40f9a26c623;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he5d25598cd2ed17273442dfa5854ca8123f102cd900eb5036cbcb4300f626bcd97cb3f0a7f025d044aaa646139d41b0e0922dd2ba11d614a46bd6b98ad2e3c311d718a018ce3403a1a2c88dd2f35941fb6acf476d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha2a5054b803b199e6ed59b27f3a4f019c3e97a4af072787e6d2c53f496dbc2902842a919089815fd8c5768fa2d47bedb4e62da6c7306d16f383729b496c218bcb9c589978df340ce6a9f896ccd7e92ad04be09d28;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd3a9f70e3d243b051b54b30a56cf23f5a2573f8d84af67407e64c099747d89ce959ec48c3a4cfe230eff90065cb838f9194b8b74c3990fa7e6bce800c0907dd8b62cf3cc40f116a887f5d8f392adb1a8922ffaf29;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h76579ad37859fbcb2197639942975de380ddcd2f5b3436ad8b21f50787ec47d3bbdc88d3c968f0fa031016faa52fcb249b9ba1f3a25426869603fddb54fbba69f463899b414f0f16c070dabbe3509ecaff6937aff;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8e23a3df22f0eb5c2ce6ef0f2f00d9173ded84b7f10672ce58e3f08f20529fee4c3969b9a9eba8e51932836517f51877acd291017db39534de7613bc5c1f941390259d0628f319c6719c80825492b37271bfa4e95;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5ebf3616dd4f5f2b0065b9b8dee954e8da1c5ca7af00169ecc3f91e667694f5e6c2baf6a18933017e09454110e4754096b8ba6fa40b71799fdadae27b77ba1f8958a996c6913e199ad2f2b4846b0137ffbe855585;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he3499bac366f585a48695e13212cd37ca839972df73bf32a142f53db53cfad9ee4cef115a5aebc83aa9e40ef2fa88653490f3e7897e813f23b2a0f1eda3aa81bfa4acc7641a9aed000852713767f791d9777f8a28;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1106920c63ee423b37a6106c4929251af94d60e1cc82e1b5e4789e035bb02ad17b156bf2aac8b583ac39bad50e6af630a7789cf96ba2504b3aecdb0a38467ea0e8831108ae912aece0fc0f5cec38bea2f85fc2e22;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hdd50cb145fd1c826babbfd574fd4555c4144c20250f17d3d9b3840471e306acda921a5c0aa2a5ef8f14c32dff68935c23ef09e472cf2aa41464d0dab50feaebe7b9c27cd1ec10169a088860a449647fdfef26984;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h670ad6ecdbe248ac23bbcc43b69c0dd1ed428ebfd96729fc88e248df14d876da19cc8d362be1f8be8c816b6fbffa01e60d7dc7875bee7bd136ff796449a15ef429b6ef798d45fa84da4c7aadc2658ca3605f90812;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6a4b71154c38846c6f67af9d51ee489f5fa1dbfca163b0f06f58f474da1330c11e4a8fc3d85fc2c0c8f379f1473d6d792b905b8009f9198916656c3056f4b3fc0da72e567463de95acfb76819a2c36112ded593b6;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6ac48efd1bf4e9be1d1e396aebb7ac02a08ded2f0c92e9efa7cfd2f3a67efa9e33c334ac51efa5718c3fbb2619befcf47491ba458dbe434f359911b263e7e72020c1faa8cb0035ba61450bc81a95aadc39c4846ad;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h387a6ed3e608292387896ca777e30c17877b4f410d26514ee78de24ede41d5b444713a95c039dcefa988c283f461bb932353389c2750318e9fee8e9553f229ebf8aac2a2a901c54eefea18fc5b2a9db1fbd604627;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5cacbc87653a5691cc121572e02a3da723d48a837a5215f2023af17205de3b0f3d398b16f97034f9bc1e1d82bac361311f086230f33ea1cf21882b27452dc93908decf60d4a5e1e9f7375f59550dd0e3c83a2a4d8;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8ce3124046a4b598ec1c4b897c1c72e1376483fbd4cc2be229a2a2e05220a517797e3646f0786bbde2ade3648b4edb65e16cfa489fdfcc5076214ffc8d0cc81a2be1c8f5fd7a2cd8d3c147a89da38a310c4bd079e;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2db74e4a1f65eb94b414af7f268fc9839d8fdf436db9e69f367f6fa8b1a739a1122ea1b75458fa2a36cb0f41736502dcf4ec7dbb6c399c10ff2d4bf8c609353f874759b905c342d834dddd19bff25bf647155331;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hdcb46541c992db3d7a25ed6daaad379b6d3008820d7c7fafe61494ac02fd750fbdbf1299a34ffbe7fa2dd6c6f7dfb5be070e53a172e85ef80bd1c6ba7ebe032d2fe21fcaa2c2a95735a2bb0e0ae5b8d21ba2385f5;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5bfeb61936893afa6de1d0a4c2165334d9a7f0504afe63f1e0e9d9fffdd31203f7539d32583cb139628910e9db2c18e55604856b208f089a1f3d0ae4fdcb0b6dcb52172eae2c360ebd23b759b123213c6629e4b42;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf81086872e4f9ed4702130f7aafa90b291acef32d289fe6b742d1b6108e509fcde932fc6ce5f10470a3716bd83ca592db21ad3443beaf1b3e2265ae4a42b457e49c0ca05d7d14c484fa21b48713eaa7c8728e7091;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9dfb282f2db46b7e51264b5e42cf952ea4fd278f175d0c9978b707453a670e04d507e580d4cbca9547f83c24ded23bb1f7cda58f74cf3b855a286b024a8023bb4049fd9f82e7026d79d8a213cdb00960891106075;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h656e3145b30789d5dfd892dd266d9b81ef8175059d715817f02f2cb765a6deb205c4246afe3b92d0c9c0ddb2746df624fa8337769826bc5c9dabc32cd464bc8affe45552ebced5d46f8e29debb052d6caa5ad1438;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha21b9a1292ae3e43b264500c2824c50e4c96c3948ac8c541ab74a84b0c76359509f02a242226b43a7e706513ed43357ddfc792c424027ada829e32d62d3005f4afa87ec81998f4615bac26a4602cd56f10afcf977;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3856c90598abe3275040508bfb8e9f5ce503eeb6549e01912e2bcfb0fd7aac449139354f6744cbb351dfbb4303a4c09fa1bf9bc269bfac797e975cdcc1bd0f3800bad15b49eeebae9e2ed2e931ec3c19ccc2cf3ca;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h933a6fb906915e24b381da9e548a5f174cbbeedcb8b1aefd7515b3caa0093392cb6685bd6cfb95cce2e9075beb4f62787d7425d6ae6cad8ddb6b5e0127e95e813725f920132c53d67e2cdf2304fb2e33fb8bade3a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h535b4cdf927d7b743d5208ee02524c522a1cce4b3d3baada00bde7d52999bbd8b8c82491a43c58962640f33527ead007f95b756669ad6cad274473ed2b472ccdb7dd0afe4d079335b0f4d5cb5b275b32369934734;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2e0c0859a253baf2a73841ecd8ca8f2e2efc9e985c88ccf5e139d2615ba136ef492a8a4a65c0a1c51a6414e072d0bca5151b5205f14283668e4ebeb9bed5129a2a3922a003c405a86dc54f1f2e8f3fdd3b55676e7;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha411457772765e0b280ba30b4bc696fb959266b40878ca52d26b1cf9e019aaec5851489b0261f81688e1d964a4083ca13d47c210a50bdb55449199254984e06bb31162e95123de27bbb9d5611b6aba0b66fbb2dd2;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd16d48be8fe44b1212e9309ce7c79fb43276a711e46391c8aeefed354c24900f3e89f8d1946713aded047b6e8bf1c7325d5debfe1bee7b9cce30dda006bc0aa9c5b99ce96308cef438bdb8b6ce7f9181f6b04c6cc;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h565975080dfbfe9b04913e6cbce6a3e354b60b24e218907083629085fc4d265115ca230186845fc1fabca3bcbe73ad217b2c8ec3cee98ba6bd795481e2bdb8579e49118391423a40cc0c07c75324bcb2f146f1c78;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb5a26fcc15af7bad3757d9d3c7571274eb9367180cd058ffe24896f0242046237ff433c0fc7eb4de4c9686ad1360b79b51dc92b9d615ab47c4cab8a7f71f49b3673bcc0a557bc6e0ad54a272c8e20a8bbf4afb9d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hdf5c7dd7e9e1a45422602d31ee4ed3fd87b4dcc49ef7d36a69f6af233f199f8a6570df2887fb6037992001bbeeada785de0e6595ee791be250defd168e9193f9a771ba306ea9901f354771ba65bc02167713ca04;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h13f4090cb040454a472db654aaba2c703c85d18c91b5e79a037a4c53a42f7f12cb83177efd6c043032f4b9c992342a98d2567e642f2c05718229553253c10da3c431ee1352b4c80a9cea745af79c2318acfa3c044;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h89a77c3fc348fcef711374dd84be17f29025a2e4800b7030dd863c544daa7e7ac469fcc9f712bb321d4aef24748d07cf92573c256f6a9e9ef806e65403882a621ef508df8c1861ce7cccf036317347c50cc2412cd;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3b1095df971015fec2efd1543c127c691f048ccee75603a0f6fe2946a0bfd2ddc5090a2d0d58172005d1b5aaff5818277ab66cc5fca20f10697f09f425f3b14f6bb37278fc42201ad4a52a93721e288c936726ea0;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1fc6aed54e710e74bcad20128cb92de2e3a06a0c57159bbd65872841647fb6b20f9063fc27569ac2b212211a1f815d1408544244f581fc220032a72683f3b9d75c32a687d0d8cc98cfcaa40c4cca3be692f395c77;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfdcdaa1997b35e2bbbe3ab8c4afa8e60e0b88e122d97f68ab74c60ae9910b9b92745957b5b4ea998e38c7e5c73c1f10a32bf897302a010ef2e768f82abe6996a28b746f18d3b1e7f05565cf2c7e900c1c73a84c35;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd57a2959761e39b30c7525071c5cc0ac3d0353694165707502bc7383a036c01de73084b311eaedb9662f5ad4f92beea40a2948c66edc1d3c03bc27480d52dbb02eee74c1e295d4b5101beaaf6fbf2f25a8c5daa9f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h87a14bed8386564e41a2bc89958a36cb58f9bc43caf7b45edc224180163ef9b1bdbd3745ab66595539f30b650a8ae009d97f301da1a15a165b838e3b4a0319b87847e325ec83baa8351af73d346f9f97f311f0122;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1ac26a78ab89fcfabd58a5561bf95ea74d72dc8ac306eb03f7291a989c6a49832f85a693437baa77d2bdda5d9ffe58e86a2874cc1107d1f2633f23c261a1581cd08dd75bfd515f9b3f1aa91b766c616e4844588f3;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h20a4600d3cfd4f6438cd2f8e728afe127eec8e5e4ca8b172959f089f994235c1b6ac0f31d71b71ceffdf359a27841e80338a2209a4adb98032be5921b2ea84604116a793121120f80c34a8c9e65a6c06cab7d5760;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3c990a5461b000ca3b59f3fe81c4f71ec14a50a2c3094a9eb60b9d06e6f319a77f27a6123c3650daf2b06ce7d1e9109e75508db73a5d33fd9f391cc11ed35bc8102d1b29dbc431f3a5b23878486005e74bd9cf5c2;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h14e6880815ae5e14b5252229d0ed96d1de97fd44808f87221e274ba22c98abc85e7e68e3a8ad8c6cfaa675577c5be253610d5ebfa64a8ee06d6f9232a5aa870a897356fb4817475897b3b7315d6b790a4c58054fb;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he329b39ae5c4bc1c2c4b18d668fc043a0cfb0ed9156dba7329ebc5ae9838025997afe9fd3bed49251e73df1e00cc458bfbffd6a8049f8d4bf60164b43f83e91d60d4028c00fa49ad19eb13bbe280ec7c4f047b9f0;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc75ea712e5c37b45229ab5afea1bcb2241ff478f2bf4f78be62828bb1c970b929dcc0aa92dd6472fb351e4caa4d7b2398abd4db436068dd3c01030b3a4904ebf7717ab914d3045a0f1b7bb6e25899ab22ba77d6c7;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hcab51e1e2aa7d2f628811d57345db31b33fcde0d6792479b3279904e32408140902b48d014d194000e864208c8348546ee3d5335140c79621ee1db6ef8cd3502572edfd4b51e31ffa10544e5a3098a78d6a3f0810;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h951674442c0e9ceab1ca8990e02137279ebce3825452eae8a6d496a47a222518a3dad672d3638c2d006a4ba88bdab48f40c809c88b083ad6b64979404c4bdd7ac21eeca401ffe68d3be7771f502fa48be97b15a1e;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4abbc98cd821000835b6e93999c8ae881e0cc85e70ac237cded2e42a512ef41cabfb823b90dbbc43e97e39c1df0ef4e5c42d73c7a120b74c442affde2418814d5a2a9a720ec921fbf7fff2100499a98c2dac67c0;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf816b687d442c6e830144cf318bd883e45f02b7ace967ea5f2bc5876db2c88a852e24b5f5b99b85674ec46c76ebc82c0df2bdd57d2092c48aa30028571889a5237032662e847bec229f47aebaacb83e1125c0e255;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbdfdd65a418d230e51fb667a2cde23dac47d133ec530ec9febeceb2e23b51cc37b1e6ede84fd306482dc0386d502a02834751dd2c95e993894da41215907ccc0c927f7cac26748b1d7d5473dcd4de38b46ec9d413;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hea9fcffb99868541e24bb97989c24ca916f753b479da416ed0f68944a387ae43d7bc64399feed1e3eafa09efbf4d8ca437a01d87276c215c1f0b8255e98566f4138ec6b72ad2cf4021768f2262104619a5b767b52;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h980785cd48d498f86869290324239b17e255c5805641f54a7391a00cb1d7547f525ef5cf6883912ce9f2b75f52cdefbfbd21821195ef040bc957d06062abe210c4cc98c44dc67808f8b40e149223e33e08809902d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hdeda71fcdb4c6057678b0758a54002fdcb582cc1c82f02d52f5faaaaf91756de48ee400a73f13392d6ef4dd6f62c100af0d19fda6e111a02a2f78efd0669a555807b1f166ab3015fb5552e9eddc63c54def3e70e8;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbda3d7d3f2a46f36f835503972101a5347cd6a9def5d2e8555299e12f08111a652c4352b81d7b2df34dd4897850b9916a22c1cb452f6da6019b9af8adddd0d7e573ea279f26cb6a093b970b6621342d2dd57aa033;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h673662de4bee5bbd2d242759e9d2f1ee1e8a29f0e8feb81d5564dd13b7fe26debb2c5fdd2dd82aa5ac7db1d081b0467020b0e18f9ad516e67486b657c2ab9d1de795212e7a2dd214967a69a505bf7f09b8948c97;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc1ef128dbdfacdcdb0661a4dd47253acdf95f6c5db8d242f6f57d01bbe8bd0fb2fd7ce5afc4aa8fa7cbe1364a25ad2870d26ffae3c19924d121fc71625e7df5eb91dfba98c74d9255139367771f4777ed35ea9ed7;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he3184a4c69cb0c6a9caa3d9b38028bf708d27afbb2b3ec5a07196d5c0844cc6e3ab89679f59715c5c6afa57dff7df3ca010d933e7ddcc739371dd12951ba5260543123872a2151b6e4f2722cb2888b4b1b386058;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h39e67eb85cc88945f59f50154ff25bf09dec5937c12b29e5250b170def84c54a9d34569767891c9ba6ba2e37e0990953bb8af7f9426ee99724ec126eb9af0b787f004e63d1c9ef3e4042eaec68e4d541920e9589a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7c6c264b8d08e65e29d6992f4a0526d66b83ae811eb7fbac8805cff4f8cb18168cf462aa30d9ac7cb969a9a724e487bbe1684d921d71fdf25368b19053f0deb1c89a59a0a0b8cb2bf4546b50a0bf534f2c3994963;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h52d314ba2d53b62bdfe55a985b3eccb13c3ce06dcaa7bd1e9de97f724823f2bea498fbecdc8cdfdea49397f4a7caf86522d4d4c06e8f2c6ade94d0ab7e6a3c627e2282b96f65ed4ec2690c9c72e46e019d01fb516;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h98523670a82bd8cc97cc52f71c057b54d30259052399650ef16c18789801e48e224371db6036a8f76ceb4a62ea7b6b02486c0103b629fe797f8f9541bcaaf4724fc47a044c052fcd7da1d86c6df98448380dc98bb;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc88a74af6749753958754c8cf697eb75eab6aee290547f864a899bad221f8bae12c689db6da1017daa0bcf98f1cf8d3e6697258523f6b9812a39783afab7d64b4ae3c97051eeb50cf014657ef01f472afa40b059e;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4d800dd6bae83b6bdebbe47260f35eb6a06bce3851e02e556ff78fee6d7618dc120a18d39a80463476d7c659dc4b00f416e8066a1aa72faee2ae6bd4a2b69b412f44955f1b20e1d7131ffe70b9e5cffb59f53393c;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h911792500ba1a8f70ab968f2191ca31db80245705ad3c782b72423af830c228ac3222da9710e1d25058dc39d314c677611fbcc7b66026214ab59821f86bfd81e7a0694909e2b5f993b0facd1e1fda6937f5ff40c5;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbd293959c1fa06d9f0cee91a09ddcfc326a1cf22dda5a2e8bfabb8df75f647acfa3420fcc46f77b171f51c83dd6230086822519eaa822f54f39125d83342496d2f8fef9e921450b2949e4f385fd81a124aedd569b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h737c991a0a58f78cf957670d06f178b0ddf2f763d64f9476b45171f2793e7d0ba3ff7d42f403428a09bcf6e472314fde80388b68b3d49847e79940f59f619d97ba16cf479764d4a6c91bf132272eb2f8f81edb02;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h615ecd50742fc790fcf752d1111c94d56bc7380db4755c906faa16d711ccab0652eaa3077ee70ed25c284caa4ed79548bf1033cdf3b551ec9b07fc7f8bc2327c31aa63077497439b68985e99747f9cb9751d30b15;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbea00a3dc70b91d4d69ac880d7241f8a705c625da4409d7e3539a90bf2f73c6c0e547ffc61613a903177bc5997b68d35cef195cd6b868b7a1faa61dc8cadc96e4a9693eafe63804c5c9ba8054bdf8c62a2e4cfa14;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h42f87fca04409b70d3ad2d95fe17b06501cf450a5f25e70d056535b8a8b72f777b12b7b7e159139f6d74f57f79a138f67e9cb0d77555dc050dbee40d734ef1f3d2ad6d6c87b26406e7aff54c1d41e4c2d8cb8983d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h24b6916b699ed24de4e3036027bcfd0af88f66a6903fc57cf0078f89f923297c0e999c827a80797477a91915f1c772f360751d4bacd1fc25e4ea33f0b1da5b571bb70200f21f2fd9b2c4c7741a17578bfa13f4080;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb700918a180dd9d7cefb425413aa38f8eea573bdf3909e8e522116a78b3049294849bab09b5d9997fc21828542ab15f905d55ac7130b448f9ab7c4497bf07837b5b623c061bda2e35ee44b9c8c0ef57301c1d16a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h77e8c5871584c2831ef770bbd1190d0a33127b55f527c439db1e2d3737116a0db56aafa52e4097a67ac276fd75e7d6b27562535d510f6d7f77d7e5710dc6249f358ff27389ab42d1fd7bbca2541adab4c518393ef;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfc6f7005358532f548b633df3b263ce14a889575890ba95d4958fc6d04d31915f2dc1c46dbf7077a7046ee164ba05110329ce23aa5960965e856e0948e15ceead00952dfea9bd22df4bb26e6b55b5c18d91f9300f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb80691aa5d4e697a13f444825957f2be3558762db3bb62765a1939d6b6def62d1571885fc832784b18006cbc8c5c13639470d1f033972e6d96c7f097c8d6ef6b976d0ebeeb935a66a1fbfe82c7af808c20a4c9140;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf21eba98fdd176332c8e1641566208b728a3fbceafb112a0d82aa194965e5760bccc1c548eb19a6b42d1a93ef1ef94d88efcd4e4acf74c0c4f058841b49c2324892542736c1fd196d29584b5a57dca7a44020b6bb;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc06e9a23d9437ef1c7d675c9a70239a5928420218d0f583b3a5021b857cbd3ca9c5347775a0405d3313434b162171ea0132425dedd9b136af476c72adbea033d94184b835c46448fc31baa24b34774f84a7b36850;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7fe673568f6d62df2f249fd6c7eb4451560b529f6ca34911b9ed318d45542c678e81cbbe44fa19cc0aa9915a2752b71bf6fe3388f600d13b8c1032eb783bf13db22a9bdd047a31185a50a1e0c40d902d084ef32aa;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc1b12599b9c1ffdcf6c2446d5228489efb811f24dea63870ded80c878b9ff11006939c27fe37e373d1e5f9e087cb487bcfce139a48c0d2f15afc9cedac9be9db542d4bf137f4008b41864acb95707d04ccc9e5d1a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3d330c0f944a38b3bce0eaa09591c38e2a30c9706b5291677f541501406573a54e8530898f10175cd90e0447e93bf42e2431866878af191b278c515ad8da8cca35532317df3c8fc039a9a33db93fd6d5a96cf15eb;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4a4003579587a63a1291fdea958a831375e2186b90a8593696086f55b8228e0a49009c85e53e6013157c43416fdaf73999ca89e12bc5d7e32795678d93a8438e2afa3bf759b1fa7ee31912a8797d32c18afedcab6;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9b5a1d6d5f2135ea3bf5ce3383d84dd9e474ec9431138c53841ee2900c96354b33e3fb3e505642403264171d94526b641dfcbb1f318a62056a7cdeb0f250e342ac3806c6cb2c5e2583e7a54cf7673df2cbe34c743;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h29b2efc84fcbd22bf9bf3df9db32c540a4b30ba1d7f33a848b1a4e471d309471911e1c5b3601b2f9cfa1b5b568ac3bfca2201558bc1ed0cb57eb91990e132367fdcc17a67d21ecb4b5aad16118efe3f6087b7b14;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb91a5a30d3f8220b438168ed9917c40970e153782efff1e088fcfad4fd3266a4699269f00579984e993d6d9047c6d1514bb557900659df94777ece302736e85b6bf2cc968f798be9ef07ca3e2572cdc8499cc0232;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7d4de1e0ada8d58cba74814577e8e8e7325e026776b271c7d3df089b2f36ddd398583197efb200334b9b823bcd3c958c5c169a261d08d42d4967fe724445521fe9f79b46d9991f80ae57612b5afa4ff38b63d13ea;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hca554c4ec347e2f38d210a4363e941c18f75f879173a2bd078124e4069271be5d492acb627b8b4a2b98b9b0ee8243db15a94eb7fe5c10154bde1a33aa59dfd0611c4d3a6c4df682308bf9a79d9229da8d242051ae;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3850c0b8502ff113b0f8d333a7125d0db1bb2041b2c3322ccd4858ec267a680b1980cf00c8a2bd100d0ec3b81a04c06030754932097782590da2eacf7fa58b38acd4ef4ead13e9eaf76dfc9a8acffe7dc53f7cef7;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h767a38de14fdb78a670b8576f5bf8238f4e27022d24ae669932edd8efc07015609a5bcb1ee8224400abce88ec1e4d5e8dd894a7e44c4b7779c5d13e18ac75cf969ca4141ad22e8abe3b604a17f61491629534c99;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'heba1c60e33636beda1d1e3272b8eb5d5e0086113ccd4e2635c7d2eea94a544cf4611f7b524219855d2a4204af0b42ad7a6b0d4aac36a4cd79d8e53f3939100b0089e61abca4b2fc8993e53b92c4f649781d0e9cfc;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7e51f1da46077846dad63e334d13c39a7b6ee0ed13c50af7749800222577c2075da0336bc2db36883fe15dbab8606b5845dd16b32d5a11b45003e923881f708c4e7fd2579ffb5d496ae432440d9682ab7dbb90a33;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5a615dc2e2e6ba23b65a9e8abc9acf244a38d6c4d3fc339f3cd7fec187df906df7fc57b1ffa314ef45958f950533f1680d07baa641c5800d9b82c31bf424ad0f18431aa217fe988fc5cab2dd784472b48b548a69c;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5f8e469c15f3e36e54ae0646c4a1fba371b30ab495c8906c683ad68ab342b8905e4f6988dab7266d9b0256dc34aa40a31a43cfc725d644c7094d1144294566f271621663eb7b5bc9480e7edfa73cbfee0cdd05065;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9ac22e4c76c67df632a31c20dd924e2cce19ab1749ed265061d782b386e776490275bbf21331d96ef9017182799dc0d63c65b1fe760baef7730ebacc216ae6a27da42e65c72510825bd17c1f69b1920352a189901;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf7bd2b44828517130f974f15b28920fd04cf7c2e4ac29971e8f53ff50d91478b7914af58cf9d6808df26d850160a94d662ee3c30e464292eeeb7488b8dd6a5cb642e90d58d2f66ee5bebda99b3cca330bea6be628;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h840cb12aebbb9ee8a0a61cb4f16f5689c56cd1cf7649cc32f2d7773b2807dddf594f62ee9d253c308c2835c2056f4b274927a9bf562793e1da871ed838d81f43cd68cbf171b7fae954097621d00b0dd1c2996fe01;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4e432ed78433a7ac1595acc89686515bdb8e3e0b58ce94aa08f1244a911e96970d43bdac97ed4814448e10961257d5368f10a8f8e089345008c40f7a0d0514a98e3f279e8f256af17ec1727ca70c4e13f24e632d0;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h56746de05b307aedfae289ece1a1b01c35aabd6e47dcf2aeb453f09c5c5338bab99f4d5bf0cca9a3b5673bd67532815a22036c99c0114caaf7109bbe9e681eb11cc6c56f3de3d34e48227798d8d10351f6fbc501;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfa0dc57f60bdf8fa35f5827dd4f5070a619566f43ba3cd0113292af9dfe316dc6acc581bc44ef091c635d941291d6fb08633eefba522e55faa45f4246a2d213848a85eae5921ce444f12b31eaa87dfeb7a8bcc790;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc803be38672c4cdabf2f8983f11768614f48e648f1933948cfd1a17d8b110ed1a3683908fac8ede48414746564eda41d91e47c7c56bd11013caa891a09b1feb8d9de791b0b2e9fa49d0899ef66dfcd870f6043617;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9e289cfded3c2cec1bcbad6f835bd432481e045feb39be74a0d815282d79fadcb8a7318ec8b25a255d8750152d68163ae85df59acf71d0832a61c29e6c2862780058ad7a826ac11ebb038e5a1830d2b69ebb35f47;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb43cd4bef60ad365b5dbae71b55091bdcc64cc176d0e7b4299308d9d82ae318ef78816043a697c9ca1acee90d336ac2e04b30e3ed4016469def7463c7034d628baaac94acd0bea32c636025fc75a63775406329b9;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hcc600ee3ebee3cf7346fcd0e02f7c246a706075ef486733858eaf33d18faef4d8abc6e7a40213dae1c17bd85cc47cb759fa1583c0baeaae8c5fbd4242ab7712ddfc5fc7a04fa26baf3f9a2659f981fb87aa84f99e;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8ebcb1252b15bfb0aacbaed256d7c63fad2b4439d320ef146f7c58ed4f8e44c18251a8714d1eaa588e4a4286a669609aa115806ae37ac0907ce4c6bc72b13ac7fd67ca889948831186d73c42d5505e1c5dd40c06e;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h926af0accc116ace9b6c646f7fe2696185b36aebe8f1fa72d05108a8296d8423caf96b50ddfb78c060029f56b1eb68f45b79336c077dbc336ec43c21f97fecdd73633818b394add039770ecc545f91a657452437e;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hcd651dfed26ffbed1ba05462a7906d29968a4f22ca86cfd63d3d6bf565969a7a90fd38cc90890ae64ec18aa3bf630d282a59235f8aedf107bb910f424bfb1071f76b53595ef7d3dcd910593f32acfeb983aca1a08;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfa79dbf892aa6688da55a4790035d0ab41cc6543de026f9424bd21aa04bce502812697614a40e9c773c1c0946d4b3497be6bc2ecc16138c0ab3684a92dc95c197988448b53c6f3e396ef3d9198cacaccea56e68bb;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'heeb7b9ba9e49c830834b6961577b513625d43403894a463daa9fe7a1a9c6a9841fbb024b695c0dbfb90c87e1835f5ba174f9c1ea94089414868e8011b1e35bfe9ec24c29abde0e7b36f9116526f01bcfb2b88b639;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3b32751c9b8ff3f0880f4b2212558eb106620f561be3afc88d51a7334ed4576bc0971de069f4eb24cd2e0503da9e7125629024d00c9db915e2abb046cb559d0fc78c164e825253cd67af251f84099a01ea8ba6835;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha0b9bf5898c257ea00b8b1b34875656f6317df836ca6f12f93e3f6f6dd618f5f8f236ccbd23757e54ddab025e558d519f30a44d3b2c4e7293434985d4efe0835a3d0e530a30d42c2518c3e64fe9529528ddc14c2d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hcbbb9ad10ef6f9c3e56e18e4589fa7cb4e849993dfe3bec40028ac85e3a6da39e097a349cd0a4ace3fe431231b36e568a43d1d6090c12e5ed19dffd1ab78163d767125798806af99ae6e9fefb7dc922d5718f7356;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4f2a394dd7c244f1f172bbfecc45766203a60761e073205bedee5fb34994a19fc986bdfbd60d0b167420f08c4d519da9a08060f74f685124f5c0fa4a580c5c7e65de4d65d9e7f1279d6b9acfbadf87b81505d7ec3;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb0d05f70992102cd8557df05a694da9f4f434c29597afb11825d723ec628502c2dbbe9add9b277c7aa3736de237d5ac6182a752c52924a60464c8adf8d10bfcc9780d48c2dc22dc2e1b5963be03b3dc038ba7a2a0;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb35e5f828898c7504b9458fe47ec9a045bd217b430ead62da56c5f082cd75b75ea302f30ecfe271dc8f6b213aa59029713dcda048d0bc2f39813d1b231373167c81bfa2f23208a65b1c335d3a00549df72c6382d1;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3168e4a81f99c2abc3314e72f1834b025a9f9fcb47a2600030500169a5438804fb47f2718f9545b18827a270d5e3790cc75491cf78059080714f756f670cd88ced031e9fadabaab4356252f239d5be063cafa2449;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h976c962a7c8a9c24b0c0e4fbb510ccd6334a6f092dce05e273915707ed4382df5f8b0ec1b41eaafbd7470c97fbd5464426b509c40ec3f852c42bdf1db755d5f7dbc9a8db58a895af0ff70c4fc52b38563b5ea82e4;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc5664f346f3b9223dd558f5143e4efe65a959373d5d4213aaf32b72dcbb447f3c84f3736d584959c1c8233eff7dcf0f08b6d8d66d48ff2245608f36798b21bf5d3356201c0cc53b717b5fc0477f9474e0484ac9b4;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha608dab93605a7a6ef0a665edd0070c20757755f171a16dd9bd4cd302077f9d44b6c0f6b39c475d865f1fc9912a305fea9373c8b82ad4812b0d0726a8f589ef0c719498d34f648bb445229ba68900f9065bc64057;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb578be6d291b7d2d918617cfecd9890eb457f58b0f61d4a9debbbbfac5f0b6a678465105d9ffa22e205ed76d2c3918daba6a4d608560d111225018e190a86669b8f24fef18bbff6159bf7a2af822aa81986e5ab59;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h54547e6622a2f46d975a0b90a972fc12aab45bf0259e22c85fb053ecab7e67190616853c4c2215bbbd154eb36a0ad39d4db3c3f4b78afd163aafcd190bc505471fe589b33bf93c2415809675de8f8d5e78c06dae5;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'had0774b5f814ec6dc491c79fb8fccdb8f41dae4e0e41dce315c0f4b1a640dc563d9745a976edf1c9701c02daf9ec286a17e551a93a72af456dbc7d54648360e0202044925ac372f10ff1e5c2008ad10485fe4c8e;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd8d9bd5bf3aa78ed5d35a3096a0c488f5aa00660024eac264d40b91197387857a33f19faf034a5c35297118285a3270e2782227b175294bdaa6c16146f021e9b7bc7e56ef33ae38957787e883e7e278f792ab2158;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc601d59033e5b2a4a79aa007538ec7af01b5862a7554f3f16760b6ef0eb7bea4d906c1f9784fd8a0d1ee39fe7e34c1fc118db0ed8011454a18b6a374385672d46788350a159672907dd41673fadf62eb10cddd0ba;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hed86b3f0757c19f046f1068e5f1ab6b94d328291a30f6e7bd8921f6df37a48869f3a5e159d3c8ee4835635383de496e0a0091baef307a696291be8a7a345d4859430a9443cecca4d3f4e831870b02af29875eb5f9;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5bab92900c3b40dfd255a6da029d679825336a653c0feeae6933ee667cefe25b3a76c8dc300e007698c226602e5ca34af2ed44c63a65e5c49411da6cbf774d8dd3613386409009b265a04c9249a55af20a65b2a20;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6e613f1d099c398e46a086b4ecf167e3af366345c7766424e43a4731e963dc8331e4652677a12789c64c224900dd4b8da31b7a6007119b38b9f6bae59513420a692a8fb40c117ae004f7bca4d97823c017268c636;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb3930956edfd27cddd9fd63d88add47a04bc9197acae4eb04d00a12d10acfd8d8230c0d3be3ff3f53dfb81920ff0e6b1eeb8f7eda12430acde1b665d2be99567def3ff0a73e90e3150d04659bd802fc5f172f2687;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h421a3256de5616d3bf2dfb6b395a6dd43ec663f341ed8d813649143c60b5950423d24a520975620a5da287e2fc34b326e71725e8ed751f7fd31b49fd47b584f1317ebe78e6fde2c8048acf22a8f5fad48d8d34fe2;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2056e30f59c50c82a179b28feb491234cf26a41be66edd4b09b8d8250547dfe36789d32d3569bbc4ac181cea9c1893662015333dfdffece73d4b02cae5b01ba4dfcedd86b9093ed73f312a114b5a2952b32ff970b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h549b1814554624f9aef5ab839f5ecb0c6ae2622cc5dfb90de932667987f3beb32fc2f671f8140eb4b6d613bc837dbccb69cc1a99706f9f557f087f831dada1be72bbcf99cc340d23362719d55f778d26975362a99;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h60a815daef1b597557155566c4fd5eed4b9d6a80a56fe3df3fa9bd579deffc471539eec8000fe2a46ceab58500432d74dd054d8b3bfa2ba823034aef7ea72eb5e1ac27eddaef775b094bd1dd0a9da98b30fa10308;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc2f77894e03b480da6b78c71ac3764cdcec9e71b3fbacb020fbcc34304bc188dfa2dcd4194ac136e759d6f469df6b646bb0ea901b6c1e284e374a1edb4e70c7ab0008b0c5f727604f2d1268129df4c402c11d2030;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3dde268b1f742986edd930278bb8999791575cf1b5d5d6f65af8ebe698ae7b27fbc3c90d379d3fced9ba207904c3872387c00b46f2849af070fa839d7702c302b2d55f660deefaaa1b53432baa175c53d2fb7856d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8abe23085f86df137d1be3a769c1e1a66fe8d3075aa6fd3a6c2a5184aec74ebb2ab5494e525b0831bfc1d8b7ba48dd0c6952e4f0417e5a969dcebc538246eaf9a5ce3f3c6db88361b4659de43f55fac7b883b7257;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8aedce24573392cd1d27c0fb4c7d0e9e0023aa9e98484f073e5dc46f393935fc3c696a3b532de1c32a71fe324db9aa8d61fee2a784108a3cfaca6dd6382a48cd76e12f52b4b2e5ed3a3d2a2db2b3a1b147c672eb5;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha9a5ad909eb47f6a3f8401fb2f4d7d2c29c31c90464b8fce8c2d315b8a68227240b31e37db9cadfcc2ea96b295663bb8785c4efd5457f4c33cdb76650a8bdcf3c08af183f6f699aedfa4274d7162cd5c439448e8a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h579cacef21295d5cf6664bc4227b5e127807e70a9ef3f5093df52624d10f2b2717a2fe89bf9c4211cee84d84f3b19765770866fb18201b0083051f9deb1956db6305027a2424e64e1ec5c53e0068764498f22e258;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4286da491f212798a1aa01b62be89052b7ef2e34aec7c526cf985f10ac0a4de61b13f5a920accef6ff3ed65495e8e8d6d7fe2ec7a46973a7584586e15b75e6dd52b7354484e065bc52ac10acfd6acff6bfde6c636;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h94e3464d5d94da6c907390daf3bb5305552dde4e38ce8f871664d96e5e30b7bcf013b238040991cd6d32514c3875536a2af385e218d9f531c1673e85f132032ebbefb6c9dc8fba6c4187888bcf9f47467dbcc2fae;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf1732325c0e8388047be3f4cf536bbbaad65929796bcf6e33c7a3f2a670a38ec2f586ba453a2647a6f2166c3883d51ffb9d17e6a37e512a83ddf1153ee03810551793c57c5a4f7a2b5d2c1831fb5a953cc83a4741;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h90ca27badd651d8ad2191c574bd9d589cf313ded84180d148f575758d51aa10ae7ca88ae7de75908fd5c81e36e51665c326b191b2db9d909d64fbc4d6c4881660ac656882cda852b30e0b4a9424d472d55740581e;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb6a3e6692c6f4bbad2474535e214793274278d849f7c3fbdcfc3a9d7af8c84e575031d7670ad47ad20db1e7e67f5d8e7ccf8c5467e4add7c5c781062d12ab9db915432572fad119f7663bfe1df414d05066283ac8;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6b25470e7fdff5d07bda3f52818a8d79250e31f6cd1fb3bc4dcf86e116e594925ed93a17b4f268f9aa9032c28e059ac9e52288e75f3422b500f2ca3277b7c58186cd4aa8e2637e47f39b6eb6080f74b40854c069f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7005e606bec41e998915d0989dd9a31543c7b48d1eaed640b033c9701b7220920f4898bbb705c1ab72bf4bbe011c85163b20bd9e48f05d0d55fe0da44034262c5cc6522a8f8ef68cee71a89df5ae8992deda1310d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h852b4e2a71d108fc901088bb06e217c3e967cf277d5f229f3c99d4add52113efeb42aa69cc114db94ee67556212adccf5e89219194cba5a7e84859c85c8fda65bf51c20a4f4b8d7d95ba2740c8bb3dd290eeb699f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfa563585cfb3d64050a46fe85c3fdf3bfb6e79ebad07c2ec1812b416d06e9df14b7fa5e3d26a332f2cfe8ae49f222ed6f75b776f8d401b91927857d3b18e101198425f36fe2dd2a29db15de3331da1ac96778686f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'had63dd60811eb92f08bf63ced01135fd93831ae5aa4fe41e6dfeeddb270aef3c7d392b7783f72c58db86439a3fe6a8f5d66b4c18b986670b8c32c0ed8900fe3707bdf2af20065d343aa1ef39ea8631f8719bceb20;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h97e72d4bd7a09586f99d9a7546e3216ba4edd342bc15a38f4f895e388dd66e5a2e3bed956bb9035d3cb74d6beecec69554e7624af8b16ffd383533b1e2fc8761e98d329d6ca035ab1d95c6472e89e0dca87391c4c;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h82bb8c1be4af89bb0d1aab36c47da235244cb7ff2fd61ab445f13be2e07036b3be04ddf8dc90d17430c7b9f51d559623b0b8bcf4132ff7fde430e05b2f265223191c7927600c0425485115158222383e844f5c3cf;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8423b2eca4745d6dc5dbff28ca0cce1e0a3c0c68e8737b6850e646919e3a84553bac9afa81f7836152f6e2e8cb70f5d8c9ebd7864c4fba2bb93b68b79f876ee7a5311314817733df9b00f2e59d7e10be44b9f397;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hff919bc5aa34f7823d501c4468c154e1e75f0274166fa3c41cb091cd1b9546ba955fbb1c337bbd9ac86c401cf2850e048a24f6b06a465dd05606258bc846ac120998b3f7a64b52e9a6e9ee6db2690cdcb4e0d2397;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8c4e28499b781a0cf0ba93dc595f4678f59a8075f039a2a7afba6642422f6cb9d38fbabf123c206a67cf5693a07c9a199ddd9c979daba3b882f236c8d4e80e5cc9d835a09af09433dafdc16e196216a9888ba8e9e;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbe9d0396378086eec6e14f6438326009d882f524003f96b9746708763e46c2ef92ecf396b38196fe9a1f48c43ff8920b7fc54da77ce423d2a0b5b4e7ba11c18a435d22c6b9977230402799886c6202aae9331e7cf;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7f757e7bfff21305062b6307edaf206ff8c6ee33b01494a59e4b600d053e52915574b5ccb94b8bea824912b570af44aa311690fdaa9a6819660f7912e2609d57dda8fcde9b4a3be2ae2ce031d1d05d10ea2714079;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf77ef965dd3e4c86bcea68a083c65dd4086810fe033b80974a102979879b19e4370e2fdf13212bfdfaf713804222b18d5b811ad969787f3ca3469c4df23e9409b6b2c1d6cd7a2b788a80373c429b6483d80ce30a0;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1a45581e60f5cfa9104d63b93b64cf939d70c9cdf32ddf8db43361045e12ed7d9eaad24fec39476c42c8c556982be350378bbf8ccf698b8953f94515ed1b649af8573d5501de6925a625a06cbc5b53808ee7f9a36;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8f14b2b6a9a84a0c83712495b7c18007a4877db26fd729b3aed68ef513620f91a0b7661db91ecc2b18ba1982dcfa455e0a9745425866e6ad6349f62033e418efea1a30e176af7f011d31841761f5ec3e342aa0159;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h483f5f3f64d926fba6a9ac3530dff6e1e3a4c23d3022f6081d75ef72f102bfeccc3d79e194380ebec32aa955181e532d302152ad364269956cea667a5d447aeba32c006118edd17d49bc64074c4b75523b5dce277;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc70889f1601e1786f0d48c772b84cb9b4cf4c850f485acc6bf6a9a9e9f2d9eb60accab0f6330fb5e80762996dc054014ce5f2bc1de9ddca50c6f2d62df4099fda660d46af70a1d6c9a7544b851fc219178a3e9532;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc56198637e17865ffbb1281fbe9cb2bb3f7eb1c9612eaa2eb7fb12b8b9950b435d98995d3b44fda07a4b90781c1c6a04e0e21920ef5d18c36e361fc2dd41bd5bc2541ef074d7a70b5d75e5bb6cbc862216fd6b5a5;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hcabeac6f627982acbaeda01801557dd6a346931dad3659cbf0fb7ff6da127e047b0cacbc2955b0eed9fe42bd5cc77b49c61c0d0dfb34496c4ec02a0e2e41221f44679031dd5a304c6acedc05609796ee9b11cf807;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hab460071b98224c033fbd8f9ccffe65b1766ad5e0379402c4e0ed434aca15bdab6846ae90eaab732e64e59e783d6bc9fbbcf5fecd296ca813c1f09c93fb75df8656a414b32cd0259824b36856e11b10431696960f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h68bf03b9a3ca80e9035f11f4c0cb043bfdde0425188a45cd89028adec6f81650810a57b0a101d4b929ca1f7f0d76f91c38a1f777d661a31a88d6875b25367c5c1d4ea1bdd2fc229b5ebf896ce2a65f337f764d0e1;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hdb37f8b3536c65aae30957a2333f61c89792c0ef5ebc1a21e7ebbdcac6a6224186ac4a39e0ff99d381b40c4a423904483f2440db844f67796a4c736ed672a688f827e0f8d2e94adef556452b8585397e5c1da896;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hada055ef90489a7194811a8fea5fb27f5f95ce37e1fe2939ff48c7352e05e781302de664f56875a18c5c8b7f2d6d02fbdc7c692c463a1fe0073129a65f9257a72925bc703ce29cce6e83f26521edb69c42759a550;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1a9bc33e954a1b4956e8b866ceb6eed32415ed430987e5e64ab354df3a5bb2e9673c7c981f402a6b4b3dc032797a12e56262ed673175038116b4f919ff41d762f514df3c43901fc27418a9ff178b8c98c09225d81;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf9d580447513e4ff99c0b0f3adc0262fe6db48adfd42939cbb7efdabceea7062e8e758572400197a959485fbf95e022d11601a8dd856c1c651bd011836bfd93484821c25444c0c9a945d9670e5383e3da755e9dc2;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbb4f80c69731862d15ff89a516d3f4fd80414344cea3545165fcc8cef56560968f7b6880f5a0db01e2a58fdf3955dfc376bf90d4f1e161526d17bfcd749456f7c3952db50a6b83cfdcaa67710b7a8056f97cd43bf;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7f8076d4cb997f2f7dedaa616f44b517e5fa9bb7c01c4bdfc84063cf9d1314439b314269fa1c4e5abb122f175391afd3c961ab606c279d1c580304b9baa34f42b1fae3731b483059f51c7bb4b866a3a2405115269;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3b6f5c5803d721cd90b1ca5eea9e437e2cf59ef756723b6645e259e73c90ebd57a16ea8cb0333e709b7164f37d55bdb58b60f456bccd358cb204d1256307fb560a838dad4905784e561509847fd087c5355e126b9;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hcf8883da426c1d7168aae6b447b401205d5350323d80bfb32b67fab311a34c03f580aeb5383dbac4e835c242cd60cbe89e47bef33bc9c369dba351a4a992748783e4670f61bbc40971e31b0aa4c6a20ab22aa08f1;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9a5f24b2fc2c3da3bacdfc3b28496344727a809195853db9362df324c37fb65d5bcd1acfcdac2f0158c5116d268c10d77afd7423c4ee98fd109342412e645f08c08739678943e8ebb7e84007e835e18cc049f41dc;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h58ade7a2fd660df378a8ee8f14052d85df4c150aa222394af1c62dcf6ef548c43b8f45e9c6e2164593715dba752d594613418de6659ebcca28b1af23c6e9136690430339963fb2a08acc7a8fce5a7624eb820d6a4;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h29791871e06f7fab52edccb6a236ad2f47c3abcb77e2a60ab7aeeb140ae1289ffcbfc0f5c59074fecf0af92c6010203a74aa3645cfbf3f3b4ae6908410f000b75ada12d28612996d3385dfc62fe929bba1ef3c7c0;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h29cb7bc268f25966031e573b440e335c8a91bdecea3bdf63d96c6a892b2d78c2e9ef2d6664313086330fa18795458f962bb488bfefa1eda242cfd4fafe7c79e9b42b713ace248b2b8296b5f4392110f899301f7a1;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9f716b750b2951b6e3744c7c9cf76958b1d3dd1205605af771ce61b9476d67c5b8f0fa2f3aaa383e411a7c3326b34b2a169722c39bf33783fbf02c6c28c5506f8e5cff948bcd0049b14454addd5d28b73352be29e;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1115abeab03b1d40f7d6a71e85e40bdd45982c63b96b067a6d2fee2dfb84b31329399bda2a4d1aecad827c914330d88f84e18778c24e66590fd64ee04e3fbbd967162b14f79c58bfa6d806eda95b733d13e3ff900;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hadca0796fccb873e443579fcd02dee20f07d923df24b8818112d64bbe3f021206245500e727c55bb0e6c984075b520e4e9ffb71fd727ecaee65c8478469587a2068a5b9c6f63486819cf684dd5182a4205982c9c9;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he30e63e4b287a0b6689962e3106e03920205b46a844c272284dd8d510f0e03d8cc12a511fba002589722492df092557e52b871663751259325b9c92bb1161033c55f9a3ad188a2c7b7cbf8b8ccb7b68d3d5db7b5f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h27662fc10efd41c39669e9dcae7f65e317dc2a8e730afc4846e165acea7dd332fe9076b65a8059b666d34a83eb882be935174184f5459717cd6e40a0c6d5b3bf6380d69550eb48b9a6354fbf9014da5b981218d6a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h44ffc68cebaba28d1df1bcb735df654e19264d679297ffca6c6b28811aa36eb6d34fa3dba214bc9e582deabe1c7cb18d8010b1e7b659ea3bf790a0b239a6868e83732b8d817be643b295f1043a3b3a3fec1afc057;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9130ced59b92eacbba58cf677d9027d4257a7bafb80e7e049f5109c78ff5fe3d2b95252a9d8dd3a1584983ebe48fac8de0c75ba1ce49cbb1e3f00a6c81c25ca70ba3cd66a3c74b7091a3db0fc56134f3d864b22c1;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2583e507a1ebc61bab8e465b9a8485b081d81c7a4cafb922da2355bad2c909e12a076113fd737c4407e552f50217040079e1ab31fb0d46a6f6fe205612039f97cce18697df7ac529c11a7082d59f252c3cacff2f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hda2a41b0c788f29a5d05e1a9fbf7beb2f3d0d4e4b0220b690f4b919a1da955597aebc80c8b968e12e68e6432dab4848ac513cdd72ee1073bcbcb3e2de8e9ba6839be35c3454a38cb107906dd19321159800fb07e;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h73c93428f08a26d5ecbe2d25dea39512e871e42f8b676bc4c12b15e34cc18dff1a5ed352808ecd0e2bda25787dc453d822d66d5697dac739e063fcf72994455f5d91b5ef4662d25b9bf59e457c7c1c4f9fb226645;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h14c731ce61a0ea7522d1b805020c6b411025b2e4590f9033431f503f00eecbdc0b2848dc122a1c12c430a2146150cb3a975131285f3a0c5dc9bf96a88bec535e3d10958ae78ead012d2169fb44a7fe21536cd3dc5;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3aa38b4f219335e70edc707010a64c5a3c7753abe48adf586a4ed452fa393303fe3378c856393301817fc4ed581992b8a13b6f8a04ffd94c4efdd9782261dc50d11a6f969de5df80e1327c9477f9831ee722e276;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1ae69d53a5d36cbb1dbe72dfa079c833e69144722a7a82cb8c3ff1c5e93a1bf4be47fdf7d2aeb1122bc2555dcb7d340d7d3285b1a6fa0c4f3b3781a92aacf4d4e8e2067b5b4d618fac61f645ce0abcaea4028eb54;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h26520f47b9b5836e80211828779065d4db1564dfc77740d3289733438816568ece2d8156e634f44e88763507fcc603655a6d2287bb41d313327056bc66512a137d970f3690246b69d15dca2e41734049ae1801153;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf2791b979f5f1279b73964a172e2345eebb836b3d893334946b9b650ad8acc4d7c73d8f835269372bcf6b069bc8a394e1378ca57bc0599b77bb1ec5069532c5a27730e02ea02b2609aef4aee5248c6511edee7143;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8f08267d3e96498506fa9a36c3a5d90fde88278328543eb0bec89b61ff222dec8d5ef434cd25aa28b6285945facc979e2d213271e82a8ec6780e5fcf4139d980ef348e719c04a1cfa0630cd4f2cd20bfa92a0e097;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h20fe4f5800af0747d97f95ba2b5cfd04469f761c15419d417cdf4d3dd169364c666e171be9c0f79de380d1aa0af80bcaabf0a840dd4d894753fcbed34cfa625c5d895d70f60e65e49fceb0a1bef792ae8638bac10;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfe3221c58e3caf4b868ab322b68129b9302ed416f5c2e144de5fe5ab7e258080bdf0737e2f42b1e14416bcf8df0d07678b7c286d2f4e55f52f77a83319b4908820c10560dab3cf7af7245734d514916a394ca80a5;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3749042defd89f70ed91f28722b242f5ee8a516a067a5ca44e4189846967d381d4c70efb880485dcbe191fa8ab45980203c9a4d35f74b2395dcb6d34e6391e5130c8b71fa87700de07e5c1e7d9de58d9294670d28;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf3fcfd9cae1c27443809ce03c4bbf59bdde46509732800043ef9158e2ae29e228a0194ad07cf0778b729b095d3e3e67c9aa544d3b36b8bfc19c01b07ea8a0d53cefde12990c0abd1f01fb84a7b578218057786bbb;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4de6227bb662461095be60a8ed518c41b4bdf4eabc1f408f7824886d066427bbf1a9254d0526312b2dc1fff3f218788570dda09916afc9cc5b633790d2c2d825a8604c450fb60ce8411514188a07c2fa300793b21;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4e74ef890c6f3670176b964ec99f3b1341d05020716ab4f1197004a126884664e7556e42d7c1cf5ba360ba1d38b0b9aa4fd2fb3d905a34c8995779ee7fc6f3a41cb8d31a7b6e248a49eeb832f606d013b4af5130f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1522da65bbc5f9ffb3dc9079d49eb21457675ead703db3cac94ba6f62e9ef7519811abd4fd02c9b164a416ef4bafba6957e49a4df2085ec2986481fb32d273f063e43789d9923a6afd439589d0de82e75e44efd69;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb2c94f0e4fe4bd6f197868bec17f36bae7543098dc78a78e392cf6323e4c962030ca7e14603d1c0c30c2d2a9081b15edb62c0833699db8bd3975880b1f2ff56dba95d62e0369ebb51623f6ddb58e9b9c5142108f0;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he45ef97ac018f2d72952f04e870d0213f9dbc23668c7f2815fdd3cd9fdd3595926230555dee927a2b2f2b6495df4a218e8898d471a95b4fb7911db8446cdffde58f79e2863ebd4889c9c5d9d7ee3285cb37ae8b57;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf192c68eb72de176d88615a22697868d60ec58141f984b55871a55438a85a650fb257f3ab0cae5987af0eaee31b416160aa14119c9fa32605fd356d07c382ff8660981777b7ba8e40b5528323697e79f41cd2db8a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h539287146d1530c302cce528275965a42eeb565751c8232e7f9fc733a406effb4b90e395a1d1e42e53da13fbd16ac940b10162a3669a193ecafa274a9d61616f258a2404e1f3190dd4a6c28daf44ed3a1fa4a4897;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h867a352eaf1ffd5d922157beb06f25717226f2f50abd99d422e0802a9900e4f995041ab5a74d7788ead82df99a8de20acd7c4c9bf4a9bb1bd81cb31cb6543dfc877502b64525bc9d78d4f33db74bb9125c4ea2a7f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5bf911e4c2ed16a54bbe3e90a3fba93ba2c58beb7081f73b433987d438f89bb72fa80751861fcd8e7b8f477bae12608af96a00a23ca4f0821acc4dbbbd95e5fb1f988dc0d117b43be912ad38fdd3c0cfc839a867d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h31c3e42f0f20e9b8e9fb88cfcd50cf615ec25f6281d564e91eaf1deb2a2614d3d27054a989e2050c82303b6f9475b08831171096c3c807afbe83ad543dfcd45bceca18cbbc8750b5639232a99e60970a1f357ed73;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9aeb54ba4ef76be77a5d926d0f990ab9692c724e2ca41e205e6403b7601e84b5f036a30fac5e766e3a790f3d7d62988746aa44210a06ab8c2bd19e46e0a6b4ca9403a230fca0120ea8ab86b64547b8465de1a5515;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9aafcaad9d8088916746e8812f6b6b9c10f127ed76acd4ec8f6b2fe15415225f4009ea450f620254a66154e5ae17fd4926011c04477038f828b1439f896d8f25e9a5851cfa0124a386c394d55118213a504e53f1e;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4b515c9744741b02fbcb1b1fadd3c57c6dbe566dbb9c2af6f71a261756bdf69f87562d5e1612f7ed2fd91e32384ca5dbbc3f0027b469baa53405b4b8bac4b406b36356fa766f41e7b33bf545895252050379f9ba0;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h73e39acb43926d46da0427f6291922300de08d3ec14f2f6be68c6d6961d78a629893ed674a6d9e2c44b9c4ec68b3dcfd2dd5138c35b53b5934a9e3d0f0b97275cdc43a94340ee75ee7e52a24aea0684ef77df4259;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf7ddf0bb6907e3e05c6f3c8bf7c5d90add67df59339eb7ba628fd853389a944df0eae858e3fa4a0b1ddc10ade66c4ed117160c14d91ba51ceb55b5280d1892cab1f5e6fdd30d1c3ea06785038cb0087ccd1f52f36;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h85e896ad0f4d94a55de461e0d20258b65127dd0515e77061ea90dd56c71935929e1edfadc8cbfb2144a6f93b70aaef194900203fdb1a3d8d80c62afc720dafec2a5619728515642239c249f3dd43527e6b4a29763;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5425c32d421b9df1e1e7c60c736178331e7ccda97cfdf2c293129684575062e1cfc9192724c0ab3885e11fb6c7e25bf547e7fc09ef127809f38f2b70260c65a1197e8500bd87655e14b2f15a7fbe3c0e8b74db07f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h302c3555d0d40141551776d9f84a30ee3feafc7cf54db641f0b4bd827ae089784101303a8e012ddd20d8bfee3ac138af2695767546686f66da6d4b9fbb4fe76ecdd7eb443a63208b859b5b2a097938bed00bdb76d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3ea87e90c31cecc53458bd8ccc624ca3b18adf2baefaa30c2dffb4005c8080890468840ba20959e9e1524594f1c152bef7f1164d260853db324a9c2c2a14360d9b6516fcf4022c7d2fa0ec9b614e7f9fcb53ec835;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha6cd7228cccd3dc7c0f09e437f25586a8025b94c7aa5306b3aa6c7de7bba2a89b877aaf8ad664fd3c0a98a21887f385bff085e672ae781d4016ba21d3fe511f2adc256624fadc505d794a2449eb7f6637439049af;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9ff96ad38030a07cbdd1ab930d2b43a708abeaffa94e992a3d9bab78f646a8fb29b51f5e0176a19cf4bcd0aeb1380260515dd672f8cd715240c717296ece2ab43c25b11e3026199486496ce2378b6533b9c0e2587;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h788a538e56f6e11d1a39a340d007d46b7c65a2056a99879be5424c7892819159001973c02e1fea1cc6862d3dc4fd36843c63ae6c46191b7be17fd426d9f4ab172e0a5d25cc88bc096fe27270b0a1a42fe24083a69;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h43334cd421d3994ac7346106aa67bd6537c59d512e0030ff039a533543d302925f44517c019f0244099ba2ddb1fd5ee8d3255ca161fa9e76de4c1f933e80dd275b9760f5514bd60379e24389bdaf4ced178abe18d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h55446e4e43048cdaac7c28f07e85c965929d9f44afc40752a2625baa64a7e912d76bd941b8a67e7d4006ebbd4038c29de815fd171383cf951a446753616e0eebd5d402007035a6e2fa6b15505a16eec54e27d83e0;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf3bd697f79507aec113a541c4583234cef1fe0bb277f459331a79781dba5326694d07fb96b85e8fd55aac8c1bb6485c17ffdfc5bafb8dc4cd9f2d16d8e4dd7bc2c6aa16fe5907f43eb5252e86925f443f3b443067;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'heb56ff0035ad03dfca3c449c9e0bf1aa59685e7b6bbe57219243bb6a6c3801679b329114dd6ae28445dc6cda3cf5a651889b646f2182a9eeea0fb1730661781dbbc4b80c0b86850e8aa059487986d9f4534cb2cca;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9276159bf1f9008051d1f80af92a7cd199e3bee179d60d3374cd60d6ea8403ba55f3c7412b62e21c0a55ef1047b78db5a2ba47f29521714c7470c3fcca6edcd122ea032a721a1bdb809cdb7414b118ad303b24f97;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc94a6d82d298d6f4bf14f871e9a42ba104392a5757c1d43c40b62d3e21fea9cec503f558b88eb0cc1a1a106434cbf3dc324e717ba1c964f4529833124322c298db00c1438b2bd39bfa6308af9eb97a7836b9df90b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9fef43d073d59804927603c298704bc9b24585362f2bc7da00809f48b8d41fbcd48299f169cdfb9200956331d52f1d7292d9de9977971a441e0ff4c5045c5c43316bf86f1e3bb7e4fde7b8355cc9f8db997a7f9f5;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7d957fcb0de481d99a77dad13f363e6ed7263befe5d2affbc3e61bd9c1e14f2857e321623c0478f62ff1f85894333e27f6c5a109b68b17848e710e3ed6ce5290d15de538dbd2c846f9e362b9107a55b6ee88d6b83;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1538d5ffa12f0686e9c303863a830624ff8a2aedeb642acfcf186952f040bb95b20eda1f35fb29d49a97829da9cd7e0c854558f2dad989a476479889ce1c0c354dcfb4f77eb3dbf50a9e3d39f56eef734d7e1ad02;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfcfa206e237959d510a0de5aff981ffe1222fcb375fe54a2298bb186dead9551e20c04d9682f20344f2aa71c103079990085565d1ca008ed72883db7fa47834639b62d44e3aed8e220b6e20e39a03c6b49faaffd;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha434599520f68aeb7eb5c940c42e5edadfbb9e2a614e1c18bcb4996c21a19076aa10390450680c53f9b1cb0dff214ca4de7b894521c7c77181664154960b565e339109855e5c2d51f29eb39a955c7296e122dc0b6;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h200897a6ab747b5758acfe4b8e700e2e372209fcde67943923dd1eddaa4dd8009726b395780221af7b84e4e1b11d404a024ce5ee02e3ab5e5b4735ebf9a158da4cee389b94ed306f9e158e4b7c86e29615e57d873;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8e18e76f379ff581644671949b4df8024d51654e9870d73c37385c79adba18df29e0c24c822d696690886062f508d34a26a91b4220ebf19d87fe59492f7c4c7a78928f01aa504709a478a1c28228a1694124911bd;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h92a10d3fcc152b23cdde833712f0b7845d951084a0553629d3079d82e453150d32800f3d1a5509d28fd8a5c4ec04d077aeae303fb01e0a5afe3925de8b38f76b7d4b44702eff36b52984af68ada69de2162f7c2c1;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hff6437ef9569053fbc5531dcbf4da93175c886f1f46b04f8cf6801395ea699d673e2513b778cef5ff324e079278bb54b4f1d94d665898b3e49bfa549010e1c828f85689d5c5c902243165b1e5436f266518abd614;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb796af5fd211b17b096b1e12a2c315dbf6a021c533d5599cc9eeaf4d068f6cda4e98024fe99657832339de19b040a9e100f5e03f499e6567819f5396c0e722d0860c3e612a606a288d7259bb7530eee724b6af9af;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3f98e4744ac18fa51261d9309520bf0b50f54cca54d089568648d33f66fa74a974d23870b8bdae6b4f2a3f5ffdb7d83599bb8734b8c02ca06c3e80fc0d82c03ee6b1db22f9eec4a9c96fb53feb42c89a3959e6971;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8a08253e8cf4b0128258e29e6c0f3d154456dffc95a305619a9989a489a9884cbf84c6d4594fc0225550233a8246bab3193572a2c697a23a4bc5dae86f48f5ce36548ec0737ded7eb193676812393ade6d830368b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h40a2f20af04c73698d92988f7b5ce48258d07af0b2e4abc3bd2950f0c61b0ba07e408aa27cef8a74463fd5892e579e4b3370d8ba17b0bec7f36f92cd4e3a0b253dc6fa363aae9ae0ac045ac952af37be798077590;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h37bd548667260ef030f7335def538d2c2fa09130c64c517fd566ec53e4b24a9c2b3fc7a4d55d81179983ea011fdbce43d213869da9f2e114bb014d7207c221b116dad6ba4958b9c00045d9ad409f026cbcc6cd65d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h124ce3f374247faa0bcdf23edfb770dbc17aab1f113d8ea569c33bc3071d2efd324ed5ebd6d7dd2a399f0495bd545ae513ce3be5f436cd484c24fa1f5fa04c6fab34ec0f4271dff1d7796f400fb73ef07897508a3;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb606c5f51e22b42ba4da87be4514b748ecfbfaf3fc33baf44bd25cfe9b520249efb833f2959c09515b85ddebf9430c82277f10e86b6759d95630d4dcf04041e7dab8407ce16fe48e5c6d3a7c40b1fec90fbb3f367;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc4c2f586806e00429b2fb342659bead6ac191e38c380a18ca736a08274aeb10dcc38a3e4ac2fa51c482b351a049547d759e03784d78cb20f20ad2ca73b3f9bf1244c63af29196c744222f57b5d219e57e41ebfdb8;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6e50373476dfbf9f688352fac917804f1ed188d5c4a0155fef960297c609d910c3a73b0b5c807ff542b3a0971e16f01ec25cadde7c33646e80bf09cb4d40e4d5674cb71a97017467a9d3b5e722e426f61d85d4c65;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb9e6567c345cb47c353f4d22025d93794f60c0adab57a7cd4b488145538980a14b41054094ac3f47c6bcac8cc09a923e4a788313926ffea95a792e56ed6e7d651a44ec91abb62e612f8944f92111428bd70556743;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he0cb980917b2b979c6818aed613e13844620c6d127b67c97312c2b1db5bd24d5265c696436179c40c446b2d758aece4a9e1eff044c15bcb114d6e40ac422e01488cd90a3142801d89652fc6c2239cbd2333d799d3;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfb4c81be03ac63257d932f8978311c16a10c16854456f44dd60414b81a37f5f3a4c28bfb93a137349d41c026733b5038636424c8adbb00c0b21b3d8667a2613b2c6940a7be2caaa4007f0fa7cadf6562e278d7681;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hab6a55a55ac8c6c1cba7596d24803e108b98b11d5a43486242aedcdf745ea592ccd3cc8cb79733c7c55d228501d25feb0a39877a4fe113702798e1cafd3e5b468d4f5ca4e1515803f694db7d0bc5485a16cbcc60f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6c8e48f501fcad3de0cf186f4976489969dca65c848752ecd7f7cf713603c49dec8daf11534611e1f48bf1d4f1837d5e7c0c53598083329eeb20597b7f1ae36aa97bceb72e8b4e27c537d52e8fb2c450625564696;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h965cf1fc167483e9713cd7a3aec6712662714fc335de4c605f7ab927a65a66aa6c752fad834753f5cdbcb9270ae7b8d7b4a0e23288e37b2e312a6b223b4a90f85ba7aa183b8287a82c574c8c79217208a43d8f44a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'heeac11f9db68da0475e3d91263895fe587ea70ee279fc473b71582c15680ac5780463231f0fad286c869eeb3684a5175255f5bd8048bfdf314eba4ecb1a88df4369bb50aec60eb08dd5481c9fd0070d7caf127629;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h996ea3ea54ebbd88b6b8f54ca561992e0c118df9922adda60a5ddeaa5173e019abdef80a1ab431c2f261c3c8243fa94a15a92ec8aea927de2a1529eef459724a67be76575167181dc788d95b5b6cc5eb5af2407e0;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbc940e2dba5533bbb45f29bbe5ef58a9afcade63b9b0e3a2c0a2166cdb81ad1f5e7715f4b99c09932c54a37846a04976404c387268bb427a3f5afcef9028baf61bca1d09c7e0e80c7e94b2d271c637f750b82839e;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h31306c89142fb0de10d2c48d0ad48f6df56d1175f360d05fb4e4da1d09e04923a219cb63691e78d23888eae282cdeed97d2a33fba152e8fe9e029548d77710b38cf01984c50f305d63cf962d1f02e110f1830889e;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hec772728fea7f0317e04c7643f19aa337b09d18b96056ba7dc7ac16bd8382d9905e07691e5a5df5303aabc9f3e3ca98ac9b392b4b66618c86ef814fd79a76f4e29eb331e51d48cd64b255ef8ef230c45a342e22d8;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he360adb7b8b0a6b12a3e70fed20211f7f7cdd57e4b15b3b5f8d639d6749e26288cfef445992fec1650bd223786076d4961d7e0099846d5def8d5f2e9439fe2533fa83dc8dedc311c6b97ae2a755803e23f17afad0;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7628526947225f8d1cc43b825210b554660c3c145912b3e0e0977e91aca14f1acc64ca3ca38f3c400f1dca4665f23d904ec807e9aea788d0adea60806bf3d435c02c471b0502e6bfcb78fcf2490bc976de04d3598;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h474045172dbb886e34491a0b0e108071937a6d48f5bd185af7ad04359d62b217fa96625543d1deecd834bac51ddb0fd34dc66ea1087c108e5b6f444a49324bcc66832ade37e5c969ae331a9298e18d6a68c13ab1f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h20202a88086f3ac7b75e7b86cc06c49015fa242ac647559702c1f8b5afa80d73f791722ec197ccf5e35b519d2b41882478bc6aa868754ac455b35399d9327f5167410ea9724bce8b45f732f2558b454e618d1507b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf85398256377cae1d64b75375ce3f540cabf10796ed7020cb138aa220edd386b538de1be3547e43627300e49d1823502552ba3e395ff8356f8e9d4654f5a8a2b6a3ce329223285d3a6d5b50ee3cf8bf6cfef01348;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h43ac4a9224ca3a04758835c81c3f40be7f25ad3da86cd32b764bd3e8bcbb2a98c0b107e85690299a03c4aa20d3d70bae6d73db5888ec8cc2ad79651ee809270c074ebbfa4109a72d82a2b2c5faf201804997ebbe3;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf1c67e4f177ff620060b5fa7520704c86991f6c85f766a57b4ee158b07be65d1e82b3f0d2c04f1e3f06f2bbd891e43a33ceaf473705cdf3968bf9dfd328af6e897b9febec83d8480495ce6409f375704bd4209c84;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3282e08d06ae041235d9ebf0ed1436ea88af85cd1bcce48c21801cebf90f3493475663c99f21521db424b562f4f0a903f6a251d04a68eb12ec6a4e15d101ab91768393656bbf86e63943aaf9c7225b7bb21204b14;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb5b1bf83ea32d0630a77f80551f3c96a451d9fd8f15e60f7162a894558c8a91a285ca5ee4f69d8d4f7e2cbc47977624464268107a3541bec407a8c6a01b0f3b86f6f5139644e476f81cbebd91e4a8e6455551bc7f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h54cbae8a9ec8e6bcfbb503ad0230d2f8207accb36e2c6a69418bbffec4ab72e7e481f5376fc44f0e4c98f65efb2f4159f84d2f042d944e7d206ccec5b3c2d558a8cf15b40683fd113505f4ac54bd00eb7b25e6e21;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc8d8286f3d85b56ab076d2ebdbbbc20caeb7d5621615aa5f42afa8e1d93278e16746e9840c0e85051423e797a1949028ebce98252118d0f106c2a599d0bdf0abd8d1ef2ca0457e4907e8f188fb80a137cbc95dcd6;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h10bce4603d29828f20917bd8c947cb038e6e8f2da2873193ed8dad68568249543131f6beac3a28c19a9df865d9086686510858b71bd759b49b5e1db5725d96a31d665767c35d8a0de72ea17712adb6db9a45bed69;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hac16b6ea70d5141fb41b58c8badbb5f925890d06c69ec111f57a6e2f5a01299dfd4c619f40d674c9f45b3db1cb13d0196115d0fb0f0d192b19500860fbfd1db39571d37c418fa27528e370659f98f751b2f887414;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfc8c5d7d119cc558fa276a920993c03835746e0577394e3099e9247a316edc6e803881a2787f50de30aa09dca1359cba3b2f83f38cd8d769c96196c9f3e4bc7cc2340afac94d422656396a2515fdf7f4460dc3cff;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd859443b3afe7fa5b59e38302a417404ebbfeaf6927677f9cf8eb74faa230d4533143ba8a73bbc0388308c53aeae5b2a39a0236f0af0c5f083092ca8f7943e45f453fa6c52849a0efb673357178ce4de94901e50b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2a84fc2718404228f1153eed0e44210fc9351731c64cef9e474f8c97441aefeb06eaed3e018a1186ee3d9020ccc87b9941eac2e98f5b558d5a5bdf106c0ee82624f40c1d4caa9d30fb9c4f8ebd539395ad3afcb58;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5f97c06ae1ea6109f57c20c712be838abd55ce3817439eb5365af512d54fbb4930625f5993ec12af72ae0d1bbc3f9ab267f5b714d911955f9c024ac10e365da4541e302c60a7fb97cd684f7bd7069f0369b20f105;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h63025f58606f8053841a56bd0797b1d8beae1e909026d16548a8b6108c8991c579d176181a1b517094ed9a38daa27533a2392defe1c9aa0d6da8b8ece62696a3b0019881d8c12d0c1d5d8878a1da07c8f424c896c;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha9062ec02a46c84b8d7922f730ffbd306da7f638ec5251fe17fd024c1687b84c007face627559a004d04dd37de0ee40b08d93d6f9514d37b47c657158089830548e2625832ecd842cb3416b88813098a811d4385b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6bc9dfa2e7497f52af7cea5f31b8ca9491d35851b3e48de2d9ca7a2f0155c0a429d6f98ae923f18cb3b7001158c23a8b3d83bd01896511401121dd0413f73282f5faa48934b1920df8045cf4d01fd43ed507355c7;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2b019c2eb36dc3035670de3d1bc93f8348ad12597c3892d1d1b8be543e38216fe57ff1de796703b8b15fc870b2ec9ecd5455b67ce98029596171f5b3f95c8897a3121c60770cb8a0dd339179eed72e5f8df2bb167;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc3ce85546bbf6a2b0b8a855c629e173d639195eff0baf3ff5c28f76f952b26d7e6c3c4d579b691f24d2ea16c20d496e1d2fb8c849e0d1f946a4c94b5396a6fdcbcbe55cb6b7ac820af7cde6477c6a9de8af12d80b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h68d5a9b06235bf1bcb53777dcb404422d5a593e964b132ae173995b7191c0660a61a2941968ee537c6e1faec9d048902e989f495a2c0c0692b5941468b78e36253994d1542ec9e887803501d6c03522023b19b94d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h97f211ec3d4c36c8b44bb24920098000f0d540e2c238b64ad10b01a2a392a68e60b6e9eb44fa189907c6a940b8bbbbde699123cac4aa7bf16d75a53a62806d8909e21fce6f493dded41eb57a0c38841502e0e01d3;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h154bb0e172439b0840e3be78c050f32af9add957abaefbd1647ff0ba6213f5fc4a65d5157b83b7b7806feb480343affc351621e187280a7c83beb18d2cc2778b86dbe62377d2c9301149c54c51f99a7738e9069d9;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h49bfbbbde4d08ab648ff4e95887a46314f439b31fd7a5ce94ff84915055ffc0c87c1e01fbe52e7ff8efd4d519827881221f550009f65759a08be100f9d81793ab4796910f157a742767986a7f78d9f3c8efcf1331;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5d4bdd80376e0864b1561230beefeddf5a8fa5afab582efb3551eef6e6e4d3bddf8353899831cbfd545ac941aad53a3b0434bad89252f69d366cff799f3d18fa43238ed6654af6255565fdd71a36cc60d020c236;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hdf98dc48d62b1a5a8a950eab5e9a3dbae037e72ed0284b2fe41352fa215abc38170f4fc6dfc89831e4bfef13c2fb2dc3c64dde6df81f49b6cede59aeaab8afa6e4b35ca7eb3818fdba9d1e575697351a6d76e0e33;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h84a4df802bf60fb34a797d71bd6c1913a45d5a17fc440f9bec5805b9c3ab04aedc301d2a9cc1b4eef7488da0c88f11968e563aaa31cbac15a0ce138a7e77b71ddad810a8af3e4856f9e6df08769167c7a80f15e42;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3a6b4f9e567dbd17cf22ded193367f37c03e082a37c127db522c6ae9bdaa684addacd894e0527676cfdde662cc9453a46128c235255907964a937a40ab36f9f40e761ca3477ec493151301f73c7cefd44f5f515d8;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h65b27894e5b2e67759d7e929a9cc52a7604af9a809f7d94faf2b33ea872fd0a9d0e4d0b3c84bed2b6908682bdc6267f9a424c2cb8ce737b7678190ea1b760aadc834bac6f28fb9a0ff31dab36e6c46e6c61d6f4ba;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5ac9cb24f2238e87a4e1fb657a3591e32b705e0d8f8068a5057ae84c16ac552fcf3a84d0a60923c11368ff9eb5ae7012e0cd611dd494e003720e020cf49c0d3daa4f5d1be977f074f81673ce7e68ed2f378f1ba2b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he19aa1cb4c129d4263a7cec31c9ff8d4ab07d564a0b42c89a8c8e72811ba27800ae36dc470b74bd94bf017372c988285a0a4e114797f4d8340262de4d687baadb99a7f0f2f69431f5291e219ec9537ec7c5b2ec89;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf333ca05e5bfd6cbae7d052d90864379ea0f65ae6292f25aa126fd51928bda4dd30366939747d257e8d34d9df9daf972ebc8e4b7c3fb07c848af8030bf9a79a91d2a5ee1f8e19ba83b6308f43739f6c1dbc499a41;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hdb41e127e2f8eb99d6579121f4ca99f92f057ed505192d8c8fdbc7a59ecd1ee314a5d2e773bb8a37d16fc5963b532174a7533b04ff453f569edfd829c9f3f41f9a3805a931d7dd28b6efabdd067514af01a5cef8f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6ab13467b6d688acf8ed8e6faebda029e0dfc005fdd0c9dcac731e9e1c0882170117e82fa7bd0a777424440e1390d267ebcd21770311f1974c72a179d021fcc9d0915a026d3e3b5ebb6fc44991af05c5bf285de6b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hdf8765cabf1e697712f84f882fa449d97c205cb50a85cd717496fb730383cf27717bcd1e4ee685331976721015d0cb009bf5a908d6a19671b99e3bc674767178905520002494e8587fa0a6551c5225ae93ebf025f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h231e2c0355198c8c34bda9f09027861edb3fe83e6a07bc5ea925eaf424b5d71fb6307674692df313cf4337602ef3c3ea66a5b9ffb399d6ee65ceb099f3e168057573966e809ab802a065b13d52d5e694ce72d6dd9;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h303f662bc8940d50676c1f2672e725f70a3c35d43252d9d6c3a918ac3d0e61a3e8e68186ee88824bcea9bfbf7d6da10eea46157a11e912e7427f7c2fde9b64c81aa51c39cdd918ba55fb1eee159d9c60ae120eaad;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha7e17133f0986c7d53e179f55e177ffd0e7a91e0cefd1decee1525ac7df8a5877443ecfd45a2b6dad59a55ec5b1ee7a2e7de70ddc4e38bfc3f5d8ad5b5410697a796eca6455080bcfc1b723f7f33855b3f8b9f38e;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h617fcdf0f36e837b363ec5f6b966151a8cebc2a2db40494bd75392762468671e55a2640ab494cd723a1cc6e44fb5e9c964f80ca658f2ce007d11764d1fa6a04a08ce7d39e26da9f2a0e91017b3e6afc08b97cf412;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd878dcb0490a713edb72c921feaf49ea57ccffdafc3295a33b74cd461600b7f1568cc4a26144e92a0d9c8df75bda114c72c385ddd4417437259a6ef3cfa8bae0fe04d7c7d0c3ab47e7ba5b7185acc6b8828df6a69;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5d6b9757cbb73352d1f263206eecd52a55c76dcdf2836b38c7f7cf807ecd61b86f16a90835bda59f2569ebfe98ae52254245bf73d0cfcd1a5a88e6dc3414683ef775fe5a97b802f7c987c77dc4410e719e2a85d34;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9761c6b820209b9c88b057344852d6d3e9ab07776da0b078357dcdf6ebf971206245a37beace842c4be0789a5d776a48f6ce9a0dd51f95b89cf4174a2d7bc4e4a64a7a06253d8550cbd1cee96b882c9f81f9c8a6b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf32b3b1ffc3cb0db8dc5cb5e06a800715db585280da0ec3555f79b183052cfafdfcda2f9fcf1fdcecb83bd603b22318318ee1ec3a3e55ee7aac2553a7930c4380d865fd542e2a0a1d3eacf4f9bf9de0168f6cb09c;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hdb1253d744f85527e4f2922ded9c338cf7b1995350fcdfc2fba92a3c10ad6fcb3db192ad09d0fb2c4484b7969b02c489e17759c4141fe59a91fa901299c8d86be6e6bcb964e2850fbe23c5d229cf488146e35ad27;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb54e4467c9bfa0b28fb1ec3d276b11dec9b53aa95e265c85e1590164aef309bccde3d06c3ea3893e41c1106dad741655f9f4ab9a5d2f8e745f66ede306d84b0f16d080a675ef50a9b7ab7ceaeae21080eb6041f6f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8cb02999abdccf3849a0ee1ca0499bfb74e657b2c07a467cf7240addd69053aabd7c54a9876a16f8c7ae591a733a0541e36b0c3c6a247b01bb2753071fa02218c828c714d66fc858b1dddf6dff6cc630b24e7b98b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf2bbb95f37c922754978ed9201d6b8e152b057bfe27c037b5df9d2b09ddfd8e2f10daeddc467e0c1b0d5ddccb0adfbbf5e32ceeb3bb6b4810475b44440a566805150a64d963878d1e2c2e2f2b0792976cbbe5885b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h847ae5530efc9ed6f6780c6b33373345f771e900b7ac74c19e020c6bc043c92b700bf06211ef70eea99d757c310ec72a04e18b151a24d6357917e63780234059023504c6ae0449e9253a8b78444a47e3a820bb535;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8dc8f20567b14b005457e84a0dd1680f75baf4541cc8e5370f35cc1eb54ffcb122f2ce23aaffbbab995cf06bf96db59d5dd9dbc3813e5ccef19f7419712cc7b5825a3903459ebc181feac3520f2782bb4c0de4fa6;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h52e38e8dafd93012bd434104f511d738d616948d17bb23127b50cc3881e076dbfeabbf9034cc066cbe3292607e3aebd4c408f0cdf99f09fb595023c6ae95bd450b410210adf88c19049c65d3d0e24b17fdacc0f4f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7c703966a162b710fef097ff5e44f43b352aff6dcf46585c6a8a94ddb9033fe4115fbb842d031b44435ce164e4babd5c7bc88ac0dd9dbe2fc887cc244296d8e472634d61cc3079eaf284dc7783ff2302af8d37eea;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1ee161c91f9198de439f49f968ad5442686e7ab5de5268149008d6309a6de648cbeb22a463cd09cfdc140e1708ab7bf11ff58ca4bc9ba04dd1a508203cfa0c5b6dbc7d54da7273786e66ca8c6dab903c8db564831;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he548e3b4fbbd4cda1918733934c01adeeef91528d0c9175a069def406939ea39707baef680485751b728487497a54b2bf916bebc14f42d95feb7b36cdfdd4a4a0edcd8795e2249be5892b2b05455f18d243aaf821;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he47423200e895d90ea3a4c8772a3b8e4f25871a2413ceda1e5f10899fba6d9b8f73447710e4f3e0d15d4996f803bc688d216a73fd3cd743749d28addb767736497fb18dfec609dc5651d4a560a0a3613bd8b14028;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h18780069788621a3183605c23e568e430b48f2fe881c3be96d23b885e7fab536cc28683929a7266fb436b78149232e7421644ffe20a2aafb2d9e701ee991970356a66dd20012a9647dd39fa229f3610def1535fcb;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h10e11ccd50d316b834857e0129fbe219fd390bc207196bbf7363151d12ef605363f9ffbca8c0fcfe9d597f8de2d29b36a04ac5dff7edc4165c0eea4425f30828b86a9f34357039f6aab24f5ddf0c89eeb5c395dff;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he29b60ebf2e095a377aff8a627c48b988a164feecbe31b537e10ce4f206faf884d9e806f8b9ce047f7732fb8ed2e2af118ebdee849a02ade86086fd1cce8cfb3e53902adc9d5aae2a34c7fa2bf0f522c67a7b1049;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h51e166882b432d5403af50d7bbf4bf54536b6308a4da9c42f0efa1c72858cee8f05512d781df8b13a7ab6b06efdd5ca4f61c63092f0615b601fb1895bc386aa8eeb196f1d8ea72e7e349b8082183178ff0567b37d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hcb6c8ecc48148482f534cbd6df0c29f718f347b11004242a86662c024eeb743b5afe7d8c1d28973f414c81e730ee04bbbd99d708aba09783aea0b57b16f65642f2b8c0f637adc94967d85e9d2e86393d539da8a9c;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha2600c128873358b0c3ba59119754267051036dd99ad7f7eed0b141e1b3bec441976295c3ea092cae6558b7982132298d7074831b41169298e16fce5a75206b3271ed6e5d2aa6e106350892fc89b88c3699c848f4;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc637bdcf084be4b206769e336c855055ca3bf67007be693b684770fc00ca6faf7780b8c70c91f81f30a2403bb86a6f6d5f5f0b462a3f9b0b0651ce9dbfab2c918aa24ba19ee9c1d940dee89fb1a82acffcf45d7af;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9e263c686b90958e8c734f905e691214445bc438b33ed1484af4674a82d90d54e06a026680264ddaf54f6195fe799eec56cdceaa76df1d69682e63915b0eaa1838f32ce94f2e2fbab2bb1b7a861d71aa8fba75b24;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8f626b5c7022e3e7376d075bdda04e7c322f312f1f8da83d514b1bf98b2e0f7b516c416e03af318dd2b6b2866ad80f9269f28e0850e5b514823932296e13ac1b2135f575f06f9e8d08dedb98a938c9bc1585530d3;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he4292408f9b78ff2517c30b21d025eccb974e440bc61cd89c4c75d057e3aee16adb834ecc8afaebdfbdf78b4673bcef38d1555f49768bb886ff314528a7585e89ee49de73e61bbdfc7382eece16ad1d1977afb120;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'heb06357cccc63097f5ec1f9f450482da80470de7188f6823e2537639c54530b82b90fde4b977df8b2092ef9821ae2264bde190fdde0c2a4c0cb85e23bc53ded5662551ec41cfea937b3296e46de9facece9b3f752;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd82282d9212da1384cb52e6c5d702989f041faa19f9fc2aeae3ceb749d53d59a3f71b007fdd8c6f03a3da5f01035c81288407d89c41169705c48e6f3a642b2782d83d9d2323dc8034256a1a4cfd59ca381a81852f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9752abbd9633670cb2be4dc89ff6fa34ebeed859ad07700d305570df513f18e1fd1a9ed425272f91d5349130545e3ad15f9a7b15bc75b6cedda6bcee178857e9e5184690d7adadf02b4e5571ff9b4c2fb33bec6f6;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hedaa38073c2008b471170a149384367c3ed9ee23266d06d8564a14752774fa6fd1e6c08e4b38bada439498085009dec707d5411c5ae9bb9d7ecdc270a4f5b4b35ea34759b0e80b1a33b085052dc5a9883ca02b039;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1387ab4e0b12dcda2151efcc0b8284a7c4c18aaffcf9332831e67925fa81218e8a043fce888d5990c0ed8dbbc78ed0e590aa06d834764496be77d82f0a9a05ca0fd0e80f9a4037afe29fe13c3eab4ce2af0d97de9;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbb79461b6f7747e058b21c23e9440174d2d84518032dc05af44d96f32705518a898920f7e1c86a37c785609c9e0fe8596ffc431ef01b668b34c4ad77884926417540f989fe289e4b54c1ff85f03d51987e3b618f7;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he01ac6f16f34df7e110a9964986324aa083626c0b1322512b16d91357c25d777057e7c0e26eab61e285391c84c5024a49de921e9f8e64fee5acd14e10dad9bce487c555609e17c961fae18e29b014f26da9100ad6;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb9f2c9663f53b8cb320b1586c4a323d6181b4f5cdb09af60ba9f36822c7f82a2beddac2d6809d7cfa1448e2dc98dc82d4e1596c29a32716e8a6ef85f5798287af469e62424b666107b218c23a568f0baeacb43278;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb72d03853ac4bb15c1dfed3dcad34acd9e78b36aea20498554b43d147d706382a037d108fb6a3b364ee97dd713e8f6d4745888a1b29dd327c135411d9a0b70ba0907c1ef5199a322ba228bc21476ec6908a14ff3;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h14678015c988fc27547d99695d0efe7333be412d12fda369f36e7117e65b99753359f5ebe4e9385fac262ec71039489768cb324b91ea21575572618afb2b25faaa809e9d89f4337d96ae2ef58958c897054061a7a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h235b960f3cdc7c43091c418c60f46c8cf5deb39b016787b301fd57e71ca2b81f3ae0c8e77195a7e1937c139488968a95b39d6b79d34361d1ffaae5471f716c12f41c8774b12b29ad25863964606713b1b6f112e87;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h54b4d38c60c56ab8c8dcb94871d92fe45eb65391f346856306e3128a1e21154dd8a05f7e3c67c4b8c723fec5849822149af8988b49a6077c9aa5f5f279543019ebae15ec23bb9316d3f078bbcf8344f267da6a134;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd1e3f2935231c4a1251264659e35ea865a10c8c114f34ec17cb6247b1f24924361826da21dde98f86e164324b395b49f85335ad99187f9f6b74032821b3a93aa781cc81874ff27d5059e07a38f882d6e0d8563cac;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6e4c05c7cda52319e07d5c8078b35726ed4157862c556ba3d79af2a93ad3b0f1c52a2603a9124a767e9f95ec2c5ef735abf8a8e36d0a538fba3a02808d5624a04f74851c8c63a60cfa23efcd6bd937bc626ba46c9;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h71ebab0e4ed6e742957bd88b958cc35003db6947b62683ef98e6424a329b26c013e50a4b902e10b0d6b7441e917cc588592b8e9ef2c1776f283b10e70a18a7ca453c7b5e2863d0bfe14bcb9321047014643ebdf99;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha7314eb48452d41a82563360ed123dc7c23023a4b1890f4dcf767b2089307dc8aa19cf0fbbb8264b2a7ab182b06edc2e96734391ebc6274fc2cf30f6f824eb690b6815faad49609c09dc0b5ae822d0837d941a260;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8eced0bbeb0cbcfb67625bd04362dc51cc32eb8172b6d65952fef0b6a0cd52d1a587ee69d085c4ef01b421b216e3b0b5f654febb20605c6915b474e9b4aeb92d7e89b1252364199d2688440d546173daba53640c3;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9bba2291aff2c5a0f23b211c68642f8ace770bd06fd44455081fd83f4178786048ea4b943c5d54c2250abb591c4aa5764e6ef1bbdb8a92e50ab1acca00aafc8046f250c1504c2c70f2b9582d86f9ae11bc19c675a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he1a3f72f654f3df69b0fce89e96917dc30a89351bd86b555afa96a35a7d8890d42aef70d03c59961c3fed15d208b65181d7f2d5ad58ea56118c4e94dc13479ef29e736dd95f334bb1b79ff0d3301349f291533a9d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he948912fc933176a904b1c1bd178ae195a150323e50a2d521f47297d6b2e5374307a3c60c6585d3d4027aa040520b7183832d6a762835e134388a0190c987f3b772110cf4825d5d767e10c10bc58f0f94e81ea61f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h66d887eed30e6f4e8936a7424162c61e4ca5e6398358b53039951fd2399d77b12c20ad66810b858e41eb5571368a34530a94197dfaed783fbef6f82852dee6f3ffcccd4ffe9954ccde443007d3f43992bea55b77e;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h999d7296cadf0a7d6d7beee169bfa69c85aaaeeb0c15b23661e55c7640c4aa2d64df5e5dc0b2e612683fbb16f5c340b614d049d82f2aef6b4928f717e9957060aed86c79e50f846ebcc07dfbfab3bfe44245a7c0b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hab3ba226d0e4287b9fcaac58fc733e0c60b865a64b312b4353e42f0428d5652a31bc3eb0c862395c92ef711c5b4d734dd3a8bbd948b44b9b8ffde00d594ffa441129244cc8a388763ffba9653df6cad114539edb7;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf0cdb68791d273a1e937c36c412ae12299f12b24c80c39b30f3eadb4a44331f5373ce9bd0b9f161d03b74f4cab753f3bd89d480010751a2e46d61efe7b17360c4cd411eaeeb68450ae4c91d9806713031c383e01d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc093f6575ac2d1a11b8bdd3c3152ff32ef3623608123c7841730c774b39a412c0dfcdf1aa11b5de7d39bd59289974996c9500614946fac102ea3a3437cba26771923785db9b1b8a83ec234aa96b2b86f467842627;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9238e706b30a7645a30b1d6ac5448add00c7ffbfe107375605d2e89b85777b5a03e18f61bfa390b238632a524d96adef1a3633af62149936b9e0af98e7eec9095d41b5c2fff5bbcdffc0993cc7850dc3af3946be8;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9be3b279fb03f9cc3b1c7bdecd00e5679977f77fad58f77abfd96098f8e19115d6a39bedba3791f10c4f76f52158090b59b3974eb5e74cf832436702c8851082b6e46fda6679296710491ff6d8c4beb4e1475cb6f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h93e1475507508c3aca78c57162ed346a03e204fc7f234b329e5bdd88c49a88b4eb2311e65a9a7f920b9858c5078666a164351bc80340f3d774f1f02bf8eaf97fac56d3d52919ff8c321bd1bd56ea07482185476f0;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3bbded5949498960fdaffdb52fd19076f8d9988a14015477cca94cc4a8e59cef4ab5c39274642898faf43e5abba705debd32be024806eab86375a52605726f357bcaf1c2968de319e3d309111ed5abe6f04cdfa0a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc566a9d6c28ec46981702427b14ad6062542c4232d81b64d1f5752c84581e0f813f5529e3febb20dd0e62f1e191e58bf6e6c75f84ad1da5c9d3d64c7975e9b9be6712f50c3dc74ff22dbb084995fa6b2ca3f0508d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8ce6f3c1ced6b84a232d20f346db763d1622a8c9e801410aa96f4660af3ccf4247a46c12284654cd583345abff2bf8399c436aea009e24ad7eff08132a53df4ef7b51b5cfd64f6ab892449282cf53792f59c2b0c4;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8beecda2090d81776fb3b2edf3b1344435abef0d3455bed949a5c5a39d49c6df99fd6ea1c58aaa699736656e70f677a15e8914581986aa1f84fb8b2a73403a077f9658b020c315c8c2a697d4daf1ac0a20a50c376;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8b2bd027e04ba97469e021e00e5c646af95b3b0700c989e75643a482f2868ae444ac1c7633db77cf45b99d4a3cc71d686c2a0ff80d63677c90001b91e62462c525643ed2153aa1f6cf19eb067b47fa490a296bffe;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8c78a29628613d56d8d379886b28402d38bed22b1f26c2ad6f3c9ec397c4fb95c6f9f01405263b3845284084ad57ebdc5c630f3e2167e54c97ab673911130a0c907c9a58272874d3dcbd38aa90f379c2d38c1d11a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9f7373c99912531d34099786359bba04ecf79392c60c08b66ce08da6260ff52a0dcc99c47de4c0e2e6d300ccbd5f373fd556cd451dac8b2fc0f413d08e14ef3f09242eb8fcfb9d25c87c844d27d3e4297e3cfaa92;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h75ee001ea585cda514e76cc66b572bca05e4bb4dc837f13eea6f550da6febe79f49b6d7f5179fbcc1ecc990932fe1ecaefada5e575654d74cdcc44d056c67d1060a7aee37f4f0c4ff23673f92a1e486c126825737;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h70a59922f57bb6f6d23bebbde00aab42852e9b02c41551257323b17ef75c623380d0b3dab0d37886566dd6f26f782647e8a1e075bb64e2b35930294547408e52d193bd0bece49ce89b92226cbb13585dc5c67d99a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5d14573dd0a6d809dcdfea59628f6b75384aac0d6e9449f7bd55fbbf97bbc726ce3d895c964a8af7d56aaa652e0a844f986d2a4e49495aecea1f0cd1a9b0a8afc8fbab5d73e07cc561b5d3f8157f299f704a44daa;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5fd76cfcffde11e96c6bd376edf9005769f741fb909d9401a469d06f1fa46f68a66af0d9be43ea59067d149fd796f31bc4982b81670341048ebfeb0dbac8a1ecab55d43a525ccc5c3f90bf862062db49a6eb8a0da;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he80171ae92cd1359c38791e3252685559abdfe1f6528351be15ebfde4f0ea842e70f26eb13f97dfece3d048f61c5e53c1cd6a43941f9d47bf898eef2e79f216ae8ae10d5cf76b35d19a91496140b6188cb06cc575;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6bf835e280608f639a75a7a97f9eed664592ceeb71fd0320e3819a550765d33730e8fa42a34bcbf5d0a292c8af305c4eeef76644ba4c68c1fa49423b45b42c8d718224b760c076e6d80d70a34a4a46354ea63ca9f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc4caefdb9813b9f9319dbc1f3c9b46ced057043053899e8d0a9c4a9ed9809422a0e74c0935608b07f40052a48631f205006a802673feb35025e96eba20463b702aa45daf88887a51d0fa1bfa9d67d16839987517d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfaf58eaa511c7438241b568cd3aaefbb25ca8cc7105771e614e3c7657965009298876130ba51389ea9c6fd6c3e824ef666c9e07fb7b66da087e1c455e85ad51cfbd34fd2e4e4b264866a432034545030a68bef9e2;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha5e050aa92c25852fa9268eb17ff958f64f872860abd57c7a829f86db2ecc577b2f96210bb2f3de810c75d2d64f0b555d28a53f9fe0d00aed7f44e2a3d61751f97725ec7a0c50efa70b00a2fb6f6023046bbf07ef;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h830ed6560b59590545492ea6410766f266b564010af4a426c6af5b0c731bd6cb9665b2c07f92c609d5452c35cc6bc2f466679aad47596df1fc31132258f6a906caae78054f7c0ca1ccf4e43df58e6d3453df898c;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hacff8e7b760fe459eff6f74b6e50fc2382de4f9bca0f3a08add38b3facbdf607e126e4f3cb3cde940b3b4fb155c484ad2399257043a5d6a93ff4dc8dcdbf25fc5458a3bfb194f88de1167fda5dd81b8bd8913745b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4de8bfba1153cf31c98b7d7988496ccd9e6fb7415d71712e4fabb33e25ac7b2f74bd39ff1f7756bd26b766f368f1e35e15fadea665679428cb9057487239bf7e933fcc0303f08e4a784cbddfb34505306cf83f5c6;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h79059556e1e985718269d994b4250679e0708f06f6619b227b04fdc723ab15911c4f0b6fd43ac36fcdf2b969462b71f681572a8dcecce0a3662059f5dcdf46ef5809935a9a89421085e7d2170380db313fef73021;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4dbd77a22979fc3eba00f01a1696efbcc8600c2caecb442ca3939c9249eb0db1439d61f962e67ea0e133f10b341ab45b16aa62cecdee0cb75fc185531dd029613b11af9b2c257049deb4bf23db2ab36b022c66606;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7b244bc9ccda674c7b0fcf88fc622b74a83353aa03d69b40e29c7c5da4908cb0122f8f8013e9e836e01db866b2053bf85fd7d98c9dfe810aa1279623536afb67972b17763ec02fdf39c528b9897d261c56800ab94;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha451651f7eaa6a28bec76bef4ecd2715c57523b76aad88eaf35f4c91c5b38d1db14b979919c2d73861465a7b5b6043f18fefa1e762532a091ed9b4b208a29b4ecd02082a37033f7472d150b9ba9fe8d4f68b90bdc;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3c349d7562a0504ffec245ed68021c8f3c546ea1eaf940a299e349746cc5a0f95074ad3d8f992521ae9d565d2e6aa46a989dac37ea4d22d404296a201465b0f3f42ab3aa8678261b0d023fa8d4bb7b5469cd05a5a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd95d2fd9890b10dbdc92ad0b89818b36398bf070d60d72c86de47a2db1c198b4ae90893f050429733745a057a3e81f035afc07c1a34532731830209fe5c96fb2160aa4886c6d8c17c9550fad724d1894763b49370;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd17831a904cdaecc3e0d96203b769c913081ea83c69f4efd9157fb1ee3006984c20ff27bacde4549872899c8190a225ecf737945b1a799be13ed9a28f7434ecdb8ee9015c9f49ca204ae1dbf94f57d25510e5e2c4;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha6ea51b1a20273ba21ebbff98fea821413b672c72afce8743d9205a747dcc31ed0ae32c135cec0034af8ac303fa6bdffbc10767aaf8899b4182972c80c354bec43b57fd1376e7b2668cf6c59d59472dac98e99081;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hba8d136d5a1cce9083d613f280e9667064a47a5640c4055166ad5dc921973faee994f0d3aff55c459b62d7058935b909bef8f4903a2b377e0b9035b15b88628bd1c5dbb39899eba656dbb8287837cc0f6722eb66c;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he1ababa80a976c566871730f1a4ecc9de96e5e2f74731af0673277b4a1360a0df5afc1b53da792e437b34cf794f7b730922a3b7e69761ede9c61a39901fa69a7bf69922c8b66e50e19cf7bea88bb2cfe01b2f5422;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h51d4681c69a9e01e361937ba48acdd070f35d0f16b1af9dc5010e7002333ee1a8e7192dabd7a9df9c836cd61594c905d7e6139fe8688e99c323fc0f5c83e07de7c0f69f02d75be9df275dc739bac3416cc24cf2f7;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hddc9837a06a2645c578915e2b9d5ed2b186d0ac8320eff447ec468f74174be19876be1c9f31b54d53da7d77a37d240858846faec31a5b5fdc4c4e2068edd08f396288493baccf392722d1ef0f88f2ec1f0f0a39bc;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4df16a0976a693b6aa385875c8ce9b7bac8650bb202386c0a28eb837ecda5f6322bf6a2e299cff26746090f255978b4881e273a17717ab76599beda1529c10027c8a92c9a041d7d82a636a375bae8a661923577df;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hac0d56f55e4c73a435b30a573b074c152f2da9bfd628f932791a26172230d87c30ba25c005a2780764037876638826ef5c2470d363f27f2fda1f3d0e62c1acf931b31052de1d24ed681747ebdcc8d0b6c91e3d255;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6025306de56530f331c2855e0c21c3baeaebd808e6e66bed6c93fa2441823c5251c55080388f0f22acecbdaf013262d38511d454118fb679be084222be3143468a23ccca05e41f690111ad642efe8990810f88e54;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hca8beb25037473cc9181f3b0423e31b91a1416e2a425a1d073d5a8cc3fe1c9e2aac587d51e801e03e47d6984d50e781745f28fd0f3ca52b4e601c134fc63d79cee2aff22ef4c319d63c24069cc43d69b9f7ff6e80;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h61993bf0a8021117590b8c050fe38b860f201d9acbffff9be3ff07fe42c810e4275639f1777b61c27df92dd9681f4a05535e72baa47e63b97883e03e0f2ace69e212bbb3b2db9c91ab2ba9609f0cdf1ef26640d3e;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3220d293f412ff73da21ef5694878769798fdad581264e311e4575339daa8c935486fb0ce5dae343f1e3687f3c69455aa19945becae7ddb7e0fe5015e4006ca2cbd6a543ae1c1a00bc395da4dcaed27aa25109ba7;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h91215b2937d2a9b0227c4288ddb6fe0d97605f4bd483a62fde3380ea2ad0d00e39b3263a16c1f882de9fb6727cfaf29e769fe8898069e0142c7a86a4bcae985d86a28ed589653626b7a224207dfc035a7c536c83a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3a3fa95321eeef12ad25b6dc5d68e5a5596d5fa3948cb4ebcd9c280f68ec74625efb4dac5051bfaad8e1678da0401aa9a0b50543a817d9ba3ac5d7bba4d8c2f141727f4cfc8aa434788960d97cc72f0537894bb8b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd49360cf52cc612d23d537f2233c7e58ff3afbcf5063bfa706bebfbb4885e97e53c81c4ddddf32a8505b57e6564070563a1d0d090d2608be6f560c107f6f69088b2df75c743a7f3636d8c1638f1bc8346890d2e4c;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfb167cd47b0a532304f27ce6b1eaf61c60c0b384c0856ba519e061d130da0a4d4e589645b2d6a30f279017b5ad088edc111fe8a7b0f23f61cca21a5693f2ddb5b4dd5b0cc1c6ce3c24e485b6cb9ebd02cc82878d7;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h653bf25a263354f016d4ff042be02d2c8bfb67309e1769df2b48cba1039be21284c8340926593c4725ebf7705ea0200d430d2a0f8c9ba4de43b311a4db9a09d1663f5b07db671975db6a974d72f2a49838b0071e7;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1a8cc4c58a77dd7146f0a56ab44a4b4c03855f8c6dcf44455df3aab361b8ba123aa72f2384378b15a52fdf8f4bad2eaae1f76d27fc5f774e94fc04d0fe39b8722254a9ca3b1894153bd61abac8e3c7853b8e08a1e;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbc128b5c525ee9a9443423d03aa584a5741d8aed1acb208804d4a7581186d322fab2145886d2d446a502e0cc408e71f1fc9ebb0ed27cecbf35f1e4c7a25a682af5a1fc1c29d7bb61ad1bea13539ac243dbab72898;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h73983c66b7bb63dcfbe794e2e31e844f4be3a51c32fe4d3e2e2d4f7564407be8209f656591318d087a62549c29c3501dbd80a0ebe3354168c9fd3f628e8672f4d4a4fd8d2bff722cefb5e6a0193a6039ed650a256;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb51406f49aa7d9eddd818ba9ca1225f0f9d815318f4077beb0efcc2f3e58fd634c207e745af288e9c2798fe43fc317398ee8380976de2d1e7dc73134aab2be762fd8f3b0afe7f5f2e00c70f6d74e0df4068e5adcf;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha4f740b7610581b3cc91c024eef0b63bf8b13a211a5e4e310ac45a8beedc24a8c9879fe06b58de96f090ce1c160022b29d62eed5ab2d5aa64bfd5e63ec29642799e637b2325d9c07d300e56866e123c2394c7f96b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6d55e53aa265a71a25af39f22e65a4765161b3d8a8423748cb8758ace69be4c56f736d101adaf259ef572bfc9f3b16b8fdab9b11f7fefcb98eaab401a6aab63e834751f2e79581ce882c06f1935052f8716c3619a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h77db924805ae2d19faba0b703884fb843b4fafe3ba67bac31b9ad4c62994067ff10fb6e86dd381f2255b704cb356884370c5cfe0f51df2ae380327cff0958706950d68faa559f2cab2996b88acf45ae132b6e8db5;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h40308b6d713934a230ff8e2691ac79b6f0ef79e8d0e1a8a51d0c050d37e404ea1557394684314ebcf0767a719e9fcfa6a71d7bad9016a43e731200a751d52ba076d3128dd33411d31147be65b5d220ed15cc48b65;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd6897e5da1a3160a09afeaeb79963aafa94856064cb2f4e4a4ebf4163a1a34fd41e9fd7fe4e894e55ffe761a04d128744229d44bd46e30721645fef06602ba1fee2061266daaca95a5d89ae18d95122edab67b04a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6981b2617592ad0eda072c9e0a4668303fdadb571bbe42e035353eb32267f70139a83af5e00a861f36a765f98ee07e98922822410662dffcc9033eb43d1b78bd6e1871ec9e380ffeac2345281f85ccd503c2d8010;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3877eadf310fe5298616a5d43a9e0c65f78c17456138759ca683385ef85a4587b2f1d2f6337ac8b70a99ac81bf17b9c155ba705a580b3fd0dce75f537acd75a461dfd743b77b3e24ceb48749f263d91bd3330b34c;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h977f5d6aa59ecdd960e9b7b4bf3570d1266a37e3cd2e7984bf9c60419a927ea9cd67d15c79ee4ddbf0380f4d0be1fe727de9b129075cdfc61e6d24b148b1be4e6256d4455546cbde5f9d358c177b1f1ee010dee93;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha5cd62dd37aa2de336d37d7f083e9716c4157aa604e48d04214e6079702233a8d9662c108df9088ab34e251f08f0651d53f43d10176036c27ad318807f11ec2b089d28cf52164802e6505ccd917c168845d9a62f2;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he028e8658dc918e8459d49d03b9abd0c5d5aa4432a91e9e1c5a5c209d0ba0708a3fcb915ad953bcc69e0aa2dc28c6922d16f20c42a4485b586d97ae818c2ab24b95e32b4831aa00eef052797cb250a958a8ee2c8e;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h98c07bd8792eafc851809a292abdf6ab908c1a7835305d288334833356ec349ff5f9e918933d803835b8f8f6eaa192854d0740e9a6195e6f956390461d1290ebff1a57ac2444c21a93fba5024095a7b71b801dd6e;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha325bad21c414c324238d1cae9a28960138e3793b8de4485bbae920fcd2b6fb537baa95451fe7a02c73545a201e8aec0635e013b6a9170d88ae26eedb6fb77e50ff26830bc93fdb282519a45d18879c43e6ae3d0;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4acc8fa05aa2097c2af0067c8738dcc075fd2f18849b50a24c39d6ad8148913953f5958677e6824ea7aee4876c7e2700c2199d1090e63c3ac17e2e9a654c27567c06e5df0672b7e67012ff56e65f48a09e96c7783;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h31c771df9e1bfd3a1417a45c5086d001ac20b37110a6a38fa0c4f24a1eed8282e94a3f7f2505136e38fa25da869147587fed456ce2de53c7925102a4a90a3ab03d25fa74ea72d2efb90633d56536e282e80f8d08a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3cfa82ca58907f95e65b8af12e07d07d196eb2a522978fd3c431d8371ea18d10dbb2f87740f3cf79616aa99f0ef23edd986920798f259631553e152114d8435061116aaaadf43aff280cafe2435867d766e24e0cd;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he19e910727c5dd28e7ca8bcd8f8727fc35b3a977dc8a40a948c72efddba5a8b8547a7a8163b54c9ec347baea8882ca8472b3e8f500eb81db0d7163b688110cb4011af569b6ac81d41df88fca7f71ae2a052efef05;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6182d94ac3d71484156644b3095fa99b626dc7810806e61c7117b92346b7c2799e847f00b52170bfb2285dea2c50af4e302dee1556c65736a6980cc20bfb86690f88eeb573ab3a98d8d0303e5d9c71dd0f2774c5;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1601eb96fbcc72d47812353d47d9b3d6e567443c51f6bc59221761e3ffa25c80a14aad8458487334b93f6712ced38ec159c4076db874a264cf94c59950717e4cc04feca2df5d66c271c7c1449cc5a08a26c4d9069;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9cb8e7e08a52b0239ce562a31cf6b38dd3194ff89351b91c6b1db5dcdcc5a236a7c67ce3874d6451860e3af8bf1724e71859cb95221d3ccf5e216a86290d8daa5ee27da14967fb378d6ecee92f8d73164820144be;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h10a1f25c3cc78480fd447da06392ac86e8938ce41092d56d909cc60fb5b0a16d0313ec9f45cdef766ee2d3a3401ac6d1bcaa6086f958e49759176b709391f9902751504e4c4361a0ad12efbf24600723c1ea3eb90;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7de824950d5db5bedf740734cd494d1664681b6ea6bbdd3c3c6a97189935e3ca8350bae0184bac2a270ad0f6eacb028ecc9c6e67f622800238f86c2d47a1ac5254f13ce9ded514de55bcff63985cb8526d52f001b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha7541e86b7f93c88f523b9c7554c5baa70841ee9bab463b109b0a176747cb2315c3a7232c0ba87d69e797ad955f4e2d4a0dd4031951b4bacf96e8329f5c8add710e9d5b148d1dd89917ac1e936f294bd09006f6ca;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h77f50738aa39b8c5fe01c8449a21f4d0d89591155547ab5778d2a8eb6fd39926f8f190aae3bf36d4e354a4a7b6849aca2433ee9c0746d5bee49873f7b7d6a057bd43555ed65e31ed3608bc8f719449dda4741c3d4;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h75aea6e06c8ffff831640b021421d317c4e7f766c663eb57ac0c1fee9fa5892562a4a7d5626d179e3f05ba5e9ac3b79a19225e024e5d0aff241b9f79999cd3f5f231dccf312600b728b0425bd2c554be1f3fa4bbb;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf5dd226b91f8fe4df253e65e2420bb01ef4b6060edc850322cc380b63dfd3d1a884e23202f15056d11911b7e13fc27b2448ee2e8cef4484bcc725cc4a7f99419ac66acbd80dc2c7af19868170f1879e0fc8ec7424;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc91b3621ff3599b4b68cda627102db63e113a56b02fe411fa124e7bf186694fbacc6d8a6d1e2a60d52940b720da7bc1f87e2cf38d14c6f96d658258fb540d0655b271b33f5ad3172ba7fa0127e8dda5779dff005b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9e801cf730efbd65032ea76097298a782449c1a0e9f4d392e1618a9a88b9ea1d50e212da6f7a2c617e735a9c936936c71af79b777f549878d3e4143eb5ab6da74c24ccd0cf3add96da004c11cca7bee0fa5fd21d0;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h84bf774194ba87cc50d393c28e7696edb3599ce82ea2da0f24a4e03f2651f4c309633fe6d78d89638242d3b8e510812d30ba72e06c36cba4684811121cb71762b8c3ce18b1f9a37e194ae3d5733a88707095440b4;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hce4ba88d597951bcaa64bf97da45b8341586f6665c1efc33668b61ecc009da6b38e6aa205e53f6f882f578a270c60b338d45d36d4f3a1f6faf1940dac288b7189183eb3f84a4daf4258ccf64b924238ad407d6557;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1dcd88e5ca6271f9f377949740423e6d216a468013c5082be39175390225b8e352972b956a97e2add173454ef3841cb6836c747519af7c1bc11718779c557a98eb09114602c7406ca8ed31dab97abfb84c424d546;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9db5131f333a5bdb677c67e5aa0f4ba65e2526d2cf4a386f90ed038c8d4b4b638ae9e79edc44cfbad7da536993e45b117c5e7acdbdcf55ab76ff87e44fc0d2ded093810cc17acb855bb31b8cb64a49f23e3dc2413;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hcfa1a3896d82d69675a75e73d263537cc2268664f02222221e71a69aa0f729022a49d88e1a7bd485377811daede1cda1d081668e9775aa2225c7516582f3f5da64bdbe23d9e00f71f57aaabcce2df54482b4fd6b6;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h12e4fbee824aa7372ce2cc7a8d7dd19a80731e1768e2bb82ccacd57aaf8f6a9191d922a76bda092c612326b7af0ebc1c5349a32cd8fd26e4da9076f8febe7015b06260d71356ba8606146564e185028a263081a1e;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h188786530ea5ab12f93e6f8e7fb48a1e53e3c63205eea6f6e476d05d459b8ebdb21f0c42b9be15c85f4b08a49cb30297ef840a530014488620abffdb8ccc67dc0bfdfefa0fd62584b7ac2381e67d9711f8a143afb;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7d95dbb4db64fcd8b4cf3923c4680343b8c0bd3c486c268e78852f1d59ce0b91c8f3d7ad0e6368108317bd0b10a4e0cc3b5abfb2527b7867cccef1d3bc1105e40ea3d7e074c73958840e3fea1c7e3a024bdf4bed9;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3a7061aa9ba590bea699742c12c05af15d1b28536c63fc7779376231fe2f21e9fddf4177c9edc5d1d1c0759d11c4f62741d5c9f5ebdaec245a9ccbd37667212df95e5d59c83be194c5458b19e117c8794b8339fc3;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf656ae4b1e0a81c5e5ae18bcd8b9da08c84971be0fb22dfed835c85ef9ed20f4363e3c3124b874a5c9eb672bd2b77363fb7a949dc71c09ce5d4942b17d7eaa17bab22afecf056011af42256bf8703b68100f308b2;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb47c0f48a07e43e5b6e2f1d062614abc2a1732f884585831bf9991fa8c14f5e3dd0698f21a24dae7fbf53f45bbb26892f2f46232e878d9de8cb9f8cab565968f9d352b1665dcf06cb51e26b05b5c948c8307a6625;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h773fcfae5024ff3afebf8cb121ff6dcfafe1842c497f73f94ba8de521e9d0b0c1c288c8dc35508844f663d3d9218579dea6a66701d0671e0ed22abdbd78630353f9bc36410c70ad6dd5aabdd740171eb1b6f50780;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc92ce05871d64df7d6679323dd2f5eaeaff1d46edea594e13ac6bcfa519d24c794053a23bd647f6083c6899c813b0ea590fa70d95f41da378e61401693232a53265c6885eb5d2a90fdecbcea2638710ddd3010a28;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he817d1d8643d171639c5c64fc543ee8fec0e2d9aa2133cf8a4d0e9b0dabe365b5e68aade5a570fa55259917750b5a691750fc1a89ce314f6ebe651ba495549c4f07ce3a58f6d7766b7fb170389de0db997e1f1803;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1a44436d9e554587663f50ee8d2f3d723297da05e3df07dcf6d11855f0dabd9bac680a7ffaf6be5349e148e0906a5032ba030bd840ee0df2c09ccb2c5e0aa6883e0b198160586255a236a3c121eb47d66f4a760f0;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha3329be05bd7bcab41e10ecf36b689fd0e7afcff9f47624ce7d00cedaca9352f9f2d1356ab330b92222ff8a7ea0cbbf8109f7bba9569a7635a331e7993ca1ed62547345a217cab1945836567e947ca5189884b93c;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h205b4bfa7d900ba14f23cb108c4e24ede67c57a03a10e6a9d30c2d194050179950be3598e771628070225c3770f0308a72687acaa576e3ddd8dfed08ddc393827c0dc77b391ab8ebbd0dd1e1527fe48f770cdd2a8;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h443c64c05c9c4fdaea0c901847d8e08bdda2057a8a282ef11fb42c56619bc6c2ad2ed8719a9eea764f05729e773e691f931896911178e66f699dcb826ca7dd38debd5ea363fc26ecc4ef667da7e1340ec894e212e;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfa167d7ed3d6eb96c7ec14324f19f2e5361e3f9e343b419c6c20917d76d7b81617cc71e24c878fe924b71d2a31fcf3a6550c2dafc1a7faffff0369493b1698c1f7474a13777b82df3fecddd7fbf8161a9b1516786;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3b2157d11e50fbaa183756d5ef6f2b326d8087071d48ae95c4a359bc64a8c43193e014eba8ea1c710fa68defeefc23dd3a27ab39ae69eb3fd2584fbd145a302b85c098027e40edc1af647f0eea41e16330f2ecefc;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5f3bf8d3b87396860a02a0800a0df4b5764887c85878f8a04e6c5cba705e91c2c0e7da1e32f6c59a3cb11c0b080bf95e45e891dc47bb532483beff1b48b5b6c54678a2f9b51ba2a9593908d9ebee1ab43704c496f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3f4d848cdb36c2919451418412ace34a2c16e102f79bc998bc1f511ce6b27df2df8fd2725e833e1900ec4e83e72ecc40b937959c0b2acde8d15fa0bb547831c465d5b4acda15a428ad5952e1d1280ec38a5fb105b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb70b6f04c40a135f30f246d4310f78d6963a91ee6b8824f6575d785ac4dac36428454b7a02510fbf95ee9a1c5bba6bc9e1ef2068be5e9bed9b2f44c6294290bdaf2e98836b470017c32a2d65ad37e465c6dd25cae;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1d6c65af499f1357a9bbfe446f0858a032035573ae19291b6582cfcf6213dd7454709148fb577ad60eab2936eb85e2c29ccf7380009afe0640b2ea84ce88108b5fcd3a0aafd18515a6bb916d48abeec2b6e31ee00;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha2437ab8b93ec03b6da1b70e700f9dffa10ff0cd2d49f5fe5c0f6faaa085e9cbe620f7c3f4956e23b1b626f5258405b858ec0872b576e1c3701d1b8ea408c570a795e40daa0b8d3fb11baf9b4ce1a0b3cfc98f88d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h277b0f021d627bbdebfb61b6916bbabaabc21e57bd16fe0db30b6f87e77a66177e4d9c8756fc3b2b0213f7b69e371adfbd9ce182faa02c1bb8b0e4ed75d6f22c536f12a4d62b12f51ca366bd526580afbe24d18f5;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9a87598ed4374efc7635caff0953a2c751d174f85622136437e1809897172c7fea02ec4e9b3db7db0a3326dc8643b210ac8bb48453aa84490aa3d7056a262c28ebb4d5182ae2423166fb2116448c6bb011c2aca2c;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he6f1fc3ff54341ce1e430cfa02089363b3da3e051f2ae6a6defa02837cf7f8c38518b83df37ced84fb785dcdf1af99cd8bdb3420459647162bbb3529e3103bf88e8d10dd9409035321463902f12665c7d8c698b66;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb71b409dcf2a1f0745dabf077129b73a6901939303c5139037f2a95b57037bfe331b8822b301089e51025aeb88b2a355058be772144e72e16764fd3c93dddd748e7a7ba373a93db47a14971905bacf42d8e717102;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf4b9f712d4a8301b7ec59d6eabaff1973855236f1201d4e74053577eb347fdfb5600ccad4b5079f9c7031c7e964184dfbdcf3f247746e33959c16591f83b73d02340ca8e4767457db452adb57236dc44c0854b52d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf5f0da1f1f38f74f5d592276b7b979684154ecea7d4fca4dd46d237ca041083a831036a24fee521fcc994bd17f925145c1d949c38dbdfdca3070a0d19d5f37bc4bb685800b128e094e7b1757aa874e03c12866496;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h782995e6cd315a897a301d1dbd898a03ac95af2f48e388794cddf330a7a2b039cf64418906c79590ef396c0c71b8a021ec275d95a5e6ad034ebe70a8f1689966d9b6437938195d7d1b17c41742a37b769f4aa6b05;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he4200217edf02b73bb9bd55092e2375f8121e37dd8b1ae4211fffc6c01d8c40e8698ff109fa94bd3bf04952acdbb07b3b005eaf935b50ca772bd9e27a5eef465df9b0f60dd9164a3b61b87ae25608bb896d4accbe;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'haf6545ba0b7b7f2def81378bc45edf2016fe0c0893ca6e6194fb17f04b787fbdcf27584583d0cf43039cb191aa59d7ffee6bf40f94fb12bee95dcaa96e08e154b637ff60a5dfb0d19ce027a886146fd30dfc3c9bc;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc6ce1c9652fa85d3a50822ad5356aad4112e0bd9936b95bf9fe2047ff892e7075aa1a7911ff457a9b8b35fc99b314399f784bd55d10f9e77a20b0999cfd98deaca91ef61aa5770ff67f692ef1ce3af375bbdb4eee;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4511569bf9205796faa04136573efba00ebd74daaa19309083ce6f5b3df78e3d3d1160cefaa7c19d69fc78eb38cf66023229c62b5d594634979d2e51f0aa518c4628d95159b43da60faaeb58ca61386410da012ef;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h779cdec2ee561729f174d28bd3f50e1d1e4d875f42b90b851ac15587c76977c2cdb2f73c46f3aa0bb1e602b44932ed06df4be6feda9c5a426c40de643144c0f03052677e368a52768a454059043d113605ea7d7a5;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3c1792b9d33019de5ad2babe1a96bef9e81f39296565d769c2d236de1116d4e72e740a69413e96f4b08d70f00111b583ef8b817c1ede2e90a62eac46c3bcf39d6636475049e552b33d921fe0ed0c11971a9542eee;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb354cb6e8d56dde96450731985ab73b7fd51552469717cfd724dfc3472e9c7f7b37f9c8cfcf6e0131ae837e57ac76381c31b3d6328a070fc8aaa21211d7fd2e186720bd5d0a25570dfb29abf392d6b7f9def6acfc;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h759c136327f6c93ccc7a8ff69a8252d9ae9298b7cabcd93052f04f193be4ac2009276f7e37194508cb3146db5fe7f2f9cc271ecd710059589915ed56ad5b36a147b43a4bbc10512eaa314ec614e4d9a8a3ad31d75;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h382ca3c05ccc8005fc9329389b4eb0db7dbd87854e2381b4bccf29e7576dc395a355a13d032b71b21dd34b83d7305396c97d1b3ca4cf25fffe07b962bd4faaf0fd85849d325515cfc281f2b4bf2db27fe5030636e;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7c5e205719986c14f5521bd9a861f5390ec6d2e54084b9dfd5e9a56508f26809f320f1f4be878b533eb5e468bc8669a4b0f2ef77d57361dd89455ad4b633994956368d247ea271418e8536243704575169ed1605;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h35374eaff9157e176ac5cd1df932953d8d822510b2ff3aa2215f9354a16bc6894a810fe3bb1004674ff03e7b02946c45a104cd84cd3081ee4f56e37d23b4094473c0234d41796ae19aab7334f2f2ebbf57fb2be40;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hee9488b22a6888ff44558bd34cde4e86a8e9c1ccb93c122d485ed037e6d0f3065bd62ed18013d4426aa4cb84c862d306dccfd2bfb0117f39e9486ad492158702f7c68ce9fb8f2fc63a1b008f1658f49d6b0f5c8cd;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd3aba7abb92c8e44e095c78f91a29d5d7c88f38420d62825656ba8f72d186755c51c1585aef3b57e212ca9881b314fc2653a02b7c5527c969b4538dfa9da62ce4a7289eba111515e660a7438abade04999a43b631;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h644aed29c6f0891854ecc1719d346a44b17d7daa327c229ecfeda293e78e1732a9a48351a3aa557a7fde714e38e36ca869c0689aa37677e1f19ec5e0ab6f5ebb9eef57822e26f4273efa1dab979e63b3b3dfad780;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6e3249b2166ff225b9a8b235322f7557236a8b37328d45681ac13ef0df2ac1c0409fd5f6daf86190920fa78dab617e183115bc612ebeffef41356330d7619a373cc89b5813f8c0e88ef196b4bc509895fd06971d1;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf02f649195be0aecc58655b41d831c11f18889604fc15a274c3d26f392db5f075d85379aff7225d72b15ac9766a5bf32107e7cd7a915ce4befeef2c785fbb82935b6307f06490ad6867ca57c14d705e8d6d13464a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hcc7f69fb13e4520f64be9dfa1d6abfb747076ba694b594869f44b96bab5ba79a9abc1a2222bc0eeec729a86031ed3ebcc62a691c890a6d36b9ea6a9a2a82908463638028ce92d17f0106007c7d6f7b3271475ef61;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h306f049d013f23a6d9b29e73463d9ca01f8d602cf3d38b1224b4c11d71c0ca53ba5a82ff6a22c349d1229350f62bf27702aa98742af265e6e6979002f29ac896a72edc8bc19b9b17576478176c44d8bb4577684b0;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha823f4f485aec10bd7d8e292313802435f8f5049c0c17416196252d63e7eda0b29ab770afaedca8deeb36cfe5e3b80a21b78f7ce2fea0b17825bbab07ca2041e5b96b75a6ccb436e3789f431bb15f6bd68a3fa975;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha5136091bebd7bb4d88ab974a3a50042f749eed846a93e0cae79fabb38ae44d26ec9b2f7ef9ae3ca2ab925ba905bfdf0136bb9daa64e3483af8c85a1af83ce6f72856dcc1f7bd32f3c9ffdeaffd64a610f35196a9;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha59edf574a646681c3d4aea153c737ce45cb65a7da2a68425e3a031b257a483888d9edd353dbb48b65f9c5a4cbe9a5237c90372ad1d7e60342865f4840c55a73f97942d9e769c1f36683b6a6526d5786334a0f629;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h16abddf9ea24fd99cc6b17fcfff7e0e6dfd0da874df11eaf65a2a518ca0e53097089a6393b52d29d3b8574adf0175c16e80878689ce90a0f6c289f3b437702bc4a74461127fed3c329799c5bcb8835a4b4b0166bb;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7c18362df743985eaaef38d1c65ece8f45ab8f4cb26a83e6c1985e6ce14ce60e2710beded94a3fb35885881660dacadb8ab3ba2d2136a006ea63f6c687d90963a85dd48f1f08a82cc5c34410e6cc78b00fd9bc767;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc8bf954964f6448fff71c24d2bbc39fdb1c03d703fb0e7cee42b60e60150ab2dff7c7b2abc2dc077cd2af1b37fe2417d247388bf1ca73043cc72e779144c1b7952928c056fc4cbaeadf29689ec3ec1467ff92dad1;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1160d695aa4dfb6ba01be6b3c67357a9a8d7bef45162b20a6099277a8906d4112de8a8bef26167809122bb2d9d7e4a6afe9f3edef9f871385b71e2dad8fa177e24769202a236e2fe7ac2907150bce9e05bb93bc84;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha6835ed054621ab452c3f6399cd9ef5bad56d9b84e654d35be05d5a4ce130b59379db57411be6d795ce5ffc9ae7c1e57839c88bac0467be3d5636e4b3788e2e4832ed70129c7809a88ca663c5c52a299a156fdbdc;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h384824548218a9ff4e92545df700e75acc46358cc665dd3a6b5248241d20a0f2e288999432c0c323eaa9e780b5758341c9171c2e2cc054cb664ef1859a871fd49b9bef2a9adf95f80b6fe6ea3d8437bc3e35416f5;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb90503aa550f98872ac6a00ac1b2dd1dc7082db7b5442f624c8ce2dc8a48c3ab649ea57c6a8da83ad62dc00dc55ebec41d43b5d6988558825a7532a231c6fc80f9eb912c05a54d90755040a747faae891945d49dc;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hca3caa3c44928f37551d9ee46c1dd7b087c0e0bc29c30ed88a6907caf64e36dd7973f05ca35af3083e5e3742fac525c2f3b0b6610ac054549a20b4c5d204ebbad70cab997e3f35be75028e6015164bbd5356ca117;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h30e1ee2dfe80234151132c7c485dc1b8c40248eda0dca30a852451e937c6ad888f489cb5b089a239cc30dd67461a0f76c2fa1cb0ede098f9952e7fe55bc9681271b62af871d127f5c4f641d71ed75475d9a72c749;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hdc32ebcf5d3ee9e01e69eac2b86fe9f7871fbde1918d9a0f9b1d831f74d8732fed7d41376afe173accd2bb9e782ebfe886e4bd8c37097112ee6654aa39d97b214758f77a6aed5b3dbb3fee0c7537c1628a81b6846;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h645d67d0cab6e3327ecb539a36a987046363fa737c11d69f73efc0f8a460fa8f2cb7635c2fd136c8e684a9d8b3b357aa1b93d4d65efec4c927b4cc033f9a90e245c82773c00115e35985145d04b0a59b28ad5c007;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7be08783a70114432d9dea49e535abb9287dd4c0f1947cb29dbd35ce74e06b59414bcdefe2e53da60a07ba2ce35fac01d8725a83ca85a622d7d87f319cbc25d2eb3107920430e4e8cb03936257ec27e8d28e7f537;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd9a6de12688d426d4c6485ebbfe9e065d410e22c555a4c7346966c98e1131209ff30a4c34fe1096da3df56788ab94a83b712697ee7b976f59843f51e9e6bafe11adf6a7370be31639bfcbc89e0bc920fb1ec07054;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h81f62ae536636f2c1de9cf0a542d659c81ceb709b80a500682d2aa3dc04f1431b828f9724eb79d31126382c4dd352cad026db1fb699e51c8b25c0c94f2801f565436e51a36fca78b56ab3a8d1e9b8c379ff41531e;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbda2620dd3f11316b5d01fc576686c836bc7af74c7c5f9e7006a79f777ba75f1beaa2e0cd5de281f2ffee4227a68a2ca492283ed75217c3bfbb233fb4dcad6838afc6e5c7d7f23c52357d629542672f319887c7a3;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfdc5e7d3d215027590d9f370651f3f5b5839e33f3a200e4be3a5475e37865f96ff9908c6199f6114baad8ff38f1fe6945106f63889a3591dbf6fdba3b712c16228de22243183709666543f82c43db443548af3ed7;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb8f42362407e86b3cf0ad27916cec491a19fd5dfcec88a690a3524fb503691791a1fa83c6b50278aea99812def7fcf95c9f15a2a08b8801ac7324c1af144b69be0ed92f356b365228e416ded59efac2bcdd37f548;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hea2c7b852a979f2bfe8445f51174e1ab07b5a29b0dc615b5893af9d2b728fc42978894bc284e684b9fa6fd60b74f81c8c5e1f4822ee28867435c51a9bd6c5220e78ed577f8f9dc883c3333e41e3031c10519d1d1d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h68be7a56d0b17c4b2423762f805f52f2e3df71176a79904d4ac8f6a8b6acd3ed0d8a59c86a98a52406826fc3583188333bb44291102e30fb9faad60c53c94b5d4c5ed096c50afecb1eca919c2ec62c39d66d397d5;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb385215d9b95014de5d05dae71aebf5c8218d7f1f7b8336fb679b95270944255992910c39a29794d02abca0aebb2df94089832ce8b0306b85bbd74c35500cb9d3f09d1be743f16a2088dc858e97833f1de0a928e3;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfac7fae323d1c3aff4dca3bbfed0e00898c294882460170236708d546b0e591b90cd3f68ef3ee2a9c612237ba6563093148e3183802bd67f8ac40a009697508692e824c7add9fd1dabf9b90e996d47eff6f75e42f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3eaaf1825b643e07eb29b8d83f33a2c561f9b5d8780fb396d5714f53437a5829d75cb498f21b7c8b8972c0cf5fd9e6459aec7bcbc9c02960460fcd1da7e545da40036e716284dcf6a20cde4cce439303a6d1b933a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4abcc5a327a4983019706ca77de9b210346c7c6a2ee3c843d10ab40038a2b5adac4184b96d19312ac9468cb83c22ac0c70e74b7af0257c1e2867a932d0ce8ffdad7dd9a333dc76c163aeca739fb19c3b86a74bbae;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h57fdccfe90ae028c218765e0885d80df27b52e9ff9fd9879dc739ec749990a7dc70c2875991afa20c4e8b88b52f81e05017828cda077bf1e297854485ff471a82a613676bc0d81abedf95cc2ac07384af15609e84;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha38f9a8bc0a21ec0c04691a9ccccf402f1ba0cabe482a7c1c6cc3707d1db566090b6c2dabd852f1b4801b2105b98da50b8d79ccc8ce8fd2c95330a34268c80d8a2cd44a5f1132a8fcb30011a8467e65a26714c2da;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h99ea3cecd058294536a1b82041630ad9bec67d9e19e1eaf41032e16133232511ea91c2f44dde5abfde05905a828cea514e33f4e5e01f62a74ceff31f1f00e77a9f83dc9c4592ad0e7eaf3ceabc9eaf3d6fa79f14c;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5728814584b9dde6d1dc579db17206e748d1f36a6a98ed46562fcd9fbbffaa291be66956da97419fbf1e66f14aeed1b9a6796ffe717ea631e1a0ecb27d80e453157a30338df7d68ea9749af5c405154a6814e421e;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4a1d2519621bbb7b456b6eae354b5abc82ae053466ddb706410534eaf6059cac2b2613b1a9bc503ff2f657461ae0d309c5e6e423286d02611567d74a3270fb04b36597a69aad333b00cf76a70a3130063f20a7f48;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3cb405b2cab3a3e5aaebb465581cd7d09a7bec5d200a50c2e6ceab1d6ae3895701717a135ddff6c58dc39524ebb94065e3381ed0c3b549cc9e25b91591f56a6660b6323ba08c7c19b0e11625db906a900925cc37c;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf0ebf92f881e722c3b20682c57f7f276034c6ce4f5414504fc6b538db3c65fe22c39e681b6a5018fdd0408b46655ebe0fd440879d076ec37df7adaed0305eef5d3d83a6ab1ad958a34e6730bf55639c302b584a24;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2c8730f5aedb430788d362ef1a542d4082380fd08bc5a033ca231177ec1276e7c3747ba3d21a3ad375783f99c2736ec1f63b6651efcebdcbad78927e18a6ec41cd1ad1d58b77ed754a0f33a92c46626c86d95583a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1a6c8939b5b8b6a65eb528b79b54e280dbf22c50f4e4efa378a51742afd3a004858df83a59034a86403b6caf1e7b8786b337e93e6989df32cea6bf6b70754d3e13d9e132876f0e7d497c0f67006de8d8da4abba29;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbd3d1e362c6ab9e9b73438a18eb56e2ae8b7b99fc11feb58dbffe01d28ffacbe6f58eb978069f21819cb22368410018e3987d861f1bd7614335d9ec2c7203a298d55a9124789137d5973d0135042416f5a3913e3c;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8e82781224f9d5169b661f49aa473d558e4fb3ae1e3011a1de806c4ccc1417c90820ae81f752ef26a0b37724d9e22190a2dcced1c2ea9aa4a0ee4bf3d07d19374360686ab0af101df09a0f8e6aefc54bb0f00c68b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h35161abd0e1165181c94010c8c8f230b9feee30f57191971da354aa811f0b937a57766a79794e0cfb3c94e83d1061ef3f2ef00848f9722ce3361fc8a25b340b8d45c073dedd9ccdab214365a0549a0a479ffa4356;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he9200b0aba3e0136b76ea8be007a342e1a8a16ff307df6ddf3c5edbc348fb4746ffed28c855ef9d4830b58f1ea68f3220b121cac15ff903b7d015c56dbf1de08ed52a270e321e03e1abbd69d9c2d1aae1ded56787;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h37780cb6f15a23ef3810e18219a962912fcce849def959d6420b935277b97e76c5908035cbf38693351c2347c955c3fabb9f661359c19d1c9b1c0f306db04ec6c68f32df63890351842baef874666fd542369fef2;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc00f1d6882f6fd5f1ca9db51e1bf4f9e92cc30248f21ae4bd8b225ff6c63d12ac920c916bfb338fff63f798cd54dd554a6d64803de646a2dd02bc9d1d3da2b9b46d9ce2d5a9dcec4d8f74b37c0268e750ed8e813a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hcc13f71770ac27c5ba4e4d0327631df9dc2352adddf1c9a334d7ee16660d4496e3805f5962a30d9ce04554ab672617c421f7699f5764eee872b111f343e18205d52e44d98d1e02fe651d77c99d8607696f1654867;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'heb6756cb00674f73305ec4c74f6eb6f690ed075cdb4c1b05630ce2e45b8f0f2873f9b4464f6c7ceaf47cea587305efd0e5c2b7fc1fbe72d764fa3a2c0fa956e85de8c780fef3a6dea0a6b0fb476dc388c33a93ee5;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h753e29d45d90e3acedf7fb6dd9cb2557106fddcae4c1c598df3324881a2112202a3a96b6121305e99400146a1dfee7901c09d474dbf969f9f7437a58574a871c007a0bae427603a5a8be85b3f924b17c2cf9dd194;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h19cf1f6a9199f5621b74a26b510a60f3f91791e174ae1a2fce598f8bbb9724de5d690ba45cc633914162b6353eef2c8b975571ca47a05683aaa440c381acf06582539ec6e3ed138b2bbc1186f151e90c0b142cc01;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc3866fdfb68306a783b30a491d92e9b736f5a7d8a470149e5260242e0d39c80b2eab69ad6dbde7ea697a5581b4e6301844602bdbd50e2f0e0262162627c09cd82de32b0b67d8cf614cc35bd4034e1b42ac92f8c8d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h58ceb88cbddef9e0c2e4669a9111514309237f66c4caebbddcf7a9107db57a5311f96177b93fe106995bf7fd922bd7cbe5b795775583c6fc2ee2dfe7f2f8b65490b4cd09b446f575a5fabd0e344202de641bd3b2d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h76bb367489d70676243b760ab30ff5fb5d18bff4c8dbd06294c59a35dc1949762cb09c09cf1fcd578e3d0acdefecdea609b1a64d0f581cbb6ad1875c10d48c978aba42c1a141e62aec7900be528b5aa29efc59564;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbe197880976caa7b77b1d6faf0c1fd2d30ef58ef44eb90d57b1c1acb623fa00d929cfb228d6a05c638cc9678ad2ed1206334add43fe9f7df8552ceeeb8410679a4dc37f37285be0caeead635ac8aa38860af356a3;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9d6ed82f59dc2c6e7ffec35d6ef4adacca579dce57320efbb9423f4991564802f4e7efe9da2d884f87e1db033f54f48a5fa95b7435a7582e77080a430cdab6254ab000f1fe3faf7f7a351e1c7d98a34a3d33ef6ab;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hffbd99e07b219bf8369e90fb871c971483f7932d5243c345eddf79f663e1494ea9684c0e3b2cde62cafa221cfc03be8b605f74a6393e815ece8f7daa65210e9d8808b206b5bc59088cf76aa8fb1fc54e4912f1545;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb7097e01dfc0ea45706c6532b6c779c7f3824b359b4597dc5ac7df34a27a42b592280e7115823058fc09323a9c88d443ed8aeda7aa3b4afba4f25629ab4deec4b89c7cee405d25600cb5af7e8d28bb0641c58161c;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h18f344227260efed702015775473e9138abe3e9720623a7bdb1ca848a62bbd135161ef2461e4a80b0648b7629715a5373be0a4208aee059fa9c373068a2ea17fa640da177728db2b44d2e6f102a026177635266da;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb7e7310cc95c9be4ecdd2b62224e2bc2fe37b4d55dd00803c8bbdb824bb22fbac45a49ee953af7a941c15c6c323a173b6662236cceb591a538c023151b65f2ade7089fb1aabe5ee8b352b213f8b20eba919111cf8;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb7c4f623a4a3dc0e219370c2917f4600a8690f2d179d73d597138309855b254fdd836d1dec0d682b1102e9754006d30f72bd2b7ebf4a75adb98f9f391b6d390b5831ea55c6323d078779b9ad6d8e323196c6144bf;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h17e6f203720280c4dae68df2f4b92bbd3cab524a193e18cd38ec7561a09761e82a826d9a053efdd7da605d6b9ffb1cb1c34c26d4a9f1a0e78487148a13664546235575236d160baeb5592d6f9772c3de383b7e9ff;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6783694688c55065d6e918c250e32b72d11556a8af53ed8efd0ca04f8aab895a00bce8e73236b5edf5e644fa7a140a6a829c585b4825d75f53ff73a3b72a7b5c6f3aa7da0cb217242d482813de0b65aa7055839c2;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbf3d7d99d289c9f5d1829a952e4ab789d68084053b553dc997cf678443be09595e451402c2ec6e7791bc007c8ee481d65fb22ba7d071f690c2bb92b2b746599e2ed1819b11e27fc29bc7c3d3f9e15e2f8799f52df;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h340b81516d6ae4e4abb50140c3c0bdf222e5f8d6878031c4c26ed5488c989c6509dc9df18b7cd021a8c8600bef3d9c5c7fe4b017f8efee66d3e698d28e9e0c12f92796f94d458dec1cd3eec71421db7a74ac9dd0a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h169832f2555719c6799c6277d5be2c5553baf2608d9f6526f78729decc78bb7eb33adabe8f69f7326abd5ae6676e2f9b441903220869d6d1b4d91dda965acf62fb40775d70c995096ecdf18a06f9e2b6ae67e6e37;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc19c4b5d6d8d7c5e823df7ae5517911ad8a4e72cfcead63a7a120619548b8b28cb284135527acb4381ae152743af1c20a2cb331eefdbeeea716c2d582d979e2559fb9d3470f2b23a8a862fb2095b4967f1a135c3f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he69e9f3ceecf30cfa8dc58b9ca31360ffec0643cf68aa43674b5617d71913201f00dec978fa0b9ca019cb343db418ca04198d445d18cb9cece4bf5e79d6509516245b25433fa22f41ef92fac607c491192427b35;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8900163947240adb452def3de8f24f5abb88ceb8cb86b581e9f4833167f633fce895558bcea172965711449e8d175e53194586bca45eca620ca6c977caf7ee51d855f7da7aac950be449e6cb2fdfc131e138a4844;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1e949c485652d855ac341407f7ec2bd202e3c7ab7ecdc52cc354b60372ffcbdc5c48175260be1e01f2759523ec034e736c25e3374be90df34964077694c545846d414b946e10f4f76dd2fcb499582281270d3bfe1;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha1fe26da821b54d4e765c6fb5d8efc913ac73e657d8d8947dd820643fc4389adb68948c2a1c728cedd4b91320e7ce96de6778749ccfb5eeed3fc3e20e341ca8d355ca0f38d7586fb44b38e99d9275261d99416c77;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8f65cc225abeaf71fd9cca6fae30a81838eb2bb792a2eeb2165627cf2d8a5135ce8a5116ba3a688a66603cee8061fbc419db2c4d632570cd1b4ed7315c28d1531c7b22b0b77ae7c0c34d70b6666a21dd7be0264ef;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7753b997d57ad6b02df11560ee75fca4d41dd756c0ea53124bb291dccb99079061ec0e5ee0f3cd4d7d8209f78fec82522f5a50875caadffd60952d8a34f2a51d0b60cc96b6fe56bc4e2ca882ea9a88dd10ea6b6bf;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha45e0d70c36cc33f695587777567c6e3d5b9de7907d61991395b44be2a20af7d71728c335b83177c3611195bde236eac9ed7f4cfb17b1c70531e136fd18bbacf85f7d9989ff5bb7a587c3de1e133f7f9f7ead254f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h28abef34fe9e8df9bf3d3f726ba3a3d44b2c55534ba3e9300873880c03e939416379ae6493fb5a8ceaf7ca8a278dee4f6db35ed1d3e7c16f6e4fd92de8b6cf87312fa9b30fdeb2ea9737e9706d8b572c74d584e41;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8f98528a63e6d0319d9b61cdd7fdf8cb5dd0fb7e375b76d3cf74d79dcc0e786362332deba44c2b44bd5b77f7ae9dd975edc102f8b20b5e31c4a75b0003e11ecc01f7e9994e1f0b60cc117d45b94615256675ac1b1;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h888f601b5453a5734e6e41c0d7e33e9210b1ee0b9c3446765b910d720a26ea32472ac3c25b6bcf95124c373db4831434dcb4c23fbd1e7dcf657c6c8f772e330a251214933bb577c3e4986946bb86099812383eff4;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h68baec8b2425a0bee8b50e35aec5682de7474c73db71e5faccf37c92e20700711b63b0d8cec0c6e92a8d0fbb6365829cca5c99d0a0358e760ee50fe8862f37df9a32012665a633bbe4e7a7cea36100f810cd1bfed;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfe5a22d732ac27f46a905f9cc0974ae3b841f5d76919ec5618758c44709ebd39c861326251d78f92da53cf4b09aa873435113ab984da1c58f5a8899a8d4da827c6c6ce0641a23f98746dd50f33d3989a26482ea71;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9862b4ca17b0c11d9417978c9d7dae284128bbbf2a6b3744a80c72f313d9d495fa46c2e91b99454ee2698385e1a897a2d9493fa5ee0ad3ba9f36cacbf77761ed16f3c8edca4edbe1fa6b87fd21639c98653dd9c1f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hdcec73d74e63f980be652bd6463bd53f0cbf7bd8994aa6b4e80ed3acf44a046dc63f4e277bb687897d4c768a9b63c8054eff897309312903598dc4cae49ee8d075a9243bc94da12c1728fef7915b8771d8bb60f44;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9950cabe2448ca0909762a6e7f38e7302be48b4f6cc1fe576bafed61b59f7691916f64b50848cacd1f528384d9485d2225b5fafd68890c55a0571ceb0644baf2f138416ef80dd8dcebeba3c37bef4082cee1f6c1a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h391aced43a96b5a02fff022aa200dc8d1ea4a80a59234eca0239ece00bdc6688ef93047fdb5618e6b3abca3aa408250c42e7af44eaf94c6fb9580d3b08e193ed50ea07d655c71e920696cd25a728b54d9a6388bb5;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h120095a4d7839775ab54f01fb9879008e4bc0839b987569add2bcec024605868a7301c2eccf28f72475c52de30bae3a92d42768528a4f6ab450c56eeecbffbd96a77d7f0eb36a358984cffe5631930da3520bfd2;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5ba13f1360a14053fc310d467e10a10ace73936293f2fdf5f56c5b082855da9dd71d8b8dbe3a4c888cc2c6550a87c98d56d135a5e73af1538f8abcdc1c63e1042f642d367b3fb551cf0c212c2d5800ffd1110aa16;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd595ea2e7fd0ab85b2a5b3bc12eb764f8b5a66f41123a07df4ac0647db38f27dcca4834ab148ae814dc8c57e78bc98c11fba5081199667c997eff40504f0b3f869dbaebf97bf93b87e1bb956503c9a49dfb2cab6d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h69030ea27cc32e474123435dc8e0ec54fa9e245225c4452512e29b206abcc69fd193b91cb06654bba0e44d28803afce90e4ad21f100d9107935820e62ab749099a9ead00b136b8185c241a2c4a3ad2146c66d1425;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h99a7d0271dac945903e2088f55e0aad3f21fac2e99cf5d084df26cb06d6322da360674524e6c7d91505e13e5e39c727c65bc0d3c07be8f73337122e04c5222b623f7fd99ff59f8e9915a94368c56c806fd9c8be9e;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h23b7b3817e02ff2cc49aaa8f576e0c3b704732eb2975765de4600f9869656353ca17dc4fe0ed3b91ae24eefe42e619cf14539d25cdf768b64935ed9d12061fcd619301c17f986c5f506fef74ea31e12034a27ffbe;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha8ff9d77cbba45d09f9928633fb992fce0c55b4f385da346b5819071f70e8c07d48f6f7b5e8753ea8fe75eb813a92090e41df0d57c962ad74953b5d694dbd2d26aa883c020b8d395e2ee9aff80681fbbe7ba0415;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hecd25e7cb6120bb2598a3854ff994589b83fc1cef35038fa42be5e612f6c35a8f99350ca99a6115bba7ce5e1a61fd8a9ef4f19a7dc397395b8220b73674364e573b149c05dd2c7404cc4b9afc7f6c4805dee9b378;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4353273cd9dc51791fab2cafcad32bed1970fe6e729bfbfc6a7a35bfd8518a5539eaac75408d60568bf7a1bd8d90d71c7ae0298f3e9622f39ccb8696a90c46b059a8ee6c1d8c0afe1786e3efde72ff99b210c3a11;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3671ef5d5ed75cf9deb4a983d56a375043807aab42a8d740dfd681b1de98abd1b9ad1093f479f1096cca3e1ac0c08a768001c3ae7dc063b821406b08ebb4e4c8bcc5b9fbe1366d32dc2de22b122b41174d2292249;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfa3351d6b69d7075e7fb96b373ce0cf7130a03a3a0ae68766845febe414e249cd071862d356ef4239f6d375956b30732cb31a07b875fd9019e4e085442dd81939d0174c747c7c05f63b7aeb528181d7ed46acdc1c;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'heae4ae7db74049234b8a5a05314a34503b18a72b8eadd4357d1b5db95f2733103186caf2804e06897fd2b8e1b004038f718efc918bc1e0351b91b6aaa720fe84c58ccc6a6a99c1fcf9fdb55f6785e27fc12b3152b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he0dfd2f2d336e49cb40ee463dc9a5c8935a427c3a1dc5e78b194e1595fd13365ea60c09f0a35bac358b6bf9f3df148f87d6b5e3ed379b0e0812a2fc750e562eca0c96d92d5e1cefcb5a4971ccd5b1acee2b3ac57c;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1d7b34ff6790b3b8bd01922707f5a7a16c0598b6cce8bec659d2998f9565c7df2c114de4a6bc381fd0b6790045702dfdfed4872c1664cc6e7412cc2284e51461c1efaba8be473966a20286100647a51e1f605d4b0;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4f49a49f6a8e6e1ec1acdee19d22b3204293931a74108194f5322ac72f0073d3dd1dc9bf57f952537fc81e5b7a250f57c8beae0fa29d8c8bc7e08bdb522b9c152622b012d6ba360c9c71119c8ba0c9736a71f033e;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf643382b86298a0104e5f45fe2d5921c189e95259895c95430e5f866116fec99a1fad1144240e0d7837b0e03e66a70d64523bf5a11b6ad2ed881693e920b0019a7ba4d3e0d5dbf34c82337e398cccf0bcf8254f7a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3b238f7095b0d1efcb1d921bb0a2d358e302247daa5f46fe630e16c938a4830ecfc951bb227a5e1fff0151c6c340128dac4ed5d2bd8c6343426794f43b310bc4cba4387cb28a5b64f0a95b7c62e3349a60ac75b26;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha0cf942f5a1781ddc1f1305c9153f3b528a0f0d5fe5cef980211c1301d6afe9193627f4bf955f38b0964b90732dbd3ac598393b4d20a97129d31efa39a30e71ff4946c8efe8437ed4d897dcf25ca99c635b9e544c;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h61b92d347b8bd3b0b8b1ed6adf4ae4f1ec482ffdf89c896b6824e1b366230d9883d4550a1c64d991cd35335e2b54e3782fcf191d5aef8bed1a31782b6eb1f203782bffee188b8974d7b9c976166bc18f824142ebd;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2e832504fa3a74f89a281474a7d5c590c51a6ac19d24e963f7be46b8b71df4979e09ffadf804a82aebeaf786546f773f713999acb3e58a671dedc24f2a7d6c44e59a55b5fb9ebea4ed0fbaa456e37a8314ee7b196;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3590bb39779f7694e77fab4d2399a1e4e3dd81b0fce5e39194cd06ee7a9d20dc0e703ee3ce569b4c865f85d3b87314969aed4b236cb52246964b3f4da8e010219bcf1bd4c523b5f2f3da456464c9b4bb59f408549;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1b99663d7ec3fc3978729639574dc59f963060bc55a0ba4c0a9a2d1b8908242ea169580f136629ec410feda7fb8ace4a045769971e8657b1760888374eb70cf6cd686a139ae494a8a7f408829216db14ff7d6ba72;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h361be80e418b83bc88804ca227c86fe670ef1e84ee5a64ee5a4c657dffdd8b5b03323b61040f880117248aea7a5ff8294a6297b9cdaaaae7bae79aa64c79484be44e1a1905d371c75a16c742fff8ccd1ce187372f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4c00332edac867e65603ff4b9898b217eecd40ee61279ba3db495bd799fc41a1921c12c61314b7ac58203e16a20f69ad4dd72e27a3ebabfe4e2f1114eedf89ad421c2191f8efd230891e11e731bc568304869aac6;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hea155e740b7758339de5ddb88012244280bea7192983e194e530313a5487f3de3302e47920e2eafeb5bb0d8fa50ffbf81728e207ef3161648932c8ca557bc4bac8846ea2c8f245cfed30fd168d5f700a95b41fb18;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1cdf1d471d6906fea3abcdafd034499d5b7c758309cf349217679c689df04cdef8faba4cb0d1a36c1b885f2bde9358dc5041446911925a9cfb85d0340897bfe9295579ee55d81ea00da9b2b4aaa333f982765a3df;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3d6782ffd88cb7b50787cad285e8f155583a6749f527fd6f7e1121c68e1d8c8dd9b72184c61c64fafe87a7f865e3ec24af5f6654ea068aeec3d57950b478691ebec75fc0d0f64021bda407f45eb982a04bc111f3c;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc083ccf0ec201307917a5a1cafbb767a340553205bce893c90b24c7bcd479c3ef29a5db952cd9b25b640d4458739d98025e78c2e8ea3c03b7981568c1c1cc92dcad25717751c725d2479fe5e3c711b7e498ea8763;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h70e1a5d2ae5884835f124c27343982aa91a269fd80d6e5ab5fbfdc7608aed7ab4fed18af27b32b283956ab0af4f267e278742ccd9f35dde899ac5904848e5102cdc458a4279012a9263f544cabc56e47654738945;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7a2f637dca60c8ed0489a5b4b8297e79319d53cf68df79ea143056cffa7c472a54ea8ff682f739c90644e79107ae07fd6533e1b2120da8bc5698efb89f57e8d6abe9c24ee3741d727da6deac40e47ae750f16efc8;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf2e16ba79b63516d6da6f6df5b034c721774dfac8a7fce69f983f21edce2ef14f08298fb6fa640e492c2b1506c7587e64d4557d6cda11c7989a6f7aec687b44fbe6f784a4038b1b4ccad766ee680bb5a76c0e78ce;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h26badaa643a7432639848a29eb294a6ee0f1f530a1f2543cf85b67f01adc1b0056eddbbcb255cad3d0a9c6ed2283aeda0f42ff7fdf622ef4ed9784fb937c2b361a31e263df4e47b362fdebad59ae5d2c23487b8cb;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfc41acfe1a916e344894829d2e4b58166e5bdae350b708de21eed61138d4a449fd4267f04642eb0279e94808f68034c42c0001af4b7d95c29d24282dd6c3b61e6a715a9df2bc42789d014d3e9a8300ff9f189b17b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he2eaf31135eeba59369dcb9efc238ae05478023b642e4d744efb53c5ee4752d149ddfcf12a72059b80f86c4b9a1e1feb5cc7daa8aed12ddd53976f1cba313a904f6bb42304b94f0a7aa8d7423fef711832faaa4f0;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7ccf7085215863695c765215d218568f8a4286e52a7aa48d5e59051b957fbf2a8fa9f05f6914c6e37399caa94d28b80e95c8755d2625ce5bb208c1d1b1be8705dc3eeab3d1c352281978265f697e4f0b2e676909f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5568fd4ecd3175a908d375fb51cd8655c5312ee8c395d4da7698ade4ae78b2cb71051dd7af26c3116e4cfd9102254a39942ef4011badfd38a616a53016b18ce0f45e9b831df72db5c0b6804866d1a8d4cc75bd046;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc68d819042d0e117449560647e8a65918d4bb49b83e3df5fea3ebf9a4aaf915ae587cf5f773b7d4d0e92d331f1472267f68c21c00d99abca091d65c8ba3709767ca1fe40fa53df356195c51ea5761bf8a08eb7425;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6b728d37a86d99aaa0a17e75dd924699e205b9ee7fc120ab37725d63e052c2b5515b41a82dbd8e6c788077cb2da05cae19037733bb4c8b9ff032d731a21c9f3740f5d2166fa6afa6f525fbb31b5572f7eeac6cdd9;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3abce122d677ebecbb38df10b14d0da23b6804c3d0be90e4159b4e34d90d3bec1cfc1aac04b020f94335427d9c92ff2819992e050f8ab4dd30060a4ed8708516461cf7aed9ebf960a65ad24588e1c38ff0fea60f8;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6cea22f59140abb24d98dce86c0ceed4d64ff2070e411299fbd685f27386bca627763f0dcc38df0e4089cb34d276d1421e3e76eab5de0cd238dedbc56e0e609ee27bb558ec8eb7652e733c77a8f3ffaef6b3e16db;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h12f779b78e3b184e21222f426c832aa5dd9b936d3aa5c9d52030dd41936f4cc9ff7624d3bb5dcce84562cc1914e91bf8fd962270a815921d59b6c5e2e73586901f1c100abecb46cf4fdebcc1485ff3a54f040a50e;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h576ab52136feb44fa565b1c708b46c30614a21a944996e63a6c6ce3ae0eba70909baaace83da3d5c0511ab79eb2c3a6a0f4e960f3ebb484b6f56ecc643df0cee6d87489917bc8b6703ce6f03bd3926d365717f6c3;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd0c5b6c67dffc0993bf63ca935256c8f06a1db5524099c7c738c2cdbd5213875504a41c6cf641f1af0715f5156be34126ac6902526c7f6772f1567fff17ad9419b5d697ab354ffbd45dcef7d683b7deecdd426c97;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbd0649c9dcf89ea6511ca6999ba14dfe46de00080a44c0d559a24d0a5444923859138d9361e9d10efa12b9cb71fdbc1c7ebb4ea85f62b7a64e62c90deb9d9307e696655748b54f356d70103a57a55bfdf6302010a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha68804754a8e9e1f7258a175c4ec644c9635eb9baff5a84059565f11680d446340f9e56a4c730ac0cedb3284efb9f838f1cfb1d79d600cd4e07f888531df239629b5a1dfe4db8e11e2847fd6877393c1294db6b34;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8c12a20e8920af03b451981e714864b850b59de7c78ab04aef997451ebba5e6476b4d0d40ef56fe2afcbaa062a312797aee7d9cac81e986a7ecc673e80aa6ccb58dff6639255847e6ade0f346cea753147181f815;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h66a6a5bc9416856807b8bf28d6495f300c938b1a43e5414f20ddd64a2328ad53d4f60943d53e9271f7fddbfc80e9463fefc2eadf07b88725030cc755d6769be76da648aa87712e501e068f213b29c97aa48961ed4;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7dcde6852b8007ead780c18dd38704c3f144adc041c939681738ecccc4010ec4dc4baf88e30572cef5f799950524f73c3d9b66ccd2502a1b1182b2b78d5abd92cae4e7cd85b691a08d97802ff7735b3cfdfd518de;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h279776890ccf2479954f73e113306c3ce60400f9a6855233d175f3c32e5fc2becc3efc058602fe05d8c583e7309772e8ce1c26ce168b221fe8f2d9388fa274de64a926636fb253cd7be9896916598fb5644de249b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5aa98f3dc2b7198e5fc27c199ac6dbf6f47b5b49234d8d975d7a1fcbbaf8d15deee769fae8dce46b08b72ebff29827a22f126ff0456bb30ecaa56c9a5303e2f500798b928cf2b73edb9125af0450b8ed21f8bba38;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h10d43b28321913af983b454ef0b2c2d61f5c613cc567d900a33aa0b35f08196cd23e7879c26b681e8604f67775c14f02e527bca656d908134beea94737c42e1f51b2ea89f4aa92e8000877b3a33271fde2a661531;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h91cf80529535e9ac6bf95d55e5ddbb3aab27525b76654513f489e0a769557888d5c97a394c17c926372a22d21666460474e4a6936c326a2f7f90d44ebea136e08e90e6c90402402d4a1259a118efd47781f29c0b6;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hed0889de76e5346973802ba4c1f6e9aa302bd959f3506b2ee63a5c3e79e67f06269bc2abb43292fc3f327467f09735d6e7588f4d905830cd02008bb9192ddfdb4533872cff47b0ab117d56741288a1203b16cf644;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hcbe5f4338d8f5ca0976f1c732e6a686e6b41e3fb86a1abc2eace651e00b5422197dc29ccc06a7144c2b6cb222fd4a93612abbf93add3b28d3232aee485742da2a74222632b317b2be0f1c3d22f714fc4386d5fad2;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h79ac3dd4b23502f992406289a3710b237ea2579b20ae027eeff4194fd4cf41da58da9bc36718decfc1614efd146790e30c970041930c747161539542c5b7c8c139bc4aa01bac433a4aa68e5debeb955ba61f33acc;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8b5dc79a48d62302c98fcf68e48e25a64b78d40d8acf5260ded974f157178ef833afec508cd94e3d0ff36003e7f9d1e03b73bb42150af7f4f79466969fc2582976b774d10424d2041b2c1c9a0bd4c377d7bbe7eab;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h59ea7a10e8512a319f6642c77dcc67766646e68b3fa8deaa6372cff1fd3b5b65f70c6921fca734b4e27cfc0821fbc2ea12c085b3cf524c622646f4eff83121738f1a0f7c703c860ac0f85aaa3e6d1762a7a564305;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h416966ddd8d0deec9546af4257b6f745d174643cbce52d44215b7b1b326c2979e74e4181f3f959ecde9526a2943195ceb9256d6f7bb47d1ec53f940efca167e1fce1cc0f4140e76373c08810e7033191fa86832d6;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h55fe048b91d4203bee4a90add3a7d027dee8f63f9b82652536b1b27976ef2e81b2f9f80c163b82652e098de3d6e5b390d52654ba483426b323b693c99fea60582ed24ae8f506781922922c2c43aaa7ee01e8ebf88;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6b7826ac95c057b4342f66dbd64fc0ea7ed78f3df84f2f25016f3a519a2fcb296a53e90b83bde782e279a16ad146c7fcdad593f2c1e3ee151708c11368c9548d6bd12676c396e42e7ba20cec9aa0ce4dbbcef1042;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9617b13e23021184266d879fd6783771f5e83246b5497852d491ef0c0094b74f3d4e9af7d27befd90478873b829182e69dcf4b25f44dc72997db47358436d7776bd1c7fcdef4e680ebc123b80ea9883f09df07cf9;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hef68c77ca67235f7137c9ddbce9b5d0d5f253a976fdf2ec00f88484588432284ff2e07f7c25bc8455baac7493bbc808a414f80910a280c4a081d2f679088854265ad98e7f59e0a86c5e6843cb05c1ee5b0e2c45cb;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfafa96a69d4318062461c765a27f2ef17bd8c06264d964f25dd329e09ff46a0383e7803263ce835104b867ea9de72109fa85799f382adea8294a1e68cc86767d5b83d0d78c1f42b92e2252af5f311f6661242b0df;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h91d99326b92c3dd83c19095c78719ca24f9ad3499572b80e2c2445eb9c7496428dd584c3e6fa79793cc0d5b344268cfb50dafb77fc4af43fb1a7acb9a99f3098706c5420797f95de51bd44b4b11eea129c8b88598;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha027b152f216acf0abc9845054560010540bf31d34e098a871498a4a7931828aacf3d9c0784066facbb1b79088fa786440aea67a2b93c8a6c332830d5ef5ffb5ce84d59d165ab6421a1977b88cfa9cc7e3372dceb;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3f9e363a8bd22f2727c18f6464578ddd9aeb9a590940223a19d2759b556066233e332e6cd3d1cfc973f08605d0a8f9c79783c6c6c6a9ee551d68eecf576e06bdbc5c36186ba32e4ed6e47bfd8a725445ce8b9bec1;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4e49d50cbec1c7858ca7bf53be82ce320e1a22c759ef6be39029ad395a4651a8c1655f976475e9d91d61e90eb582a32d449c5b590ee0732964eb88024d90019cfb09fc812eef2e3660562821c3df4fea864de6012;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h970d5159e155211e3e75a71c5d30fea3eecb0ec24dd369816eed6459f79e61cc78501083f498f39997045ac32a2356fe0739999ec48cf504ebce43170901ec4b93480daa8eafb096eb1ab1cf1c24d01c2443cdf2d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfd84dbf82e688a307326f1f6320dd779733c6037265ede5a7847909390ad03e6b5d023811b5a3186c48a4a33a79c93ad73138fc9a2041916e19d01d262b2790e15b7df215d2648554362d3a5c83506bf855aacd0a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2bbc18a6cfa0e8ccd5410f1b399df9430a3b5431aae80024174f6d70fa7444c3c874c3e4471f18a005b3cb3f6a64a4b62fec8aefb81f58e97e800b5938029e65c17987a773aef4bd8519e92ff64fbec2f9fc8de5;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h267e29c4f7667760abcc2634c17c59dd541bea14f39f3f7ca6d0b7e70e2e5a9f0f33ebf21facc52ca56675317e1897ad7549118593e1f3e242853cbc8789d347cbb8efb5e79aa469e974147f434adfe7bd0f17a56;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6d480808c53db0cd368bbc664ad924e66f48f096150d2861ea3d19cbf52219c7d51719c887e4795c3b0c940c5b26702c44ef5ab5336b3dca54fd8c016e1ffe4bd95d895c3ee94c12839409a83bf5cb48c78a3928;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h597e5deffff9cc9d28064792c7d06cc8fc69917af1210b045d3e710cf0d6f5d799e0f2ff0585b42b6728be87314317877f2cc090f99b7a567c8b4fa8fd097c0fbf49eafd5a68a7cee8ac4bdc69f58021ac8d29b04;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h23fe7d67c10b972251c4800485b1b2551b99f4a060592e627a49d3861943c97bc59aeb996ac2121e82208e603623f6a1ecfdd507e511fb8f29ffefde4c3e7e9eaa3a9895f545cbe1dafbe1259d1334a9471517415;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc2d683d57f65a15f638ab0f69c397a95b9e7d487d0f7786e345720fdae492c71dc19a97206c89f52aa2f42f5e2436a51657749000beccfa6e24f4689266201ab063d0b9a6b05efbd4cf0627d9a5c84b15d2bf3797;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8466fe68bbaa684ed0761ff17e4ff5a1c42c3bc9b3f14cdc0a01841f20a86d8275b8513651fff0fce4a2fe398e166a476dc1918346d3a39a61e3143f6ae13b74dd6fc8c9f92f01c527fc9082a82bdbf452e9b7a24;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1eb4bf7800b3336cfcae94f58244025bcee8ab3e3e33bc84582d8fd71ff4f440e3082d9df60461f048f18c55956050288e8d64e5a1f57ea741c209fb08f7f9bffa13fd97948ee5ea2de6cd049191f7e42d11805f4;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfbc1ad92ad443d5daad99ef621a356959484505d71d406bc69c26a0138b0f5382ed096e095b90ab2b282f803f88717febf3dac25069331aa815b720d63b362b4765c5ee15339e8790b706486de888376b42a91040;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hdee440b32fb95de582b3cd88e2b64431efcaeb6575a1ca1b6009faee9b0d91a4fbcdff5d59fad13a552efe2c14825c9db92017c9b584ca5e5cf0e44cfc8e3daef3d021b948362643c82abce0a6ae4040754270c0a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8a87b214de9d624d7326a6cf754e1afb0826e122d1cf452d0bff76eb80bda0fb6a6da9984bab80646194f635ca456513b62c3c57d67a1eccdb45dbc22c02fe62fc241b1cfefe9cd496af44ea9d23b4f391d3beb1d;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h97926bcd109564214cc1464dbbc16060601aba27a386042842eea29cd7b100d132be6ad5136078acd9d01d8747b2517cad0b6a88b4141e54b175c7cecc5c3f2f01e5f50a239a4aba3784af922baa0802a43fbf918;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h507bbcc88affdf364a5c5f8ebb8de321efbf47128fc4a698f4c8e91454c87383b1b3049fe8d88a82f136774e44a36c11978bd53c329f0b84691bb742f5086d5fefbf2abef8834d915c9c9a1f976863ed1cde59378;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc9bd0cd6b12e415bb8ddb5b3c20f9b7cf0fbdc686d12cd823eef68b5b67fa2a8760b963e3cd9bef5ea671131eb35638f441af7225df384b5d42539796f066c2d4465e43296ce929d132b6615a871cce64226a1bec;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9f5c95e751ed26821d27e3d69b6204095a7f891fc9b9d099cfbe2d62654ce25a958ecbc491906cc25bc8ecc2538ff6097d1c6bb7d15a13a78eea874f501d8d177e81bd5ade09c63740f287c500d192160c55d20a8;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf9c6027486651fc7361c6ba2f635b6e0c510f37723bbd8347d8e7cae38c4ddb376ada8f99351c307e97f849e0189b84f0ecd8ef677ec4c2b22abd54dd5aba59d9cec6b6686b4d20579e7825a64d5fe818ed30fdc8;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc13805346ebd462928b1f5fffc40658223cbee9e4f644c29dfd1fd72feb6ead5147bac23aefdaae52f4d70638a9829e1ff76d01ad042e4550c3432f8ecb4fa42ef0d255fb57e59536c109414cb6ae11b75a24b0d2;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc77db93863b24b8fd25913a80db0a2a2cd4d150b6c3af3284b8e0b5a46cf065e15203937b5b35a94f4eba9be53bf935695bb24b6bf0a02d593667d58cb80552ecbea5e6419cabe78346296c8d7c6ff3dff16d3679;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf374b24d9b457c73513118c3526b3fc7d25de1ff8ec727e0e45c6beb154f9c655e4d38b0d0d81a81436a78331196add8618703c5533d6fec35562f1c91a3dca0db6634a854ca6fc581b6f03f04ba66cc24c622491;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd7e9fbbf36a1b91bb87d6cbebd66ecd5acefa0b0369aaa05ed14193ffeba9d1eb622623b17380bc11437acf4eede1583927e951cec9fd8d5295ad6f05a368ffb6cb9d4ac8a637cda44cf6ac02f1fb70eb1b6ab677;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h898d6fe01ab70b7919eb88b00325f991ecb7262f9216484a2e098b9a6f6ae12a81cc50220c5796beed1554d0a11527ca7591da9236b32aa23093baec3b684f2c4fe6cf3fcaba43393f92200d113abfb42d0a88712;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'habc139c60341d72326f30e9095bad236012420e63c53933e7bec9b2e4fca638b2d2b3f03924ae12db5fcad77ecea5ab461c05878d45962823e2c2b926d92ca4a2b0c0ade3aff147150a4932b9b0feaa1e3d8ef08;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbe397ceac312a454b7f1f58393781313a57b419a48a74305da552bc5cfd9182ee9c49c383e27304e3c5ff97d24a90df6ffc553421808f19e2c737135c85656b2a75c4cedf2f087e49b9bbb746079fc84ce5a5ddbe;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd15f9089ee9295b86b4766c8def8cb17954711fd26386c6b72c636044501bff5428f994271a4714dbcb4c9343d685e7bcacec2cd21bab42f063a0a148b267d0ffc4c547e02564d9bf743fc30b9f8ab8036cffdfd2;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h455c6a8d0d7388f26feeeb33ee11c3490b2117a522c1bec94b893d7923ab6e11914ce304d95c0e8307700db39460e54ff8b8e4b24041973426987d705779ef134c580265e61381c964f7a932c8ab9f8d616dfa234;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc102109d319cf470a1ef8b4512051f78ff6b103850969def5973976c4601e547941605aaf6f792416afee79a291e9fe2357196acdbdbaf3b505519924f5b5e43dd36e030841bed2234edaecc0b8f7b9b8040c9bbc;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h278d86a0beb72b0c53ebdfef636ca18e492eb9cb730bd93d1215adf1610e66d092b0ceec2a20906d6f94cc858eb97e1abc1c8b1a8dc1210ba5c5ead447ea5b141728918269cd19d766edc1737d58e3e7133c4a801;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h13a47642faeb335d2927bffd17e2a6f427ee17695d8a7feef584f6df24a42d997d10a7a2075c924cf4e3a8fb4bdf86ece239e225c0bdc73daaeccbb616f70629087e91e84405d9b7660d01c7186e973bf2b5c6dba;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6df3aab0fdd5ca39da4504d8773b57ebac86555826255679a01ad26b502c6f32377db2e07fa00d9d6e11c417ef7eb816928a291285f7ec1794904b17b5179da1718d0bcb2557f17d03cfb76a6ad41a28a3d7b6b0a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb8a80273f8392eabb8c36e1ae8112e3811d0fb92f5ccced3afd7058abdde48dffda400ded8b30a895424671c2ca5c7e3ca2ce5bb8445ce0e268e94422c70756426eb380eae8c05dba12cfed310a81ff93e94b0304;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h208549d36b1e4d6d2c1edae5373ba654e79365d555b067846b22442b941999738d5d03c567425d2afe3f5df5ce4620b67fe33775ab8250b04252feed52bbe1a6ee7b88cd87e2a316a7ef7804790b5a84552d22c40;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3e2b994fe2ae9d4605ccd19539bd543a8e4a3c47a3747aad9cb6745a7fe64f41b81f95104eb2b635803be58853600abf942cab9c7b1dd5a13842526587df2c08b0703077260cf0dc45255c3b86579c2fc3e589d93;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'haac0b926e07f4685d98e96b2e28456bc77feee400ef591ab55e2d1058f6c6c331e327bbe2a01edc31c2b49bea6c7d3c3c052ccfe0880a2fb681257be4b7a4d1ebd64774de1c576b63335586d0f543c4c56fcec8b9;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9314429d36a6625784fcc134e2587b911ed515afb050cea9326ba3828fa7673ae9f65b2f33f78615108b66f682c15e5f52721ed81702f15e834ffbf7cfe8af31822293789c2611291c21040f2cf3d257725ad7b10;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6858163155cc33a92f77d30594223cf0c863c48776a3918ef3c5eeb0d05386132ad1886d93a1b6f2505fdbfd3f309c9457bc1dba5e6352fd957dbb600feda64965e5c85aa134bcbf299faf65d0a6739c2dc4b90f6;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3280deb2a45cfc02c62099e7e679df1388f63ba639323b439a30ff85fcbcfbe22ccd6380633b1af668f904091fe87e4a790ca641c03a0ea144665821d6beef9dc284440b2383bd882aa036387ca64e931a4ac8853;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h16596dc95bb1ac0669cc15d8f9c96d3b4838e86d2082fd69ad667ac4bb18dd991f26d5d39c4ce28e9027b2d2a9cfb30fe493841bfc597506345bea0109a049707380446658a1dcc734d5c5468ace190548f3e86b7;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8131a2b807e42a03866fcdfde2ae2b56ad8acbb60b42dff1aa10eba2945f3269a8715a1b9503e1a9e9be44e6e35dc03e3a3cb76cb91e899736b76e3c644daacfb09cd6ba98e494a708070ece3a4fc916acc27ff46;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h690a7ded50abdfea96471177c70f5223721e17e1cce430876d003f77e2cb0b384b094f1303d43be1872441949be6fa69fdaa1e4c5e367fdecb59419e9c771ff69f60a4a769490c7817d28e64a314ea4e674f653f6;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf807c7a834434af8eddacba619b978d794ed20037f8636e6f06aebd18df5e3e88a814ae9032e739c372422a4e0d2e6f0dcc84c96016f658b8355d3a3b9c7d7b47b3dc45955c8811924d95660ca0fc77a3a03b130f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5ce648c60227afec2ff67588e0b268436342acf3ad95a748e42aa67d7a9a63f134fe0731355e7e9144dc739eff83385784d79145537fff1f4919254ec7ccff17a9230de83715622227a068bdd9b5ae149df8c4c90;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2812475dbbcd6402221098c54f7fc9a9e1e5364d803ccb0f107c1e6212b91271f4fbc8259f526ebd1e5f0156f18e7e63c06dc69f359bd3cbc4ca94e6852d68b91ef6502894080d6a46f3cba3d6c7ae8770f513780;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h820de55502d1f05635ab8c576e518946ce4606ecf08bf974371d53d61cf8a00b8be5727ce86f06f56d5de3704c2b5df90bb34ac52c7f9097c834a8858e547a14f81606c81dcb0db24205a3755b8ccca2afcf6f161;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hac85df22744a54b3557d7f3dec2826ebd8ec0c3dad311d2c48e044da2f7d2b5d8af390a0fa7e02807cd9a1c62b6e327b101d03c8128082ab1b26a833c020f8add5471b6ead81df26276a6b98fc3240e39c6bb320f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf8a172bc6a0b1e5cff85e2f3b002394bff785ed6ea823a040202c8405413570335ad95fba5989626ecccb39d4fea2a204d9d2bd45e42272263b17537a686398d5ec72eb016a171ae018692a52ca845979c7e38c22;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h124836fce50a537b5011742eabb2cc8133e5e29dd13f96305c6d1861c4ca48db3b736a04f92f8c2f82686febaa2a2e025d6be5aa02fe108a15781836afeca05ef768d010d0188a763069fd1e2917e2a15a3f48063;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h234efaac9a648c43838d4af36e0d93046d3812fb43b87dc79aa0f6b8a53977878ade91f96688ff2148e7c4ea09c3ab7f76f445132ead9e28efd2a9c31d838b92fad56c28a57c68311ba67d81539d9a1cda8cb8323;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4ece897707b1241c3073f79a2610e5dd210b12069071b9474b9931f9e4cc5525a5cc4c5f2bd269cd120905568170f1f3b71f98a7204fb9fd6fe716d004b1517a8bf91c96a4862758454bb7724547a576fc430697f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc265bac847b65f95ed615cc6b7ee813a12336b9c7d21d9f98961f9b1e3f5a0c0b1ef8e8706f6adc72700277f5bcbbcbd9095e0083080fab50cbf691cb950c0a65bc8666b5c1e43bf6347f640dd3264f402a379e09;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd8acbf2ea66636f7ddf2f2814bc22d585798fce3b9d6937fb8b325ad5a24688bb4e1acdd52dddda35a3be5f1d57f0947d50dd99d3636594475cda0fd8ae72c270445cef65a5216e0b0c824011d1bc227361f1376b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5e5956485d684ac24c51f465d738fc166cbb404923d62f2d37cea3e440bcbfdd0f4f342f217be3ba7e7c55540119e764207bc976e737777b8e8f28f98079bbea90f4802cdc43d291649311702ee1f5f036c3b23df;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5e731d3b291d829b7cade04176c7e5b274cba560612c34fe50ca5f95eae66170b0734528ec7167d3957f7b6e4ca89d95b46986c1d79a0d4f1ebfef6bb9020eaffcd93ceaeff602afcd914e929138d7e74db0a2c88;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7877aba6e4472145adbd3fad8e2a1669181c5ef6fb3a2220de99051eb833814ed47791865c66826fc43d14ecd7be09206f2c996f5cca3b069573c5ee67f3b784285fae61ed5ee0b4803e9970f3df7635247caf250;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4a8dd0f159503f00f4762d28c75f310125174189c076583ceb2a0941c512b9df09adbc8250ff97ad96d0b591ab2c9d70a662cce149b6695fd40cefc7ddb9e89c06ff8028548c5eb706d8adf0184444537c0b7e88a;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6fb53c0337ed7ad4ec45547f3284b6c3725d38ab55477d68b0c571cbb6a75afe2292f396402151db0326222a8ac45ec73f73e0ade69056db852c7917d122ce2c5e6612cf0b535ba69012a0868ff149d7a818cdc5b;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2118253ee29e8a157499ecccb193c8c9fa5327a0c920db58faba5f9fa4248aa3cb24eaffead32a774db5ec3f6b1fa8ce195b7ef94a4b6fdb4794f8c83e3c4e67ec0bf4f4fc058cad8b16d408a39ef7b7f7da49968;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h97f8f5128a7fd3061324f4bd8b11a879e22d3fa1ab9eea1ee3007a9a047849774c8907e374b4e2fbd0e9fd314a8ffa88bdc29e6da4379130fdea50a5eb8505f6a9fe3ad3bda3fc7a466b07264189576e234dacbab;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3a1e40c7c91ac2f7e3a24cca8b80a05e0bd03f32e01e42b7761331236c425eb111cb1bd641864522c0cc89648b7bc6fa802282540b90789c2614e62382d0c376437b1431a018e3eb4213f6be901deddaac729f4ac;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha14a09057ca73baefb247bfe2de2e6cf22f993fba32b74213cbf7c84d71c3c9934511748eed7066e660de3434ddac01b21280559936f7df4a970a45a6a2718cb93c0c3b83ca97ece221e5889409104b225bb7e43f;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hda7d11e669b76602fa0a9809d4103af024e70c7395a9e418e69e8a8e390e0438973e038b83de1af92b3dc0557c83df3e2f0f07b4655bfdbe932f7b7a9b16bb596ce364a5105b258bc00e950512c8b7b3f6c8b29ae;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4168c84c8d82d5d186087f498335800ef30d07e546fc05d22076aa1ef097949dd0558f9d0073ce975765a153493da51e0060b88edacbb44f1f07371507eb5179d45109bee4fe465c2fe39277b924aa13e521abffe;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc4fa64d09073de13457dec01cde5b4dcafece0c7b0f6bcd45f5091caef4b08c95cd5c6c96f7f5b0b005a3a68d933dfe82f82453b64984c405e630c02f0cfc8fa03ed967fb2684ef196facc74a750b2a1ae0357891;
        #1
        {src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2e3ed212e1486cc83c05961906ba0cf5d5bab952fd3b8bf13049d73de045567c2968a88d5a88c18129f4f93a48bc08a73e3cb12a2aa10c27d3905c80d6a231af6e455bfefd1fe901fa2ba768e8f3e965daf9f4a4f;
        #1
        $finish();
    end
endmodule
