module testbench();
    reg [12:0] src0;
    reg [12:0] src1;
    reg [12:0] src2;
    reg [12:0] src3;
    reg [12:0] src4;
    reg [12:0] src5;
    reg [12:0] src6;
    reg [12:0] src7;
    reg [12:0] src8;
    reg [12:0] src9;
    reg [12:0] src10;
    reg [12:0] src11;
    reg [12:0] src12;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [16:0] srcsum;
    wire [16:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12])<<12);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h0;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1ffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h158f73003073671b80a629d598f7501bb8c97bb6cc1;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h156bacefbe44960f1adcd32f88bd4eea3436b8d37e1;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h153b61f3475bbfd87553b771fabf59f6d46f6319dd9;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h18847c2aa67dbaf3e8ac7ef72396bc48253a901830b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h7816151b9987c7131514fe28d37e6645024bcc7994;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h6056c945670b17da37c8253ab9eb2c2c7411ef739b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1c2b844d26dc749ece96ae6f323fbfb12c74a03aa9d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hee01b842464461db32de5793cb380716a3c2a63c21;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hafd32f148d13451428bb8e91975c0788f819db0d62;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h4618c5ec4a774304df74d6e17c56490bd81197d6;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hdd2a93858fd32bc35ddcba6a6f65e9c543af1218d7;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h17273c17254eefbdd2d879272115c81e66e6703673f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h9c2883a44d0bc59006059305736f0850a33dcec381;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hc20627fa0b6e154649c4b5685a5a52d8591eb58df3;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h7ce2260927bca7fc6318d47dabaf3f6efe4fa2c79c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h16c5c6701bab1f679a3a7d67dbc26a919c732d70d5f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1eebf55f777e6f8e9cdb86a86071e165bc48713d800;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h271892085795bdf8207cd647cb1f11034dbd959a75;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h14678adc01551a508e6e0f39b1a76df8bee66224cc;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h17a1a47a46a22b529e041fd9ef198e930533c006d8d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h6ffe69a53fe61abab14d6d2b111f0fc7cb0b72a54e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1ac9914bf11daa68d5ceb503b7d09229090d051488d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'ha6b5ea692ab3f0d66208d06d3dbe0be14d1fa7de0e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h9bf3407e9cc115b46e517ebe90d3db53f905ba4926;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h14cfec1c8f14a8e0cc9395e2dd88acc290fdb3709df;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1984437ac7b1022f20d430dd90549d2949d9fe59071;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h18b025f9cec3074478708bfbe3dfd320d69d77b75d7;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h10d6077e8570514f880a3290f903d88e5cf5b5a1961;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'ha286805197a5abca9ca09d8f84b208b25c5edc4b3c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h91b34e7f852ade3df2b66a538b169392a2ae91ea85;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h5b6a46a1112208a108de8043c4ef9352fa845161e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'had37c509e227e19d2245f5e085d9c75f4fb621ee81;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h123d7ea5a75ac55b671132668df0d23cdffcd25fc08;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h11c60e2757a9280d081c581e5f0b8eaa94dbbf1f9e9;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h765224208a81946454335d6fd5b482102c7bd32a48;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h9c2e72f542c0c0afc761d782e44f31d79cd51118e5;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h187193e7423e513580ef930253ae8e7827ed003cba;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1e3a4796978fe23710b169922d2d73a6766139afcd4;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h8cff5bc1b430422161455bdcf927406c851960cebc;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1833ba4f11a5068b4b4eef864c375ded0e28b418e3b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h9c73ab5f50de79f7850e33cb5d24eaea7291a61dcb;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1aca042e29eab6f1da90e4f2ef752189c564ef141b3;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h6861b3bb008cef9a8fb80b7b059bd9433623d45bba;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hde93f49e36ac8aaf9b54ae9049b255d2952d6c5042;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1cdcda912117df517a5d126e416e533bf8e763e50d0;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'ha355e60183e4e9ee4e29716d8ec66ca44aef5f2851;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h101f525936e1e0196d2118bf46b9087504aed558193;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h6316a6b4f75e57d1257030b2f38732a2b5ac83baf6;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h18f206b032b221bfd3346414aea62a77b32c34eb27f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1857b425f4262063b24c62ab370b0462024e609a7bc;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h175ff9715eab7917ab2fca302ec21e3adbcab0502fd;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h381e467992b2a4558e9ac466c0790dadba790afa7e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h2416e73f12bb566433e6742590a5a8fd3d65d8b2b5;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1ad35b3493b07575a81e1bb0cc614a64e6eb30a6c71;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1d6089a31369952e729a72fac2688a66186a0c0e10a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h17844dd7e6b0d31547178c10d15c77f97d9ed7e6946;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hea98fc2d5866cd5f89c3c7485f7fae7b5a136ff0ca;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h14c77f1f08c001db46757ba065861f33e80b58f4730;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1cebc376533653b6f2a3fd56dce46b15a20b6943356;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h147d1a123651f53c8d9c9c53b5befad99366fb5c0df;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h22ecbc4cdf383787b67cc817a0b56c9bf2b3d6cf02;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h6972c850ac068eb4ec124d4ec9ba8ab6713e2b5d3e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1ade40bf381cc240700172ace31a5ecfacc1854c584;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hc6de64fab23c7ddd93b95973df7b1e06994a436c74;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hfe3acd8594c0f6e4579c5ff0f80008736088a44984;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1f4e9b84056005c51b33d24e5c3ffdffe94616f425b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h2c5839574b92ace252bcbe637f3e081fa69f33db5d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1c3f8b21a638ae8192d4889118d46be886cf46a86be;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hb7f16193266c9662e73521b99e6654b768b142d877;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1cf0065171caaa654cfbce5f3c09d788e6f2c39d1bb;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h12405e4d6fdea1456c2c043cc23ee3193f1a892b6e8;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h14b5e1eacdc2eb3194aad03eaf920167f19a8041aad;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1a314c7317662fec7cdf7544c41f493dc5394c32796;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h585fbd98548c20d226db914c76cde96590b126dea2;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hd98deb0cfc794dcb03695f711d00b9b35504490d8e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1baf091ece3f1ce8b0ab9f1a2258817c08e8b6b69f3;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hff28e5ebf012965a244e8eeb116457b759caf13906;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hd15c3b50888afa72fae9f427c288e6256b7df34cce;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hc18fc95e6fa9acd72541dd39cacfeab821dbf614a2;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'ha26efbf2aa3dfe02c6f2fab700145fc38ffc455da0;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h4940b29e019f7dad9b15661f2c420a1539bf4e0cf1;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h6fccdfad6651805abaa23029e23535e873526c46bb;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'ha505e2e0f479f98618323fdfa9a571fb3f68311e31;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'ha246b69a0911a510bc051548a94198f9a6827331a5;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h161379c13239715d501fda4a6671aed56b1c0b8d68;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h55fe389cb4a0c3272144feab940efdfa27962a7856;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1209bfee099bf9969ecb4f85309b7e71e781a23de9d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1ae168357b456baf6f5eb4195b32c7481007ee8c706;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h7ca0a512c9a9ec33009d9391c7cf8b9fc1f214441f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h18e67ebb81936f021932a5cb991fb58ed258ec30ce9;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1f2ceadee04081d25972495120e131d64044a57e3d7;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1be418ccfefa0ce8ccc6aad1aea084e992d288dfb0c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1bdae3853563d7863e3ea28ef760393f08d428ebb97;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h173e7512be1e95fb469b036056ddaded3a750b66749;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1fbeeb837e5ef6fa2283790b0124070d165d52b83cd;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h16924cf03fe4e43ea1fa88d70c8bb6624db3a8ddd3c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1712b606481dce36aebda6bc5083f106b98e4375c77;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h12b193288793bcc4a56fe6ce08cd500334d4a8092a7;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1f6d165e191049a119da815655e83e3d05572f882a1;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hee02c3526c262f2848138b68b11c208010b45b1d0a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1390584f2520ec3d66715862c7605e4c99e0520f60a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h705c14fc761da6873c50e015351d97c9eb5bcc6c03;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1d893ce5e60ab2396cc1cfd82a759215ed8c3db8a82;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hdbc8b6938c25aacbde4fe6aea37184e15b761e7255;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h2f20fd63f38a1210c6c56985aa6c26ba5ff3fbb262;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hf54fc1ca4390254b8010007f3b07999ea51b178c3;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'haae4de600a7438bd8147eaca6752e4cf7499341cea;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h13f8e6636ecca3f16c8af902138940a41f680ffbe7c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1a844b325bc43c7440a4ca18585a5b75c939886158c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h66c1648ba916d4c13ecc4228afcf9836e15147781e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hc855435b25dad0b4d8ebd9e8f7ea2c3820034c5ec0;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1e5e8c7337b9e42730e3eccb682c092b8e6319acb65;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h123a344ae52d206921736da0eb524c46e0e7e12e58b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hcda63b6f7d386d92968e7f0ef0fdf0bf45519c7c7f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1f9c64ccbbd9d6eda41087da7a299bd60a6066eacc8;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h114d30f13089825569f9b7388a80b9c83e7b4b6eaf9;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h11893c1e9282588c94b2fa086e2aeaa4d8ee33f0b26;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h3cd39668250c450d77490194f314dbb8bca66b228a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he15096fc0815ed0171ef6d331f4e3ef63a632554fa;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hd9759299f957e84743139f6cc1ff93bf8b98eff92c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1150be09f462b3f0b7ee2b94b019184d750968a06bd;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h10043cf611e8fe0958fadfa2ec14ced4d83dfc049d8;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1129a27ee5f537f1ae2b430531cb9dd0a1a08f7f9d7;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1be39b5878fc2db7be5e97702e1bfb142bf38ed367f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h10de2101e539d184f59875a05ffd4c52aed4c9e80b7;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h18afae6cb86512a4c4dc2aefcb7d7b641a2e83662d2;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h103454c9824a2edd883715161503d512fc238a24a59;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h15f1e74dcf590632c4b3f5e26a305813be19101d8cd;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h145ba48e1a7c861118e0fb903fc37b3f0578089b5fc;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1034d1c242da4677ec72a1b21a6320debc023fb357;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h46651aa29ff60dbeb5ba7949b25d1d93f7f9b2957e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1a66927b3f1ed675052fdcfab37902c3961fdb72bba;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hbd4ea593e2d9ad20e5fa6d2dc7e6b6a47e531dad17;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'haa4b42f20b0e2d6497cfd7b3499077781f527bd241;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1b187ed6f05210aa0e070a0a9534c8b49160223d8a8;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hf3abf0f2dad259978d6bc3aa22c46e3d0020ddcefe;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1fcdbc2c6f4fc8339b5bad7e6bc440524b54175451d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h138bfe18ac4a8771c107fb2bac9759d1300554445a0;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1ddba08baa980bc0da4b56c9eb6a4a0c74531522932;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1cd6d9a437bd59090d1a81c37446337358a816f774d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1eea255737a07704c5d2b45eb5c1a26d01ef747263;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h148c7bf692ed9a43d56696510253284157ef0686dd5;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1b1dca51fb19b90a647b65f1aa70b0424fbd3638a6c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h57ae56b6ab60b67f015bebbb421d94bee777113560;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1e8424a79a39c484ac793ea6743b1750d4eb57900e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1f80975dc9e8b7475ae323bbed195d99a8dcd7feef2;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1df8ef6e61cc407c05b3ac03da2cc66447e1e7c0a16;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h14a23797198fcee2ac2315485cdf8e56d09c725b8d5;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1c875c808340916872bd55558b2ef58e24498378fff;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h12b0acf22cb31794b143f0027055c300bf768678418;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h20a69915342f102fd53ae5d2a8ba6ba43fd8fa482c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h4e583dba47c26cba1a3c65965ea81975b80179ab53;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h10843fc2fa02cc11306137acda74fd7d26c58cf679b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h6fbeb73ba1e8f0a68948da2e7095d0269d1a2b88a5;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1ebec6a32e5a27a3fd8c666d474a015a6e953f10689;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1789140f4ae4bc76bfee96bbe4d9d2965277b795c84;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hb20005665ff82aba4fad48ca656e2f1ac4ba1efb32;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h113ea044442b7e751e8e7b61c9430148065d45c6d55;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h29f378aa064f102193746f64faebe99dac04471b5f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h13d2db34d85f24adb9c1d6797bdd22cc3b701bc7b7f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h10c63ccfe6f93b54c780dbf92b046b3698537258c09;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'ha769e2f4b892f8ce7af8e72fbf121c99516ba37959;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1192ede7b39744084304d92b981e737b86211ceefe1;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hb50bcc1600959f55095b6907eeaf0da0917a9795c5;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h19b990b96fdddf73e4b709903b2f047ab501844e199;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hec013ff6b87715586074f72bdfddf1ec9156950a7d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1e1d5c521dc92db486e6430407c289dd9c146ffa864;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h14e32c69ed52e573efffae8cdb622069614d68f77ed;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1825eb33fe16b48041c79dbb2161afcb445f866098d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h5e46ffb7730db48b6bd747e0ab67f736e0fa1f461a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he2b311c41fb74659b5c6b4375a4345530c89b1e31b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h9c7d94d4a8199567b42857b57641f1374c6dbe71d9;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h15ba9fbbc9791a0c7350e990c6e231eea38fed623ce;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h82f8b050939f7261ad4944999e3b433667dfceba17;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h133b4d100587f5cc4b7e2df3c023fc0ee4f52681d07;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1e7e6844ca29c1a278ae7950c005d5f41f6aec742ef;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h163540af64e879de146f5dd8864f342f34e99db3272;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1d90ef2c14a8d78e52e9ae87f9a8d4035408dad9865;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h10925736831628dc28c0a1e82e268db9f1606b1c28a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h6161362582a0e6a9be36463205be10e022686463e1;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h162ee0a1c6ef8fe31afc67abe43568181e25ebe8489;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hecfe9f8f1e98800b1a704e79a5ef69a8f331f29b74;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hfc338f597d9e214673d4c10ae8e7a464d9e3a81f28;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1da75f6dbcf8470101d14e3166edd9467f25d970be3;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1e37c56d49bf5a5bed65d2171d68a12b277db76f5e5;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h19cb7b2c21829579b5ce8427c3b3e9b816f32baecbc;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h7366873d73c28f6219803b0744d8e6a73f5683da39;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h162244acb76946edde62befe295d820a652b78b5870;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1d7d069b2d060537f92b571ca878e018deee2593d35;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h50fd365378f1b9e0501f025edbe566d80a118b586e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h13901807c237f5d244df394f7d75209b78641765f37;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1634eb0767c9cfa40cfc9b76b86f110c9ea6a03c554;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hae7856abe6ea5260b9fb95ed1330e7c6085e96dbae;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h108f44a27e905d636b54645766b282666b32623df3e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hd9933f83cb45e0eef91713f2afbc85b8ce6b47980c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he5d82289f1c039688cffe8b1bf293151b2c8238290;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h12b85977a1e19ba1a0c416d18c4e9e47261f8e85ac0;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h60f874025d0c454342bfd17cbbae23de4fc2bc79ed;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hb2b151fd67a7db0693712633de381fb2f583d5b927;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1824592bd8b0c038f80ce0c94470063fb16abadece4;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h13588498fca025e5d8dd9c241291dd687e09001efe0;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hf2e168be8db3b62882fbb60065a50461a2a26572e0;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h7dc4c1ae3e0f7f87bada2898df42c74244c026b53;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1f8d4f6903fe1d439cc89c2248a08ac09ade92e1759;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he67ff3303379cc62082773dbdcf720319f45228dcd;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h8baf14eb96ebcb2fdfbbecbeadd4dbe400f6e8f682;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hbf2e487c18ef6dfa48b9a390ff66d1ed70d43cc158;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h18948e69a64ef0430dafed18e637bd943a47a1ea050;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h19548c6736feb71e01982109fe8629da4931731da0f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h71fb9c9b4825a30526572f73b3de1dae87f48e4323;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hfcd7021c67a0eccf08c2c6af95eeac6d133a316322;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hd438afbb93729ff6b27d1b40f42910d33e18421589;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h4a2e39f46078b03e03f8a0c5c70d6bdff47a558a5f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h9f706af6eba2e0945938b83701ab1f1749c0218279;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hef8ee89033f786e751c283c35c2c42d67adbdde995;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h3225be60deca562ea5a9ab32a5103902172da6aa18;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1e6b1ec6deab705281b2e9aaaaa7b88cbd08072837c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h82163f95a709d2a99f031310388a363e3487a03b28;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hbf4829dce70a11403816b81d5ccab0a3486cbeda20;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hcf38ec2d194e61ec281053e5f01cff44a3eb5c8b70;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h10fff5540d2a0192caabde7c9073e55cac83f8408f3;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h798738c3378fd3bda23c3c5fa9fbaac8eefa58ffc;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h18de252b2b5b1964bed1fb211808fa181515d7db47;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1a064c4ceda9481e40aa86f319744e047947502275b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h10180bea18b7403736a4bd6ee926289fc3ae4b4444d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hd02fadb28c47ae186ceaf3087bd8ba9735fcf1637f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h7eafa2e12355de7d23d48a429a844d530528ac6761;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1d057d6c050ba713f7c1ca3c5169fd57ead778844c3;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hd687f7ba56ae589693419300e98c1356b911abcdb3;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1c89cf492a252813d9a9248d0c7a73cd4f7878effdb;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1e73b929d40825e471c28311e6f7738b83ea997e6ac;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h6811b4ceab7130007a587e42ba7b2f7f72d31d246d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h11083bbb44eb9b7edb3a8265f23b5e818ed1cc46fb2;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h18e46ceed44d0139e7c280c8e191cc81b95995f93c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1eada1a2d2d15be245756202b4b7b0b6d414cb547d4;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1bd7abf17742e6b678413fc5b8087303bfb541aa926;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h123181865160b0051513ec20818e2e05559cb2c29a2;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h18b3f6eadbc14f00a909c7b3ac55977484728391b9;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h13c157e9120df1af501e73b10c3d7171560e581ee3c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1ede0f657d1ae1c0410ef84268b4ca1117aab16ecdd;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1e6ba940e9a5d14de4b264004c94a11beb1339221a7;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1bf24e0f977aea84f87d50bdd1b9f6c65b43e72e589;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hf19e2ee53af7508f6001388f16633f0eeec23d8ccd;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h62d773fe52aab7e020f0339da4c2abcad95f5b58c0;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h2ea91b1aa2ef81f59d482b04a083fdd5fac93efb5c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h2ff45185569ed3e363fba8c48bf6c9126af8f7dc8e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'ha8096b2c26f3a02417e45a668a00fc8d2ed194e421;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1e0c904c24e98038351c488857dab6aa7298c31da76;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hf61d2165e6f7d5452ba1d158aa88a70da0bea92a5f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h17b52bf5b97c549e5e5e728ac63dff1afaf61ebed0d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h64b6514b7e547d8055c41fa00672b8f0738f3ec6f0;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1a6e9d8070539809da66700ff6110374db5e019bd77;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h147c8d9c2acf0cc25857a05d3a8b466388e196d7bf3;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1755a188405850a7f2505f6c47569ab3a6217b8fa0c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hf5ae197786e18d3e41205df449a8d0092293e38358;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h3e7aab4afe18ba9d2baf94122513cefdfc44196256;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h7c821656ff20f77080ccc6ae357b152cae5cc3f948;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h675ea6754ba759d9bab6223f270e20a7381a5cfbd6;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h9b395ef4fb86d6fc4ab9f7ba160953b2fa59c218fd;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1d750c4618b72096bd466214bdee760bba9108c874c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h12e57271e7bc0027c3ddcd40134de42990928a2ae29;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1c7e614da82ec1a2623a8a2aee8121c5ae6df4fcf37;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h86dc15a330b609db41acb632e4a3bd020c733ada20;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1cae77c075dc220096a9ca7002807a4736a46c64e3b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1034f4d990f9f2df333d75cfde1a0cb2f574870611e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1497287d2679fa0966a1afead01e3533668170dccb2;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h102856aa51175255d20b6a874d99b34416dec94b085;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h81f3a0d03d829a88720cc122b9e5d28f7b9812e5a7;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h18d52b17a61f7f9c87f979a62446326457ac0e3be90;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he2ae15abe48e9629eac4ebad40332045df549c2e60;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h16bf69e5b57027b54d56dface889507b6b73c43b9ef;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hb0f3082f3398321a5b89817a8e025e9c098abd010d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h130d9a323a5ecefcaea162801b096f4910d9f4f76c0;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1640cb8695ee9f6dfe883d398d557783d985a7ec989;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hcd662d3adea9d94e38fbe8e755da2f669f4ca8fc40;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hf33733b1e0100436d514892e837cce51b974b1062d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h153ebde563b3429f84e492474919d7b841f9a5e4000;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h19a23ee32f160306284795884639a895d30575421ac;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h149eea2565ee542bf3a2103f605986026087655fbd4;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1a72b5a858a87ae412434a9117e48a6aafd540e8dbf;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h15ec7bdf3e4d91a9cb28fe3868f444166a57e1fa1c2;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hf67cdc6e9102f115601d12ea91b70e459cb4e08bf5;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hb7a22c7e5af9e9f5611a17f375444c2fc47905bd1b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hb82e1b0dddbe243ea9e68925eadfdea7380e01defd;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1ccdfe007c67bd4ea31fdb10bda17ae6d80d793a0b2;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h498d39707f65d4d7378894b91c3f0f5f8cadd75fb6;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h13817cae886f616a7a05ee870ea1bef5b1ef078ce3e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hd850b41310a6262c3f762bd1f55b7e7235e6282625;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hc890da54a0b4acef9f961b4285facf2a98264defc;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h969bc865b60d86ead09d703c0752e7b206a515bf91;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hfa1fb632a59e0dd26a2b226d0f3832f9a2756a3afd;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h19a13f0d9bd7860d564a363cb56dba15cdbd8dcd301;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h734a36cf1f9ef836c75908507698e882f88226a7c9;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h56f1106688b1ecba2057e9d366c8fc3a70369dcfcc;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1f3b724d6692b53f9ec60c3bdb277e7101452f45c6;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h178e7a6276b64a634217c8808a55b52be376a984e1a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h133556e09b77a09be179ea5e8d95e0b4ae4e3ea63af;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h74799717a206c15c4888cb86c3ce4a28f6e8fdd758;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h72699d354e420b7b860a6f495c4446e6b9aa3a90e5;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1464485790cc7c17f754d38ca1b14451ac0fa3a5302;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1e278af372f003473612d0f81858c88e9df27e3a560;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h63d9c1509968ea2b83d0981a1154c8fcb65aa6d10e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h105bcf73fea88370ff4a739bd526cb543fd6c3b8dca;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he9dac63259e83d467b53a09acf61723f8c4bccf75b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h19d9c0a1886cf50f512d0c8f20c81166acbdfa75cc0;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hc58b5d875e840a9be31d292499467780dfec0bc9b9;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h32bab13b30fa1b099aa2648ffaa024b6c249100318;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1fb54db8810a17fe3516098421e7a3293be21d841ff;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h14cdf598c34465a850095c035ec20658d4fd3f0a762;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hc3c3b78aa8e3419166774b4fd0f43a2a956e3c745e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h3e03edfa5b0cc48df570f035cc825ab537ff4ed925;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1b099d276105e1d881a5c1209333c83ea5212225dbc;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h11d84151d81bf9eb61a4faab0d5c71df0f048cbfb7b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1294304e251e194128473106af53013a3139f19d2de;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h13e644b434254959cd3ed5c32f93a13eda6f46ab0d8;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hd0590cd12d59c80cba19cc05cbab2aa3e6cc68a252;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h153e800c520d00d7107d6553b415158cb9330097f8e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hb566904cb27cb4ace44a3c94f34cf2a3cbd68be79b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h12f434a2b847cf7805ad0e6263ffcd0b03f6598a95c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1c056759db29227552bb6e5fa9bb330677c451d1b7e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h160021d1036841080663ae1705cb7ea19e93ecd8ea8;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1f6c80386091c613449e124221b183bbdceecaf6c29;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h9ebdca00458983ed26bd9936f21f16440bc5aa770b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hc56decb8129373cf24db707c45f6ce13dc2816d969;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hf8244a84842d3aae40645d5680097ae3093d7846f7;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1e272b598ee4b6d908b849bda7e252602248628b1b4;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h15e8a152d48a9d88007ab196535eb953402429dc92e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1cd65268d16611fbe4706466a875e941778812c3afa;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1235925eeeecf341bc5c48cc0a47ca6136d619ffa83;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hb0d7665e08c4633e88ff297e6df0b49f7385e00f0c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1e9e7a69cc57e697ae2f690e056f94c644c5e52fe1d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hfb5b5140227f6b39ada80d2d36df5150c3a9a3f308;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h2f07407142deb28bb79802c43fa7544dea6f25a185;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1a4a15d5ef597ebb1cfe1edf9d8f5a70eff34cd8da6;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h721d4e8d0a78173b7b7beba540c708064cd13a1561;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1bf87fcca974c17d3cec63e75d874c296c273b5211c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h863ec71b6877178c41dc7f7d6c0b245e1507207153;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1ffeb0987f52c117da1ec66ded774c290c6456079c0;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h742ed2eaf74a2128f6a09b746136f5059373b579b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1686c0fb8983bbe022098ef9f0f92c85ac9ebe80d44;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1fc77fef2b3fb3497478806576d373daf3ce504c3b3;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he34405bc2418651a8ed7faab8fef9978b3062cfeeb;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1021184816c41adfa12acb7e69fc05b25392dc84e0f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h10dc60c3404c68bc23f3770f739b8c52c270ea92a83;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hd8373dd6759921e54e66616c294a11e9c379b7bc5a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h689172da32e0645de839ef80715937fe20daaae146;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h197d0ab6693e22372fdd1abfcafd88e8fb942230f4b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hb8411e5e6710d2e4c9d998b016c96cd42925daaaaa;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1fa0f6ce67cd671a83e1143f2e97a7b89f82d614ecb;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1aaf6d05d4bce8e203a91f993f5c05fe0bf400b04a8;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hb4659634ddf5fb5c802c5def11baed9667f899303d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hba188412ed12949dcf279e1a72d6cde5185f8ace70;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hec092039b1f7b6fb04db378fd362e5e761cf9259f7;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hcc2e796ae2c9f1c4b3efd2ed9aaf332c0917809e90;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h2f17777b95d31c3a4f2d9ef016eca5b673d1146624;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h106cc09528ad462353cf07a52c89f9416a60123f48f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1773fe6038e19084cd0a6b9bcb9f4cd50e44b3a7bbf;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'ha2e0b617866106169984ff003b236543a7e564700b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1cc8698904ee62808b1cdfbbf85f178f2d70485d924;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he48bdb12c7fe0b0dc5e79d817b4a2f876e9e3fc337;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h17f30e8aabfb7302fb970ceae619ad92a6edebee24b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he15aac83edeb1f8cee8adffaba3db53365da570c3;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h12d520fce3773d9f34cc8e7953782c91ea7014ef993;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1b429768f85542b902fb73d1abdd9c43a27562acbde;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h157f93c5985b8ef388f452831a503e1b49a3091eb1;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1ec5a1643c00f2bf8c195bec28121b9cda36c311658;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h36adbb5e48858de53a3a258355133de719529e2415;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h11f2a1ef0f4e30e88a3bd3c86b88a298d6c8931a574;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h19b1d7de6a3a35d251d8323c32911f4ac0291e640dc;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1d2007cd71841d83b02ce4557ae1df409390b713631;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h14b3f01fcad5971cd411d07c19decd8dfc3a66e208f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h196e61d0de09d068acdea6ec403d4661e6a4efe76d5;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h7765bf8f739c0633f5cd9218655d7462a39b6a74e2;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h12e2c03dd1d2199a859e9e46163b863643cbbe973ec;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1edfb2912d20a553e28e07532d4f1581c516c77e605;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h15203733deed1c27b73f107bb509198b90048478f74;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h7be70de8d99e4e2dcc905641a8a74093b1e133039b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h479303ea2587577b58bf387e2ce6b85dd8b80412fd;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1cfb5e51e732b4501846a8af29fd6647ebe7ab2f78f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h18d4ab34ded012a356bcad4a8a27d0b54c4f36560f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1884184f2c85983ac5bf842980c47e3b8f1da54b93;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1c3c5d9d84b24220e6827375bb185d3838911594ff5;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1f1f99a5bf1d5c9912c4aaca31dbfe6dc5e1e3babd8;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h11270041840cf01e0adbdfeb25741ff35f58bf9e465;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h8adf2e30a6be1d8aad9a026c8dc7cd1be7f7bfc507;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hd00bb11758e8da27fc23e5c5a1702cef2a3a7ccb7d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h145b253fef4cb22a85fc124d10e0e61cb0f3f408f1b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h39be2830fb2abe8cf0e737faf5fbd1b5a59696eb16;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hfcdcc022cf0ca7afd561a1e18bf74011433de47096;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h4b2126d75a6dc2d46586deb10febd32c5fb91a1858;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he287e8fc5d67263b984589aaab9e88fa6cca93822f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h179b009b3004c41ad922b56743c79f655c776ca837;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1337641734dc4144eef69622289079793e944438f63;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h23c4d9a024f704506017a78c66f5ffbd7242fb8fb5;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1ba5abb2e6c1c752a674637e5abf5b22016807653b8;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h104f41aa030ac656acb75b4439f61334e15fa6e3959;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h100c35af818ee713e518346d37f72ab4af3e0cd64cf;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hd58b4d3b4e05857359fd57505546582e98dc09d228;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1d9f387aaee810f708900792d2858a34470ced0269e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h51b1ad196d6a2dd00f3092f2fccbb7eda017b4cc83;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h2a5c30e92e45c1edde349df7dd5013b31bce6065c9;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1e0931a5fb24858a0b9ca2317c83e5f69510af95034;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h86c69887833f61fbf8f2b5bc543d93aee75c29975b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1ad4717ab78684038f70fc9e4da4d64edc7cd2ddb78;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hbb641b43c80c8b501f77c3276432bfce39180242f4;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h166054ba4b8726a655c552f28e5a8222eb580e1661f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h10c173c384c18d7270093ccd460ee74e2df24065a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1b4cf9dffd3496a35a4c04daa35a761cd29c7dd56c9;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h13b922ea5113d3c1b4e8d0c91d68eaa3db1e76997f1;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h17e06a63d3428357530adbb87b3b7cde8f6f65e8846;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hee51e67e620424b97a9459ccc10328436089fd9360;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h9f331752effd01c6498648cf8ff8425722bf37e447;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h18ce7cff7b0de252db401d525d423ff82be90154aee;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1711d048d25f620e4d9f96af3cd0e2cf47ac65967ea;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h194cde1d971ac34817c6a194ce489e607d7a7422eaa;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h34292c3463ddcee681f5cf8663117d14664095ecab;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h106defb62ef6a49e8a98256b9eb17497384efe12e71;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h10ba873eb0a4816c9b123c7c3bc7f2c9b1185a61d0f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h187f270deb86fe73234776e80ffd0ebe7145c36dbe4;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h80d69a47ad7ff0e3c3a14273cc9f3f9a6fc19a3185;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h5ec023a22aa25fcd96eb39922e8e5e848a2f75002e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h39903835df9904e1152afa24606d2f299a94d4660b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h2bd65391d88c06f76437fcc3876742fc7a4d7a626e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h5e9211ea5db4a49fea8853c51963927da403fcd090;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h181ffd2b85f6e49f6d82df98ab3d4744ca46eb3b835;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hfc989a8805ba38f633f6a75a3fed4a6b43d8f51e1;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1dd568a77bee637386419964f198cfe548d57416947;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1a55920435fc968be694ebd78ae63e88466617ab316;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1e3d992568b4eba0a56fb31d1b7778c626ce48f8ab3;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1873ceca1dea01d49d56dea0d70919e615e8c7306ff;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1e3f4b408a919c57e2c3e45e1fa1b7b3e323ec4ca79;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h15e91f537f3c22f64411ebb7d1dce41bd2e2b5416d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h14d7bd8af210de5d78d56f754175b8a43cb496bf662;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h7e6788630750d0fe7bfa3210cb40ede6acafc43cb2;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hbe2fa844cf4acb30e8ab5fca0a24ca705e0bf491f1;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he1c04ecda0b4a71aef2005715cd316309b1b956708;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h828f15154fb02ee778defa19a49a23de02d4a1ce5;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h13f66026547a09029d7dccd68aae265ce99e37ee1de;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'ha18812f501e2748857c925609cd2dcc1ed99b0c363;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h10d52cf6c6d573bb9f9b6c42d034fd1fdc296086dc8;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h13f82145a7a4102dc6fbc06b7582f63f8df94532572;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h9fe110b185db1c295e70187aa4c8037c81b2ac44ea;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h15426f3de16ad1bffbc65ecd0f5a8d1ac7070c57691;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h4ed7f8fae95ec91291e45e67d52b15598e6b07cfcf;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h82c6a61c337d2facb41e6487b8dbed100dec45c1c6;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h90340ebc9b08aa3af8db0c2488e54ed327838f0a56;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h192b0051adade483821018bbbac189d068e59de5fdb;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h9e34f1a91dd8f3418fa6f37d24dbfc0cf4ecb1c33b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h17fe6cd064f1998fc7201512fcddb588e5e65ad35d2;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h221a4fd69de7412f842a99b09e2a32de19699fed75;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1aab5722d4cef18788acb5d753623399b7c3718cd4a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1c6edda9c50ab81eeeeed1887a1b7fe7002984c1b6a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h127eb88aa6dbf24e180c26f8e864ee1e01a2938ff5a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1e589eb228d1095790575d1dd4ae92b93d0e6e0be25;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h5989c25b10a321c67e2811fa93354080d02cab556;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h446e7b55b194b7b9a56444686d2afbe010fd9a92c0;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1375f67824a9120549dec27c59ee146c7d4dd66826a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1bb69ac9c5b873b1f2ab90e777faac28eef25bc2166;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he3858d73a90a5c26f526ce3e0466a8c35cfae0cfcc;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h17d96d8e2c0ce4f1e683b872d849d47a412e8ef1986;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h113ba1f244e513d6bf7caa042d33dd3332b247d25c8;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h7839ec6067bb5ba4d61b8035cebf03f50a6a10d69e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1603f6f7463ee7e8c0d585467f3c25592a4313879be;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h4c16085cc31e0a43ed31cf99dc38de4fc1f037851d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he4fd587ccec90c4688828ba9667581653564411c12;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'haeedd192e0946d5ac423bfe2e3e7c13ddc1d896ed4;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'ha0679057c6e9a7c8369e2c48c1fef0255942fe8c0a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h110b70ce49bb918b65bc37a434288d3fff51167b3de;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hd946a6be2aacaba18c26bf6bcd1e4e03e0a84b8e2a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1ad1d8b12cf178b26ec7de0633af06a9156313c7a55;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hc62aea99ac7abe7c32455f9a9dede58fce4ef631c1;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h14581240ba57483c3d85358824771994ab8505ffc47;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h537ab6cb3137c4d9aac6047991b5d011d057864786;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'ha6906d2df874ab540658ee204f6929dc26fb2fdf9f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1195494f3bbe8ff82110b0b469fd69e4ef64b1da59a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h822a766e04ce82bc1e2e3005c480cabd3e5161c838;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h3eda9d0263b3bd228d79e30cb0c9d3f265c79b6638;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h10a9879e1df1e525143f1f388bb41b7f94c210922e5;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h86fd1b61a8020864712b45f421caff2e6d68fc3a53;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hacb88fd36ecd272d9496fa3fe9c082a19bc27632eb;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h84dd3c861d49cf258638f3ce4b9c754ccdaf48841e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h18a8368f926323a62072f6f764dd681a6bbca4ce67c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1005a6dca728eb3bf08d0ef61ec2781d661e4a34a8e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h18c5587c2c280d327bc5b6ea8c2042300e5d7ab4a7;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hfad5e3620f8278c01660cd8a52d5307909f1b7ff7a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h184ec7baedecf5983768b12fd5c2838bd99d498ff33;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1b72dddd5fbc6250cf68463dadac0302604be8c5841;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1c091dfdd90144e95eb3caa9c099c6a54ebfc85abe6;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h833044c7be9c5af17e87c9003bf549b70cdcac0a23;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h494c4d687e71149c6ab4779a8eb6d3d878203443ac;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h87f370f2f047963252a07b8da0e73c1927d9b6690b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h4079efd48906384707fdefb526a5e953e22750673e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h315aa34741541f5d6b52180948c1ed28db59d97743;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h6466f6ea60d705356c48f2074f81d732dd1081645c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h11f2fecf43864e0b895fc09567af3071a7ee0f9e446;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h244f7464dd43031a22578f3b1137f8ee94641344ba;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h13cafec1a4d35b844cffbc27f8d75fa8aaac8227c95;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1730164b7dc7f29d7191497ce40a3f2106421af29a8;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he03d5784d900d257cb94c8e4c7ce597d3caadc9051;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h10f56c08216a174b8f8eeac3c76045f359e8b6b88a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1a13e67d041ed38eed9b3ea00ced3e85d6185e76f5b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1cf2b829a77cdc0aa057de3fdf74081545be22033e8;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h140a425206a56bf6f14e2f0d24bfaf60342b326b07d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1401c0b24360f332b2f6ea592cfdc05711602cc57da;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h8a18c579ae2325cfcbab5e62c3fee69e67a6cdb1c7;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1df2ef766b4e4b9f44ca67f15622ccc75914131c1c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hddaa1a11abcf336e45b5f30f7c91d34f56c2011976;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hdb484a911923c8dfeb2ebab8ac9d874295efc78d06;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h198940cbdf7ac7646652fb70d722db621e7e3dc4f26;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h8d57c0a50594cb5acaadf7941b6d34edad0ac50a25;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h4999b14bff8f0b5dce36831c81ea517f54cf3babe;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he038bb8bee5c2f36063ca8313a6452cb74d7579d42;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h4a3ec74f7180ae8b1aceb66267d4cb9a90f7be317d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h9f57b542ac4ebb7d04a4c4e68f5fa320f3156d31f0;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1d96ed6bba84e21917ee495616c533528c2378f99c6;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h188f4330bfd6fa01d52b27c46a9662c2a8c068e2ca1;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h56aba7cd5b928018f5c4ec409101a347b17d913e7d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h273811a20bf9a6f96aec842d040c0a4a4d3ac45fab;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h17ff61eb8e5b6ebc54e84525cbbcc28125bb6dab8b0;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h8d178658fe9a2ac0a766bab8c54dac176f11eea76e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1499508b9a3ef55f9bcb684e4d9f9f6b61605d1425;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hd2c20bb20c0c796ebdf795b11aead2a13d3aa94f92;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hc23abc7d89dd579bb8826a86bf47d0610cd9c185d7;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h6e764045f46142d7b17d94a657ca50357f221883da;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h242abb7959e752ddf9e11e7fb3c4b8694a11c49fed;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1bc48acbc6f5eb7e1c395c04cdd34af0a3b2e0e63db;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1cda2c6adace6175889f35599c899652fd2b846ecad;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1c84d9e5ff54e9760510ee5c5e655b5011faa17822c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h276d3f7835106685ff2b2a2b6a710a518dd34c4d04;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'haed11d603bbe5def0392027413ff6168d9b9d55ebc;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h3828d45d746957ae73181295731117503a08e4ed98;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h17a31551af4a1f57f3470e58d524d04e9d2b9e37db9;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hb343ab616a443fe6cffd0bb0b3e5569ab416da1abb;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hd9e94be672ead049db9c465d61af8e4033e8b09851;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h16595ba4e2d06ea3ffee862e2081c90a09d32c48c98;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h16e5eea72c376a00d20c408d384b62b4756bba95507;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h10556860d7c6e3425f476e05a09319fd526da58be7c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h8d096db38cd44d272aa8d64c37fdef0d2df4ffea5e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1fe6b187122d648544897c84632e628b7ee078eb8fe;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h179100c33b0859f72055ecdab0f142ef8c3ddc50fa3;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1860688ddaf61b4009bdb59e8ab5e02094736daedd9;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h19db2bcb47db0cb48b298dbef7db8d2db39c4c9982c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hc0704ccad32b088ba7395134e5234d5c8b51c18dff;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hb2891b7324c905e64f3126ac6428165ea2807a4f7b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hd111f073d43715340c8be6e8d49e81bc01c5dd1bef;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h688c4d43a8bc1b83b71833a20a1bcabba0d6da957c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h3d1dc28cb321a65107f6e7a49d144237e15e4137e7;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hb15cd8acae2072b416f7e3e32d5f14c05583c57422;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1e254b3cb70edd021be4e174310c1ad86d2168c1a68;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h7e4dffaf0f251061a68701f63849c15c9728348de4;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1bcd1119ab6091de89779c32ded14c2fce05398ad4a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h2480dca621f106777181b02d1bb71ead8bbbb7f266;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1e6b5c95f21cc7bb4b9fe376c0d9e5a5fec4741c2dd;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h59f6ee127dc56113a8e3af3e04d76482772205237;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hedbbd07b1f7315408a6ba8a95c8b4f3cb955415180;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h555c9beb59352dde0fb60f2fc0477c78110aa4d9a5;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h5ad8987e2efd1acf6a64b0f6079c27c66de4764464;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h16f25cb49c0b2ed0acc1680fe15b7818f20e0d05739;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1af67a5a4a324e84ddc7612d3970b4a2eaeb996b1fe;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1bf37abe046a28af4f4ed090d595ffbbc3b8d2a6506;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h8947a5d2aa0131b26da408bd803e9597e51a0dce46;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hdbca8215bb2195305566d4e55679db680bf5d4d537;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h13e13dd104012c7a3622f7e6165ade11ae8e90ead93;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h9ad6543b0b5cf181471b7cfd8a456107058048ff1b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hbaa8b3f88995c0c535871ce58968e685dc67ae7cb4;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h144c8e9aefdd6891ff7ea91dacf8ea690c14d004f4;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h143fd57d3cedd6c38a352108407275a329aea9ba454;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h2c49d7697da953fdb22da2d4ef5010b567302fa1f8;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'ha255e270cb6c68ae0c499e6e8b342772b26b981340;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1593827c44497f53a8e3cab110679cd0cd212909787;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1bfe12c44a2f27413cb71e62da9bc5e624a3fb2a5ca;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h58dc0b799b9c378181bbfd7cd7f5e1ed82be2b1038;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1537bbfc4489d52bc28f653295525d1341f4329e49e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h2f6d83a035076a9403656ccf6309c49ea05f9b2aee;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'ha4b589833e2aa8c3e77a1ef2735c34d01eb3a3cb5a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1728e1297ad0b689dd6b8db5efbe264cd3ab01814d2;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h10a8a40dc49c5e217f38cae99d39c11af1bf8504963;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h4a0ecbee24a6604c4f1a2199ebe16b82dc9f714b5f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h117f7f2e78e607bfc93caa3710f23972ba9574d4996;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h121bbbcb35bd39ecd6d352593e9bccce8108100b3be;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hd0b60689b0d914f9e85bad5a8409c996251e58fe45;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h673faeb1e6c7801116d256851289d37e5cd9caab;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1e8af6a448d40a023006cc57eeddb3959cef999e2e3;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h18b5a162b79faae5395195713087ee3fc59f6092cf9;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h8c49511f5172e8d33f5501908b99f9e6e771074ca1;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1ef420096754143950469a65afa35abc836357340bb;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h30a3cd060dda3f03fb6e7aab692389cc4b2cc4896a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1d525e9296876fa7800bbb02e3dd97745a0b623c501;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hc1aaacd77973d170fdd6a0d53c57a9e5ed3ba30560;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hacbba2041c76d4b9c7e589207f5d5ea79a79d14a60;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1335f6e44012dd3ed079d88be86d088e6a7d96aa958;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h620867b0e5a7fe24c5441c3ec8f110b093e39d260;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1ccc298ab1c4976c7882a73980eaaebefc17e4fe091;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1fd984ded50185a166058a48c233896b8ac152c43e9;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h185cc8940e6badc6b67eff507864621792b9a843e26;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1b8b3070c4ca6f89441794b50dcb2233d67548fe64f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h6ef519c9544d1adf8609a50f25e0c309d115a4eb0c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1d864e07a9910b1a7e29d25ac20cf59393db2aac6fd;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1cbd7d610f67e963b0018b392be15f02faea303827e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h4a389fd28df4962082949bab76f6940ed970918531;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h134513aa32616862265d52ae464d98606f85605ddf6;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h19677326fb65979e23e2c8afdf9f5dd705402c7cdbb;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hc641c5dcf1983aee6d0ece5326946a45a142a94ea3;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hfa939323b40cb0e40732e51c94807515fcfe871b86;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h6823fd2274dca77275271a17b272364defc04a0d77;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h186f207e27d8c3960bedec24c1a8845ffca536ae98d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hc6590eac24d1b062880d39a796199cc7ba745d54fa;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h924a60ce3f634d4f4060a7da398261bb173ea569f0;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1dd822ca3c6b8d0d9888a328543219eee412c72849e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1590cf0f42ed751db7c714aed6f4249d448ff1db2d4;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'heeb5576aab7f63c46113e8d19e6db31d2424f41042;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h103229f36b95f34854d09fac1f516ea44c86b1190f0;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1f757df3af9b88bffe21a8f06228ccd79f9bb49c00f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h12c5011fa3ee5befce22771e263d468998533b67a7c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1a35dddc97ea7db2a62f81e053adcabe7c59b66a956;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h17786311e462f78b3bd29f3e7833db9ad0e9b85ee9;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h46ffc74c4db54d26bfef3a5768d59fb45cdb32b1f1;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h5b631d2caf22b6b1f0e289323a1403eebe67b76b36;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h3070add603704759f46d9992176e6282377aa06297;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h19aab40a6052e197fd19d1a77f6a5e4c003b6d61345;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h3684d614e3b79cc2c1fc376c03d5d401b6d468dbfd;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h9120ef421e252e5bbfd12e7ce50d88eeee190ccad2;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h16ad992835fdec85fea199e4c7b3bf055cd0d39a13c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h15ef73bd90525ef9729af8d340e77eb4479480a949d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h9d2b000195ced2e5feee3879f63e2b7a9002065e6a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hc1d01f9a4b59981a2bb70b6f98cb77ba956b54c22b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h393037ac4918f5e3faae149d8bd939fa08aec5fa2d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h11af1442ac5bd97db1a95b837269cdc60fd525d06d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hbb656cdba34aaf4a9d02bd62a291fb5a9bc475aa55;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h152a7081f2da17b381c4d5ab6ec5f0c848b66e9e478;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hb259c8d031d44ae71eee5adad0e482b7b7002fe407;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1ca4cdebd480573fa59e02bc5474aebf4c54b0d73de;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h3af433ad41723e8e8711048aabc13172de830bee25;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hc0ac5ee919ef1d6f35b196b93e4c3948f807076b41;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hcc5d8c68fc72eede109892ac209c1f1d39a3a1960c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1e8c940b5526facb77d0f3964591e4dcff28dad66b9;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h24409c9c46412f8ca4ccd5e5941a114153c06ef221;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h7f4d592e1c2010f2b39eb13320caec63524070b97a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hd0207014531f6fcace2a8921aa1ae64221457dc9d2;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h157dfe7056128ff9919e6502ab411e5a8a3ad0718d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hd97fe27e387e1dc2bf9f81930897e89389571c916d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h101bb3f2f146270ad45591e8b3b8df6ef2f97e47c0e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hea292c852431b41b25332391c520f97562a1d5adfb;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1dca6f38f11aa4f09d501685c9d33608abcb5b1ef00;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1747dfe313dbb09474265c569f49208c895f0948e73;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1e565f588a8bc9db9241a5d8d371be7436611e281c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h126251be52850525b480cd09a87fdf49f1c00845b23;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h9e19b74c5cbd3b565aee30f6d44c226af0c93ab3f4;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1de63d80d7b4a81ddd35a3cd11753593f9455d5f0cd;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1a07c6b6285e02152d59bbcfa03f037b43ed9aaf61a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h4d83c550c89c61c8cba9c633ab3efdc9aefcbaa2b2;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1c1eb450ed6b25a97f115fd3d1a8bdd7cce932b085c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'ha2a3053ac0537d292512334c0afd48e9e8891c8dad;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h194f391fd9448941d5741961c5861edbb1e2b3dac4d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hdb818407a5a6297dbdcd563093f7f1ef39760b7;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h15186e8ead2b4a855474af4bf390f164b31215a1ac8;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h30b7153caadef33778eabdb417f7d70d3ff6c89e2;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1039805b32f5cf0759148c1a8783be96b4a937b962c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h17edc8690c48876841663adade360452181dcfcb302;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he726cf37270bc471ff7a2fe825b3a4314d25631adc;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h15730f3fcc0a4bbdcdba8e4f92350516c9dbcc31e6;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'ha6b4a434f65d71c8f82b571e90004c7b94b6a772df;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1fa12669f235213d9b10160bd06088bc685aa17d961;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1cff3b4f1b76b2a123fcccfc951b694431c1ab74775;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hccaf3234b63c1bdc2bea81d2fd16852b8093b8c375;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h10ca337885157f8689a17336233b74bf895f9c5caaa;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1af94b5b7fd7534bdfb2e965d85fdeef9263836286a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h5a6c99df1cd60a23c403e017f2dc5974d1e12ec234;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1fe93b3624ac8ea4a1b6228007ec9da1b96fe67020e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h18b4f522e7a9cf1b9d3b0317ca7d446e79a3a860e4d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1fa60f858a6654225d85facd4dc3a1ad82c85d257fb;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1e2f51976a7ab906f26dd2c736dc246548527cd84d7;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1e5af535d52c6219c6d474899a126e724766a9a00c7;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h14c7363cee139aa4f412ca36c70628581368eccdd34;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1403152d31625a77f53f7827f61ab0e65cc3b88ffc3;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h6534d061bdcdfa73202cbae139a0fccd72c4aba553;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h7c92d1b18aa2bc0c27f57749ac4b02fb9dcefdafa;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h18ae04f4805abab6a01eea4dc4f5433c1a3c3dcde9e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1b6542a20dbf588e94b6a0d6a2705e2b06c59acf513;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hb84e2853013461d52bb47fcb6b57375596f05871c4;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h95ad961625f2f53b93f10ade1eec44280b9ae7e97b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1018c92a72b5da6a91028961bfb28ee7316469a697;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hfdb5bfec18069ab70155a20c96723ca8d2429d32b8;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1a27f61e586f288e2fafba79bae73eaae20dbf53a36;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h61037988b4bff2df875b75f8352d9f17302fff574a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h74894c121d07cebdaa708315233a43feae19a8b871;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h841488d8dec04fa2a10fb157551a3f464c76919f23;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h561a370461fc0ff0af3a23daec8f5e30f866a079c7;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hd29add958a179da91ff19253cd21cffaf008889e74;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h15212197e5cbbf0df6aa1bf981b94040a617e8ced5;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h7df3c4799aa1117c5a67a8b75a2a1b0ed9e5f6ed79;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hac58a4b7e7fa1ecad0381d024e1d92cca4e4d693de;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'heeeb39df4b5fe2504ef08e3ace44d047566afd9161;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h11690ca7d85c10c908d69a8c444eca145505b74322b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1e5c7102a815807958bb1bff07673c5157240b9ce76;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1e4f4a127de83971872a82d3da369727dc9bd52b08f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'ha1c7dec529d61e265f5259d33e5f1b6defb89adcca;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h2cdb3efcf97df622102b91ba04f9f40a05f54108a2;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h8c5fc69341fc2ce138511dd792e7fef06a88cddf99;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hf6a59e5ed9d335e4d039d66d25aa4d57b19208e4f6;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h183ec284207eb209cf4f11bdf37e7595e65cfc635e4;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h18d3381e82f2b7651e7329cc306edef62b5f1ee1480;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h6747b6dabc2bf5334c375eb09d98226c456e50badd;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h717ccaf07d715c90bbad41029f3c562798d5ab9d23;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h17314be87e5c746bda9be66da4eb9616cfa0dea7209;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h561c4b61920d24e0ed3de0075522e15e7c52a03d83;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h18236acdd6616e1cbd520053f365f7f229c20fc6d63;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h135193e9429d62c53b317c25a5ecba76a2b3f339b53;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h489c87910d3043d1d75896dc954b9e25f6d47d95fb;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hf0a4a7b2edfca1e5888eda6e271fe214f2cb71927c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he805786adc3af74b2bdf1ba9bf719c1a641aea6435;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1811b38d6ed6a2ea7fbadc6d514860af6dc26e4bec0;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h53e8f8cbb9ee1fea575f537b2aca0d7cba32a39b45;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h5f5d8486c2d300b527c2d9dcfef761506605f93f92;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h5da8e1c42831e48fd38b9379234d017b3f2ad99c07;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h4a854c2f2ac316c2c98e389964c5ca8f68f9debf46;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1b11a63bf058fde1b1a48738576f4237255248dfd85;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1d89ba4c6e29314eb123fc53508fe1e6334ce23dd5f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1f83cd5dd6af237c36ebc9224d9346360f692cd2249;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1a5c7eda3adc9729a89e02c50965d5a5fee7867f5c7;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h14fd882db21692fa76b72f82b1617bfad9fa4e4e3cb;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h2cc45f579b5efd74d40f334783d81173cf86381b74;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h55bc593154a2860d6d0831211efb791dd8f6e0529f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hba21edf0f21aa901eb0984f054831546cef67ed6e3;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hdac491b1bed8ad17330cf711e6cdc10332aeb6b3b1;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1f011768bc55864107fbb0c9ed7ff4436ba8bfb8ee0;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hdc1709516978ab0d12820f187bcc445c172fcb4022;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h773b91bad01df61f74adcafdf1bc23776fcff1b679;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1f4aed715b11fff1afd8448dec29be7b480d08ea0ce;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h6113cf614a53aec5ce09ad31bcbf86a37d7bc0e46;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1fc059f1015cedf2ce218f02840cd80b4434c1d68f5;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'ha7500a4d0184b00b7baa9c011beea2f89af08a701;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1329238f1ce93f48018b0ae4116f1a350f979a64b24;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h7b3690642d7ae38516bcd0feeaa97646b57b1e1801;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h93f1b0f6820392ade40bcbcfb2783f54eccea4c008;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'ha149524f00c87295c42d0f3e4725e832062e66ae6b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1f833c143acf449823dbd6c69969fe30f1d0ace8449;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h42a299f5acbde89e5c30c19847a1ccff4838a92230;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h433c22eb787500bc71fb404d5115a503c3a99544;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h724d15ed2cfac9c04d8cdc7bce32149d3115581d87;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hd374f8f2cad6a20e9c579dce30e93b4d9296f2fc7;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hee4901ffcbcd0a99defe56f025e0d5b1fa88d92df8;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h6f98dd54d364faf6f5b74be136146913c25520df9;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h341e79434cb9c7911eec462fced39076cd6bcea19c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h8c4670a97fc88cd50a63bf458c62e13a76dcebbec4;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1d71b2a382e317eb3405edee65061749a02cb6476f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h129e6b4e1535111bcd90459f3d3add1b24aaed9b56e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1cb504ac1dce0aaa305a82a7b3a927d235c43c0b1e5;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'haa40f2410772ab707d28b9cbb0601a545a54dcf9e4;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h8b183dc27dd68563f750d4a8d7f546e08d8adfb837;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h12d824fc06f8c1393e22a5938c30992b5ed6fe29842;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hd8a4fce561b88f1a6c8656e425886eab745e395136;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hfd69d994f6d34812ddf4ce6793d4d9f61eea8c60a1;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h19be45fae103a00302dcf85e3dab30a426c504fcb06;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h14393475ff16c923ec7ec0e43a515cae01e6f353448;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h165560d6c6a1ef373467672cfba1f883a9d07b3ccab;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h46a58a91d97e23165d0e9536afcdcc2b01dfc61f91;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h9e42abdfd6884f83e5fa0edd1bb3b28379e752bb99;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1d1bd9e6c7890c40ae72bb123e9799a478b0d691ad1;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1363ae17564b2093e7f5860a210929fd6b26270e7e8;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hf6e7ee2dd695426847f0044f073a61efffa3d33c73;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h17e31765a4f1beb346eff3a69a0ed05b0f8250947ea;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1cf0d97261bfd15d28dd6fd1cb43b1502d140b004f4;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h125e2cec6c3c49a5bd32f7653d78f7a37e552259cc6;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1841cd4b46588c314c410ae2eec8e1eb203ad3195d4;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1eda97b19d0f3f1ee76f2e67d244ff651f22a1eabb9;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1a4c1b8fcd86fc9f294a7a4c57f4cc12d38d0b22365;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1291caa0d7ed163d210c596f3305c2e1024e6ea018f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1fb348a11fd2eb18c1da21019315cd0b5daf9b52b69;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hff7ca64f84cd3e7d2f393a66461aaad4dbcac8d632;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1edd80e92d40b4731a95594923a9b7e445414e7ec20;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h74ad25ba11168268ef0156d4881dc542852bc46139;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1fd7948f29b28c43c14f69151f8ddcdaaaecd6a2519;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h14b462ed533eb53b78d3be5d3fe4ac3fbb2a8f07115;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1f43f1b39abd464b62a5f419e282ffecce58559d3a1;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h69d110410d62c19aed24483c7ca5536496680eabe7;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1cabe0613a179cc1333a41823d980f7541d956bc217;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h14818f8e7f436e0636269f077b356af6d11e4a49e49;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h8dd50749f22a4575c2e76b7f0a443ef18c16d2f4a6;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h56365b4550a2652b4ddbf1d8ba8b91f546dd422e1a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h8f1a225d77b0d8ad1e5d95d4b050116ba11c9fef35;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h6c56b82e5e59ab62e6c0725a96c53995a08a7503dd;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hcdd27946bd52994e10ae8cc70a18265eb8fee4423d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hd410c38c31d4c22b8fa4ae78eb127577c1ad79bbe6;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hef36e31332e2c3fde9607ad77c8693130772ac09ff;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hc937d090ff51c741501922bfeaf9334593f6951171;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h167a16fa17fb6ce1a11b212af4643326044bff4739;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h19a83672bb2f2352adab4739b8fd0f04bacc3b6870b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h5879b1e72517573358b003002cfbeba880e9690bd;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1a227b565b763097951188f655b85f26c340949512e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1d9e13f8af9ee45fed1de9a97d9fb0769c9d2a27917;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hde3934a9f56aef73a3af79bdd8f0ac20ef810fb24b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hfd2f51b335fe356d46d2b26e428a8bc1ed19237698;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1fdae83adc0777aae528b7d014dda5031dfdd3d3611;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h18f9bf615e792cbf83ebe141dca5422408c52bdbc06;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1e0a055c1e2d21de0d004f5c56e1a8f597c08fcfa18;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h152e34f241101ad58561d8ffa0fcaed8874693b7cca;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he147c00952aca8f3c8db32b09ead8e664e577f1b48;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h70e049898c157e7592cb43c019a319a152e73abcc8;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h22229b4a054825e5899e3e81c5604bcdbb5c63fdae;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h4a5a8cc4dc074c190c2be65b3b70287fad879b4a80;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h5485c669f3f7b22bc02dac97c1e0add9111ef23620;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1fcdf162b75105b26251554f6038687bc2ee7c3b994;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1601cca042009709aa15bc8dfff797da77bd1f4d0f3;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1d65db2594ca97b2e5090ae6dfebbe853fd8ef63828;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hbb35c68ec8b477b2d82235ffa456ed1784df287551;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hee5cab98ad088d4b7cacf21e54e1c63aefff426ed8;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h16e4caf2c66a41bbfaf420c9f2ca6f44896463d68db;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1bda44c4a29d298d9d80304ccc282911969fa16bfeb;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1cbd4544494f91b510bd0c53180dc88b42dc7e67415;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h2700bba5636e5e57592fc859d43d4fd850e6e403e4;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1028e8a0af15a2eddad04c58c832860405b63e6f172;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h2042fa04b8ddd031d06625a679f406ae8599803aaa;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h762765e217c2ebc03c81cc2fad0e3a4a9e92d1fc12;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h8453c31f932864e63a355368d50d999ae01c5c0226;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h2e80be5acf0f0b09f36b05149333da3e55202d7208;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hf5580fd713450018385aba4c1d03abf56bd8297ca7;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h4f23d862e424b915b764108e4304c30568d9193d16;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h16990e3b97461f611e742a16a69fc233d69f83cb71e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h18afe4b6aa9c940394786840641259554744154bbb4;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'ha423ceb3ec393fa771d920710a7fc7f2c76f6c3df2;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h184e32e1b9109768f4f1222cc7ac8863feef459f20d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hea4b7a275091dbf157aca6c310435fbe8f142ea154;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h5128a7a2bcd3d0184748b014a26cea36d65f0b74d1;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h9e4ada98e5a48e52ac297aeb7d9f868b941254579c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h129112ad68987399073f4a309657a061e47014b8dc9;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h11cc06297dd0b8378ac59e9fa2e0a493b29e361f6b0;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h17881e24fa73ab7c435f952381eef1041fc2d04b428;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1a983eaac3a97898fdfed1ec3049a84ba7e773247b8;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1c1dd7d856ba7cf1d6f4275dc888b03dbbb4d75310f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'heb2c312563a9ce3229f6a8f41305ad0170ffd04c50;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h12f2d5b5acff112131762463a94eee351f1b8e239c1;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h4a45aa706bc28f094d3fbb83ce8adb745e276b1934;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h5b91723f0edc1ed7487c4fc7afe368597b8d0ef5fd;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hd01e6f2712d29b490497fc7d5905b91a6289703834;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1f3ea6980965c945a64dfa2de7f9fd4ccdd43c2320;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1ac1d3c32d70b7b876a1cd275358c51fdc9654804e5;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h3326dace7f59468f95e346426b0d93f222bc9035b0;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1d0bb3aa767c1716749123ebbec891992990422db31;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1907f932223288ea13dea0fad9ef5ee0827faa9adee;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h181b7e815c95212160e19d9ee2d7a207b0e7d763c80;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1d78226c7f505c738584085e8812470f274f9e6dafa;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1c7998456ef6ce65cc600c1bf94e73909216a7875ae;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hd38e0c1128b55f56afcbc589ee39b5ecc9a629062a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1de30bbe80c527f9ddb9f23254a401d2b9906835d09;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1e185dc866018b3be700deb7e105efed7ae961a83aa;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1b287f33c1863ef06f07ca92fd6c223ae2eb0b67cc9;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1d7271f4e340e9ed5e68320b3080048a49a0f9b489f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h12337d32ebadbc13570c64fd5211d7aaf639fc1722b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he2bff5247077ba34e924d0eae0cc5cd4ed62452b51;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he045d41a3f3e886b5f4d3169b3b44f8254d3a453c1;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1c6f38e66199ac977090704983ac3063ac1a9f79f4c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1afc9879b29eba4ebd8aa0efb3bc993eafe205a198b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hab184d57491452aab956bd5e1c3b575d4fab86184;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1b9f06373767543094347a8101fdf73386ed7535b08;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1aeb012a50dfeeb23f0a64f3b4f9657842fe32f1c0e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h9ba39c3a2e32f9fdbfacc3548412703aef4b93b5f5;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1c19a2046dec6f2af322a35377e2e76c633c47589a9;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h19296f56e16eaae694437407844b9b934d2a1b2d830;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h5903b44aedb1091462c87c02deaba2b91e5a903e0f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h13d8bc4fe171ff68ac8671aa1cc32c181c23aaecd36;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h102b47dc4258d433a97ad164fe021eec31748f0cbdb;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1f75e7d239bc170da898d4b095fc9b813e612a2bfc7;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'ha96f00c3fc983bfced3c7089668b500a4afb0faad3;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1ea877e17160767c62bd7224b229602c3a7cd0ca9c7;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'ha868a8b877ace0226943cf6bdffb5a5a8e83e8716c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1dc5701f1d140cb5f1a206bcf451165ba38e984d9e6;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h11218401918570b746f7a0155e8a6ae716c1a457406;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h2246b8b4424af76b60306a9e1448e7ccaba9fb17e4;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h18bee3bea5dbb713801f722324a102e30ed8854335c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1b2b26c60e09f772cabfb06b6d91ac9c5c9eeed3ec5;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h178b0656a74b530f669d1bbe67b7e81a85893ce5588;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h31e0649bc74379c66dc9e165680a7b9cc8647f071b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h150fca4a1d1199e6fd9bf83441c44e1c519f5dfc9e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1666efdcf636d41452a88f757c016a390a206fcda9f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h166b687546f95532a50727e8883e83dc0b716f4c9bd;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1ab6a1a11fece107071975bb84357282e7c1499d0cd;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h4008c131c9f432f20053dcc9e304e15231649ec3c0;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h231fcc2e7229d81352a00fc34762f5a2cb742eec7e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1619d38cc33c74092848957d4feeb8a025a19eec79e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h726c4244ac55271a9ef1f69ff111bb613e6612e107;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1fafdb448df034a829fbd26eff69d2e391e61fedcce;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h229548fdcb0bd1c23c4c667cb0229f26327c101c35;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h35db53cbc03b4d75c15dc63d8d3b90f2b508fa4f4f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hca44575480de77773b4cf5ef3ee6aa3e529017bc9a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1648cf502bd0a6980f2a7c315d4b09a46f39a6a048d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h2ef0ffdef92fd5f00aa2c621bf7d06590f323ab718;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1a3c16cdefd2b30a4386a2320d8df50bc4ce75b3d4d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h444322d69090435f6dc664917c4f4591c1610606e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h10675a91f1c41f7f21772b151ed1f190c399a71f1f0;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h37ca6153ce8902f7f0566c1b20ea90291855538555;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h141f06727e3d1df45646664e4b671d71858407da10c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hd6d280baf112ca3cff2c659c14847f3a777f5ff8d7;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hb5026f5de53bc0f299eabec8c824dbb5836c5ced23;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h249e0eb7eab0a283b6d8077204844e580e77a660d2;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h107de74c62eb6a1b51aa71447ced7966cf46037fff2;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hfa1970933c3605bcea379f61e064207dd163414190;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h78637ec73330fdf348c0235472c4388f81241cdbb9;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h82928d7c43c2aa08be784e1382060d87c10bb9b583;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h19c6b31b9dd9d95368954dc23c168a1980b34f3cdcb;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h19dfb2540207950f1c8f191addd9b00ca1ba769997d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1ec499cffd007024dc965111c04aae5211832b157f0;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h16e271c4c506ef4f3ed84d2e5b6793d189248d441b4;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h208030854ca4620998f00b66cb56640679b1d05ac7;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'haf787fc08c9627315750ad29163e42d3f38cc1abe1;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h18f0ac8c1873ddfc5158c871370f3b1bad2f8a709ec;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1200ed17204f2cdf3bd00eaec75d0147fc9cff5451c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'ha5b197a6976c70cd264812ed7ab952e088d0f64d03;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hc50a80b85e0acf11868867be5a4817816d81a03950;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h13ba854a53f8e1ba7b6585f96fcec2d703128d35ddf;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1fde42efbf4b6a22d5162d096dfe254b9d3d1095dca;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hbef4f6406d243a2f176fa43418a47d8f94237466d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h16b296edebdf7ecf89ab4924d30666f592dc3163479;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hd842e7134681b33306c5752b12b536d306edf6554d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1334d78945b716e2332f0ebb0995ba87d69e59114eb;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1363ba0e2f58af167b0ed3de2a012439a3a305ba2f6;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hdde5972eaf410f212ebf6c39d1881c9b43be332bbd;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h187b19ec2df9b7b66fdf076afc364a153df4cc34e00;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h52e879292488e2862239aa3609a07e705651bd6c02;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h17e73204d9497bbfea964021434f57e6393e917d648;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h71ef4652541faf702aa8b962f5e1fe243c58266f1d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h5318ddd828a44699e4d81eca1b92df30f14a9ba415;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h4230d94db3dc0a0fa22b6c170672dc09e369d05a88;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h13efdb740b62943707e589c851afc5a5728fadda752;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h6ed4b13783891ae2226394a51f8611f1c8676627ce;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1e575ec578cd69cb6d697aa38fb97916ee99278e788;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1ec12d4bb771d695f3e77c7257394f4231b37e6c671;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h2d210bf4bf87e74d29f7e626da0df3bfc9111f8904;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1d7fcb7d0670f2e45fe20d7e0b73ca2f2fb89c48db2;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1ae1698ab89be9d16eb69e84bce8a5977fd5e50758;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hec1938ab85aa4c43b5009354aa82b422996cedf9f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h153eae5c962975b8fdd7ef2ff4603beb7266d6f41f7;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1c75338d8040fbf3d2c77fc83da039b74a1a8f23f34;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he534bb17ccbe3bfdbaa94894271a8980a443cbe0d0;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h499afb5198f7fd0a260eab45af6f733ab77938a365;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1e633de35232fd9527d1a92ccc33e812a92747ab250;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1ae57789d3b873bc234ea6992fd73c8b383471bbcec;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h79016fd2712f99cb586b777901be1668441011debf;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1ff032eb47d135711b76127c026f88b778f31924cac;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1868fac4a9850f67e965395ebcd075a28c01bfc9a9;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1dd44fd87f335f0faafd900150bf534486fd813ce54;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h10b40bde13dc448ec2c809624796f3ed0f2fda0274a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hd0f69be1f15cbe79ec51b74b55f36ce3d43de3ef23;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h6450349efaf5d0b533a4036450e7d433b1fe18f68c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h21186ed768c8bcaac45690a215acefe93d62a4a1b2;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h106841f61f3cf9c4ec25f41b07e110db2c81907484e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1f902bd69edd0546caf1bf2f47c6f75c7704bfdb519;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1dcac0befffe696dc0fef9ecd5eb694f7b435f55d6c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h18c717e2985fe53d81ec36e2404706778a50b2ff5a3;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h5dfb2271d36c8cdb7ee4236b99a58a9c597549b265;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hb18b992aaa82e6a10f0dd98f94e4a7afa87611b857;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h2da32fcb78905760e1e4432e3532b456e46ad0c055;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h642b75116d81257e969a9d1f04083b8aa81e32b490;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h6e91512b1ed2f7011144c168200e877f1a147c80c2;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hcc846bdd1c7266b3ce2be630ef767bf6976cec46b2;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h16cf7cd35b7206fb0778542c983186fa7554436963f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h78338559d295b62f225f1af76b5d38c2125554d722;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1c7250323433637af137f65fb2b083d41273ccde4b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h40eabb9557ee9d3fe00b96ff8899b078a50c751c9a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h80564f188ad9890e9c3b2fa277a05df4052763f93;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h4ad78eea84c50ef94a300808337e43ada15dfc039d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'ha46427a607ec4d2f2be0b46f8959e71d2abe5565a8;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h13b1e36cae27e917610351995dc1edd10d7074c0bb0;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h127a9a5600fc3de6c8f9342f9e12e996b14e4ca9841;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h3c8e48b436dbf06c8d1b6b856b0686b9ec6ee5ed69;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h2309827cddc90f881d7e0591d47cc38a21159c56d8;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hd6e66e486bbf04c16a0c9829b21509cd71abe5e965;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h20f44b513175b47d597d4d96dc18849d0f66048ac9;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1f16dfd41c91c8ba356b70e78b6c114c0c5657e3b82;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1755e359dab6c689cc78ec36f2e02555bf852b69130;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h113eab837e864aa340251535170d0fb2f98674ad3e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h106315df4e862cb74b9151283f967e25d4faf75574d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1c24d340d5458542a0b049b0d3d55967b422cf2ff46;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h171659c61ddc3666c15dde69a4345c842b5319b0b34;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h177a61d63d42fe44116d10dd508868103b8d587beb1;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h183c2b3080b3533be69554ca5a195f47505a9af9e68;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'ha26ed93ebe54c39c874b3c50160ff538b1996eba8;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h14f737d0922cd1ac85989aba277770be42b484ca938;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h940a787acf0f9e130e8b45437583ccf1d60e27f9f5;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h34f9b6f9b9364fae09bac0c45b256967c54572f220;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1f6f2b322bbe932ba55cc6a48ac2aca8524bfc0672e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hc73745b7287b486c5cb0483fd0fe3b41e2aa387505;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hc672152290d0f89c7086f9dc29e08a99708fb06e3d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h8a3a2c260fcbdaaebdc6405ddaa3fec5ed65e2cf79;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1546dd3e6458ce2673dc12d07e14e38fb453aa1ca33;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h12d8d636c20ef9015233426a1834f60d8e19bd02f52;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he345d4778481b473b47de4131dbe5c5236e03c52dc;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1b5d5443a09fcd8d95adb67079a4848132fb9f1daa7;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h175f411d6168fa2995f140314101a9469a4ac0d6141;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hb056676491499a1bb12f35856f4c3769b19db98ea0;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1f6ab2e6a307aa6ee26bff560e808f0c03f05a15f89;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h339777230706eecf2717133639d59096791594f281;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h106d61b899d19f657093e3a15ccf3fa9986dd872dba;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hc3ce23a3e1645a0494fb2f52348f35842cd38e15f2;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hc7af290231a50429427c85c33e1d0bd59fba14d88a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h18b6935bafb17eb3d992629d34934b4ff3b089a1fb0;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h75141423ac5e2b919891226419abca6cb3744b9af9;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h190d59cfa63bfa8056c5a48f96d85d15b9a3b046c84;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h4c200a2624ed8fa1ea2da68499a0c37d5f632acd18;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hfff9241f1682ffc98fd1326fd4c98f377c92a8e22c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1ad5b16fde0ce7871fb1bbc14cd21adff46aec1d235;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1c0f67c0da9fff84008b65e36eaa2f30d31a2b9068f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hd5815485f4a2bf0e9d231be6964af585d006f7ea33;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1dab4c3a42d203c965bc95f368d4267936784c041db;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h13fa8dd17f3dc61f8473d7f68e7e3f451bfc7e63368;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hc3630027368959aebe558dd5eea8d63eb6837c78ae;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h12ef12f5943b0d2711d1edf1115d336d623ae4f6c8a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h16143320ba14210092658e42983d649996a4570dac3;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h6899dbaf8f358a26377fb58cef7706f7692cb6c3f4;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1360073aa6e1d2cf141d149ccb996a672c26de6c74b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he4d2f55e84a135d52c3a8ff050308ce6223b09949b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h7d72f3cd2a7108260411275ecbc0d1290d648547bd;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h9d7c7a5469f6663e538f4d83a226cd366a7a52399c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h16e31c0dfb4df381ecf96dfe704af65b35d2b4f8140;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1cf987615fc1bdbf1ed4bd3e7f32c27004b5173148b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1fc59abb8f40186dfaf8cdf3cb14314ff925f21e21c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h102a4f2e85453b3e35851e45ac75aadec61bb3853da;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1e703c03d8ba3dd4f9eb306390886364d465faf5fef;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hafcea666e5829551788b7aa03bd23a9d2323590705;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hd60879851746538cf1ff80d2be0d2eacc286dccb81;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h17a19be3ad7876af43d5c0cc53015c7e041ea906cb1;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he4437032d2508011f7248d06f79081c76d886912d3;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h2400a18120ff80d9b4d531266d06edb954cf920dc8;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h168dcaa7bda3133f968db0bc19bfebc67dfe1a14777;
        #1
        $finish();
    end
endmodule
