module testbench();
    reg [24:0] src0;
    reg [24:0] src1;
    reg [24:0] src2;
    reg [24:0] src3;
    reg [24:0] src4;
    reg [24:0] src5;
    reg [24:0] src6;
    reg [24:0] src7;
    reg [24:0] src8;
    reg [24:0] src9;
    reg [24:0] src10;
    reg [24:0] src11;
    reg [24:0] src12;
    reg [24:0] src13;
    reg [24:0] src14;
    reg [24:0] src15;
    reg [24:0] src16;
    reg [24:0] src17;
    reg [24:0] src18;
    reg [24:0] src19;
    reg [24:0] src20;
    reg [24:0] src21;
    reg [24:0] src22;
    reg [24:0] src23;
    reg [24:0] src24;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [0:0] dst26;
    wire [0:0] dst27;
    wire [0:0] dst28;
    wire [0:0] dst29;
    wire [29:0] srcsum;
    wire [29:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25),
        .dst26(dst26),
        .dst27(dst27),
        .dst28(dst28),
        .dst29(dst29));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13] + src0[14] + src0[15] + src0[16] + src0[17] + src0[18] + src0[19] + src0[20] + src0[21] + src0[22] + src0[23] + src0[24])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13] + src1[14] + src1[15] + src1[16] + src1[17] + src1[18] + src1[19] + src1[20] + src1[21] + src1[22] + src1[23] + src1[24])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13] + src2[14] + src2[15] + src2[16] + src2[17] + src2[18] + src2[19] + src2[20] + src2[21] + src2[22] + src2[23] + src2[24])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13] + src3[14] + src3[15] + src3[16] + src3[17] + src3[18] + src3[19] + src3[20] + src3[21] + src3[22] + src3[23] + src3[24])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13] + src4[14] + src4[15] + src4[16] + src4[17] + src4[18] + src4[19] + src4[20] + src4[21] + src4[22] + src4[23] + src4[24])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13] + src5[14] + src5[15] + src5[16] + src5[17] + src5[18] + src5[19] + src5[20] + src5[21] + src5[22] + src5[23] + src5[24])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13] + src6[14] + src6[15] + src6[16] + src6[17] + src6[18] + src6[19] + src6[20] + src6[21] + src6[22] + src6[23] + src6[24])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13] + src7[14] + src7[15] + src7[16] + src7[17] + src7[18] + src7[19] + src7[20] + src7[21] + src7[22] + src7[23] + src7[24])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13] + src8[14] + src8[15] + src8[16] + src8[17] + src8[18] + src8[19] + src8[20] + src8[21] + src8[22] + src8[23] + src8[24])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13] + src9[14] + src9[15] + src9[16] + src9[17] + src9[18] + src9[19] + src9[20] + src9[21] + src9[22] + src9[23] + src9[24])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13] + src10[14] + src10[15] + src10[16] + src10[17] + src10[18] + src10[19] + src10[20] + src10[21] + src10[22] + src10[23] + src10[24])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13] + src11[14] + src11[15] + src11[16] + src11[17] + src11[18] + src11[19] + src11[20] + src11[21] + src11[22] + src11[23] + src11[24])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12] + src12[13] + src12[14] + src12[15] + src12[16] + src12[17] + src12[18] + src12[19] + src12[20] + src12[21] + src12[22] + src12[23] + src12[24])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13] + src13[14] + src13[15] + src13[16] + src13[17] + src13[18] + src13[19] + src13[20] + src13[21] + src13[22] + src13[23] + src13[24])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14] + src14[15] + src14[16] + src14[17] + src14[18] + src14[19] + src14[20] + src14[21] + src14[22] + src14[23] + src14[24])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15] + src15[16] + src15[17] + src15[18] + src15[19] + src15[20] + src15[21] + src15[22] + src15[23] + src15[24])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16] + src16[17] + src16[18] + src16[19] + src16[20] + src16[21] + src16[22] + src16[23] + src16[24])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17] + src17[18] + src17[19] + src17[20] + src17[21] + src17[22] + src17[23] + src17[24])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15] + src18[16] + src18[17] + src18[18] + src18[19] + src18[20] + src18[21] + src18[22] + src18[23] + src18[24])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13] + src19[14] + src19[15] + src19[16] + src19[17] + src19[18] + src19[19] + src19[20] + src19[21] + src19[22] + src19[23] + src19[24])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6] + src20[7] + src20[8] + src20[9] + src20[10] + src20[11] + src20[12] + src20[13] + src20[14] + src20[15] + src20[16] + src20[17] + src20[18] + src20[19] + src20[20] + src20[21] + src20[22] + src20[23] + src20[24])<<20) + ((src21[0] + src21[1] + src21[2] + src21[3] + src21[4] + src21[5] + src21[6] + src21[7] + src21[8] + src21[9] + src21[10] + src21[11] + src21[12] + src21[13] + src21[14] + src21[15] + src21[16] + src21[17] + src21[18] + src21[19] + src21[20] + src21[21] + src21[22] + src21[23] + src21[24])<<21) + ((src22[0] + src22[1] + src22[2] + src22[3] + src22[4] + src22[5] + src22[6] + src22[7] + src22[8] + src22[9] + src22[10] + src22[11] + src22[12] + src22[13] + src22[14] + src22[15] + src22[16] + src22[17] + src22[18] + src22[19] + src22[20] + src22[21] + src22[22] + src22[23] + src22[24])<<22) + ((src23[0] + src23[1] + src23[2] + src23[3] + src23[4] + src23[5] + src23[6] + src23[7] + src23[8] + src23[9] + src23[10] + src23[11] + src23[12] + src23[13] + src23[14] + src23[15] + src23[16] + src23[17] + src23[18] + src23[19] + src23[20] + src23[21] + src23[22] + src23[23] + src23[24])<<23) + ((src24[0] + src24[1] + src24[2] + src24[3] + src24[4] + src24[5] + src24[6] + src24[7] + src24[8] + src24[9] + src24[10] + src24[11] + src24[12] + src24[13] + src24[14] + src24[15] + src24[16] + src24[17] + src24[18] + src24[19] + src24[20] + src24[21] + src24[22] + src24[23] + src24[24])<<24);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25) + ((dst26[0])<<26) + ((dst27[0])<<27) + ((dst28[0])<<28) + ((dst29[0])<<29);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h0;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h89c6c9fc0d15b34789da47b52ad9c525ef219df2e3f9d095f1bc85f3ffb44d5c67023b3d8795fde33d6884dede02054ea9c15f1e545b51ec525cd4cc9ff2d2f3f808abd2ded6c6982bd99e61d893;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e35835dd1920bf57f90c902672b330ec8ef5a83a3a56d875f99e2fe3d8ae029eb3c4adaa508884e19f8636dc9ef2b3908739e6a3231a7f7174ea7e4ceeba1e276e819545b0895f76ae5881e97fd;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h12cc79ce9d91a694d85ae5d0434341c9eea1a3db95dee996bfc6ef7a53b56df34b751d51e2552f9c972eaf299bfe58556feda06bb133eec341bef0e0d7a0ed95e48e9e8656c8600c97f3ff01befba;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h93a60d5174279553e4e4471b0f41aecb315e5bac3c55219878210f292e728389145a38a90416d9bdf6132d7d8b8576bea4db46f0f77429a665bebf42851b36cea327cde656d19474c3b9f3d83cee;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1473b15fe300121a08314d20f0bc263e78a6a434db0cacf2b00352b08a7e259379009eba4f0ad41c41556d621615470728ca1bfbe2e4e9ac7d4e0cffc12d769a5bc937cbb02d1e45a1c9cd65844ea;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he0f752107ce155e7806a171b6cf0cadda2ae1008a014c7907c4282a01231e0f6b5129c59c9734433a9ae432b3127ec2b0e7d53a41a9fda2490649cf63748ebfbc7d9188679af0f02066c6ede94b3;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1201385a1961071b2ef31852981717fd9cc27f92d1c18bd45be3a8593ed78c8d3472704e871af6217fbe7a2ecc536cf3dd9922a55cce0cda3e0380fe3396c3a3cc377d3e02b2d3f59d14bd90edc4f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1125b806460c7c2e3cae08482ba2f01ccf9add450371ec85d12f59396db953732d9f87b4dccad7d99f31c3e1468e958f4559e6d2d8b7db550fb8179e905cbdbc0205d288745234fec2705a244828b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h8eddc9e55128edf99382f40b4be6b8b7d9aed067dc8e59a6fdb96e0c30aaf032f32b2a6a374eb17600df03f0e6ea5b0d4a236f3d1744c849e3ca2497419859965b454c8fc3bad2f0c3817c39f1e7;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h6e5e175d26e7a1509e32aa2e8323a41da25a9421889acecdfb0ca10d368e31c536da5cf7288d07c7a9bbd6585037078befa31e822ac49e3aebd15356ef46ee52e723074b752f5df401ebd16163ad;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hdee06c06219203bf739b5ee1516cba34bc8cbd7115f7fd7e2454783f92249aebbd3d389def4b1ad6536eaba66a8553050104e31f73fd5a0646a4fd5599e5d3ef9daf3cffd51f3f069320858957aa;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h192c8b8fb55ae2850098391318ac71df0ef9da022e9d82965e0ec330d7b3fd39cd068e345563a957c6c5c4dd84c22c805be8d3993987afe63c033516bd14c160b7dee9c02594f4c42f86b8a42ce28;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h3e3526f9e84746498af0190040a413b2619fcdfc49913f933e0b015845532ab46914ebbe4f9b5773a80e51585ebd97ed13dbf2df02d07ed918d28af09c0ba43afcf13991e70885ca6ec15696dc07;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1eaad1fc499672b2ce1fad1cdb37d750705ad3387f744778d7ebe1920f0175348098bdaebf167b36ad99d310fb146feb2d0175df56ff031036e590058ecf02da25ed5e9e18d1c19dc14aeb3fed722;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h172b23216b8973c01c56f3f0f672345ebb839b4232bf1e79aa7daa9743ce37ed0abcec3c157b88a0305783ae76442e52c47a5e152420cf18a9447602ca7529563f7760cb0c896227f4bb9153c605e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h6b4b97bf58f50cb6e69f50bde8360ae109f99ae6d3ed46abdeffdf0c78735cc9ae427a07e026b411c8534a146b6fe988dadccb7dae8833a6ab8f31c35f04f7f01be1fac9e2705f7e4afffaf9937e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h18f9bdc1404b94f2823190d6b64a6efd27b1a7337fed3830d21892794546f5b359d353e3838341b050da9b043ff36a97ac6f248090da721a67d1bfeaebc387cffb996d9ef5e70dce57e9a72f5fa4f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h7352add1158b66fc5586c93b0e0d7ceded2d2b52afedf83ea537fa99436672c51eab545a60bf3df09e28ea8d5c059daabdf36be0bbaf2169715e846e435576f692e3c4fbb6f32acd772d1c25ae47;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h144cff6d917fbd538d38765a25eaf156cb199207cb1206e12605d359edf1de8b5660bea46d3b5e4c96da297d8080aa0cb0d4874868839f79e525850b6961115fd5232b0b3beb484ad69197703e5ca;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h469505e0152332edb14c0431faed7e67e63f4819847bc2a51cac8758e810175fc02c91c191773a564d413186de63852131dd7fff7ef8305451f9b048019fef453640c1db174b042ffc5f0b49c847;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1be354b789dd2d7499192e725731841af8706e2227ef3646f1dea9a26faa92710c1b6f63509700980b1146221709edd6cb40d9358ad46ba0910271ae2eca897dd9f70b0fe478e45af706a87931251;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h183a7f07090a63a5b9d921c73e4dbbcde8e15041eadcb3224d7baa231ebfa7886eb5f1040466922c78b9b6eb095e23455e5d924b2625a27e1911832f995ca216b3fa393f21005d76b0906cda8dcef;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b178e03c850a62fec0a7681cf95113536417a4c17dc2cff003d00dce14e84ca8c430253a9aacda6c16f885fed3611aca8d5171b836d6421a1172eca32c04c32f06ba3b42cc3996cb401030e6d4d4;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h188f7b48b170c794be82d1bc408b09804a22d784014b82242b39e4d06fe4ae66edbe2f18f310f5cea1cb332fb88bc5c0feae4dac3f7ea427c468dee5a3ee5037d421ccb73f93becf1347cccb7d45f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h6e7788f42cf962561d6c4015f8fe4f4316e6c7a93141e821d74eefcee14e686565fedd297f39e518667a8adee7bafad17e7ff81a08e70d0ad1b1e4a163cf89a2245685d885fa84d6e69f234432c8;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hdc577f0c4362324789bbafe7b50aca5ea60e603e37b2f3b45c3d3e20c5f0ee98e3f8b32b1a747abfdee46a016b4a4fc814f4d6fbe239cbd03cf06b2ada155602b4a61006a6440f92ee9b3b5f92a1;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h7fb9f0a1ba4c357c2d864595ebe0164e176e21d61183b5572b8328b59cc1f2db8fdd0467b18c8f51207451b8eba7034cea997c2a888abdf700ab757de6ff4dfcc5ad3e12dbc8943305cc374a923;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1bcbeb44c469f49d59bc68c9c4165e4353ae82a42b331748cb703ccb35e8d8ca9f0a71f7381c9df816b185f802d51b262407058e05b67084e1fc448dbb257901089dd3bb3706d3365e30fd149104f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf4e38542079bcd75b2e790318f309980dfa343a904531452668f9abe679e7dec52bde8608fd80f02c702f2937c30164ca900f9b146982cb5428747cd018e6500a4aa969653233c6f29cc7c06f65b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h19e0c5142af7a61384a0d12c1dcc9c2cad11bbd55d731176080d5d079a4e2a15845d0f63eecb8e26634ff5520c7ff4239ba21f3ea389bf898d3d88535ba631ae732b1c3d43f2f8e81fb45a3831256;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h171e73123338ca4bacad1d7b887f92aff16bfe39e5dd9aad0750537c78526177fbd9dacb4eab2995ace12ba9c4c08cc2ff09fff0f02d134d40020e2f8fcd4703431512901d54c9cb2db1f8ae1527e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10db8f9c4b81bca6d7d71f4e7e7861010fdb5ebb75377e1332a558053ed478b3416443db59e759d272b7c8d840bf620e8d8f4bf1c1e441d09cef8d7acc9efbdfd3cb78057c3db4305db1940f3ec1;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hef2eca54c1b1c9224ebec17bfe4c162074e1ed20d71893a74a6c9ab469588cb3c738d106110e3aed5e984957f7b05da2128622315b223cd1b9f0b7e092bd63df1cf70f9d73551a11b03ff2443751;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1be370cde3439b5fb01c3732696f705f355633e01364655cf20ac74c15a2edb25ada456b7ef7bf9047bcfcb570ea186589ae3e747992dade6017911d561d7a4a284938709b19b60dc8ed2e18c5953;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hffeaa1aba9621a67c625e0d0017b0420ab70a09cdc638f4f410bac4d03edc3ebfa6c88e778045cff68570312a9fbd3001c6db1d911e68ce8e0d024c891406eee3e467aab792b06b5d760d63d92f5;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h152a595a9f273c1643df583ae5e6f85b906d3541a336482e52e960956c5988c316160c438091b5b6995a76739804fa13e810e39bc39d99e7b8f5e95ab484608beceb968b75d2cb0868fe39f076c1f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d3f3678ec61efafe35941a5ea5a299a2f79efc4651755238aea292312d237620bd201970ea627f2c3546a00a976ac82633c7fee4bb6f9e3555e146a3cdd71ba1f7359750914e65d4b3557cd793bf;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h15a900734da9f749911fec4dd2fd6a2b163c0af846ca5b402ea3d12b8953385ea504685c65802682348666b000e7c5281042db015e08964a65af41c9f40b9b8289dbfd6ea3baa34016eb829c342a8;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1cf6711eaeb9d49f3926303251f15228fdc1419182b00d7a410d9022fa69e2a00ae872182ecbd82a09c4c2469ffcbd624ed78be8d6ccb30a6e8cd302cbf724ad0c773f70283741042c91d6d086ba8;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16d71220ba83c8f67b71ad5972ce6262b342d0545da15527fc9923af62a1dace9b34eb39ca5cf51b5e17f8973391111535be5be55d36ed03a05d2773dae71525e6dc327196eb118b7186407c7a263;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hce182a10da403e53dd3ca70324c2e162f179d349fa4cc403946930ec7806070e9a7730694c0b100e60b288ec814f9381e260487c3dc0d351666996687e546bf2e9d0080bc51a5d777a3b3e8a00a9;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h11cea380c7da4cbae41de9d6e4150dbb53438956d1bb0178a77d7fc3df14c6ea80b65e5fd86d0cbac8578bed96edc526a4403f06ae6fd43999f63577da81c0702e14eb428481b1b3532a7595a6f84;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h320345a674c6565a27dc26720f6c0eee49e402cabc05065936053061b197ab80953456ec052eef696297b43be1933c8c952a9079563616e2ea5a1490ed4f020a66964e749bd216cf04342af3dd88;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf469eaeceee730f5989a8b455b4ee6373ef1c9fcbbdfbd16bdbbb1e7946b34524d80120321e2a0ca350761472341a151c2e4455135aede281fa41ac28d78afa3321c23f8b8e90e28168b1a3b1025;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1eba0cd9aab8fd6d52b8e0d8e201d87c097af1cc8478ad1901800148d1f352e697768d2c4bc32a4282a69ac11e239d1e87ef3465364a4f7aa66aef9467ec2fef1f80abe8b1fc5b5d7f0537490e54;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ec73cabf14b150e26e57b7cbd57e45da5f828795a0a16f3f758a73421c294e9457ad907f98e25ce13ad299a8dc90df36f332e01b30db8ef033cd5425d0fe301fd0d8f3337df9f416fbcef4ae720f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h623ffb0d63ac5572779dcde22fd8e0255749682e40d02cad62a3417073103557ee2f49b8952048fd2df1217a090652fbd12a5aa06d62db966b7ff302415585ccb18d35a5f1c4565d77324d6ec535;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h684ec48ddd8a34e05acb153be66b9d5a94b2d8b7959fae3be1abd3549c29a690bdee474809702a5978931cfd0c784c133e8ecf9681d630f43f243822a86e3d0001be1506e658a0ced3999142ad3d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1270ef94eb5c79e585243f076f736e2e8aea72e6a79c8a23027f337b28017a85c1534201e73e731c2f6c0dddb3742f1052613f231ab5d5ee5c788db4a6ccc5235064724c1e73fd12f50df48555df5;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hce1eed0be97b05076607171dc90d0eb4db11df47f110dafdd5f2babb3e560d68a711bc2e752a2d87ba2112a49ce62d6c79a8698a8654365da252f42ab06e07ce22af36b32d13c82e70e2077f063b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h641dd91bc17b2e520221de31c3b68aa730646da26710d6be5fcf878e02c4b5961658f9d75cd74e9e686ad3692a3f558c41eb917ddfb53627661c8c13504a1665bc7bb59810720c8aa26c36740d21;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h8c2dab55b41aeaeffa0be9f2ee772bf59a3c0d379f754465eef10887e886064a84c6ba0f9f8edbfe5cae8ddfa19edbc1e0de68af14c785b1cc50dc3b1e7394784db867ab0e9912aae88f486afa0f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1902c126912e8d615ea6cd1b5df10c133a72c41fa47dc06a08cd5914411348639037c0058ba536106965903248379251df16a25ea2408ded9a27a62b15b96a0caf1045925a65064fe6865a082fb21;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc6868da8e8adfc046e9f2e743c117e0ad63e9b9f56ee4f87d3d72c848d5e67015f0db89b074a0005ac4a7a6fcd50032c95be93ae5b833ef68f163c95e5bdab0a8c6d1c876fbb03405d004a6f3ba6;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1aa86002d3cc6d415e24e37b1326dfcb035a16b804d86139254a1c543eb9bedf884d6645652e40c40454c5de3c5d1553041fa4e8892dbfa81f89ea374c0c51bc2d7aaa28a23d987a42fe3bf65da82;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hacea7d955b45856280a811af1955d4b97c43c02ac103261f8de67d64ce5a12e5993c63e5208b9069e18d7dcd86f94ff75a5d07ca92a70b648a9f56bcb1dcfa13d1da42d75bbe8d3a0168d8c2bac1;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ce090f9dafbb5ab2a44e94f213dca526d22f382bf59f8c192a4b30d33eeb3e74c10bb5838fcdf68863c7740eb54e93d885b6400a59e1ada93dfbfe682af2c68b4266d19333a2723c9450d0537ef3;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb7a7d6a3f0c1d1081c6d67d8c976f1119cf706f35f1bb2be66f34a92e01a18067f5abb595291be7b663341bbff0f223f2b3be41c1b6a95a0d8ab62f75a5cff220991bb3322a0cf703e895ac65878;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h672ae9a1c7025d01e4ba2453cb5473f360c24566f8bbe46ea656b49df0816d833d6fdc412dc869f1eaa898a62cd5f845aade62c61257e382a3d715497b956c77f860d00fbcf5fcd446a471ac74d9;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h4d000ef4f743c34fd6eb49eb4582a8cc40ae027373910dd916ca2d4964e264206eb7e86e865c4b0f9c261871ec268edb949be5709bf787e8e1115c13855680415091adb626949915c1269ebff90f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h12df489584d46ffd897096635b30599b92ed73e16ee11a966af4e14db2407f46f493deb1640d45020702ae183a6b899f51cb2b7e25246c8b496fde1be20ebb333f53f63eecae8204e10db10f36f41;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e3c5e0a9894eafb856d780531a507619c78dcba9ba9c32383164f69a9e61fb27862b410b2fd5137f506eb536e8f3b13c159f50e360acd7e48623c081dfa32bbdc3b52d421a96c5e7fe1535acfcfc;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a47142965cd3be3eaeb3dfad5f528455b2160734b79f90ea6608dbc9c871f98acb613a747a58e15e9331484e33592d2cdb531fe520d02512cee5ccb0106934738d02d359917e15ac23db8ef6f30e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h9d3b0f9526dbc876070c294dcb7dcdbca7f57d5021f4da0334ff84821e43cabfbf82ec2ef0acf18ae81ff305d2e2f0c40c63229cc438c7eea9934a89c438b8ddadf18c45257b04a79680fc0c214f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h24887da91ecf9b6015d79794fde2be9c4e9fa482aa64c9b2b8b1db341b60f2fa682be5c5350a03a64348ef588771d31cc11ba008ecdd4e63de6d4b2c5511413a186d48753b842838cd9ed59cd253;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f0fa41bf1692b7595f1eeb4f06550a84b46aa06de6717887e55ffea73cdc1bfb59133284199942a738cf9cb22371ab5408d46f1eeeb3d81b33ea843ac93deb5502ea1b942337803ea9dfb62893bf;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h124af80956f02be9d6a310357326e973a68dde9e4ace6c0a90923c91078bb79deb796b685b24bdf2c7dd80d33a95745b5fda63953c486479a699fc182e4537c18c87d0e60da7210a5c696fefd0282;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h407fb4321874e7ba65965b7ff21b1ffdf8124c394b247f7765337ddf3307e7975c860a662b9a6c5b5fd7996bb8307ddabef0c3a4689d493793d6ab6233e5a202a9d40c0aaa71ca4be0d1df6f160e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h2275ab63e9c4a7b7568fcacf2b3edb6b193dbd601e585abecf0437e4d2d92ff97970b226f292ef43fa8302ff6a0d0fc88d4616d4f1d2d1a43852e642b5e5713301eb7e86ccf8aa9ac2c347089743;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h198dd6b7847954e1552f3f190925e0bf815ef29ad4d916251c4b4cf1b18d6f45416a3130eee534ca7884dcb1c688bc4d0074cb1fe4695f4a6773cfc7fd03dac69ee3b1707c5abe2fdf22d3621086a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h11eb9bee26363bfc5b76658118968aa8a071b1f623f765ff2a41d111b2c37ccce8355a0d102bf1f211bafafb85254de6604860e3f37eeae8676de70a2577d7d2cd605e4b1f7bf8d5522fac55c4f31;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc412c774dc57b6f726187d2b145640305b75c6a1ba53f901d82068969f173dc1d247c6b27574cc4a328b4d4331eb8901a690b84aaa607eab4081b0c1713566b8712d35db6792fbb47aba2b15557f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h14f3615fd54b80b890c00f6f424b68aa6bac1e9d562dd816aae63e64f51148d8975e75912c8e3c90c5862112e464d1b9cf6cdb4e332700500fa05c546ba24779b54b8f6aa178644a57379b1999dfe;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf09017053f2b748b2ef2cec96e151dcfe5ed47ffb5726d3945719e4275c16ed0bb16b05d226cd3b784f859e8b02ac14667337023124089c7cabcf00faf96eca4e25e09cad86d21102e12e7af84e7;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a8c1dc0f8f6c2ff10778a633c8662ee5b027294b807fa22d744f7c05fe01a8d34a7660d9bb39bcc433e485c8ed68e38e6f88cd3a364e7a26b0beef06a41067a6ef83a8c0959dc54ab255db139dca;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h20e25a9dcd4dfaf9a5f43aafd914ee99b6b2ddd5e9958df34a6281a153cb23291094909ec09b01584ae5d3a9fb384ba7dd9b86b01b8eba9afc184b600d96384d6779c29f6b9657902162950aa956;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hfcf0d6af255952965c8fe32c5f27c4c713a9a4404931ddb7bc5d583f3a75f008bb110810026f8507d4ef301a653c18903bd6f3f302c5d1d019d7a7b0d8d3c641ce29afca0d04cef622b3f9989ef7;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h55952825d8db7434e267fdf0b13c5bc43faed7f82d60dbb6a69bc5f55622a905c26c064a0b25fe71dbf4008f21de7f3bff85731108d471fb55e23c19bacc44e204b92c6698986ed6adef78d09d93;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h96b20d891fbc1e31b4213c0d96b1a9ee6cbe76d1b09c9c194db21c45c0b617e1cdba16ba2963f599f5649be41e44287623375cff001014de6869c444ead8812390efbea8019ef55afe2d9d1339dc;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d1e49d7a7d495abe69d54916a43285c1035497cae630a0a0a57f0142d3278707cf42255a53d0fb67614824db3dcc1db818ea96eae8f7829f79b2f5e7e24e4542470c772470c17f2dd003e7f3b657;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h13dd4ddc693d7766ed490085cc735419d778032763f5bf64fba8ed6210017cf4353158288b8073a60fe3aacb69cb451a910676e1f2ab645cea8e0eb2cde0da9e46f3fb4b91cb0efd42b468947594d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h118efaa7430dccc7f5673e7431ed58746e0b1bbb2b6cf534c1401103b2099bb89a34a58d65c1d9a1e7eeb08a0370fad277e7df7f20170546031b9b5bf3330195ff303567cc2c6ddd47ccde4d9e53a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h55896ebf70b7dac0865f87d2691688f2023c2b655576f0613286a1e18749a1b8016039ad0c08d801e8fd5fee81189da0ba219cf395863caa44c83694ad76f4eb7ceeb3ffa5037717dc86530f964b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha34203f7177a7fb57ddd7e4b2060c16aa3f000e5c4816387804df31a8f70cf7d7135f5e473101641460a41fc4130e09fb6e3a7e715ac99b5f5ee3dbeae7fbc70b5bf78d00f101c460622ecffc9ed;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h149f16401be8a529f325ec1831e726b7026a000b4841559fe5018a0b9048b064e3335cad05066cd2ac5c2dd8ef452cfd6927c240cb194f34723b03aad3369e7487d6bec6cb532d79c5307a93d9fbf;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e800cbcc58eb4d18c3cccc1148a5773ee5b5ac8b037d1c60616b4dd7b9b1a39f30dad0d91e171e2107cf6eaf47547da121dead699c6da6859023cc1c13c48063a0681f9f81ce7743ee4f32a9f487;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha1ae4fc48dee299940231d1a3089b233b583e9de64f3dcff4915f08ce77d7073f3ba70b50a1ecda3b671abecb3aedc2a51e2f0d342da1efdf65b2186d530caa6be506b335da89f3f48953ae851f1;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hda90935d1deea701fd1194d03ea6fd1986c6d2b166b33875fc093cd82760bafe82ad8def451c0ce7b9576643ce7608bb63b976c0cf0f6cab180642b6ad753ff27ad6c0b39faf91b12887e5ead3a9;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a1137cf6384f0513e3c1513ac398fe3c6ce4b94433613113d61665a24d5a6510a94d2305f4cb9c5be806babab7f4131a4c2d72f83011948f48da43287ce9d51b99e11d9c83159219d44c4b97596a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc7d9f39ac127ae4c2fbffed263965c439c9b6098fdbee51ce54926536a7574db2f844307f76d7dfbd4ef626f3cfe1c850923ce0ee8e616e9827d9eba446903a86d20e971cbb6a0432aa043b143b3;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f6a4c3b43835a3836719e38d57acbcf90811b791d20332d081c13a15b45359ccaf810f41f9ece379e0124861e72368fb64ceaacb8e39ca26958252bdef092af86ae0eb8148e3b59dd73d860f17bc;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h30b9bc78b4717529f5ceff50aa05964120ca96a444a3d4cf263da1b7f2038262d876df242737639ff7ad4c63d093dd08dcc717de3031625bd3f1b0b74927dea9ddfd82dbfbfc18b5b6cab6a909b9;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h898682d75d34bd17f59006aab3c08ca599ebe9742750fc93ff0cd93e0cb6febb27fd3c65303fa827aa28b3a79b7b5dbddec72f08ae8431c86a201db9cf1db436955c77e0da78ef200eed0c3e34bc;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h6bd0cbbdf498777f8142b90f935cafa89f2790ef6ef1cb13a6ef94fe0b10d7e6d95f3e42e89c71a143a842b1aff12152cd38bea67f3213754162a87023829de8106fe3a6482845a246edd0d78f28;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h8790a50ee951159ad4d7f43359e9cf23e50896630e85bd84d84e53380e3ce10dbde901571ad264796195719c627dec6bb00c2aebabbc8f33b6454c766ba58b3011ff5255da7ebca5d33b2b6bb0dc;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h15fc216291cd4d1c74a463c05e9bef305b4d36e5c8800c7070ec23c764a2f1efa1732c0cc2760dd4bfec4523b467477c83737355520671edcb75346bcc7a47dd27cb3c7ee2ea3db1a27e177ba3022;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1df66842f95976d4909c15bf048b4800ffef31f4b43810834fecb4cbec800c1e877d161c478dc6582f27ace0f2138057d7454920a643c37d2f64f5c036f61718c16efe6c7c9fa8e3d6514f0133a18;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h53ed2d46b1334e5da5612528289b8b110f5c3fe1b6d8e2e566575675b0762fdb1cc9bdb3a42b61baecb6af70fcc8eeb89fb60e1d3b679fb58728feda4e767b69637982a87f311c8b84871ccbf511;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd1be3c495bd59984eb47762fb3ca51aa1fa52c20f422400b4a7ce7de8562a40c8438591cb0afb6944e565cccfe0f4bfcbf7da34a44cd602fddbe7d8d974ff1746dc498959b6980b501a67ecead0c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e5b5173c410d4f8fe365ed6acb97142ecfbec3424a2073554264539339efd28e0d51f7675a39c49f154bdef2658b6a57c2a23b15a0734d48fcc6a207ac1ae2c96aaba84abca08a17f860e6deba2f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f42f65e3fca3c32622ab8566a93e76fdeba27c71723fac01c05c0589bcf1cc501ef2ec0cbcdd31b2880d48d1471cf668d00befdf25ecab79b29956514b119f2f5510ff6a5da68c53af3a9dea173b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h119cc059c152a6e7901b2ceb7b104f929cfadbac10228c9ddaebdcb811601708a2fee9e888388800b6f64947b7074329cde642ef931cbbf4f19b79f7cc8d7e5e302cb413030a575dd2c6e29594f71;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hcd1a8c7ede6a98e755bb3d99f219c2cbf5c31a168294daa4368f32d75c2ed022441998dca26a083bf7598195fe1ba6b2be8f74695d89e414e6fbb0c16114c66cba78ab078aa5c909aa71e4928a24;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h938a51dd635df52ec515bf430c3e40e589aa634731b5d6f5f0de78fa57b8513e9e5a4c4612df3fe159bfa6bf27527220eef4ee685ad025d2e7ae09f511626d32c6bca4d70e04f0addc4be2cddfd5;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h165eba7e480c461aff7baebec54c2c1356a89a613e1db67393747ff945dca20eca8c0c9a11044517d5f7baafa74a2e533e680914e76061256272c9ebfbbc739c5a62fb6601c796e4d62bb0b546a40;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h11e87b1c2efb9950a28da890490fb654608d817d82e4d8a25bf7eca4c5b327058d0f8c9fad2304a03c283c700a86058d886d37f4168ff6eeb04d383f004fa4acf10f8471a5ae39089780d355a7b86;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h11e1285398b9cce302b102c32731f02a84e8d5d0e687d626b93e9caf1a38cf8e6a74f4736ae22d066db76094d0a4a0e485f228c610d0f3bc119b021656de2302bdee9b192bc1320715cfa5916feeb;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h56b3a81721a8ee514e4268670fe819735f551a5fe8205dff50ef56119343b861bffa413d632729dde57dd86d48811ca4d4637afba58c72477ed5590ed738e43397761dfb31ab0be9b41287c54d39;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h924edea500a8111515e8a0d94b6472344eaac2e4ca01e4bd14b3d5b5e10c099592088912a23e23d4a1d304493dc6129a657950f8e5abc9864f614c72cdc6df9bc3bf7f1d1b5e9b6f051a2758cb1e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h180c7ffb0ce8bd97e724e50dce676734d796cf5c150c89257803f1b974b6cc8e8bd39bfd240045f080fe17628108f534ca879021cc7efb5162d0b248b78171ddcea6aedc48ffbcba934b85d0ad6ed;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1cb9323deca30c2cbf57b963f329237e2a5a12299e75f7d09e4ee00a5a3c59affec7d4d1d910752191be92098de8d3258bf53e57f04056ade7d10822d297a33985bfdd52a4bd062145ff85c06aa0d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c7eeb0e86ea0c65cd4166f8cbb0a89d158b973bf71f96ebf4cc200e786392aed4e5d4acd668c2d8ce5202ad68d403846e6a95cbbdcab3ec870a733464dee4067f5912469baec3ff17dd3cda18978;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h474229132e1b60e17fd26dec8285a7e9b7f59c7d117b97dd445e115937cc2026c6d057c229ea5e372af1a9c2513a3d0accb62f63db3f334aaaa9f0a3015593a7818bca697c2b8af4fb284d432011;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c5f940327bfda0dccd720132248f1370584785332f26a7534e1b299f46ba595738d8e386165b6dd610dc90a5342f388284a87cc0898b670362a1937058bcbfa80702689181e736bde4969b5bbdc7;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hafe886cd00788ff5ba1a1638fbacd27c1b3fc135a4902ed951e3c5f63401296dc03f2e8159a77a8c42f1e78efd4666962d0b7dbf6050df2145dde2435b2b628ea03a36029931d88b9567e0c8b00d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h9182b92fd0fada8bc4a8ab6613b2dfcd65cb8a758156ba7ca765df57a8069f730b4423b5a8cba31833bb00aa39b2486aed825b167a7a0f036fbe7d121b601d3e9a8770ff1a0fc81c7b15bce3225e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h86b5378667b012f7a80a2137ba30aeb0f37bce1b36bda22e10e499ac38e14ccc394257503acc0fde1eb06bb99851ebf57b74c94615baf5125b1c8a4ea30b687de512df31ac92deaf07ef20d9724f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hcfdba2838c1fff5caa2d38195d94d2d5e1e7c1c998140e4b5c303732f9e88f23f82c48b0c1a35f300906959d0678c574d964dc9198e25dfe49f15f66b5ad92f7cd4cbef1ac6608ca2c944ac087e9;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h477d5b2782a015faaed329b71e7f65364d05632639f8882ceb657f7a0c595a12949c94ee85c6da297af3a2e588a4c0a4fba4747f7e51b6e0cfce9cf20ba051d347def046993ce7b71d809538e5f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h13d64fba121162a62dc8a71edb3e7aee3e82410fa14aff0da1fb4f0a0532e5dcf0aeb8e36fe3b1af47acf3c4d079f20a00eb3f261e7805f682a21ec4c4a3af5c92febfd66e6360382a61c2438c39c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha3e826bea42582c073a01e5349ed143a5af61632c1f2a22934974804aad68ae3afab0a9942bb952c62df246ad8094b24a7e02a6768fc3b4e1f87d6fc098c279c89a088655adf3be8b4ae9272bf5f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h713c742612320089c6a1d2552fa6bf266d58adcaa3c303bd21c2a91649680a651971c0290cefcc12adf24caa0383433fac2b7a4ff4d8c870cdf47b6554daaf12310ca224a2930bfe852c4cf1db4b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d0bd01e123c7c4c4788e1a4fe726432755bdcdd0dbba37aef974a2c9023f42e0722387ef5c50f2c30838ca84db3528a721173cde3336ca0479b9859b1b49bdc104cfab449ea4f4a542b9e1212727;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e6842b187a4a10f64c00574db962ea6c1dbba4c1538622be40f29f0211509ae696f31496838e79627081971192f0c8f2d73f60e918bda7fe89583844a5bb23cbab5e826c4509f16831d66a2922c5;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h19c2ca57d4b5ec1e216801fbe501e736a02620a5b1b25cd01c71274a1350da7af3362719c38ff3546d0a22cc7016348f5ca4442e5f41a19946687f9392c1130e50f488968d04078a383e0d9453598;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h29152957d4987bac6f02fd58a24f4cde2cd83c803a69890a5c1f49ec00e0a696f5ffd939ef7ef88d2b38994a214e5095cd6c6a33bda771edd7654cab4dcaa80c0acd662573d2fbe2a4643e9eb3d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha29f7524a0de89b28cfb05abe62fed97865d0e60c49dcc87e4e8a5fd6307d5e63dbf277c842e87e9103ebe7b006a29c51a58140e2f6e741125542f259871fe0cb741fb46189e15c209afe2b059cd;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c4a57fbae790114b2fad472f22afa9a41f8704f21cd0a6a270350731088139f4b03cd3e34c309c20e135bbb64e4a789ec8d960a07a191195b452340fcbd1e04fd2569016d9ae164b0ebe64880374;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf95ba6c541748a17e6598bc2ebccd0b61486878e806985bd9a7cfafdc5cad312d0cff7efb4653a9631682ed0916f5e28738ff78d33400e66e3ae8fabc1ecb78ea8be1af3398b183aff81f38c8b5f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h91cab7a864a6435fbbe5c4ab72bbe5e66c63ddcfeb8320b0c15896e42337151da0db712a55c834194097835a575512ab176f76afca456bea36f0e4ee12f76ca7abebcc1b7570c3c6afc147c59921;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d187b4e02b9d4c147f25a1d8d33f8abcd1cc0f1bf2a041aa321f06fcfeeb4cc693d97b8379f98971e69a6e35e1aa4368726ed25414e5eaa0e485e46c7a50e15c88de5ef950614f013b3a0f65772f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16abf43a7d39240bc7be292ec0d23cfa32c0251f7d2b61a28f1e043e73cfb2e71f232ce041b81b78fedbe95493b9a5bd4aa88015124153bd2196856e0ddb4817191de020bdc65a3bca21f601f371e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h14f5c2923953a2dc3cca4da359b8cff04ddc666f272f8b3ad969a039d17a30abcb8e919faa5f80cddbaa48768c9736deb9c6fac034b2f25d43344095c4cf8b4e350cecbb43eb91e780e47c748b333;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'had976b9be765918618cfd8ed673f4a3d650edcc12328c82b88bbedb92f43c31f7d5eccfd2495a51bbffdf4b9059eb1d6761c404957307ea788bcbb71a4118f39072bd9b1dce08b1c5f0bd14f4d59;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16c7f2bedb8b202930a4cfac40027ef6704a3489f9b53b30b73857e68cd42f59397e2f60737067fa81abd01f64e0fe5402f26e315da12c81088e475a7dcf6ebf6a7b3bf0f5b545f50ef4689a920de;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h785f2ddfd986f13e2b5e77055ff4176933c1255686189a254d3d228c7afc7090e2913fea8e6ecb41cacf3adafb82bacd5c8c502d926aa3d08b2ecd71f13e3fbc55a27598969dbe1cb53ea3fae62d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h7bd6adda48038a14bfb403971c5f980c09d37e12dbb9d2f6b52fc3ffe6ffc0b149cb6ca8e395377bc76ec623d1db28923040cf896cc3a64f14a85bb1152055c708fd298e9f8d0841559b7b6dc6cd;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h140dc3c54bdcacaee9554e0c4c270f8675ee8e23316e126238f9d12c6a76e6ca060014f5e3dc0fd94d2286a864bf4734d5e51d6f3c7eaa488e0342ba7a2c764173d7a445d73d71bb0ee7f97d53252;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h14c491d571b28aee07ec6c2b9944a57a3887f4616d401d5ad8e740f2f10a178a55a009c01cc3abd387b2ee35c3b1743dce632aee3ed301846c9766f59864654380021f632be5804baef9e6daa48b7;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h50a5090509a7a206eeec113e8119cdf9794bd3352af735e02fb4b9ce9535804dbdcc49a85c5a1bc0b4c8acebecfa11c8b070b6218591e38fb8a19fe3cfe3c483efe774d402099c698da3d2a7d4ac;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h799e065833b50b69b8904ae20220cb6d4bbbc7a2653cee258ccd3ec2d2e267c866ecd05f6662dd8db777749161c134a0dccb7870912046da64a2123370c240eab348d7a60c386159fe05b3ea06d7;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ab11ea13111acbb1d0ca1fe1a24d7b84c637c85b7b36eaa6d0ebf8b9bf2d8d725cfb45b753bc2406bd3c3a171f4391bc68c396e6a0ca769c9d8e75b24ccb4403c058aa2902f4c6503bebf3773a8d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h17560303ed1aeeb0fe26d1d09b1ae1f0d99c305b4a4cb9895b6995e67bb03e9074bcba2a34cd74281491a1a01520039be1f044c772c5852de6e173f3be7486df5b8219faabfd3da31cf2baad95d4;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hfc9d68f53ca68156695408385cc567e8fcfd99c4f0f4695ef60fe22a8f09d821705b35770b38dfd56ff73356b0e93dfc5ed50c064d30e1879aa739a5588fd5dab4b3873fcd56014760f764b4a015;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h6e3f1ecce0416ab7f9d3bee16eed60b7d604f221ad9ae4ea432eb70a8bc5158d4057fdfc11f0c3a2fb4648d16a58ca316150a0f14eb97fb82a1453ff1d55834f5a969c0b2194086dbcce6aa1a17d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1aed9bb6e802ea2a63ffb9b139cfa237831796c7f1b1d3e2c8d02ffcf4c580dcf46fe84463aaf982bf61dfbc8e286e0eca0991ec2d5348227c68a677054b3922f7875f0a273fe10bc3b50027b25c2;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h11d3fcc39cd66d3f58d9ca7568ba14d300b2ba2b96f4aa6ab637a60cc68136de6306f30c904bd0c42d735b4f27132608512515764b0d0c65956bea81c8c8b3e9648c148c8715d6b81df659380b604;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h11aad8984a13bce67329d4d8a9bb56cf939acc6749a25a4e63276165c77c556bfac237706a82b32c7a58f35a0cc386888549afa4e5bb70e41b4a7dd240cf9118ad8afda642c8d35d29d7278dc4c6d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h133a9ab3d0075112517ddfdd1c4666597b2bd1586cbc9b659a1104ab33e631dfb605b2ea1b70d6d965014883c6af8751d89f6195acd7ce4d112b21e2870a172c22e4ce5fa693677ef658dfb11f9a4;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h11da3fd4c1e5d4b77865966c715a3bad71070afff3b562b3324371c0cb3debd93eebafc6a2e32981ec0ed25686a7a2412fd84b3bb70cbbab1779ae2430d153e4550991c3b38a98403827ed87abcf3;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h22efcc14dc91e9513b3e0746cf78c89f9ecd04e7f293b90855f537b81e24fdc184769f3520f7e8dfd93e127b4e003fac3bf8f5aa1593384a698f32df5a335d46d3c1e89d439bfd5fb25625c52221;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f9ef3fef9c9932ec1db3cb5fde299fac1d3e8c6d1d695d9334a5dabe55dcff6a7d644896825614e26a99e3255af51755dbda9ca3f9d6918e2f4b867bedd2a483c8f344f5c5f2f31f9c9e9a1d17a6;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1746851508cc4c735f3ce7fee20feeb15de0f36d133b1a230d93282cbbf1b2f462673e0d4f2e2f14ff5b36ecedaa9c644bf5b67ff0c438e600c0d9ab7943f8f078ea50efb05e4ae178bf50fdbf3b2;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a7e33cdff2b134a555dea5beece1152c7316444e53973726637c1af30ec8a5d60bed9970d9820b4cfd76a30ec5be3ccb83a054f49b13e05e9593039a0241130dfdcb3774fcbb5848ad851396c10a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd98e9c7ef1bcc0d643a17ae77626cfe8d276eb1c5e121495d0b6936c78c108c3b4ca16461278d51e85ae7efe7352b078228ffd6fb0c24d894e3f31934433f3078b4d70cd8df6d4f20a8ddee2bcf1;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d1e5e47882264e70c841f6ff383a592a22f8122d13676a22989d73dd43a6e0da860e013a905fc438fe96a20cb365b575431f81ca9245bd9f3d6c0e54d53c5cc6d0bb5c604b1ae64f10721587fd22;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d3bfbbec1a3f5cee336d62364907490dbda76b3f872efd0cc59aabae13f3154a19739ee6c31572a36ff88ddc4f455b501e474fa570e0c34ac6e02bfa76fe4993f7b66bb13d8f959e990f4eb7351f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hbe1bc627dc45400463d676aeda040ce549ce4510724c256991f36344b902e3e99f6ba1a7d8c6c5aaa747ec7f33bca504d5b2fa0500a116e5003ee2b3acdd2d43a2f08886eceb4b65c142048fcbf2;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h377446951661be1b0b93bbfc8d94a8a2abc8774c442589be09a273f20f5eea9858402838d32bc7d6a481f3fedf743a925cd5ae6413bfd7502af645831bda18367aae205ac4ed786c53e6b288ee28;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h137baba790b833b4e65ae52e2d6b7b025e33313a160462a9e15585fe26bc4c6b4f471f95c57ce48533e5535cf982ab8ee76a24e9cc51443cb528794f165cae835a50216450bad94bae22c50a6203c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h15560fdc5340c57b2c1d821d11977c547951023c58da8b432913870b3b60e0439688b9aefc93aa9f848eb89f01c3f5706e5498a0e9c55a32865e4a815d15c22789d812f7fd6d68e70f55924264ffd;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h135d8bbf71f007988bf2e7819bf4dd29a5ea5fcdeac8c09123b09e3bead6735e47d4f1daef400e1953730ac257f0fcc27acc3aa25fa9c0c518183d3fc1c900836e2f358937c7efad1a70b0c084ccd;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h18707d3103c075dd0aa303c65b3977bf06da378e5ce891031293de50f1a5bffc297431a50c99971652e5f338dc2ed6b249f1e70e6ad14bc241d218f0d95d20927256b10d86e1b595eafc9a28d738;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b8ce6b4ab33aee5533ace19ce219bb39ba1c8d9c96327a618aad67c676dc4b1e5a6fbbf1c072c598b8de2cc301031e1b50eca2891353108b297ab9251ab022f926b60fbe14ddd53c253d906e7cfd;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h186f0006cc00f0401c78a20038df292fa93588befb82f115645841a752cb4820a3af1d325b4e666ba278b8c465d31e503d86917666ee70fab843e997b418d1df8ea7f0d4fe3aa419198a89121ca5a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h830d3029498c450a2bd872b08c9c727d3cfd235f5b7b04756636fa24231c89f02c4ade6393458a520576913941e418c38b2aa6440e4b083eaf4c050ad6473caf2e6f1681482457709c371971bc7;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h91926fc5d8fb65798f2fa13e8fb138dbbf53dceebf98dea00dd55915509f317dea17b3b496568c0dc2ed19e06a8f3c434b86d15acdb687d52154bf2cfda73516715a0909f87e9ed827fa1431319b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16d55233ec92b777ef4acd9ff99f47837183d7939cb23902fb175e0cf0b4df1d23c766fa6e412bf666c0dad0d11297c102b0471edf1ad0dfc07e1ddff9f55df4ac88f80019b6dbdaccf408e8e31ed;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h17934feb15836274291b02157c7164bc2c162cfe1072a0410a1ba72ebd7943ef0d697dcd175664bd19f7052c6df84e2105fcb8ae768769deb6ee3011d184b18122b6cba934006bd45ee70a7db080f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b51eed12a8cb8e7fcd53682b7ce1f835ad04864c43b524e1edefaf3e30059f0d18c483dd397f76af440eb517dfbc0542512508374862bd65c7afb6be227020d468caf533a075a8d1b434bd88025c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha2fe424c20bc7a0728dec200205f5c6bcd25ff6b0c2c7ab197fb5f26d826edded0ca38a3925f4fc7f27fda0386a06ed9ad0ec4be7451ec51e21f50a67d677bd6a74a8f16ac4031457bb3ed891dda;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hed177d42e9b00b9851d60d9a612c26c263d430a3e163e36b90cfadc34549b929ab8a530e672ff66bdb28051a71d01f215a35aea3273f9b4f7b8d273b73e900e6e16056c9611c9c7f7e013fcd1000;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h9af3e5dc38aab711a712dfffad2b698aed25d152ec3533537e3c22ac8ecabb1e2b3d1b2945c524e8315687b783f1abb2fb01b72d9dce20d339ebf37c0d83c3cc3444d4daab63777fc8d93a6d2f9b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f6d151a2fbd943d28fc1e6d629cf421bd1b84c1377c0a74bd83fef25a3963e551bd7753b6be030f88b168b459a9fe2ec61a1d3316e37a3e9c1c88976b72f48b0e04bca39aac8c4d4d4f5e196b099;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h42e38741c6d0376a887ca3122cb2509f81191a882a802671c48a278fbd11f1fca5755f340fd363500948cc59f1a3e1b758723bde0f42dc698d2b46a204f69d59dd8afe1c4e5fee457eb232a93d29;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h13080cbaea2ea7732be749079af4a7eca90a93011b12ba80bf2a981928fd06670c838192f5877ac6947b7e685717df9f7d9305bfa3cba3e793a404043a2029157ddd43cee7838c1bf3b5f49f47c44;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha90f01eef25ac6e303100d6d3578e4778f70aa5039c0d46b29bd46dbd952875bf9fd7c88e09d955f102bb3974694ec602e6251f9402d034e99dfdaa2e83a511f0569a435abe3316af1e6388ea790;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1deb4c4cdafd3f0dbccd2e651d4352655bd9daafe880cee38c02ba0bc61e218f63d62f8377a365ee4755a418375ccdd9299435fbc1b0ca100d44c0bc72fab84387aca6d68eff16900d0b6cdebb2b0;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h18ac176164ca88ee70ff030249ec9ece2046b93531dc99f348d1437461a3e9904de991b2728af846d43d0aa667b7868d7ff896ba23f26448a0f6020333e5ba5182c505f47a31a9865e5e29fc0bad;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc761219fa62b184fcadf022343a293668915d59784367813ca6aec75fbe7576d7949001c1c34ec7394d500e8290e8e1a20878a21ad04b5996621bffb3d572d58038b1f639b73251619cd09c304e5;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h103b8ad8a06dbf7cee320eb959b67e3c3dfddb1611aff97bb1fdc598ae0fea0459e6d7c855a5f3a6c67806e92b53d6e40eb435b54d1ee50f1fa2e80f6dedcade29d091093ccb19bc4d00f19c8c584;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10d133355d0383ea3ff7dc9a3f6533b03ea0bf872084d81516af04415565073107345af81454fe466fabd7bf4f54136ee3bcd1dfd3574b23ef322175f28b06b451de1f2d54b0d3fd33ae2db495f9e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc396e974b023bbd48f3b293bb945580bd293340344532b521821fa2af0759c15f3292a07ea33be2be70af358b3678b924ecb2f42a87b69c1c3cc51a4d945706d50edb329c9599eba9885a608a519;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e37d4ba4c1dd346081bb4768ad1bdeabd7ff021a2951430f5841638c7cc625cd26801dfaf3721debdfe52a2737af18ea30bba91bb9f2a15206d42f411095c023b585177d1db0c4c9022c7587ece8;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ca67092d094b6552a26846fcc97160c3004b2150a84cc8f10ded073b88f19e14f1dcb27d95b45e2cf0309dec4ff6b1dbaac20925f6dbdcea0b0677912200684d79e459328ac81fd6f3e8eb5b4f35;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h2af5b71e5cb02a7d407d7aa105aac5c6eba6f23e943c989aca33bb0f4e0eeef61ed096ef541c0c22d492a71f89c567d88eb4f1c912f0f9e99af535dad5ddc725440fea005c6dfc7d288973d06176;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h18ae84a08435f6b06cbdb7057bbf44221ede73774fef8215ea2e7768d8fc47a6aac8693ae0a8c0dfe64e1a4f98a368631a02905c99fe69f2469a0cbda23d8e5dfdd4737cad697cc9bbd6db9dc5726;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f4c63356e0735dc1cd986aa55ddd9b3aa054777bd23c4cbdb53f8c2fe9cce7b8251e06eb7f65985ad5b97a93b9010a7e3b3058553cbcd8a599dbd8f667ec25eda9dff1bd6dfcbd8a71c2687bbf97;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc5e608afd300b43dd25c7d50ba253356e004dae1661aa16901ec7334f26456c1917f8977a2921a649d6bf71ba0bebb4158669f96bc9015535feff4750418100d06b9fb05c3068fb2e8e9bce0ea5f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h11c91042cd200378d975a71fd3021615b3a4fa6b5b6cc378fe8627bacfa05b41d000a0cc3c67b613c30ff783c69a4e47ffc48ca89dd6fe04dc0b3bb10ecdb6553c5db55a007889c8f61d968c89e9;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb0fe780e9671ced8143a1281a7c59df27e919d25ffe3ba2a4796ae2a51d8271b1cca510d0988b7712fc542f7bf32b21092767837517cdbc5351bf23885526ba0bb58afba7e3b8a52791b4fcc9924;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h17777021256404a288774ee81e02a69d748b2c34cf02f1968e410c6d82380d3e35f5893f70f2d5c27b98029595affa93950b0d7ca9c22d6ede19a5aaf835c6a5a06151cb1b390dee451970530792;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h6e4705d1a686a1067982fa8f3540e22733d2a7625e3d77ec2c5b0673543574da42d8f88e443937f1e1cf0d595faf8a518d4587730eef2679eb207116f836f7e1269fe29c9c7ed13aac3e8def3a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ec39a154a3d72d53034bf8fc4416f6e9002d3872c58c49ded29657c6b3b2818217faf13f4026762e2bb43b9e6fad0acd05f9247b49badf6a6a9d58782018e05175e2ecf782aec519e4d083cbc4ea;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a8dd85146c66b2e7262c645149890ef348b015be93bcf20f45c5cd9cacfb40376723ea5db0b2f38a07e2e6681d4e8d83ba91c5f0baf4ad4696dc84ac1cee00dad12e7a14b82fcc0a4199cf8ddb27;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h84738dc773880ea301519203604ef24a089b5e6a664c6624052e7ee13024e9e18ee139f663280e0e47df2d8c1959f465593f094b0468d407243a37761fe0ac6e338ee86398f56aa131d440ba42bb;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1fa91db81f2f5f89715b83032b15368eb53cd77dcf1d88924aa0d3fd55d135ad19e7119a72328e0c091bdac61b919d2917b7ff6bc8db8b775633af47ce79e6a52eab241020059f7ea86c1783647ce;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d73666e19a9f6f759ec2a6937e1167d4e32c43cd001884a17b87f8653b372397e9e28e9b983e3ebcd5926ac473387a017e270145f8f3be86dfbe4a2f0338bea76aafbac5f23241c7c71198a59622;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf481f0f72b597820e8ecd2b384c1dda50b4e4fc3b673d51dfa06dfff1b63f3e1e6cc1c5b95f478bee350d169dbc5b58fc3a32e0a5f2110f9d2a9cba947df8367a3e8dc1370c5d1168e3a6d26968f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c5c380ed0782fb42d6db1143b6ae2dcea422be45e3e259a0f883c7408518db3f02931a1b85397278d49e229d3f3811efc9c82d7f03d7482fe359f851d7b90bdc900843790fd2afbb2f138dcd2b2b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h34f8141f179d5f4e1cb332d4fc1d03028d4b643a0ada992bccdeec0cb99315690d99dea208ea0d55ae7f7af87f3b45761f6b06c268fb5e5ef3572e1d5cd681366d1c39c85f3f2e9de4ad90a4aa59;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h3c6de46ccc263e01e522cfced0e5bc7ca6904eb71cd420bf41ea7501ff16d73ce12bfeeae2987e8808a96c3a59761699b709105364af33256bdcaba4ce379c4cfc86457272bc89b5a477ba014758;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb2d50ca012cb39f0434aa0b158c4d3a5834c2d286d95fb3c1bc6121a00451cb02292b44eaae36a5268e2fc8f45dc1a5db0f358ba8de8d6763c2d214ad042be37b3396ec06f8c8d2b1175913ffa94;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc46c180f6b0b30aded2a91a2a2b1ad15983c2f0c384e213aa869d35899fcacafded6145bd548225fc56be6a966183a2d57417f480f4ad4e3b5001a681b0074a482a5e1bc9b4c3350eceb831fba78;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h80011526b4127fcaa04acc101db776dd612da3d8f4bbc13ccc61b70b45b07a9e088987feeb36511d53a63135701e6a1d5a149dc5264b95b14862ca52c0b2a6aa82b420442b95d90abf0598e6960f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1dddde89c122a643d49ebe2190fb09cf72b7e44ad868d29212ff81f81534294ae41dba03c066376938e563fc36a3dc3ec43b961b69e884b43787dffd8fb13a2981dfdba2b91a14d8f9ed9ced3b16c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf5011c85a393433defa9104a99f6dcf67dd3d1a56af605ce1c448ae69fdf51091e1a6982fdb217faa82d12bf3268b9736264c107ea04611a5711b7a3739f3288c9f86a14a312d6fdf4883f2dbe69;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h469b2f9d71f72887dd450a7b982dd8c74a6d3dbb3ec475aab59985efa92b3bea6f024606131827035a9ae12819471b209e4e5e59744a3b370b2aa185c2ed5aca572afa3a5c98e734ffb90be8cff9;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hfb82ae8de686d6d62bfd52fdfe278f263c7badb7c1fab6d8aaf858e498a1e545ab526313b5b662d0b26221eb0b17160c7a7fc2c32817c2b2c5ad8ef398bfe3649d458085175f763b9ff5c08eadf8;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h82c374c8da5b52f5c8e41d8bbee2a1a45851f2e869efe3c8071a59bcb024cd1f0bbe14048fa425e5f31f0a7ae15463109bf3d4e929e88e33dffd63bb7bba9ddc1a6e54194df69bf362a7bd5965d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1315ffd419b90848ef3700ec5d9eae9415a53fd79c2151476eeb8202cd7c1977929ee25915e5a6cc7aedfebf68eb885ba2cf73505a63ff2cedc7ec47b16739be5ec49bcd44f1b46df4ecf6fd9805;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd1895273230573224ddbef97dadde04a8a6b9bc071f8f3db2090d9dcfb2ccff2de64614fdc0d2fd17f537d03c1d03bf4a7c4b1b6d4d89fed5c1dfcab42522c88546bcd5f0b4227cccf1329fdbc64;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h117fa43a958770fc2f6f718016cc221ff5097b66166eb3a8666a136e557a7fa165c7fd281fa7938ea8f92dc8ecee4435d360169d05644d1aa8da7acf5c9ac36aabc442bcda2a95ac090cd1d9fc12e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f9ea9b62367b7d5bb7de43ae757f8d55e2fd321d71b2bf1a2b72d0a7f6becbb9dff4d322c8b074fc55a783001cfac6c667b2a7a012dffefc67e848aeefc84deb09de13c6f815065d19cb61ddee9c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h12dbcd901c3b4d3a11511e0038b2ad066591ca9ded189645da58b984e3fe9940f8b09ac0e863eda2b33576d2c087d5b9e6702c3884566dde2e64ffb8835de782b1829ceb7a66bb890f2418d0b8ffa;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h19ceb2c0807b0203711ae3067181aff961300aefc07127f097a624abca21a657f2d35abf2f031f650ce194f1c94d846b832c661a94a102d2c82fb47f3a66780338ddc4ef8f178e98e67e373304e8a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h15e6139836ac2cec0917236cd1d99455b785f7d16ef97380b9aba3cb49e2c25d06c78dd4538d4af176db6e5d8172442bd30e26c799e3fb6e7eb9ef5c64cb0e0c4c9f7ebc35244d55d9f99c703f12c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h83e6470d21001377ddd407449e3d2922287543ef9c694b4a1577352b8c982be12c065ba9f7a0787d22bcd1105a61ad40a95900f5faba1b68921944756d196c167fec0e638592fd7adf1c3d040983;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hefdc1118f12550746424046f667c48ae1cb2b7e2fa35bb8cdb335e241cf18033c49672f5690d76778e31a85970671736121127fd2a8794c485c5c7b9af126804dbfc6cbfa67721cc8c79c505962a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h958b564c17696ed2fd270d175f07d12efabb2cbab3154c8c594ef4a4443ba0e1e88d13f8b33ff672968d3ee1b96f288559446a1a15775d045a56f4edf0193cfaff78c57205f8c513856032903d1;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h167a7af566f0ac45db35c10ab5b3d5ada8fbcf07ab8c89ee65d25fd13f84351c160b234477ca4b268e210ecc47fe4a2e5c5fbb6d97ca110769ca66d62e4b64f9dfcf6f1964d2e4927f3ec167c8f30;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h154ec23c74a9af5078d62a6f5f17704a44d0fe00a2d5e80f606cc00767ab761eb26a8eafc730649e91e99ffbadd745b8a2b652eda32f6d34384fb479ec8f5d14bd87654ecf34c09e6fbea4c60551d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b029a0e6c7798c9bbdaa70da9687a08841347355dab9ec6713beb15bbabc1cc3f1973439c3fb744347787430af2579128a7d33a050a28a518a7486d30e2d28947f179255f6596686b08294787852;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h187ac3df8163166f34d5476ffa30bb212f6d52e4311a0ef0fafd37a000f0a234978edd6ae73446c25e4824167131030897156573b573f2e27debd3cc2a69005c13fd82c4192796a6ebd9962386c51;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hee8d1e509e0c8100f641a7a7517ccb098264f52db3c20cef55bd1dbbcebc0a25d6bf3347dafed53412310698c14f20f4401cc64ee1c48d51a1b44a2bb875f5bdad1c2686d24926f0817add79f234;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hff3c6f8ef731ce5b6c98dfb35e60588086b0119a9ac9f790f60b44feb134a33dcf5c9a52e44653a44c896802bc333a114814cf143ae05fe6315a176e04c3b7df4b60aa953cf85e568a3bffd0f0a7;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1cd8a528325a29e4f6d4cd76b2b185b42bd16b7f9883e8afa462ad7c2c810c8c163faa11ab00599b7951cc8af4dc6d5c161ee3e1198d3646e36f63cceefc1da22ba14d3262465495fdefe1ba5b74e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h166f0ba3864cba65a9f33b1e217fded0c540a4ca045aaec5ebd9b7b0efbc6873a24d8b32cfcb7f33569cf02311bacea282d26be3a4f3ada0fbdf77ad2d3722ede83ffa1bf78ccf137523ac60fbed0;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc8d5c1c41a5b09436f09d56d9d46ffc1ad550620a92fad0d8e550097118abbb7bb176fb2bac7b990e4f523ff7d7b08c50d945945eaefef349dbe80987c5778b48beb5d62f4174815158471275ffe;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hfbff7b1f21a36856bca5e2a5057a24b6d63702734118a2fdb7454c36100f9854dbc67020c97e2435fe6d711984c1be911ff8299bcc20886e180f13c4428dca5504cb096c6e7af4e5eeeee2dc982e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1cb8aa9b48de5ec740db8e9680e583fbac347009383a5db74fdce4c820b89d2557ae98a401ac9b334c7fc3788b075b53e431c6ed12409065773e0aceb48ba03c819039a77571845f54cdfba66bd8c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hbc5eb8e58f3b878040d99abdb323cd2e00e891926b966528c3db8150fe5e08a347dadb393b757f6f2660e49a92f61506cdbcc7c67fcd8306dca451fce33e57df430c9ef346cee9bb4694f1102e3f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b82a389ddb9c7297532a62320ce5c5650c39a19ac688c8cf24e6f989f632ed8192362c65ef45a48a581a3a624c8daebd532c39515d0c8333be7fa7b43fcb92d980a06e3e6b8af13324c7aeea0550;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb0dbdafbc2a56ebb60d31853601ebeaa693a8bdaf31f7c7e0acc1b50cfab83d348a7211b8a5d1ba113fb2b28ac389ee7b06f4b106e2e761692d1c7da521f9acab88fb58e91365d9bd677efdf0c90;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1728432b23e38a8305d44badb83889d0f13af95664c6450e2298355d51b2389fa4a68a4aeed4cd140be6d001abbe31f8e61f8a3d017c280e0930fb642e552e5de2ec7723c27c0e1954a61c18b910a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h11ea9688be7dbf26887f0242e739eda1315ff1bd560180b89c3bfe8f7f38c75074c0cdf5edc2bd03e783490c9a6b5ef61c634d19459b4bc452d5ae9b656fdeb7677b4959c7e6c5a819224575b7f26;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h234bb8624ab9f216bab14b1806178e2a43220160fa78c99505269c8ffe069c215171d652118e91aab176d6e163e7686cc3a1882632e016f730d3a325bf37cd341d8b161dc110f830aeb12b3d07e0;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h19716da712542f493d52fdd97e3f7f197e327608328deab77b75adb3878be424fce505379c0433a95b1642152d0f475ee8b788fcaa1a95bd0133453e263838da57547542b920f2920ae3c29e0c0d8;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h4ba7e649bb1701cecd9e9c9411ab437724c5ff6e059c38d100d7f00d703c2c4fdc4bfd17a23043425a33929a94923512143f526364d7174a99895071bf7fdd3e905f1c05cc7aceb1e5ab6cc4e438;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b1b33417c061d6eb2cb17ef8dd171bf82a3e3c5f0c04e5b0c925b68f1bdfaaddd7143bf2256638f8a48496621ad5c27e4016acd70a73ef98baaea6130eaf0ea15038aa5ffbb3aabd1a7d14b95361;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d3ad5aa78f6be6b704fce01d3a3a0566bbe3e4083ea51b2168f9b5dcaf2f2b8e4402e7d2fe871e2b41c79851df4428c4a1075e825035530a6a3ba8554450219bf81e52935420cf65d03857ec5a0c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hcddeee8c55fa9d8e29c8ec46988c2e15cb7409d8ac04058e24c558156b27961b2475388dfb325d9cb1ce94353dd2a96044944f72a7b881fdf470b0de8c3c2a3e2f65fc2eb29089ed396680cc969e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16fa132b8ed46fdd99c8676ac06d18fa5d459d14034276d73043e93b553b4c7aad3ea8b83e21481531aa6335dabbd628d1387df7fde50605fbca94fbd45adc1cb9dedad3aee584991b35bc693f1f2;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h661a167778301a0d0d8e76edf17d0ca2e9ac880474e757eda8fea1d03bcbc1ab17bab81b297ef48ffa64b66a616fc35b519a242cf72ab2c12e8e7255aa3c6d233061502bfaf31a417d9da587d896;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h351fbd336631a51eaccebea95ee18b83f4214a932d81b7805f9d50bd760ea7df96fa932db48f4c12a261330e9b03812269994f2963163811203411159a59de9dd10ad373de4d5930ce9791d23e16;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h703ac42903e0622fe1d81e71568adeaf6fd19cf9fc41b5457a9bcc21e8de5a1f49fb38dbb7db721d4627a76e675207838c57a1c6be6e731ccd0f4bcb20c782568be88648f8c79181bba22ebb3565;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h49ff74493c5811d3646e0ebaf47ecce44dd7477b365f4f8a428d8aff8fc6567f16082f877db22a8c1e8782bf1c945130d0fb5cdb433b41dc68e2b27f90e5117bd5a98797540613e7465345b5570c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1bf88eb0b15486037078a72fa6912ba7412b841063ad3e2109945c32225fc93f3e971a67fa36476f66d02ccfd1462d6e7f1e0ae2c7f80374db4d70c88fb7c983ff01acd252097c846d80e096e481f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h14707570a2a4f919c4bebcb8d7aaa5f91a8df72cbfea4256a8b309a9deeaa63c9cf2a6601801d3ad36f0db472703f7751959a95023a8c5ac6f1925a7921050b4a900c667cd0d1050f56898c687d4b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h19ef08e9a4180a86bd98138982645fd1faa047b4af6936a2b36d08571ce958aabb5518e57998fb26696ce8372aafd2414a372b74c381d90374f16414ae6fedfa49136236d3d5bd22b0897b2dda8be;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h2962dc95610d314052e5270c6746adf5533dc68a25f76f078185c55ae3f1428c3b938ed6a800f541e570e48f5c358dba9544dcee78833a2b03afb948e007120cdabfec605dc3cc272459e5ed60ef;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h63d0415d6620858396f5c14b40c303fa888f1d2277c9b6e3f3ecddf983d9e73ac9dd0bc12e0fa67eae75ef1eec4e0ab7f96cfc1c4ecb0fa25535f7b0b0a7921381cfdf89a79ee07706c0b0d214f0;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1788e5ce8409c6455efa1e99c574861d5db98434da0dd26a0515df2323aafbd055dba4f5ed761d2f293f0aa7dba5455198815365cbb4539d9c6aa449f7843862d2dd98539583758738400e0f50f16;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd84b4abe4e98814469c041d25b75f674b8da1e5e5ce168f1fa0f2814c522979275bef75b1e4058288642eb913909730832acb6eb53cdb5987bb305bed979e565d92d57b321a27587ac308a5b12c3;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb3398869ddb5f80d03e92b25b0f7ec78247d64d901b8412e0fc7b7120e459b9dd67baf7f29074e18f01e53789db3832a166ed681a9e952114566d79e73b3b0477fa5c5fccbfb76569ab66d8b7f1b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h18431d37ee881c9ad73d5b4992b5b74bf775b90ed5462e3b89ee14bb6e0442d4466d8f6be740548b580a52d2f4b498844eec968aab576927c1a7bb2900c206e3bf065bed1c1e661333ca1aa38a13d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf99416558a6aa7dc1dfa70cf8e6cac9e7fce8dc2af78e17f8692f03f6769a9b405717f533367578d55bb93f94beb016b69d61e1293bf4a1078ab30d899fff479987de0b2af517623f37fcef102d9;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h114b7220dd7755c8ab0e38e54ea93bc2af18a17133f2f05f0863f7d88d80de57e5986aa6806004e6282c596291f854a9b954092f8a78fbb832a201caad2c5d38d49658a890da5a0baf6c7d2cc92e7;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hbfe685845acb5ac0323bc24a3bef6593cffb7c3e76abce78d40f15ec78ac084baa51814ae72c6fa2404eee5f78e7b9ad8f9d7c3625c425a75aa64bd2975f1cef2bb751bd4941ac608fc8703f063e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1126d45d303bf47a60f84135343ad6cd0027c0e6d5cf5c138460acc581173d6efb3d10eb7fa02c3d7b1bccb757c53b4d5a6c19201220cbe885f0f577f8b7d54288d8eca4e3eb75dcb67629fba1131;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h19b0574e080b9ac1a4914680bf918ef07c7734802a708b58f8286e4678f97be3e291b3383af2ef7ed34b15f813855ac4c8f7a5947cf8046265b3f12be9902c9624ad290320f2c8300d2c978000f9e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h6053629e216c414a9e4261e7e07a203dd95b22b2f6d55f2b672aed4d429df612263a1298dba236e5b4bbd38149db218d858db0cdbd595875d7c721b13c091e3b188b29ab841d5516ac01d71b11bd;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h5a4c898a30fc5df0df7cc96b8d4616ccc2571356f5a8b5013c756f2962b93910c5382d5f3296653bf8bca2cf55c3392b944eb46a3a761191133f0ab7c95e4a5d3efa39c70163a66dae5489a560a0;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h8023914f6ff5f599cbaf54eeea4fc36ecce4db4705c7f518a1c779daa4e1bf4bd6e195e3c463fc1edec452a990f0e0b55d48580b892de02f73923e8525cf6ee515da3583d622b3ffb5ab3e7c8765;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h18a4d1de956cead4dc388e7e4f99cede5f2f64d08e5a855e0e24840935d2409d2201a51f63d30b94210a53990c1a4842c6c1711f66587a63eec5035089449ca8d11a1bd75278b98e0686f46091ea8;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h4dc548a93dc396c990ffe1c6866293b4428764c0f3c63c278dff1e881541c01afb07845711bc967c3190f4241185c187e19032d7da0f9e8dc1b4b24114213b21aef01ad2a3b5dadf65df9059ea1f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10d2400134470fc88522e2a6b89f1c1d6f7ceb873a06448b4762d168d44a7a62a8b801a2efd96f8ca85f8a2449750bcd0a042ce6418b8a3e0d8025cbd8097501e1d479839d3bc7813abb97d320021;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h101f4de86e142283ee6eb7d9172a7f6c32f4198a30c68b3a35ba37c21ffffc111cb48efeaf0b52329fea185be43850c3d3440cf00142362cac6061bb1638f4c92b3d5e6b5dbeb0b0a92812531d1d1;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16a8cfb808b2978849c2dc62fb43d41ecfa88e2a4032ce4d7bc23d864557a97da2b43eaa9978724085cc4018be93ac0c72beb136402f0904efee0b91b08f0d0e1488cacb273ff2e311a744cd0ed81;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h4b9d7403a652c80673ebf23081dc4d72c4fb487ad8f3ff6d54834cbb7e34354211e87189b452632b8ba9e1a18e4b515adf0a01386d98d5176fc6dd851eab8564b77efd00f51aa5bb17a9d262cdbb;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d8fd90f8806aedc793996e77ad8b506dcecfc1ba3d57eaaff44a66cab34be22b4b609820629e8e1857f355b843ec36891d3da58b8fce1a10c58f22c03dee6eb101eb4b7a6cfbf94c635ff8f31384;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h17bc1abab7ff902a40b91bfa9c742d84207909562ccecbfefb84e9bb58964f51fe02223d8550092c56166cf71455ad5683a837435b1a3d251d4ee12671331b3258f56a753ec8788c2ebdea47f506e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1248be8cba526d84c1909e86f9fa0caf5df61334abb6140048d1626869d1233af8a6b8c1d51dd73f4c1dbd5a064b969339efe557314f6107710ddf082ff066dfd7945ae5f7c55f04bb8eaa4e9faa9;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hed9fcf9122e9b20e75f5c55ed37b5ff1d66f9239553fc2a6a518c702ac3b3fe14e45c9d5ca8919505930cc114379acbe98c7a162ef0641789ed4970435cc7910f91684af094efc81dd62c131e091;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d0ae17440fd38561c3386c55fa0bc2e62d4742453e4c58ad14767f1e77a858a8a192394a91339089d8eaf745deb046c38154056eed51e5ecf1e915bd0fe511d446c74311f4747c90ea15237c9f67;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h18a4ca6058bd800581c2b87f08aa3a46df27db2a6d0066f902bfb9dd784a529293e600891d81df2b2c583438e5c1cd9ba32bd28895adceef232989f3d28140a39c82eff690a585063dca30cef137f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hcb4ef2ec49c84a8758bc16612928305b3e92d3968ff689cd171521dc3004365dae938bf6d5c6890ab03dbd85033ad4a78986d4c8521279f8ff708b9fb73f9a5d38578e946abfb699ee50e45ae5f7;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1161bedc6e698a6b20083b24b49ae9eb4d82b3c3bba853c428c4adca5c5538ac3cf6ae3031443918c3f7c20f7158b708cf97dca3d12215785dbb0c577d0da55975f455ed839bd656c9a7401bd668;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h96e0859921e597e60c95a4e7eea31f968ec5cb40022f67a959b12594d3aee2216c9ea0bf5742c1bad3761d376f688239414925ab32b94ab175e1d68858f2032049388b50332b6c2b60c5a322bcdd;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hbaf71d71ee82d554f417ca9947d1515cebdfe34fc9b2c7408c6f1a50ab137502f842c46105d3d26fa5720bff3813f0e79f5b86e45c0624926e846a1b4e3d3157c568e3edba86c58dc39423049c39;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h8cbd778300f925b807a56ddd6e317a2c4684e1b68579b17d8b5f5c2b2964994265d371fa969fa20977e8ecfce86b96c3c7f5b2259f0c996fb65d82a266f3f0579701703f539af3c8c86c940f32c8;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1efbc8d83a3891838776028385c1e04b082a6808dd7c59b9c248627f4cea8eb12e76aeb15924f718c96537b7c2b7d3437be71316f4ac73f5b48e79c55b7887788a42183ca9b7c734ff80e57d6abd3;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h7a3a4ee8be64be0cdb5ce9906a49ff0e7581bb5df4939fd246d0657d9c365bd8807c247db91ca865b45b2306ee5775aeb77e625ff0fabf01054024679929f01a2f5f4c80c4a5152c7b0e4b04475a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b0ac2969a2787f607a6fd036aa5cb5ba641a74e4c586662f58dfcfc367effa967fe3fd23931d8f983bf6e5e042b31c950408d94dc7ac3d634a2ea27028d16ff1fb3d430086b6199fdec0a0be0091;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc410d2a102bcf7c35054bff1c5f49e70f8da897c89ac71ba270c8b97755fe4c7eb067b3c333da424958f163db36e12d0eda5d2718a137dde160e24e85cd377351cb361e55c24fc1f9a08d526dc0c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h753e2580f871ffe4d628bbe12f31b27b77722b86b6d8825cabebd5b7501a63426260ceb6cc9a734f415117e14918d9d48e2532e2573380d2d6b37f84d549d594598f364277b7c85da77d492ed1fe;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1be76c22c865a2e8814c757a4d03c21f9a141b56a787b5fec66ce85a24a2b3b0fba049b9e636f5e0c40f67e43c75b2ecf45f3d52e10534274a2d676a28ad9906f0ea6e63598b189aec9f73915181c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b47604085cf9c51dff7610a8c5ec539e9575013ceb712ee830983387143a0fd641eaf58ad3bd222c437ad32588296d984a8314c76ad9f0bf2c4c3a1a97610626c7bae70adedfa527f66e70bc6ec;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h6ef324c1ca0d239d949db4f880c37476965bcf16309e111ca306eb03a431e62644697b3280da03880455ca18c3bf440e5ea24d45f4f090812d1a83ad8fde57d484c07f382930b595fd8523b129ce;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h6e29b63061e9ff60f95188ca105bd00b06f5b4ff3a2e29af291650f58378f65be35327d064ba36c3b4d91b600a73be049d59d69a6274e574820ef36b37f4f522724539e03a9a32510c3d9c851669;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1dfc42d3630f8ee38f766c0878cbf13e8b10486e833576d5d1fbef6b20b8a839539b42442b9fb0a95b3a49e8994fcd88772a10bfc95ed942c1b40fb55935cdc18bce691d2720892226e5469c16219;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d7b406219d3474a7b002dc7afca8c3adf96ad52307e4ebc686ac2c68ecb7d0fe68b583b6fb66ed6aae01db00ff85acfb8786e08701ceedcf7e1bd0e102c0a0052ff36767e1ae05f5e3c22f16647d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1bfec8c25a79970c2f392e451aed996b2d5d46208c79a6c8cfd08e057167f620431c0a9ef1095a8a48621bf94308a9f9ee6b145e5bffd7176a5672f921bd8bff358c132c2098bc3c73d35492ebd08;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h4fb40791bee2b96014aa190737e34318698498e92e47b98515ae169b86f3016969acbc4aaa6779984a7d02c13edba221132bff02914d065af7f9df3ab79567c02b98bad56474ab633d4a0da4059;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h12aca834220247589fa34da068972973c58ecf513e191c348d49687c686ede6054006a05e1403858bc0e80d5ca559b17a3c630cc4cd663d4c3ba5253648a9ca57c6a5b74fc7a8b8a88d0908e706a2;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f8023efeb7e116fe7377109b2cc2f4a1b3fa2662b2f7cf7e7a82a9d878a94dfde75dab652c381a016eeea251efc8f5abbdd93bdd4aa778c55ebeea7050b127aa94701e7f7407d68f37e588e409b4;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h15e4bb6b2e80e7a07b9decab82063703f1886de963dcfa25ad86a2766a1555a391b565edb845d07d399d3dc87038f6675531a34a3987a67fb53895e05677bbac3948020763e422c2f495b2a238966;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1337d430895915be41d84f96deaa478077fa80dbe005c035bffcf74ae6dcfc4f99a94c768d70b3cc3eb276f33eedc8bdbfaaf9b476352fd64849a4641e4162f340d50945720670b0ea535f19eabc2;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h2126184b914aad277ddd6a98c52ec6654581bceca4c94a8f497b01a4b973be2f4a6d99bcf12badbec741a97717ee84d88bfd29778639ee1288d7d66385f596b669454d5fb99a64609226d5c93631;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1073a2f92866f7dce745dbbc22343b18b9c86e4382e64e41c0395b93386eb33f83f4bf2e94c347b5572e005896d99785f02cbed2cce02aa8006658fa8ee2601967271685b993e9a68937d74f353ad;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1cd7f8a4299521e02c31cf5aa49a83bbde474e51cfac2e3328230db2a8d5836ac623cf91b6c74a9adb5514861b293be13f0416c9e9f5344b88ea70e9555be305d3432060ccd676cbcb245e37b0b5e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hfe9b2c580b56f3ce0a894c8e554e5520c14b94b8ccdf1c31081b0121acd719e35c8b247d18adcd9624d7ec1ad4cd7bb53fa49ece042089fdac28176b447f659143fc7603e1197474f34ffc8467fe;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hfba5d9f89c6b191d92ca42caec1b0eb2ec8e5f4b0b9ac6fb6666cebe9364ec0485be13f04a49bfd447826f2913f6495ec8a6725db29f46c8acec83f5507de635c9035fd9ba8bf535cbb0c53a169c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1284f0342fb29e7a97db491fe6713212c0d3652b45368cd1e49714c4c4a49044f51f1cd0001125b05405fe11426a1617cff81cf51e0102c5655ed023de23e4782f0f791783048e1018010abaed15c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e13d0ff71da370a42b0473663dc49ddb682279191a0ff408413a09f9a39a5a365574922133b8bd33f3d68c54a5824c3787f1c1deae992b9a48ad6e0910a0473d52c2ffdb7072e01bfee16fb6b97f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h142dc450b0f3764f6160b20372aa4cda0d60efe0578b6b5572fffd03e35b1200dc7b905da82a54b1984cf656c7b95e0ef2de25d4e6a8a5d3851114c9e9ce8a2b7b67ed2b98213bf29f53ae50dfc4c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hbf240e7111371d9e4ea7de4f76b42913c65be669f08923c89962a408c31adcfc43cbe6b6eef0f5f9db3227a1eb13b429a2d20155c3166efe4657b3a0d5be5a1be96165084f3deed60b4cde4cf915;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h11a8b08393839f41d6c960435e7a553ee71e8d6681b662c8e30a05bc78a060c735a3f6d4d34e48739bb8f5167d711e1dac3f9e88e46efd2424c675ee6a4e6bd1648e9368e0303018a5c707236a14f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h146eba5498a599055e7792baad8d3901ad304766ddd9d6b548768899a046006b780fbab93076a3b1579b2b78de17d6a0228282926164d51637395491d983ad22ca882650a9c1b1cc6d8c24bfd936f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h14f7d9c8baa9d1ef7629782fcaa6945a42a3656b9e26dca05119066186d556e9b4232293e0eeaba2c5bdd9ffd412565d83b42d448841635ea64ead159590565d0865f3676ef177f71a9eef3a1958c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h6142638f212f602315c78f90dd626726d32127fcd7b5fa06de82044b472b1d91d5f3abc0876761d02f542135ebb788d90c5645c0be9250c7db9554b4ac85752709c256cd39b731b1114d8fe6f96;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h4f9efbc825a71cb118e025e9f7a5d8c0d57aa6eca5d0c79c42bb29e9a255667c86ab84423145cafbc237195f07b7e31c69d6f765ce36bc14eb49c0d02ae65fab36f060bb783844c10bc415cdc628;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h13f888b692838e91af0a4f7a5736677c05a1c22a08959aa1e9621abbe21e43016c1e237ab8fb57d03f8c9a9a91f7bde3c341da564ec65667ba4d96ed176f48661ef2c311d8985b9a3d56302cc1f81;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha173c40ad00cb7cb4a8a4f383f854bb38c8f5f258d196e6f08300cebbbb3005d0dbb78446258c21577acac4ec4d2d995ce5c1333ef47d13c2bcfd279e565d8d70d76dd56d58d7d18ec2171d926a1;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h6a833b4891831aabc4b302628298f56982eb5a0e7cf2b2847e0dd13b2368df7d0e1b7af4532879497dc280176c580142368d94cd132198251398de852b56e652299543656e13c29e7548b4849a80;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1892668fcdc23baebd7ee9763b2c53fbd6ff3f2d7af38a70a7c9f9e4afc123f1190fb028daa25ae6a4950d967a7c9b63ab831eba00a8856bcb458b089d1272ee462ae2e062fb8358175174e223204;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1387a718763405ced17f61cebf538974a93e650da744bb1a60c5714ede04d8dbc953596f1c379943a2c27bf7c4ff521860b4941b55e4fbcfcdfb66789a8a2a023276a832b19ba4021baaddb1c689;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1aa95495cfe030792479b4f1be50e44700070fe4cfa348a601d0abcf85a5406c4c2c17bdfd82bde948566d400064740bd1dd15a37336d5d0e324a56d22cba00de11c76dfb8ae52825f912f6e30040;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10ce6a781402fdf3aff1336fd40775abf6bac93011aa750531c2626131c7464cdb0fbf37bd89ede382e04286675ff54b7c388263ed2f1825601cb393b1ff37f66e9637eeb0539c1a251857592df8b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h15ce4e87eb4232ba456104a35459b7cfa64dc9578c2872cb82cb157bad457aa2625407386549419ae7591b0372c3d999960fbd2771ea7a02c6e73c111f136b6636944bfecf7cba7b389e502af99b8;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1cacab59485f3e51df3c3441afe1b02482b450836778c64130ea00e33b6ae7ca0c8e516550e243652071080dcf3d8490677710a3ba3578e92aeee1fd3357af20770c13d0f57c39321e35b27cbcc0;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16a33126721ccdbcbd45c10593d9db8b7c93b1a1f4df6dd4e2b998bc91d0ff007d71d7d29d5d9a160f0b887c8517d7f2f10de3192254cb46b9f25064bb4e746bdf0237f0bec646c7335e5a7bc8b12;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h158753807c56f37f7274561c49cb464fafc9144e55a58ffd1ce7e8272dfc0657d966aa04b1a2452cec9c7360c8cc0985589ec8754cfe132dbfe330b179f0e99a0aaa3d24bbe3a048ed479cee7d95b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h12eb607aee62253eb54e8d3c5d66db03b2adac037cadb931c3af7ab53d5237f7e2c3de5be2ed847ea26bfc8b8301f77ade2bce820f573dbba116e974263648c8f2b37d2e61848003af0d01c50f227;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1015f2a68e3b3fbea8fae0239a923d8e8e981a6b4f774bb69e54a10b5890ff7679cc4f19a6afb939743b7c96c5e1b44204a1a0345cffe2975dcc458b4af5d79cfa627895860a5a94ef6b1ede94640;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf1de77829e9372257d3b95e1dd19f2b0628aebc5fc2eb4a40f131a20db9c1dd135ec10c32cef13913b8975b7b61594c190ed7f26e226eca20864a51afb3e942ddf01832c9be00d031bc17faf2d8e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb12fda51ecbeba825ae678dd54c4608866e88c006be5ba366fad2dfb749df236e06cc46d7578efa5270d249bca4e007ba2ac4eb48eedfe25d697e894d95d33c25fc2d6c375901c0a12258672120a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he88e88cdc3ccf8788575c6a0caa7c80ce04620bf3486c5ebe104e21d08cb07ec8cbf9e5a9db040c2e216d730cdd2896103835dab1953f44fee3a6eb2523df7cf27f7acd74da42b639c7c71d952e3;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h14f5991d661af7ed0002d1ad6f7f5bb574733a5aac255f5dabab4db99acd2bf50a4720621cbd13608e8d0a66af653db722cc08b5bce787c51436bedc4d866dadd7f64617861f7ebcf8a23b56572ea;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1159e6fb03a92cf94de8d5cfe0c2cbadb76e486d2b70d1f680d03992eba7e292813c361de5acb5d1eb87164d3d763b122f3e06af03891193026aa9ff59520b605ae6bd872ca9cc714a08d164af682;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16e63ab444ecede251a51c0290ec2e7ce72baf0ecc50c98357f375cd2428ba987e497c81d567784ff5315a29b477c644f5aece9dccf121c2c78ff07eb22bfd8625435e2340ef2e1bd892a729d1dba;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h825e7057d232b3e6474bf53f2bcdfda5ad512fab2892a136d266a1b5fc1341a239c801abc4c2e5caccb2068cf4ab5ead94c6b055b6e30971f7bdd390792b7dbd46629b8aa498f40dede71eca006e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h90b11a12811231b6797d810e9589b18f5f9229361dcf643b1022ec7709b42c3575bdbefdd2aa76fca6a4511001fe5ec0ba17c3fd445e0f6001e4326d3c34260e04a16cdad1dc3ab93ed61d07dcd4;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc083756b23aa14fa035646302c77e31dd570c59095d4f12d02446f35cff1cd1e616cd3e16b9910f3fa095934b81d96f3288d9dfef89f810a22e35a9f9b941affbd3b4b05e75ebde0addbc9b9bea9;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hfb6b8b5e9e5a90dce0ca0f10f9333f1e11a1ac1a8b52b6a1f9ec65e7d34c5b2108b1dc76689c80d2bf58e6d22b53b7a3850b2a91276eb49f28979b868412fce8204e226849d813ba85b15414924;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1141bfa28987ddc7e1e1b8131dcf8f33b00efa652380eb204cda3e4fb7c8b5e7624041b269d645b646eed8a445d1f1f3ecd87872bfb061dac7bb0b3bfe002876a62fdb8aa6e061307099971bb7701;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1da706eb23ab7473334ad7c5250584a1b36eb85edec49149016b9c62c231b2380ef52f041825a99b4583189eee787370bb078d35ff7361f8c8cdec579d1d0f0ec6687ff41a3985ba051dd6f1621ba;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f5b433981b8179496cad21bbc4db95e4a899d57060d876442ef4340ce7d9b8b583bcfa28c78183676e67d16a70e4d3bf60354fd245529d4a6754d40834dc5dbd0a463cf29097237d53344196c42c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h91c73e0ac9881cf0d72af1ed5956c2bd7386081a768394e3a94c8e789c52176c37e4a8b4fed5e68abca11143fb51752fc2d56e7051e9469c320e24c023d94062cc90df691c4ee8a25f19e618097c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h788dcb8d1f101451b5fab5e0d9ff85e709d2b00224a59fe5354063b9c08bcaafb288b7ea4c7a377ba924baa6e6fde784d5428bc449b3e0fa57a2e067e16e3c15dd1cfde07c60cd5975cc0116ffc4;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h19decc6542111fffd0a370d492fe7daeb126c9e30580a7c53ebd6e3b3a31e511bfe8b6eb3e4cbe4f4220f2d363c5085589fc8e8e52d54c1e2bf65dfb046a9d1c5f619348e4de0ad9a6dcbe4fc8911;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hdd84311c182fe569a4f6cba251298b5e19e830df0cc19dd96538f25f515ca093945f2516091e1f9669d34e781c0da427664aa8fdcefc14c49693b7ca5dbf83e0a977f05f25eee1dbe071c3cb0933;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1640345eddde8aa047792b7daaf327241add10fb5c0ccf6fd4bfc2e0807f414dedad687d404a92ce0501154a0a91fba3b771562a06645fabca2c1f0e35663feb51bd92e1a07efa77f2a36290a72ab;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf9d739f2d0b2bc8275c77e61c32ec2f0fbe0a87c5121f428afdb83755af7df776607514c68acc6f7b71223e6882151c4bed77555c1736dbefd8e31ad7ca6c441645433f5d3fb8db47795e6db305c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h664e67cc02bc8dab0fc8b219e932909a2272222aeba14198d461feb5ef083d4c64c440f18b1fc51b94b0c0d9f73812c376c6731da2a621158321b37a20b64f84176efd5a405372d230ad4afcdc1a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f25e1de85eb9bcea9169b3975a0c4a7c5951381bd21de33b928e2a53753296a1e6f143cb866e300e72a309f1032c2e0b769d2a219cbad664ada167ada81f99c27706cde8e3d9f9e00cb5ee72eca5;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ca684ac9090ed6a59396be7430ab25600388958716627f83f632a02f4fcc80e8227def4d4cbed71788dca13f5b5cb0a668fa6b1cb40eda2da426e05eae3e749c8a6705b3a277f59cce93f89602e3;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h170855d281355531e37f09ca1f65f2234bd9e4f551ccd58eda95aa240a2abb51cb4cfb3a71ddeebf7aa0ae020ca002ce9c94bab5445a101509ca68ab72fcaee3ddf6c8bb07e55393d2e04c54387f9;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f349f04070fed3f8b04096855e08e2d9189d57e6324623aae797bd7fad3adb95b638d36dc7e923e176a8c3084960dfb157338edca494e840a7d514a9cbdbc76c9c89ae36e449017085d04e85734c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha03ee34f2d7ba07919247e76f6e58e6c1c9495d09d129d5f5693c24744924d0000d6e8df8ce517f216005e2b134df70122a22db3257d1c7007f6dfc8f6868a3ddec6319080ff4325254ce494fe76;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a217948068b2f8a75201505980bcc40602f1762fc2789fa2542faf866ad665a99aa8d818be377063590c9581148b0b2ba6253198f45fa15a0eebd0e68b855ba91ef2d6b167f3803862213a0ef53d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h31d2ba0923124a4f57e49c95ec58c6983119dd9503a50fd5f36a4767a4ea1817b580b316c69489089c759bd0d06efcbcfb772f8daf7d4fc47a6245df072fc585ec5050fc58d7d1a9bd12903cbb7e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h140a2de1c18302f6f9a00f2242eefaeb8be6f86bd89ccff85248397bf52692cf707d885c51cf2b924a8bfb94b1260b2917cd2ed5875269539ad8b3c00f789ed7ac8c1a5e108051c6f4440e3cda085;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he82a73938793183e236d520044cfe185ac87b44be6175bc6487528c9d77ab27a9ce0aeac25b18513580c46ec184ec30764a9497add14d1ba29478557f62d22a144a1e931c73e0257a8b74fa3dd7f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1675054ab9dc168e49f2c91bc4614b043ee9f9f2694c92fe3b7cfbde8bbf2488e1e00221d228189fee51017e2ede1538b04e0c63f7b6674897243ab4f674e86f1daa51c6eb4da459b8db7b9d35be;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h49b971e37bb84115c2ad34fd1f3b8271124777a97083fa5e3fc4efa0cc06c4c2c4f1f40288c7c4b03becd353056d3539419288e62934dc039a2acbfdc1b604c55b5ef71375ff09eaa3a3beee7fb2;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d85c8f68b04777022a66e2b288ce57e4c91cc4a8ed0cef1db09067f018d94ecf96ee931184e56ba58245dfca2bf7ad3dc53a8863463a173bf9e560381b7d460b80e2166f0f04c9c46e58ae0c190f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h11e6118f35a148a8889c89402ec81b08436449c8935d84f97ea9eb4f01830d36b991c3e64c3b12cb946c0df315751b28357147bd35e16f5ccd59f434949473851da2aff95db239a4786309f847797;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h728ffd4be202c2982333b6986243797c96e5c945c07241848aad8bfeb636da92008db074eec3512f935897d886877dfc766ae8d3244d3025d64f2c66131fbcab7e21b6f709b121cd9ff9cccf2084;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1761340adde588d06575086bf7974b2d0ac6441e29e14f428ab165b66cfb473a7c2195c38be0e2ba407a685bffc14d9d3f99d7fc964983b36f04079553f05249376542d30172cd6786447c5249cea;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h92f82650c521492e705a360ce13e5d03ce02483362b8c6696fa7946f5f020020bdad52df641380550ec51bb6d0ea81befe31b1725cb0ac0b8c0d368b04fbd1ab6c8cb25450ef3a8110c0f64f2486;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a16a5f236f2681ecd20859df663432e7e10c411a99a089055a763e73f41e6cbbfac5e4bca45ac043e09c97bf039002ec493ea0c047d28a6aeb5973740d00d5f50e45c20ded35be670cb1b9db46f7;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h18999ce07a0f6417b7c63e39736c3e581c4770fec9d8567f60dc739f48864ddb243513328ec586dd3f69b8df236ae2f3b2776414a5b0a253fe9498e23ecbe1111ed55ab45997ebfe8bde23e60d62c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b2013d500c07ea0fdb66c4819a3aba42395e74139394cb2970f3aa540af3686b13c30900ab11c5b292cb30c3470d9040b3be9b3bca5dd6c0dc408fce55f6449fdf7a61a10b8e445c8e7fba928a62;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h164aff67c03762e6170945db4747478874b80b48834f869651542ee134150c17e2d444d3d83bf802b747b654784ddc3d874fc93092f4b2a3ef9559e67bd0b0e1922cd00190bde7704f0cbe5f44e50;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h4db82c15172be7868d65310486717b6e8f99e98fdec75811eb32d200f1ba7e014b9a2dd064c6c51ac63dad0c17216ebe404e5548b9474a9fc59ebb25969c748767d3fdac00efac3a5395c50f967f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h18dc6dd48e861ecab9e0b52d530b8271986d54351856e36f9a90fc57ba5a6ffdf6362b944c538f6023d67faa89447c52e000c7866675b6b3af5e45f5f3e262e66b9faa138cd43eceaa199f42234af;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h164e6184a02544a65c4e124928245e884c745e7c236dc901e89fc9b33bde7db6a1f12a2f590cc10ad354bddc8d8137866f0ba6e969c85494adddad2820998d5de3632bb2972ae6b0ab1a3cefef422;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h12f671366cd1ab9c1c387a5558e84d043917f3329a037d1fdb86c25d693266d203a81900a716f3907aed24dd6d6ab5846cd63ebeebc159f3a2f27632c4d9a63ccfbdfafd99fd453cb981a6ee6e1fa;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha618469610acce72bf1cba9902d54293ce19417b1ec27a0e69b6f1500914146e05075d9373b786a437b72e55194e867041d9739a08843c90e0529f5ba1a856df1e6302b46c365949008ad1c98884;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h154ec480e2e683b27bcb537ff4a9887bf6085a1b7234d60de7cb42234914733c5aa04bb7bebcb438cee19b4beea3870fa909d8279aef73d47c86e20f277a146dd518e7cd49d84f6d98832c377d1ac;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b1f7d1a33fad4a3c2f49f36ddbf931167f4ee3776315516555f02a625e5b0ac0598f055c843965556afefed38d4a3d70de81a4e85def683431eea50582a4ff1adad2514521d07310380059580d55;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h3d6006c449100021157620a3ffac36f08467dbca2f5b5d2800f6a7b15724c789fb39027b4c54e6c18ce454a8fecc593d1ce08859fa7283b76091848ba4f3f70361691b99c95ae5281aea3082ddf1;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h171de3182b7e644c54891186181ddb03976dd55f5dd0d6df33ce44f3035fc68c6e7f9619276325b29e06967ae3b123ec13ba15a2524d8d22f7e1326ede891260a1a53d65335f7f516faa2d271788e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hea977eaef7d9eb25a401d960e475cef6a371aef53ad3f2020131466feb9722d1481e9007e4a6b287132b901180bceb9c6f061bda0876eaca02be5a05ebb8f59e4ad01227e7b73a35e394e18cb507;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he032dce22403362729ae9729ed27cdb1f1bd1ce6686f1a0f266f236989c6b95bc4f109f870c71e382884fa273c9950e8ed162762ae20878683946a6e454fb6f365a841eb2be87a72c394af70e662;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he978564fc86c300482dc84288e74d81a80be0a1e37dd2b25eda9f0b6e88b8f3a569cd14a76c38f5504c97ccc739b2756099f8c5e322c31a70aeb43b31bf607ff4fa0be2454507d4f12b0834e5b31;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h42be9747601ffd31d1d66dc1adee1a181526024696c3f0b2de5032511b70000d9cc8a16379d8b8b4e6132c3077b110b9be4f559c0c8ba9d3c74f7ccb04b12000c500f64f7bdb5ff577364d03cb78;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h137c3da721ed762492c359fb2a4bce20e5b0fb0cb9999494ceb0625b90a23ab2cd5952b28a1af1ea8d8db2c6cf09fc5f8dc2fe9224e3736ccf5a53ca381ff3a4595e110c1883a92052f7647a4183c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h7f25fe7738ec5b1bdec20a72e803e2eb43d44fff4a6f9b37554f640a44e62ff5864795e861b0ec214eced9f95749729de6d31ab4dafda4a05421b572316dab04355efa86c0d5f82ba4a4bb3ea75c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1534fb5774e2c8faf069d548d97aca8f61069f85eb0b2453fc2e3f330b92e6c2ad90144d1af095288d363839e54bb294133eb8d139bbffb3e8386d4e55b3c2b1a3814017c51985a0c0c2d37492f1c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h156d49d3c7ce5ccc7d00d1fae0c8d083cdb27b8ae130beb906eec51f4bd0e9ef839a178cbb4b26d4dd77340ba95542f42387107612357695ccbdbc57d4bae42dbd35fd4dcf9cbe0de5af943143b67;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h935608dddeb1f02f89c93d8182fa1e2b22f14d2ae72fc3fbd43442a37626bdb5c0a7c00d513fccb7d44a641f2348f21b05411f198466118badf19e0a3ee870e3755973cf6259f041c033231feb5a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h14a2e66d4503eaad8eca8e7fa38c28608daad1fe91325eecd72b38042679b7819536e658e16faf7b3d6f1595f9cb1399cab359916e7a4a15cf2702fecae1b0b2e351dff5a6a652edc4a84ce82df14;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a10edd4c9ccffffe197842a15b055807f555b094460379a9a12f2ecce8075d1244232331c4ae414244a98a55bd2ce3dceb39c30a119c452efd84977a9f9f5558fbb9ed96a2eb3863be3f8e9da697;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ecde29829a91993b5890489c2f570dae52a98003f95d115869f1fbf0a1a3ad756da58a733322daff843257fa9ca8efc66b4c39e8d4964a7c07e0adc22aab0dab565982aba678fb021d1fa88e7b56;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1537e2499ae5f627e6ab016506b7963fadbb755eb7697354fb395e169006aec4613dc2db0666d60c144186ca08cd66e8cd9f0deae5cba503c357f4b68d123f9b293e58c1b6b74ab51f5bfb783b535;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h18357062bf28767be8e0d633eb260255f43cf145c04cc13015b11e71bf8ae83c8da3b4179974a11e15258eeb12fc5129bd5f57c79bf450ac0d3035ea0bed1ca5801ded7d3ae29cb48ab552df77049;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf279a59f39c19a9f31e5c2ef6321aeabd1894db6bf3e44dc7cb3114bf7743089667d14c3562a5dab8010101948ed8eacbb23f1b96329308ef70358d28880109a0a51e3a7aed53f755e566806157d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1fc859eada9d907d9c63a73e4973bc3943381f9f43f81da8f3dd2d9fde99091be499d2f4b1fbd3c33812edf03e114dfab86bdefc1b923f3b0f2d482f5c06a15b006b924f284065343281b7afd25d4;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h33c101ac51c0bc14467a18f9ddc7c2245b71ac8c61a5917ca6ddb285f29460ebf0d6a744f6e8bcd3954f46bfd3c2a5af2362031b434785f2e421219e0e591ebc4a301cb8d53bb22d074598cf5bc7;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1782fab0c2522add5ce4a76c837ad74bf598153ed393bdf2677c7d50966bd643f357e0c1705db21febc5ef3a11c5cd8f8c2a98c312e52550d9e3abdf573d60b38b23524369dfb86ddffaa5bcf5751;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hfd4b6c711aafc225a2b4ca08e075f347be1ec4b2762c03851a3f74ac718c649dedd2495f68339568142ad1dff53daa00ef78c392f6aa12c8408ccd2fa470b35c16f564c19d6a40e7527d4f22b25;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h125fd8bf9d435af237c24c370893b1ead43cb9bb30e8cf5963e8ba977523bfc4db5c3b6dcb89f60cabf17f1a589a35a21a1209929837887a1d6c7fe55adfca6658694730c6dcea00a3d8a3aab653c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h77547b91e1c5d3a15430b9d85fdb16665c922248add8d94eab620137b886ca1587d851b94585649bfcd35c1497ad50971bc020848fa1918dcc7c42c4a2913d44b1c6ca0c7b90a26ccc22576f757c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h2c645cc84a74af759334baafa164b5ba2c1a843431c1d82d0be455b9fa6d54c82a6f62c560f1c65e5604f66a73ed9563bef334802064442632927e855ea244e125e6d6e1ab15efed4be1f98cfaf4;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d95e87d5eb0a5194d7270d41ffd53c1924bfb172b702e6d9a091138187ec7ef800b5f1e918b96fb54e807b91114534468f006fa52b53bd475d6493af013a0907644725057a043e78a80319f0dbde;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10f86cd92227d45ceb43eb87fc93691e7e28c9d2a888308558299a772f761518135b40860895ec12586fb939f16cd6f2e4fd167f8a3b89233906a9cf5e0e7242daf8838f43117c05abf760df0d2cd;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hec851b8607f0837362b2111ea450c0363b94d0df3b5ea3c69e32050b5a0d371053c93022e09da65e3585777a99b67a45b298f0a134e480b8c04211888456822df0f352d25e3e4afe298909cfeedc;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h71cef8124e975447639bd199ffc189b76bbb0409b25d052e4dafb7e9c5b0efb3e03557e1478e13700e12021e6d49039d6b69867ade337c8d6d40a309dd606ad866f4d5d33cd22678d8dc55892c11;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf3c0957a75fc302d687d0c1b657a136ee77127c7563872cd007de1aee60ebd5e2a1ec254e963982739488e1c63032d595a0f1d3ec50a754b707af3d8efaf5517b72bbc0a96e163c647f25c612578;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h17b61548601223760b456b9048f3aa8599694196aff5c4ae55f7d293bd4625ce0dff1e4c57890d0e8b1ceea150764ce9867d16546eb424c2b991fa6302b8607f5bf1ba567619bd74939f9cd5ffb6f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1050843665bd7693cbfe8f59c46eb71a4ab7ca1b0c75985a342118b3826a217704730c0311f2a4e4d843b73db4a3b929ed1f98d8aa4ef1890283df42919a43313198cb1a14527ca0ac440e1266bfa;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hcdfa5a17715321f5e42bf872d1aa444735a857aac58c096e0705c76cb25c4add215ab2300d79035927e51018b25c58d57db76f75610845ce9e2fa5e256720ec3ff809fb7dc7068d84eea9edcd02b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h741d5174c7ef16c40cc56fb36e5e846f12807745ab4fdaa30073d75ac9eea5510bf363b72900196e559978f54db9f55fe87e20ac59f2160d6ee0c9d97e462dcff1bb3a21b008b1bfabf2fcb0708c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h165459cd4a60030e0495adf0ed3f66178e7e514f14974ab5d0e517a2ba02be35137e1d2b82f0cc65a98d47e1504401f5dc17068468329f794f4445a4096814e4c635ce38b44e037a4dea2a1c70436;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h4a73135118a6756a01d5b5079b6eb0228efae61f66a1afe3cfd317d759bc6f535769bfad9061636977f3cfba7cd06aaeef8dca0006cb27dfbf464db6b5e4a103416a6b7a83ef3bc497e2e1a03cd3;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1500569d54dc14ca9ace0358848d1b9085d314b702fc6ebae631903c7ed921f0b734c9d0aefc6646f049ac79fc568da5412e0be25d998f35f364e9aa726d49ed319b6e373dd3c1fe64660216747dd;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10d2c98d3811088a6c26fb71c64824fda955aa596ca5f4e0419d045aad4a0591e7d658871ac339933dc403843637b5bf9fa0426e9dd0d4a4df311a566d5bf5833e7f11364bb5f431862c3b6048d74;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h9495294911cec3a52fb6a28cd69a1e211e252044d3427bd2641cf6748fd63b492566930ca81bf0a69b62930113412de20ce72d6e9e16aebeab675965e3aa11f3150b60e484a6ab138559401e6d8b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h2af0c8a0166e1030cd434669599e3b3b77153f3ff9cbd515b85eb2c5c780194f17d7af077583c51401e4d0fbd1cf51f1af5605d37d7453aba64530494f18becc3baff3ca9df5386153d40ba5366c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d3eca4096a7dca8639aaaa01738b37ed5d7846e5e05424972ffff0487b764fc45f1c4b64af3eefd7ac49d0fd72abc4476566d95e77da371039dd7937f71481a548c719008e782d3bfe833f0b08a2;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ba3c8389df6765d4cfc3f876791a8a21435d50498cc9c5b5d8c69775397a4ecc873a7d08f67364a4e86ec4b9297dbef06cf72d44f01171c50f5f97c2c2f24cd985eb5055ce83cf3d05f7edffa0d7;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h62968483b5ed806193f689762eaec9d7f8038652d9816d6d70d804783750f670ae21cf3b21b62c7d12745414e3f9bbb6fc1dfc03873e0d9719eeebbeaebbce709b4575f553fe3380ea5135e1f4e4;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h958c6ecd573417c89a046ff8ded9f95e689dba4e2f30f41d5917e79e5456eef3e1aeea6556d3964008fa49ee8f569fb09dd59acec71379ba5661bdfb0fc6b52838ed7ad411de22bdae7fef9ba93a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h17b9f0b51689b6c466523682ff2f4287971ca0cef6f45af350b7cd94c56b708f0b342a3dde114de771819c25d1a197f9fdad3add6c237315e46df0232f9abaf1eef74f412f670ce6f57cbafe4e037;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc0755ca01714b24a9d499768803aabb02e321b80755b96ab8d3ea8df9505e6d2dfbe1065d7dcdfa3f6beccb17cfbd2464898b8c5c60ef6abdac5acf98e7f3099c384f7e8309df6a8fded0dab4bbc;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16ea9ed66882c5380bd98100aa06b6b92ba38100335f023bc804c88ba10654efcfe60807f7a9b700f249ae1052ef4c6b6fbaf62102ad35f0f04e60518e20ffbcbfe5c9e98edd5eb6332a8ee6eec1c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf7255b9480b5390654a15fd5904e0dd394e01342298f0e3f294dedb0908f1d2e72e78ea84c8bbd8cdf4a2771e4a221e35dbd09f661b39c9c2fab7e9b4f8002bf2c3d2f7f87fc50966c2a58602614;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1567d2f951e13567c9f0afea2c88454989ccf743b0c79eb0abaf0d2eb45f1117e27f36db858f95e3c37a814c7fa599bc90ccb0203c9d70b41312a31529ad79702760baff2017929bce840f443b832;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb50e67628cbfe06638c63a9741f0afc90352e2fc246aa7ef1a929c0a8357dde5f7ede179d68f9b8a2a15fe059a8bf6117181046f48d7a1595175ea4ae5679869a7d5e0114ee07580e29151230f99;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h9da0e2ce0368fd8a1922d83a06212f3ad748bcc8c0cabf17048374a58832651d4b423056234ab122847cdf158f5d0563f96fedbcfd4332162dc578819eb8de93ec4d5b716d2ae1336394a586f578;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h17a0a32dcfb66504460c9b9cdf18e1916e280d101d9a8b20fff07da01f0df062ec467a48902cadff83075b51d5d031aff0007996e580446c834dd4d6710386378f61c41d9b8829499c4b7fc68c788;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1062bd58c4b6be3c3df6a385a1f09dfaf1ffed32612bcb1014c41035ff906b2d137f9a1306e4bf5fb33fd45025532fed0e863646e80610af06e613255dc4d40150a847a15b60a619c46ab43a96c69;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h199882e38de99d6075060457c63ca90b969a0ec66788326eb84d4a264cbd7134fa87950f9e446706511e295e71ce7f6b7113393271d571dd906f1776bafc416809ff56aa623b400f1275634affa0e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h9ecdf6fb20d2e86780c68b3bc9ff3544407c158babaff1a023d866f3cdda776223793f45a7e2b9e7cd8397b403678ef5e25f20d16a17e634cc20e541758b76d4b6c886a923f5a0df7656de1c306b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb96c87219254304e1589070d719d0951a60423326c7b0f058fd41ddcfa0d5e4c7a976b3d667e575b355255bd764ccb12dfd1e96af0929ca53b89bedec492455a856609aa77dc54af01b3ab2fae5a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h189bed75377f4a1ea6383a67f1a16d85cea7a7c7cfe6812f9f9907218f17b1cb010a5a5f91bda3e6d0375b1bb4fcc7109206bd9074d7177bd988511e5d2a068102a91f742b76566645754720b803d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ff50d73b8e9ca26cef4484cef60be2a548a04fa94c1c9e8a08c4d6edeea20507144f1a416f633efb0ce6ab6182da2b1222861fc27622d1e0e88805b17e824d7983db2f782a774255b76ef13946bb;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h477191ccf6ef772272b02114b2ce5648e899ba96245766eb6158d72dd0c4b56d7d38752c5b2f9eb6f06fe91797bac0b3610b50e8c9331f3b8a1761bfc0bcc0de14b8e348bf21320923a2337b4a82;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h4627725889295f2ce7791f9fd262fc5783d869b826acc3736f280f563e496c4e6301a9923e6587d350947f115390d15defec78d3b34a85cfdfb43257ae7dcc8fdd3cb1db31c9cff33d1bd2ec4f6b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h117c754c8156635429f24629e20dc92411a2cf28f194df0a430202a6e66958960542ef5fb5128616549db879cca8bdc9498078bb239689f9be5d45ca4b8b5e66ab94fc13baa31c49bb6c30551cb88;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h15a4b2f1caf20ddba999357f7fa29726bfa3cef107a668363055868c60b1bef546bcfa24ea5349799898b471a6da5bdebef44cd145fb7de5d21e4e166153340ebdde31942f584826150717c267910;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hbee90ccbc6b83d8551125db9eecce801956ff2985b1b4d80c544890ff5517b79f7e9f74025ab671539528336831fe3ab59731b3a165d02c21b61e4050d2db33d5ec3bb16ef1b39ae285e0988d735;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h109cc3a666ac21edb8d1637cd1e82b3d941ea4f80127fd78dc2c56670d4c3d2cc51cbe6a6be67fc7788475502703f7f0c26591be2f27deb69908c21571fe8f0375ff4c96210a19ea7c60f9790ab67;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c51b15e0667024625d7b38eb317fd7318ef7919f0364b8f3b8387723ba2d954832da14f2166b44b41c163655a5fc818718e72c0b6e5068bba4269fb14d9566bd23b43b4e16955d896aa6b5b34200;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h13f3355b69be6ac3178ec15ea2c3569c57a3811b2522da30c97aa9333f39e9df99ec0fbc1e0cb3b0c34847f8ba16be2de266f0c63a0b5f8eefcbf3c65095a7437c4698e764245241635dac4aa5bd0;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h124de22463ba92cc408629580d4864fe86c3f28e204b9eb6abbdc285e8a286ef99ff6cb20504d28ad265910541f8ba505b6a8dd985c3a49a42e0e131a223abd7b9aa5ad7debf4e40e55c088e12d11;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h72cf59cbcc58d7fc2f61c5ce4b2ffd36db6c7f93ca3b156ac7c109104c3105c462f5ce597df954deb52c9c2f2ae04c78d409dc7628c22b4130b38199ea8c886b59c2944e7587e6eb64397b96f31;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h135a0dab07daeeb317f2dfda1599dd8700ccf6bb9f3fe78285adccb24f3f1653789b6ccb5e6341e78e7264b4fd042b86a9d4ff062c08f0383f5d333418887baff166ba01e1681f36e8cd0787c0094;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h638e027bcba57978dd55102b57820b19627d90fab78162ff1ee8383de82649984f2cefbfe623de5ae42e8ca224843c5ab6edcee5a9cf68c1fc7998afd78eb7d6f88c5b5dd9e2d6fcc9030dc266ae;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h56470624a65e61f8029ab3e61bfc90101e8b483514b554c355d3a933278ddea57db495f281612c8b261af312a8730527d0aa05bd91ab46079d87e36286c6114329fa4b3fa9818f061ad2cc2d9bd6;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb55ef0ffc870a799a3bcb050dba3acf71488d21ea07b341d1f5b48419ab69617f0b677e63d8cd86be829282e23cd3c9223c5f54a5e40f57bc5d8a80f537c15fd1b82b85603a90211958deda2bd92;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h5481b5b6dd4272de76717059e6c0284ce570b98d7622b97d03c46d37c08648d283c264300654b272b874d097f6f2f8124d33be7effa2d9a3af8f46bc164266b4713750a4c1ad4758cc4749cf9091;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h15c2a5998da508a0415c9d1f3db0fe081e0bc9c8dc32ccbdbf5e2e16b85324de9f023f808a04b3a775b1f696ce4e61826024593c2438a092ff877158fa7d19359d90a98ea69f0e6550e6ca7a7d7b4;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h5da070fac1c8060606e38e695858798080741c207f5a483c06a1dbedc32dfb936e32502bfd369f13552bba0f19b95ac7ce4daf1e7946bc4cd1666e604af8ebc70ccd03ab21135b89b99f852ac32f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1598df030ae604e11e0a93adbdabd1c21ae23c0a3b15a22236df7b52ffefb86afb66dae265fed97d361fe40c8022d127188367f3bf512eec6c41d7bf0fc17a6502963f13b48d0fe454917da48a701;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'heb52ef9508c26949dead52ebc0c0e3710dae7cfe5bd49dbc1f419a39c71c7dc6d09e134353f67d5acc1354eb3c0b26892272a9ddd43243aca9fed23e950e1215ddf9317c48ae465d25a113ccb39b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb2855ea12829b2414d56c083c6dae7e45427505e2b32a1171dccb54c213f8a6cd5563edd93a14fddcafa2b978edc77c40c05b211c7afcfadb31569c1bbfa202911caf5b00f8a6b4a08a1885cc3cc;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h169e2d13ccbc3650a7370e8722edee7ec5a502868df38e39199782068a46f3e6f42d7038fb2aed188aac6bdd3d89cb2217775a7f1dd96b84d9a23391f78017e0f041e6f564b48820f80c7df1a11e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a015cb386beb8817133a6a9d63ad9dd710fae58199317316140cddc474ac62d21c5e6985f30361899dd156cebcf28b3e3c831e4cea93d45e668c5ee69a50672a977df9b146ac4fadc6bd999825b8;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hef443681dd23d9256da0920399a03261dd64038925a66fdd8dd5fccbd41d572763cc4d2eab1a3a5fa6951b35b9f0b40a03ceab60a0f8b59eed324de1dbf8d8b47610044eff4912150e6ee11e8d00;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h19cd4ee16a103b9df64b1805ea2cd7112feae572dd554a30e2627b61b6f2af05feed91115b75936aa83ef9df226d7b9d01a52ea5417c5c5a7e7e9776a3011de60ea6e606ba527a916c833b8753822;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb88e97f270e5d558a42a34ae60556a50a184a7046f17a708f959de857474b70345ccadb548c3675f50e1395ee46db3969467ec7b82edbbbe0418f1f5935343b86f647cea0811f7de1e986e856cb8;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h19dab9952b3330a976e55721f42516f26b6bb75279b4c2ffc9f629365800922e2acbf279a2654125e61951c7fdbf3af9fbf4964e48afbe1150c5421783d1511c42c1ff302f67d8d4bc855d2a69147;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1af42b0c6838f590047ada95210e233ea1ebe53e39a86942dd87bcf8e68f41f36371d891a0b5e9e416fde9547eee1793314157ebcc89d804af50b27d9634ca2b9778cb0a875d729b235a3293c76cc;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e5384b4999a0d52c5987c5de308602da26b85d049c9688bb232f40b07c0c910856841bfabf2eb0a8b8d846bc48252a44ba425e34891a270b5836a30034ef4c347f23874d957a6aff113b3ba4c671;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h2f5f713647501efd16853d9fc35d59bbf00020ed0445a2cd30d46592b7de4d67a716f4db96955a814f68776f5076ae4c06283579179838127e759f9476115c9e9e59c74a69a65078839a57183a1;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h42969e7fab034a0eee497b7aa80e92f8e3415140b78e9264095e04646a677fa7cff8587259a013a0fd7cbe8f5bc9cdc04d0cba0f997e833dee670758d0c27f0c535368718401585821269a5d2d65;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h149ea75f3935f557407ee5aefa4f6fb61787b7a4fc3f51ecb366455ae52e1157fa4ef9d0670663a7926db59b7d460d316019c3ba685e1b2aac83a30744c16775711c0449e90d071bdb2aa44c653c4;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d43be78d1c9e8f6aa6d759ca4af5c0ab0a3046c4086e85a739bf60c91b19e33404e13cd01af32599f522fef2aa0e7e763d2f911d7172b42f7e407a32f29b88b825abaf63a48abb09e0e89c27d745;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'haec3a0511a71d144b10c365c06aaea1272c9756941146a880fa2da4fecf6d2ea74863f6f970d515502c37bdf19c85cc16effa42029f8f0c55a71dd6632f31e5e85c89e0e09b3d8c23c68d7dd8dd8;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h45601acea64ccf2369958bfb6c529c1929403a8e5e290c42a4ee6a412b00b05ee49322c046c4cc0ad0d5f238d13c0daf8c290be323a03267c98c41601de1a5280a065af629b891238757be9291cf;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ba9a3850cf44bfc7e3985d9d85311803de25296db51de52adf6e3aa93156f388c0a7a30c8c927d87c5228caa2ae618a39b4b329bdd87468beab4bba7372b3641d171af3ccaf01a50f258c5b88c11;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h69405d9a5289fbbfb2f1cdb9dc22529629d1474520a61e26d81cc4f82b17e5fd5ab5b3ba4618eeebe8b7a5a59e7a13381e35f5b5624d7f94202ef04e505ce4021736aff92e97e7007d39718a631a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1500c74b6aab431a5b72b743289bc65b8cd5e6ed6d56d3103886ca6e21416b8b12b69ab5736ed7751ead61d71dbd43337b6e309c35a9ceec7a42da158b08ce2ddaa178476747b8c586849695b176c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h12b632523a097887a45cdd6d64c026a33d19086087d8ee09ccef893baff90cacfec50f0b2b46364f24614fb3139c68395e91b6d3b45ec79dee7e6d33669ee55e54914a75be060340f6eb05993f05a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h541d65ed045cb43a9765de6c7f6adb37d009a3d9f21d2a1d221778069d627778439b3a12f3a1d9a52c8a65946114d7b1e48335d8d6ad45f31954d5a8806d095572b275d329d96ef2c624cc746da0;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h18e42b6a6a50967d0518af8151f76f759584c631ca171be685cf56e2ca47138f2936aaebfd73486406761243dfd13edf83d3d09a445266a7926983f19d984d3d0162dd5e296f57a83c01d8f6f01ac;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h6812fba96347e0ea81a939355cf3bc9cf5fe11b7b7c58ad73ccbbcf1d3714c34e1569105a16ab590715f4e5c1287b6912f1bdb40e6f6b1633ab040562980765113d099efc4d584aba13e5c1553de;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1bd6d90f0530fceb169ef15b439e52b3de37ad15ee11e3de69490f041795a1ede3e5713935a4b08255362f8d10dfff86b1e5e92d18b20d2dc2ecdd969bdba00b8089352f0e8d6e8f20fc1efa462cf;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h8be3d53ea58235b98f2825e812cce78cca2b25c193fd95adcd864d9157a277b0d5c7b1855e9b88e8abc3db796fc5eec04536ca9e7e3930095154635f44c620f449082554d811d74404ffee489fa0;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h33cd1f670a4fdeda10951442a062596f75447c57627406dde10c98ca6cd3d3c8ad859b62d86a727e8a30d978201a511ce33950a4df4dc855c95309cd03b9c9258f05b66c053c65be3a2fb7ff1e82;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha95da1becf52e7ea0376e4dc2f8c134f04f8e2eec253f0b7c0a99cb49f0e0f64d413ee42d8f3295c01c8c346c6ac14562b9b662feebc0fa1d1747fc8d144298bb17349a88e3965f6f9ab7be368cc;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1cc2545da799c3e2e613da4fffaede5736e1e600bacb4a3969be9413d8bb86d4d78995267babe14e158772a0a6bd985efe0d997ff9899e56ef686ba21f01cca02c6d0d1c156f4918e37b99c480e82;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16120e3e85a0d0076342c97a29b0dd1b02a93fbc894e249849156d570c6d8afc7a841ae1adf5caf228b7c7f95061a43162ba0a6dade2e8d9956a5576a66a55eee0fedbba29f050634b135d85af066;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d89db51331b034810bc82c946d0c180bb150791166db3905328851b74562f42fb8a3bbecd33bc57beb8e8bf02331f7ac0e63cddef2628ce6566b1ebb0dab152e943bec43c8effec075c062cbebf7;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c0cbf9cb237ffd706836166649d3edb713281198e8f6b0f45cc9f6ac4e143c54c3d9ce5fb63c498b3b9d0259afc579f7c74ddcc2b73d558a3fc7dcf35fa016f97ecc483f0455d00fc41e38fda2d3;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he30dd01583f223272a96d5c0e58eaf9f7cef7b1f950a214fbb6248126e198c6992bd8c3a722467545ab901055deef9053837d5951266459a40e26b21c0f2a57672b04d66d1ba901b94529b0b07c3;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha6f29de1e79965f40fabe06483ceea2a20cf5c76f2b8468df146c58ea3075f04d90f81a5df462d1aae38d18d58a1c7d9a9c8ede516876fd2f028d2a15c6338a44083c3569b39f2053995132e4f23;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1264094a047e4934ccb5759de4acf7146da43ad8956f1e45339a23c61357a5d805aa347e98127666202d408bc82a19d0c251f8d6b00319b3f8c9ca77f6ceb8dc55715485010383f71924c233b611c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc7e17cbb6e44e9fc33e0748eb86bf1b3c5e810a0fe3af59094de53f8ef2c1a9a1d7c61bbf7fa5ee33dff262db09c28747a43df9cf32ad447614e91561304b358f0208d3155a40ea8e6fd4aef4f8f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h47320aee8770240b40a6d76b8b7673b91f14ead7e1cbbdc00d1d45c4f607cec9498067617287a450d263a423e5e62683949e1fcd1987ab4f66b3d4076eebde26b4665d9c78bc9f1aae5b960bd7f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h162d0464c494be02dc569c11a4270336f4e22591f6b7abeddb366cd7b4fcf45a40156c753c0a959d4bb5f0c8d880d42f5f1abb252ec5028c96742c8a1ee00e4ba150faa6dd4b7e79fea542b13771e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h139382906d01244fdbefefdebb08bb0198a8a8097a9503b03d67270171303463610a5f204d37fb787df353664c619c6da8940767b51e2f301cd5e26dfb4deda0751ec1394e32ebfe5603d43fcf825;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f9e147729bedf96a191625a55d7d2bc271bb435d2e254eae33c8161e089216d9b3a3964720483dfc9af2acf4f272d769c41245584d1af4eb9b6e48b7960c5d721cd14bee72cf1fde6245e1e87a9b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h13f64054505c0d848cbf4177a90c91cde42f27734ffa716b7dc45d901a688bf6d1a68594052e5e17ad6191a161ddf8587a07a250eae6245eb7b0a97277e7b09768521dde24e9bc0a0b6a492b176b2;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha42b95a537da727139ef6ef289730bb2a55fa83aa1d8604a5183a79200624049243a319d7b999e7cb7f6f4dc177cfac2340aefbb33296afaad43257b97e19b35a49efa0dac26d745fb97c95a4774;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1501a3c9e50cbe6483c9e19e03c1beb95371b8c64e6f8c91c5d30bfd550edb3629a0da5194b470d2f344d0fa03752d7f656bf564c570450aee6aff19b6a663937e0a28bc149ea5cde6eace9572fe9;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ff5fe6a6e5222e675542842d44c09aaab5d23234181f86ff6712fc1ee7cda147f858c606eb6aaf032eb1bbc0c211f7589f61237144dd235af83d882f6b198ea23d69cb5a53c7e1f3b27f897e3441;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hdf90192d20e439d27d5212a33ed9cc350cccba0a894f4e06477f205e3b1b782bda79d428e5bae8ab31b8e66a27529ff0b087657a8bf96e4984512e7f2facc93500328230421d6613f989072515a8;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1815562abd921614e9dcdf0884d35a39826a99f427188fd0a4718f925f4e6722f267c32306fb4281e849b1d6d9cc25b4496114be7d01d7bd6334f043555a0ea89bcff9cf3f933a3f46ca61188dfa2;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1dc8b8f5302950ab7da5d071b698bfd68b74e9f75f1743e125633ce3f340d6eaf6cb710530b864eca12a4f6fb4ea756453c1c2dfa6f5dc6538a89eb52fdc5824cd32a969a4bd45d49830e9c520b30;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f4d1852232ff20d3387dc67003e0588b56876e48faff6f3c0604fc13d1f63b562ef5a37a66a9b019265a952795896316497e0b547de36a00b14dc73de42ae0f1af55a0b78264afc4849ae7b24001;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd64430687c81add75b19067dccd71336d31764abbe5fde7e2d20588e3b2d6fbf25877b6ace2072a558adf735d61f9772978f79b8f670e95bc56398f5b1bab3c815a18490230e7e1015b132f5809e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1aaa3616bb910f855d95428166002c18423e3a52ac00c6c6e74879b1c9efcfe7af15fcf5f9a73f666b816e793cafa7bf4b4d627cbb70725c6207e2c01e160fa20a6fb2d138d78e3fcfb8574a5ace6;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h169509bc5b83227ed283b8b673d5ce60d9f280c71278097f3928c668bb3ed758af394a98b48bb523f57ce6450c8abc20a98b005e68249485821a301b84dfc1c415654caaf2cd849c7032b2a58111c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h36d66b3dbd5146c3cf44eee0aa2c06346c38a001a51ccdb4bba48fa4796487a978b24027f11ad573697f1d3f985c972958a4f85183bf400f84054c7b9ef432b60ed367953aaca83367f22f478a73;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'had1b5770612e79aa2f39bdc6d5056eecb1b6d9f3e3279510fe91ffddd64cec794df43d59f2ce68d4046bdfca4da7127dd10bf853273dc5c9f364cc5388f304689a58eff1420d083d5b761380a430;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h37d6d23d2de8539e7de72cea8fe79562ddc0d2e9ce7de1fdda1e898ac4748d52645aabeda71af5328458d04a76216cbfe4b144b1083d73944cd3cf3eabdd1ae20e03f3fb1d1f4e9bd2bccb8fe286;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f3e5a1c041c31709efaff7e79b957867aac5363f0edebb7d7ed2fb2e65e1d93b3fd25177a2196a6161d7bacf32809d46bb6321a926b31cb1ffc33b602c58097865afa9087784059dfb0d2bc05acc;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h7c50076e55c5aadb0def4c636fb1bf138ac361ed602c41d04be47cbdf592af840c23c210ca6e235108a489d0670e0021fe66ffad3d1bff5c1eab09bcb1221b41ea7d3b7a02b38178003831784a5d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h9bf16bd9292fdc5d1be55ca915e2a5b0ad17831d7ec5e7e09aefaf863c3532f5891376d6db686eda9dff1ac34391971c8288e4bbb9fd049d7f7ad830f5a86c481650773de9ece87cf68e9409d36b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1607ac615ca481d08319009d2858c56613b348ee864e89aefd98b15d69fce584ba00c094f1c64677311a82358787009d78a9a0fb5956e4011392b3ba1baf0a6a7628e2102e59738b0f49ddde2934f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16eecc88051768fa825f2c585506068073cb184763ccd2c1db2d2c04bd9b5c6a9e47dcf1e215741dc3a8fb4d7c1b059d683e52fd17786261cfad1195fe82bc60d7bd1a0f791de6b2a8a5b36d817de;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h166cf5f2f414a9a1ec951023c772870cb2f816171b6286de6f30e90bc7f1b00a32d148e04f136c31b764092faee901b187cfaf43b797841df15bbb956d730a7c26578684f2577821640d56b525def;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ce967db50e3c3fd45642d06853bb087e6888621d0c59eaa13a6e519f80ef7543e9960619d4941b6707f67b12f66aecb11617eadafa859e277e4bc9c1111cffb2fb1f49a0048b5049403de8736ac2;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b690cb7f35cbbaf8c264be004b5dad497cfabab9537d3fbc450d37ffadaccb38f5e428028b47daaf3f8ddec0a92e51e71cebefbcd880fe30e931065ad758355cbf60debf79af445d53e1ec654f4d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf768038b7cd823306d48cdab3b815a43e4780715db572fc4c98fa852a039e2750decbde209b67b3657dc1f25baeb4c4ee86ebcab24bd7bdc129797658d014a7fc69ebfffa11d77e2b25d3d550d84;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a6d1d69c766420588919bc84e67aaba9ec231c0179eb4dc240b2d67e1ddeb29d6009d465938db41680f504cbcf06a6add8b7084033df47ae220a219640426239f224eb92bab0f9bc76d3b11f1672;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h102d1d52a9ad09c71b7fbb76cce3424ef414a4a76bc8529d262b1d39571ee564d7a877394b0c64fc2dcafc51b7ba09793d4d058a330cb5c9cfc3703e8187e64beb43b9a7d5ed4f13d59b11f4996f3;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha06c9684ee489396a125b7fd33ea04a3e7f31c945d2a31083f2c19ea22553773a6903f0c9f84707e3230b792ab385df62f68d73ad64ccf43fa73912b70fe16502bc20aed7b724e43ccd19e23f398;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1924ada8a5f5ba0baffae1be08eb360be7ffe52ba31d9cad490da6fdc9ed26a33670b36048dc84ad5caa0a1b3a1191c15186d55d2d920e6f0b15a633e51c04da0a5d4371c83221bd1a8c19be96f0f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc47deb8874a8a4f707bffe7bb64450be379bdb12f91d6fdfacb9fbbaf20acc651064d681e25c01b2a7154dd355fc73e6f79716f2205c4bb9f54283e01cde9b4bf32e99705b7089ed3caebdcd62a2;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hca6e28df229cc62aeb449052a62d059fbd42f53349e0ef671a19ad1e3a763b78669dd17c2a8fe8f7461cde065b935038ed20d99e80f894daa2d006c68c3a2c0907f08d679b564bc1ce09ddecc5d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d8b5841c474ae009772d6a1c61f8db0073aa139947c24dca0f56f95e2e0c9718cbf36638d3ea567f6233f2222c2f6711b71c217d6bc54ea4e6a375792e31d40331ef0498ed31dd1747051850de6d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1141eae3bac2fb80b262127d428675c1e7ca8bb932141d263ec1b570df6274ce72273cfbe0b3a0180628c5a9646a8ac182d1ae5e20c038844c2eb25ff8acfa18e635ea364fd4e680a850550271c3;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hfed045c35bc4166a380bd98bd7514036b55b51d109b0ed9e8154f475ec88503e73a9ca8f6fbf39644e1722635dbe4ebed3a6d30fb6186a935f01f21b709b6998fa480c0b4ec467e8cffb767db92c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h6820da94ad1edc7afdcb87d0ff3d5ab2c40a13200520b9830046702b3b1de73b7904b7316c91e419b6937e77a38e0514f431113f220c7718548b18d729e501df4c6ca57c65ab1348c566c703f49d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a8675a70bf1e7b31bc5ef1450482896c2cd514200fe7f3da40908ce13ef6cfb43e242807bab678e5c87d58266028b1db53e8d8bf4789b4d1b587a4f3f0205f160b2eb258a89304cdcefc56162f7;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h7b9f5f455ebd029b78fb1b24fd535425ee92beef7bfedc5eeaf692fe3f264110db609634deb9c9c6ede4ed96099b36ddaa582155e12c2a33e744c3a3ab609a86bbde2cb7cac3ec3c6797ecb363e3;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h19097faadd41d7e69770a8c93d4473e00f588a5fe77f82c101441791e54adaf509889c0f0b81e3398344c7e11bb9c15249ead33d20ba6929f228851768854ad16dbeacd94f09e0d0fa8b1290fba01;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h175989e2f8329b4e15655815003d140a85573b9829a87008091b633a0613dfb051dc5dd828b8fa681aa73e02e307fe4270d33b35ab3528bbd9ed59b8fad3220be125afe780863bac044356457642a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h2206b5b62ff240cef55f4f26f5ff6e240ef9f82249017f663c1e9a8dc5581d11b5e97c45da532420a4531d7aea3e868275964019cb4da77d971fcd7cbb77b22e81b38329fbe489bd51e8135d6e46;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h75f66b67505c331428e88404163f45e6ad8239eb41d3c66f69482ab01c7ab3a704be738dba8f8c458be0cb188e8762d63627802076e1793fdb781d4b7b58659745a2a886b913afe16011a6c8ad53;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h187efd1ed9e096075830e31dd2dd783314bfc4681377fd8948498cf21e4d97dcde07e1b6b65d70f5323857878d106a0ab5291656c367ed834b8b36e4329f31da6b66c5307f674a4a10c2a8e6f2523;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1219954528cbcc14c92918686cd33298fe01e8933534d168bf05f94505857a3284a03b8ee9a423a00ab8251a0daa4f7525b5eba9ff344f3268dca8c08f7456cc9859af41350120122fa2365016684;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h160c9f1947c1cb015d6dbab914b2ffd2b6a7bcd01277352fde5a7bc0a03d5d0ac4238847d6c3ed44a6a875970fc1e2b0fb752e3b12c54a421354ebd6a5e594f34580d5b4c9fb330cdec1060e50825;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16227e37c3b332284817b7618885206032e1045e1e8a98ae905e154d11fb25559df02b6ea6445922180f871bc669858aab851d5d4f7cfde8832928f75a4cb04a22b57a341a9423940b1faf52c1718;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h17739f622f272aa8c80087388f4241a34811b8dcc89472c48f151624c363aa380f7cda96c9a9f574442ebbb9ac91e9067f2ebd4eeb49401faee4532daa373948b2d1c30ad1ecccb8ada61f3e83406;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h18d8d723a84cdac0e567d4e9f95e8b87da05cbbb28eff6ea3013a335b5a6ca4ff5c48950bbcef6ad586586ad5da28d5b21eb59a2732a91675c4631d540c6bb2cfe237bd716e432724ae9dc8a38d52;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h997690b072b226eb8c52b2ca538d4826826372848ae41bb66a7f07ce75f8190ab765c7a6acdbfaceb6f6d6eb5f2752d4059e9f97a02f6bb38183dcc58150457aeedc6b972c8690ee7cd8065972b2;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb45099233c5c03703e7ceb523c851555f641b833af0f9eb74ce9162a0f1c57d5092dd82a036ab745ab30a86f794fc37d38f6830fa9090a7de1299f64acf1a0676655c69e64609388e0d1388ade17;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h17f596e04a794a44dd1f097723a3175e551d82c376a7909fcf8be16de503611da17872b5926e236a3fef8048369933e229eaadd3c4c9d10588467575dec4ccf6ffd9d1afb59c7b1591a2e74501099;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1325c08a4aa7086e3576037a04ac89d104d754222d65cff63ac80f5caa3f0ea91efa600dd7005cdb8dff39c320b9db43eb3ac74e424257cbf4c3fb36653da631085b7a3e8114fb17ce8ec3c5dae55;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'heed9b48f6794e553242d7ad9025695c5e18b168d96fd4ae493b1bc6696e12b888aa7a13c07cb857d45108e0d9ee623aa36b770e3ee68b91bc7db5cd1163463ba595066a175863cb7c6fe8c906c7f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h17a69f8c735b3daa9fbebf07f71b50dd3bb4b2cb8d0a136128786ca78b82b17a2a759831d28c8b148cee951b6fffcf14c53ba6ffe611b1bd92e0068dfec5e88652b47671b064f8f227a1082320ec9;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10323761d8dd3e75956517c29145804f3df6c6ea15a08dda9de46b95c3b0fd75a003ef3b064379c5283e6477e2073bf86668db4d1cd5e7db3ed4ab4fe036b950c18b4439350163c270b5a1c3d332f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf5cc5bce584608a50b07a6f197de51fc7930b0998d9e60acc01007b400c4fb7077ec763be5d1ce1a984695f104657e09a23f68a2228e7555dc86c056ee94b09bca94bf252286fedc506e9d624f77;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ba5b493cad82429e39d6ec9e3171e3b789c0d14e404f523bff06179ca5aa5fbaf46b4f8848ccc77d29441b81f63b06a115f23ea3af057ceaf648ee194519e661574405555eebacb05d0059044d9f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h641c3319aa6b7dd933a79a18929b012bd63424d6b27640beb9364661d5ffbba48579105c16b8b26d9485d765ef35f132af5fa16134f2c409eadf814ef3757d252520a7cf3350c0406ab8da87f62f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c74922bfc71f6b764f14d57c1a253c26cc73ce1dcf0d8080576d66d1c095d92078c2ecebb1a642fc06de7f7a6964deda0f74c862562002c9873f3422fd542556851f5ed9409b732e259d33b5d5ac;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f4e6fd41452aafabbf48cffbea49ee73ddd05741636b9f9733564c6a0c0e6fff4a2685ac3ecb895014b9fe90736bbbc445f439b9b2a131b81f676d53442324219cc89593032242df711cb87c97cf;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h8c6f68286833496a981b51aec1178add9b7e338206507fcf7d4f3a4677ac584bfd09fa8d082b87a208950598c5c16926c4f86c7c17593963ee3efa5cb541dd3928e88f977c961ed353a79fbcf56b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd23bf77270492806bc959791505f1fc948e01c7f93b4b40016b7130f40199b3935819d9049a90dad15bcbaa824fe89f4c1aecdfff583c611c325fbafe1faa71bccdf9cd3515a09bca895d7cd4a97;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hbea6e82288c0855fb0db0ee7f34212c564d5f202059252c469cb1055798f2e661ffecf6f9b6a64b25a010983b540d3617e5e3068fdf371eff22c77eb8f5b7b4741ef13bcaf036a7b15c8524f1baa;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h4002289076f462f0e2f0d75de11680d35c2a9679c18638b70a2cf78ad3ff4c974b656f90944ebbd745c9b9c57c25595b79d2983509a0e5c75b400bf02f08c3e38ed8bb2bcaa023bad3c1926302ed;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h18518c0edfe1d2436f84ac77eb665e2b1f156fd9fc1235431ac02f2f97eab2343cd3330cb4312f15ac018ad88a98ede0a7a247040a48397b537958bde2cf4e418844466fc889b52eec3d44258d14c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha3d252595f0caae081016d237230056d91070df67eae0d88625aaf468bdc121a94da98366edb5a86ed5760f24e18ecff9ea235757510b1bf71015afd7ed3dafaa4cd451ee0d57c7159c06d118551;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h5f8a3e969e4c5bfcb0f6663afcdcb7acd46a775b4a738dd4f37af22637a4e4d6fd98c7310c7c029f88f5f796838b2646e63265b8eaf26accc00e95d6c6cc2987ba177128a83ee5fdd8dad0a89572;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h91850ce24fdb1f16ae983096bdee42e23d61d32e16bac99182dcdf8cc5d401758505b5a04777639a436d21028086514b7bd8d0b19efee9c47120c2ae21835f1e4d6651acf50a61065947b0f6a3d8;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc4af126ed418d5a352b144cb6385e0db79ce35657f5c4d28d7e37de6ba3b9db8893ef0075779f31782d3120f5cf0395842875b9e7df33ad93afd054b05d936dc5257a181ec6482deebcbda1393a7;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hcfbd0248108c837dfb8f67c12961b98e3b471f6ce66d243d401f59a62a77c3d80af30202f02fdf2ca4ef8ddcce9f5cbbf24a5a037b8c53723c9f95d5d2f9d6b3ca454c8c5984c74c8cc7479d3b21;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb9966f408f026c02e0c24f8a5c491afdb838c55c2a0c233938cf0647c373533120bf4415f98d248586cb2b8d27a85bc58d18086ad208f1c4ba8e10bd9030e7d784c83abf8f88ee4b46745a280c7e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h95e044c49bce0b4b156f76f8e84ee329f478efceaadb59d07123d2d819e090fd717f7fc09a4cf500e4c8e4170a88887b86b8e94380764beb7e536efe90ed2848048d7866d8c89bd087fdfbda4805;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h14ecc239a5afbe92a2fc6b0d90b07228f1c0cab8186b4c340b791d53ae2f6ec6488a61ada9d2a388002ac05f7dc1c4df64622f1630ed6c5eb27f8576ad6f97cd42cbfef4a72efa4df1a1068be918d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h13699c962806f3be30633ffbde2fdf4b0ff60a2976eca605dd51516d2999a8b02d106d068ef30e7a4c266e255c51ed70fbd14c20bc38a50787e458794db5b6b11c33b0dab2d48c06fc015eba00198;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'haffd3a68437ef8be49592acd2638b03088319ef5cf8475ea0958ce798a46fa2ba2f01173841b6db68e36e2e24fc7ce83493dd187ec46ded337a12177a2405c058d530d7aab3babd0a938b20baba2;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e7ff2998ec185b1a6cd769eccda0c966824c81500a2a7b3dbb2c314e6005dbdf9adcedeabb90b913c5ad253f9330931147017b8462c61a9b108eed7988b3103b2f1a68ad994ca0d4f47f7ee22c4a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h978b539150bc06acb25e90fb7b89258e992a14c3688a62cf11da53b0813de316cee37732e76b3e6c8f7cf7e47f07295f210d09613e957d94a08c3ff761e885b07be81d46b094f7c540996eeb0102;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h8bcc398bd918b675d2c93f7d056754797bf1c59787a2f80e1d7ee87f224bba797fe22aee47e686cd7eea415b9ca09151b568635104f333676b39d4f58790ae34fdae97c5c00ee78f153aea6fadd6;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f7802011213f91982c9abf349478efcc077a8299b7f3c4725322b4acdc1d429f0865aa047594edd50859995790fe3c306da634117527578dadc764f030d56ba46bd70466d823895a5a8710309f0e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1746f24d20104a64d914adfd44c702295878a4fb82fd8f0f921e57197f2793c0aa542514d245226e44b5b5fb8b99172e629a8dd2be08f8ca94360e87d29f52f5c505db92dbd8bf6d010b13fe6c168;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc69344e7f181d1a4d48659c58820dd799712295c747c87ccb90a0cd6d25e6f27bb588cb8f896244e2946e6e31d91aa39bc17e42e9e69952a092eab43d566cb92872d9248ac33ee7a985b40bc665;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc90633c88e36b385a60c513197a089c8abdfdb60e0e6a14c57fff75b30e45866a7f22f49b2dec5253b9cd92d4b48bd0d3ea0c815c38ec332d1568ecdb8a45ea82e6c41da2ea58eba98ea18bbff79;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h8a7f0189e96c802f0b1640bf3f0d24adc4f367b72e980093f56ba0f543231803c5410b01cca14cb8c4cd1d45e6ce4e76d0ca9c7c77d7bd274171ace53ab8858169669dcc5856c7c149e04e75571c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hde1e1a3bdb6a9e6bc394fc2031dd9e0bf158c7ddb3219943b04d4038e3ee3a35a9546f62f7951ac291647113b52aabb13a2cf88d4f35c1723beed713dd5a6d9dbf4c99cfeb9b7ca504acac73d9d7;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h193282d3395b91d7832a7c5c8a163dbeacbd06fce10fb4d48d9d116a18cacfb7da9dded2b3a3ef6eb24f332d3006d4bd9ae5d82c85ada6423f23a4c9d9340e6ba2d33ff0f8a3b163b07091ccd3b06;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a6ba91c8c794973a42992b62074377922e1362a63a53b6e7aacc6df6e6e79d03769690bcfb577f5666b45e5d65b235c68c0ed26b195b455a2693fae899fc7ffd5a53ac36c256cd86cde27681f1dc;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10f0628a4b44d9afc70fbb707a795963e9a2c678d5dbba76e5a35727f0d09f3a15bac3c2eb54af9c1233a282c9103927e95057be07a4867ba65716c20fa5ecfd3eb473b2d7f96e8c8e1f517f023f8;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha6c59d49edacab4e2df39c3afcd9d5a1789b80ffe250a60944621d96a6b32719c4b1fe78475bfb9dcdf65d8e91e71ecadb2d0315e2532b6271c62e049ae6648c3e2ce6ae8c4cec61184a09d08fd9;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1329410cf3926d1e8381b2449c7834d6e622740b5ab72d280bf2b849b21301e29c192b7d3542e872751e2afcf8c3ead56326747effb2252444446f920c69e5a0afee5c5ce7e080ca301070caf5084;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1673755daf3e26c5754784f96ed7d4c2a512372c36914ff70f51f7f8b7bb1d41808bc270ca77e40cc4dde9ca4a87e0e37f86fd2048a9b148164e5bf5bdcd6dbc619a48137eca435468ce280c28c88;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h770ca00d049f045bd6d17388efb2c22d61057f4cb530294e5f6701de4f4fe5806ed91244a19f49b7ece5474b6c455dabaee94dfc3642cd6eba2f2d1330f4f1a2ff69ded73ad3811b64704a870ac4;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h171c5ab9c389c4384b7f257b5c20546edfb399744fb7cb4505de0f623dfab6facb07649164a14a0919b14fa3b90a3b7de223ab85703cf9606c4a6a9f3d47ea1565d1f887159442117440084ecbf06;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h9c6a05aa7e5ccee6a906da7da93f927f9654d94ad23a22faa478bc15c4bd26e6ec8592483639df5135b37fe980f7f2c7d3ad45e96c2f83cf5eda189ede848d4fcbe027c5edea62c9d60a89792c05;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd8a2e43e605cf4632a09059f7e352741631c347753edd40ef99cd64fc38b53ac1423a33ee74f9fe0f53a5d41597c5a67356cd55cee3b9c619790f3b86cabd5b4545cafdffddb99d3fa0e1294f733;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h612aa926b671066f3e0c801204b7934874bce2fecc3766a138d8933ed52fb2be1a76dfeeb523a4c14a5e3b7227eeebce4d5c3711cd52ce53691ffa53cfed28b4226a9711635e0ebeda2139c84acf;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h155edd7b5ac60e155361a0e278d1f10d786512622a278caebf94c8cfccfc48364cab5957c1bda32af8efad63ddb78cced953cfa3d15af8c8b28057f61f68b60986bad84841cb9c049b9328430f0e9;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b320416f4a744616075d98ad5b3ccf2884446bc7760e6273a0278b4ceec4b9cfcb82944c3623d48d804071d199468509442507e2a82172d1f189703e8a8970246bfa9f77851f82584132e0d1f58f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h14eac5d33656009d06bcd98b5f6dd66e3ae25de2c74eed89878baf71d6f79ce6ce32df285d68b5eae3a0c0d6d91bc411635be71752b0431ee9d9be97a25459f28876b32c82cee264d1cadb5c186ed;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h19dd4b45e1b6948946597f93fa7249164b544c566f904e98d2bb976948d0dac576e5b7e14b7eaf5d957a33da99f7b7710ce12545b3a2f88a4c5d712d3e3db078a3a64127bb7edf59697a509c9b3d0;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h279c2df20110cd8d080806fc3d33a1cab2e77179b8075cd15e77bd9da10517450deaa4cb252a6ccc3014a60349eaf7da1faf233b82f4ce50071ff808bd76a5038a0cd9c63cf232ce68282f1a1e91;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h39e9a2c169998cee8c89a77396923d1e488c9225a3145142464d3421ea91fd3eddfdaf85a0ec6eb755991cae8c7371c95ff71cf27df8ca8f83208ab41fc2cc7de4829b26cbad52e1ddba2a5de0c6;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a578c5f5319e00e9848ac4df8c7755eae58b6623e02cca678e9c65c0170d48d00aaed90b4a726231f34b7b5ea988d744fe40fa0350861eddb3d4b31dabce7d936f8bb7258cecd10eefd3b506daeb;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h913859d0d2cbe2911fa33757dee8d73fcc15aeef6823a95cd68e69516e933d0151367bd8f447d6ed53ee61816ed7fc185708577d927a341c0848e9c5474f7c66ba7ebdaef59eee4d0697ed2275b6;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h7828a8ee16745022955bdb3a5fe1f5bcf67f76d856f51fc2f4211d4135c5d179fe08f9568454eff1c4d5e44cc3b97b5e2bb118450f41739e7463583670702df3d5305561b529b730b3fc198b91d0;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h9c924d3f8ded5f5fcde8849bd7c7e4ebe8e33131be1d67988ad17c109a14d64ce5a39c68ae28bf94e6774754292bacefd19fbce48d54452d8320432587432269d19680e0b0b18e7d04617b3cf652;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1492f9fe7ea4b081003b2b3e1a3e0ce70ba2aaca7de397bca64d4e0c3d9c6c7bc57590d71945547da09b4af71bfe01e24160e5d0ecf98faf57f7f277184b4552674cf288b675fb3bbdcdfbe4de782;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h59574c4dc8ec69337fcb5a1404d6a2d313e694a5778ffa936ff17000fdef8dad5e5cec92fb2be910c36a6012cf5efd147f8a484738fe45c50f74cd9ca708285011aa6c631eae37d5820d9c7e1905;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h14e3e2dff6f04f9ebefdcaa90d2c2b9191c8cddef67a9ae347e61755faa5f786430c594e88446c16803798b994ee9b25e81c60a0ba3e203817b0928c6258506f0e0399ecf5a4b153b5a5e2cc83c2;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha536140dc96833cd240c2d932df25b5e3e71fc86b8eded40309b6c89e26f19b55b39f9ac3088c77a8c4536d3fb9f07040600f4d993ac6e138a8053b79d50d87ae66c60e5119432fef3df74b992af;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h57c94624709ee1303e3dbf20bc2255f6f417a1a340c9c83b5ff20b06416edf1f196735b991ffadea77613843ad10052c945d82a194cd3c4e02d89f0713894e67b873bcf48905bc7df2cba2567abd;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h93f62a263e477197cf1328c80f18d7d4d8b22314fd4d9b87f1e04e83bcb5275ac64597e05baa23b288e7bfaea59061b9740f8e0302521e95696ef6beb1bb2e7c98e7a91201a649b5d2df78e216a2;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1824980cbb414210cc23e553b81912b559d9de175eb32ce1009c303d7430f88cc4bfb8696dc0c44ecd6ff90746d2c9af9d2d9f20fd81bbf59bae9ebc4a1b8df122691d06085af09b8fe0823668824;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1bc024fd3a376165b57803dce8fabac65b93f23235b940d1c64d899a66fcbf5f4c975e04a24e45b1c079d99a7f782b1e7c64a51534ef5194ab1ec8d904104c0d0b6ee56035c8a5d3d3defdef35a66;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h4525174c9193cb489f8be6dd136f2b3ae4c0f9f7bd3b63a5af63d47857e094ee422953b306cfe6318e97cb21c96d36b42cf98ad9437fd918ac284c279d2dd76b1b69db2abec80aa4725cd058948a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1361b9db083345401583ee6b436dc1bada44f90187ea998678aad022dbbee4d0dac0fa980af25e0ad2744280020d27667951585dfacd46d11069155ec069b47060e578017cfc0a33b21c04ffa2a5b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h8e1ce0ec0edcf4c6454ad1a3ae72b4829518ff4e8c92264b2988109ab282d25ddad97a1e21f37408d20923845edc74e5baf2657d475ba444f76f563f93ccd9db8e070ada2305a0d8a9668b2af18f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1274d29c2240102bb88c3ee5e8a42c7df70500cc88c6386202bd4f348d2850ad14feca830cfb5c3a0e06e6a797dffd4b8ddd8af84859463682c66839429fea53602eaddb6483cc5a4e8529f77a3f6;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1772fdbe9a92bef2b328968fd6c2fec2b773ddfa55f7b4925c17d96925905d45d2f3097d3af9666b9dc5ce063073d277f2d7a527d06f49e31877cb9cc0f44a147c8dba976c3e24eee5ca33f76ea06;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he194a80f20e63fc6de3756e1dc19d78eea0c4fdcf447a704739eed76e607332572d29a41e3157f72470e41a9a0b9965aa7466cb346d720bbda7a3a65f2ad5869bb405719d6f2b5d32aed1fd8c494;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h165e515cdfc15e0dbecdd97585857aecdc4e643af56da3ef490aff6b10b3a2e0dd7ea44218e4d8b1b2530ff26f52f975bfcaea2932781933471624992210a1ee2204c5c9c2a462aa27481f4d69061;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hada0fec1424961361dff6bdd7cd2bfb37bdde0dd4b635dcfa74736025bd2681964e5573c8e4d619947a9a84bb369681615c5b3005d66446b4657225661e0fc3f77d5b98fc8fe091350353d46b173;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h14c6063b23defe2d92fe645ff5070711b36624dbec0f0bf879e19b2c76b39909668ed8939747ea3ab46c7abaab79f62568e228044fab131670d72db2ca4771cc212bebdcd73fbfcf820fc00e8fd02;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h15c80ed9006f2d2ddf34703e08e99f518e7078629cbbec328a7e44d59b50bdfb6506b2db2bbf2c3f7afe2e73cb861756cd1f6ccb6c46db13e5cb7c94cb9bbaacaa71165567e24388d66a396f73a77;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1cd9ae4bab73ffc5d9ee9384eb72a29768d2158f439d945c4e5e088b22fe48b85bd285c3978d1337f978c2248ff60ba579826de2ff4a6ed303c3dc23c7dfc09768d8148c90a950243ac2afce84bfd;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h445df9565219a67fdea05ff7e737369edf0d55dd2a68ce7bb866b682b8ff3a102d228ff0c29d7c48a99ebbe57d6afcbda68985889d0b4ecdd2a88420f1df337ed07fb26c72001721ddb1434228f9;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h4b950d493c33693064a65111056150c91e25136d6fac5acaf8955b137d7d1415563b1254f1db3b43bccc0963dc673b28860c2a0c857557ba204f448ee49944c427f564742b7b30038d6a270a5bd1;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a30e08beb5e56698d7be1eca50de331abc8a5687c93a2a3fefa73607ba926fa34db04ecc6aceda475cbbc37d19a5ef66234551b9c79e870937ff28b0b07286a147a4ad33c3c177fe380a93a04dea;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16579b358d7754cd65467fe4c0576b4c6d1347a16a9a74c62a7e5a1024b45872eb77bbe408281ad3cb7704f9699b7dabbdc98e96e78965b7bb988387757eeaadb9fe4c3a8b620dada3bdca10e1004;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f6176365538d3e9923527c5a44ceb3e3929be7382f6b7f7299c07bd9c50dbcd5d945d46b79f08f321e73d35702c34e01adfbc18beb845f4d9c1c7d03a885d5eba8df604693d8361806175288ee35;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h41f0df206b62eff6d8f172182346543595b1f9a79e22059a35d44f05169099276269bae2986c8978adf00730e9959a932e20aed3df59c5069575565065d5fe726b71c9eac0e7d4c4dbc9b84da25;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1553bc41aa6f326a1c54a6ec704ad911bd443c3d4df76c16a69474003f4549191c13956d2b8b99886954f89a263275268c66a6e252fd39ee5d4c3f68a4bcfe7dc92f02281cde7ea8611fba68454ae;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1117cfe4541b466b41d3d41708c536a46605cc61ae2afec6252454cb7d0fb03f0d4af44fb17f54651ade38533aec522cc2b50466b30d3a7513673ebb6dd9cd3a991b210602297bdc49f07617e6402;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h3385308dda9872db0b92f0c83194d98969cfc874a5b6aa26607e04673f3c007321a5ad6f2e21031ce1738877cad0b3538c3fbe44a0266ce6146a55ccd7bd3444c6e0d7d613cb9e990afdfa0aeef3;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10e1adece2eea859308fd0bde3a04d7cf2bf8319f754035c18e6c679881c97f55a2305f9908e76671fae2c44dda830929ba369935cae0a5bfe2c62aba9b2377098113451cde9c110b5b9c9b50b9ab;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ca56984f94ed1a1ef19bb3929483d0181ecb5a4c1217230e827b5f02cf8843d23a6ac4cf2a88145b2e8343655894e38c05db2ec3ad0085a64253e32c49af9beda2ad773e03289995f6f1216a33c4;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h14b6445f6f36022c5a858377266f9c88c540d148c54a9b574cb74c51ba31fb51d40b9ac70587c09bdabc3c3305efd125e0889a6bf5351104065eb46339d5f688652acadc651876f49516254486bf3;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h18731c781e9e73af69ea37fb356608a93019e12da7472e458ba1c11b07287c311769b3d1a5ddb8d5d9004d3ae6015ccffbf2f272adf2a82aa1c84ba3b85f754d55be129e1a1806cd7c26fa9e65998;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1478fea4b18a965032c94d4b53461b43364b2ba9a216ecc331c21b8996b29a6fb5df835662e7969a87d74f2d8323d1e6e21adc75077cb1e17ef0f2dad73ed3a95dd69724d1fb0630705e5ab849a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1067b15dac41d45b4a625bfbd1d0241a4a2454dcbb50b5740a9d6693b3899def576cd6ea5cc9e92c0e26fe4645af7ef8cf4ea6cd8912dc64fb32abe863e374540287f9bbcad33ebea0a591bd146e2;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h72a528e42d31a8e6fc63b23319a488d8f003be18ed90fd94632c08aae061cec51dbc813c873587802caf35409a00e0a23dbb268ec477360b3f4931c938bd1cfe9278f895c0b4ef23f79585dfe5cb;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a6870b36f43cc8de753ccf6d46f6c8bf24f99b0369c5cbf1b5229672d4f00462234826a0d3cce5cb05a58077ac5214d58d586f766f1771de83cc6c4fd07b06de253194c127827294d0a02e070dc8;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h14870d1d2c8fc484c8c1c2398a92cd01931428d97423f3beb9a51a41d19b4e4b83bd078d40594496dab0d457244ca1a0a29dffc62c2421d81818229a8157c2cebcefa7ae603d6a998ee9710eaa234;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h7a8d9c4d0e6af0bf0c289545aa9a0c6602afd4cf205538e5ea649282954f7ca3b6e5bb0c174185ea88d5d201ef131115e6919611c1f6481e2c84193f8501465bd5db69487718d3df98fee608fe57;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb433407e4f0311a902e3ce4a939db8cd4aab5fd3ced33b07561fff3d55b2dbe5500b9d2ad6ffdc6f138748e8903ed57ecdd562dd9bed872aed69367abc32f000dc73d1011a03c8a76c280a1317c7;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16de029312e94b87262b8a4123a3ccb5036e5b8139d365e49f9db36b1d1c294cb61dc641dad8d57892fa553472d763ee8ecbdecd413e778da8c87fcd352dbb987374e7870d075516d2266d7f4b8b0;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h11c0980b388d8d483f1609049db50162451ddb95b428de735bd157bb107c23b3e2e1e4be2355c66fd4f8ae062bd33dab4a02810f0ab8752f4b82f0d153992c3b3be39bfc66f99e598b2e32bb55bc7;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h40d8b4a2e653fe46fbb789e376d036f3ebd9c3104ddcf651500e95a6c40f2d3c9e39097516a00b2d6c78b3b09e64bd149f6a5947b2534ff1ddb238ca7972c0808dc26759f51378efbb5426a4e940;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hfad61c7d0d2d1abbdb5f58ec12e52ae9e166042afa58c97c8f611d0104b10de06d358336fcf038b98b9969b5073fc74d97aaa04c855b27d7db6f1d43d6f457bca07a88cfa3f75717622563f152a6;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1dda73d7d458b371028ec324ebca8bfe9ecdc9ce2815bf1dff9c1c9e2c869faf6dddcbe9153afc5a4ffce3a64968b30fbc3cc5253c2f2278be755c7a7911cdcea66d64fa36b2a90883c3998a730b1;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h4eb231f758a7138f45d2ec2be5e97a132bf3baac43ad28f3138d9e1248c825ddc38b0b5cb4cd5a7717a694dceba365b954d4299e0015b490f6633b797e6f0cde01d6929b6e709782bce5229d29fc;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h5a6092731ae027557cbc3a7f1474f3cc875430a9807e4f6be9b252595748580a7441ea33a9686c21e5f36589c3a7a70c96a7f06fd3de960c5304c52654950730b1eb729c1e9d6874b501e4899961;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h8ef38e194ca8b678dd000d021063d430ae29d817d86e6e996e52322cb49563324748014da9551ad9d11673bfc8a1e3db21a6fc11b3eee3c560c98092375d409ae9b69f63fdf7d2225357de6cbf44;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h7f79b077b1ea7cb221cb464f089588eaac1f147b9e78741c76c4ff67bfb44c6307cb9ddcf4626ce5ec257f6ea8fc6fb8105f03aad09b659cbacf493a3fe5d8a5947abd89af81bbc8ae80a0d25e6b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h21336e6a1649f71b11c706e8978d252e396b91f8cc80016469fd502f3c9ff489b9d28b001725799a295376af47e92244c580d5ac1c51c2f443197357fc9bd68b7c9c6cd4963d15f484821fa44ba5;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hbe5c1461e1bcf9b91d6dc9ee216dad60c732f635ebc039572babde0f4027fe319a2e7dcb0dd05c10a872d1fc3d2bae07e5edd4013371e212f8ee076f047f63ff00ce59e2bc705498eb1fc2d6564b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h11953c9a31fe83679e73eac5b28c8386edeedb54d79f8ade507989177b3b2ece811c0cf566b147bf36f9131f2c05caaa42a3bd6590d22799fcd66580db2a19ffddd0128b8aecadf72903335bedb1d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h78d7f0645a6269ae9e85258ca1d08617444cc4e86791055d854aa11d0148a32d23c8a9bc29865df6ed382ae1cf75a660886460860c3210041e2ed563c07b6c52aac5b181b3bf19fb07341191a7fe;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c10bb724fa142d17a12a16af4c6731bbd6cf1063f0f9746b8a61a599cfb29a5fced3b7f0952a38887f5c719ccdfdb8ba055152d865faa1be809856e5bea6c4c0701843c805a3bc8391596555622;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h61991ee2c34baec4535c2122458a9b6fce17037351ffd7f495d88e07e29fa7a1d1cf53366168ee1baba6276ae6dc9ad7e6b6005a93e9fde7084b134a51b3cb54bb2d829914104b68d8c525679ed3;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e79c6a1fb675ff702f8536e96da6027c5fe75b676a4082cd321d7ccfbbad817e14db97b6b419b248b62f31a381e9b6cf9fdf29f9994ac93a156243e0ca6d1eb2254056a8b7879f7a1bb4b3295037;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h19fa7a59cd251bf9030f390d26a4ae9818a6391d222f88a7d98ae20aeae54b397db2ad0d8ab1111cbd8ea83c95571370d9def482aad9db4639a42d0b81e59285cbbc94707c79f2eb2dafb6555fb4f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h18121ab75ca633e20a8e536d226991d80e4798e83acb860dc4005dfadfd449c303d6514071fdfffa453454f246473ac81cd7bbce985369428bf702f8d199d14787db85ecf3ac790cea1bd88abdd91;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h167acc8f0710062e0f92e48f83276c26026e80a958946e999a55359374ab8130463f3b5393867617fadd8bb290848878f3d3513b1a12c7cc06edeca7231a9fb08a3ac954ce4b5f282417d43ddf39d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h3764172357d49acd4296e8cec4d8dcb3b295d72346e2de993e5c1c281ae95bc7edc5a86007381c9108baed5486c8105b62f6bd9849e531edd7cfd45c31915fed81cc0e3bdf40b187ee79c2d1436b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h13d58e1627c5ad6669cd6b5d67aa79f51d557935f4d404f8c2226768aa183fb9f1f1dd451fa97b992c391007dc85a6c9e332b7c17ce530f1e5d50743c7d5c06eec38eafed3bed45d0f3c3296e9a34;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f5b012bbb7a05abc2c2356b3d725625c2e442090aab2043e36e0e1e020684c92ba0271af4e2be025f9f9750ef09e54484a8d93bc6bd5c8701392a40f8bafdf906b0edbdcb25f928903b9efd89feb;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16946f552be53e352e1b41cfc85e524da25291695785b585759da6834dd165c54efb0e6586f1eab0aa984922007b8ff616e62bc17be4e51c7ba430dfa4f35a55469d42f97d6ad0f8f46e9c0a268c2;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b6c97b8be62f1b9ceae5a937a1afb4f1afc11b4d05c9901fd7bf46ef12ea3d7b7bcf665d4ccf95c7f3851d9fa63e8afa4f549fda203f429424e2951a465692566df88a21cccd59c76ce87c898bbd;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h363e92ab1518257861ca599ea733da22a0ebf582d8c4c56e29a771afc4987d9ea7c302447c3d7ffbdf500c70bea341faea24e2dfd3c0036a04d4b92a818971d1f1366cf8675676f59d58764deb1f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f77ac517c8fc98c6d927e850bd4e7a948c8665cf472f41fb56f205cd21e66796f6a46425709e9e49e6d730f68294f3f7838be714cf23c47e1afeb22fb6dd5cd48a0721a2e52b7a5ecb35a921a68b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h5d48d10459122a71e252360db566ea8cf15b0611ad0a713d083f8f1253669a50cc9299a826c4622d0c69a54c14a94f4714c37b9b9adf2674588f1646fee0b91d3991c8436022e37d3993c600de4e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1389c015d4cb1c01bafa236590651a9fdc30589da0571f996f8fcf3ad50372996f0fa7fee1b5500569489970427f1b7678cae429ec061e82e3899960ad91ee8e87c9d2d21b1b11b9f4fca06e7d114;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1fc3230f59543b610b1eb449a4c13366ff5a116c1c3aead200ad7232ee0d314a8d56ddf774261d1cd81cc9f43c2e5aa283e591a043c2760c9c3a9efe487860addeaceafa9b73c6f633fb1cb104a9b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hee515dd073ca432485c0a50c86e5e8693e4c8049982bdbf842a53731f99be95c6f449eddae1b195e2964e2674050dbacf084bc296d1df3de7e712d25457903d99ee0bcfc798cba4658a3e4ffea60;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b259e4425bf2bc8781229a432af9be11440ce40947083be3b0f2e16f5e234f684cea51bb37a9ad1787fabf8c3963f07b89413e496876ded1d3fb5baa0a2ad8234c51fe42b6097277b4779246f21f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1bddfbffc3fecb755066d497bcc5a7c6aac62b534b34eb4a895103a2a5a26cb8b5d136f4caefa835391fd0c65f4d0344aff17ce302b37def5141ee8d9864f58d06e3077404e1f14ac61b905cd5f6f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h13e915a7fd11150f036d405ba319dc979b412705db122da1341a7c2807eb7d14de06aa4baffeead06b631323f57a72903cd755ee68691df9e99450a62ba0c900c6261f5ddbb3681b3b1a178ab3828;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h89f6e0f7d859971159e3adcb1a4f3213f8142eedb095b008a623e953921dcc53ee03f4b04b78b7ffe589ec614241abca4f18ef9adf78bfabcbc281262405cb184f176693e1b856375c51cfa24dd3;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h9d3a8746508a88393cb06eab611f11d8851765b5044c63130c9007fbeb64dbbf02219cc3b071893aa60042eeefeba0e8647130f097803e15d701b142e0acd9da930be6eddc821e606f44d73aa53d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d68deea372379d1ebef68400457483995cb0791463a32a2ef59b28d8f606bc85ab3baaf7cf099ec0a05255d35964aa9ce71fd115f6bbe7378df00265bd3bb01e7ad4a7f4667033c4112768d86995;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd35ca0f0afc1df68b39ab82b8c5440130d9a0bd69a7d3b6569e5b754e0c4830b1b0e842237a31eda37b27ad8621213ee6dff141c33376d952ecbb1bb8c8d9b03b724dca47d10cbc255179154d6c2;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h6494a4e46a009a1462a7d1b4cce6bc92aebdc5e6fa481142bbea9934fb1ddc538b46df8b8fa934b6e3c9ef43a0809400aabc6a15e771d0627f9d609c817c831d607a24beb6c5544cbc82f626d602;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h131469f6a0ac2e85970b8d2ff5fcdd56526d1bc946e192ba1ad64f2b2a0f886e55efa00ba067f6ea4fb87dad005eac5375812b2701bf9840f1f294485f9784a6fe1890c7ce5391a67e86254782cf6;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c589b48be7b93d3b39c894f7d28203e294bb084c13ff58ac8da6352bacfa7326bb6b75d5cae763ccb20b6738f955a76c02137a139fcb9f4e672fe823c1a5b2317fcfcf34b8b31778cae2a2c71c16;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h72318067aefc5d93ff9ed39ef36a5a22ef564d235b2a04794862d05e85252682560e22bec6f581e7cf130898fe2f60e2f266335d96734fa5ca704989f73abb81fe32e64a32116bc153f348c00551;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he2430a7a0f6202b74c3b21c63c542f69bece2d804f1495d373789f769ccd5b3c4205c743a56ca4fbc27d31d8c2e9e040b59399ba5f936e9c6ab7bb17e2045161e73d04fd379954f52b2f87fd4abd;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h11e5ce285603933947a5313b210e5e40eb1f6bac5a961960a3eac75cf3821d688b0337871b6bb0b17ad19056af77a6a222a145a05c0b261f04fbb0e5bd0cc39689e597ff1407f6d1ed778d057de82;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ee93c500ae02054e78822b9954f655bc7d53cafddc785357d341380304d6813211443b87ac921beec7ed9a8abfa7b3a11c537672c104b2791e91a2cb69388ccfb4db5335513d6bf0ef5a4399cbf9;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b12d7a02b0163e125eb74124603cdc54f3574d5c935b552bb85aa313c3b1fdfcfa8180d212fc50b8f8b37ab55264fc6da844322b2a07f681b713c63f2fa039b8d33fcdc2f2e3bade30b6c7d07004;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha34da7d065198d3b4dd16cf49a12a0231f12125ac3b869ea98a0b235a03af4f3048a515d329608369e6ba754c0f72adaf6a047dee1f7e0361c4901def5a3bd9fedd79424cd25d3ad41916b376890;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h9bfc53b5c9d2e8d5f8ca4029ec228cb4730adfac87745a6a1b2aa419fdebefd27544c90ce15c91a97a3f69368a8785a9aebe7a44ecacbcbe79eb4724d50d6e73fdd0e218480cdc233912d7516942;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d23d0f6cbd2168cc41739a3428a705dce5583c8e217b737a83ec8c12ac43b0de42dd120123495bbf3a546e2d2420b4ee8c34f69426de105f6e5b03fe7a784f629dfafdca70c172f20b44ed3c57ec;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h123132c1b2fe240f7c74dfe2229b8dc37d69aab215cf170e9f10dec827d47d499b97619ffbd08a736a0808ba6152f917468c67f2b6e9a2fff217644974d3bc990e60df4a09a0ebbb55d151ddcdd06;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d49a1822593640dc615a1395f05573f7b4f1a7577716c048ff84cbe4b9b3a223629f21d8fa11f78e6d9a47bfac7ba6d3f53557fa4730f6b881487f0335862ca582f184fe22b985a9a979b429ad7;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h4b976a02f1c03221768d471ec56b89e64feb5af7fa4f94a2debe84f6bb1c9366e2a0d97ccebaef5ff72aeed3a05eb89909bddeef3508513e22931dcaae82defbe511e257e9e7c337f196b38ee2d0;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h13a51bd8987eb5d09a8392876906e5ddca4bde6cac1430dc02cb42a5fc8cbece66a8fc748c0e16bd9483b885cc387993ee4ee91dfebb3c903d4ce5dd85d1e4824b7fa04d4fb7a62495339d647cf1d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd7e49760efd5932fb8665fab7a83e1a5d9a7e0601089a9c0211bd95fe92b4c453b3fcb1d1f224c960dfd5977a7bcb3d3ebd533cc989dc954c4a65d75d4a5be613f746120bf6fc154459e655c1e1b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h14d0e882e07fa3de3f1ae452485ec4d59ebc2fa87ef5be8bf2a7af0f09dc676f376d619c360162a7b6ee2aca36994b456424ee0d7b21552717c7da169ff2f464653158dc3efd7c511f48a291fd73d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h36bcac148a97f6fb2f60ddff28fc8625380c0513263c0fa5bdd6ab38f187ccc814204f795e1ca6520cb1b0f3a815497703a1a9c42057877b08cfd11decf68ac0be1e376bae9780c038eb29226151;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h19023970ed33055ff3c21c57cc111d79e2eb41491db1b94afb15376b5df9d7c9d4b66abddbbc986b179f9c93ac7dd3c9e6fc31ddece89fa9180982227f53bcc7e40d9ea16ef810885f4314c2a523e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10a1ce52b7b0a5c02d5d038b236e4fee585f182b1df7c9ad918d3030c37387d3079656cd1eb0436288d9c4d50b2ab7d5fc28fcf70d65f1c02bf5fb26270991172efbcebe2d7464d050a263a704a32;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha0fc25101eb8f7faf07c5591ba793d63d3516e6f5beb030d61decf3779fb60aca59ea915b6c76e20bf23bbd3f1e288c7d7e26c416064b54d65a10a30cc9279491ae992d79ca57a795bb614f7fe4e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he2cd9583d0ce49f15049b4c158849c2435d163b660bda9a762397121c410410ee95271239597eef93207fdece4a60f9d0fcf553124b4e03d65124219e62ef93eba10067db3d3d1107745b81cdea5;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h126328460ada2d3a9f335d8b0859e9dcea51123f0e0cbbed3ca591a3660795571de234b91c64a34a268ad4f65ae0a9800cb5a7f64c35835604a326239a8255cc02e7af06db3218bccf3a7e2c4f898;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d643688a37a904b8d57edaed8093a4f901d55345c6e8794df6adb7e6ea8e56cd4eb786f517083572eb4eb879a234ec184d8fe4203f0f67ebc38a65ba822815c1f4ef3c6deafc4e901e80f0ca9796;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h14f6547c42160205140f3a943ea64c177404fa4d6776dde1542dd41439324c89f8faa4c99e2fc3c4324c4d3bfe3ae9e1d211c4afb3cf09451b3bdd6c8e2d860e72fbad2f014cd93812fad3ba0c705;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h15fcccf4a0463385295a0d97801a6ef574d9631b3b202981449e4d33f67f02980abaa345f4cef143f8773b1386cf139536f8b1edc00a7d31d3d44394779c52b564910d34470a789e1439fdc2c92c7;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c2b0916c80f81a4d98723eb0550087c3a025873a990c1261c5351e6abaa6adb709b1681709dad11489c3d421d7678513ff87129f868fa028666db708da55e527af08df167e7800559c51ac7c68c3;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h13bc15d7f91bbe8736e8bc2b2f9dcd97c75458642386695eed7607ea3adce9154bb4750e94595192bb18fccf0db3dad37efccd4bae167296333039e2f760411a94c9d96735b26ebed0322118d02eb;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hed46f9bbcb18f2f678a27bbb192bf9d2ec5cf7dc8ed7b165efbf7b600fb546dc2223477945e2fbd312cf75eaebd426ff8228e55d7a1814434e8c6c7ee7f7cfd59b7122694ef4de73af4f0a9af48f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h18bd37e5961333d0dcf0bb31b784158e423f95f07844f174f63f4e8af2af318ede78cbd522edcb799288adb5a810befb6b20a12c40dec98ecf31c4f1893e25823375b08340197ac61a2956570232e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb1fd924ff89781d7097052e4eae0d42f09382d0722b41e8564940bdb23b8849eda5df4e91ba8aa6997ad0a25f48ae32e6edefbd3e8af4735917f6c55b5d637adc339a81bd16a7054614e93c031bd;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h8d1bd04ee153610b7efb61996b4c8de49485bd98f7910320048f4ad2e16ce616188479bde9138707f298aadcd636d9f96aece4cecc0f171cb1e285e6183cd0da8b11a44973abed6119887b566a69;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f6aaecf67e2531e535b3f6718e3c5c980cfa37f161c50831476e1f0f275fe8831ae0261aff92015fb79978af31b145ac6e62bb4903e17c2b4f8bd53e3d9788692c2b385750eb610f27766182cc70;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h41dd261933910f12dfa75db158357d97e0eee5ac65e8f4debc37cd9806d3fcc922f1af2948755db75243c0e989ff3a7b78136c5f8e9c67468e8670549f0c37676bedfffb72b44600e156adb55b2e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h9becd445d36a4cc680415bd0770d66961cbcb0e6a7910fae87f4333cacfe94664a9fb0d0b8f85dc4a5fde61d0709ee50af45237277ae93deabd6c73350252e303cba1aa7302a14fb5cfca2e955f8;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h12000c097e4dae6ff684bf587eefecd3a475e958f36f44ba2560ae664113580d05946109b5a813653e3eca8b87763f27903c8813e2c4846b31e4ef140729974333930b51f99831fe684e2dd7600b9;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h6c97ae6df02a98ab8f77cb017b9aebdbe13dbcd6bc6a599c114ec519b246e99ffe21738eef3ac552468f996275459a09d6b6a1fdd8ca42c6fd946baa4e841351bcf7ab48e183174713203e8f35e4;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h18bddb68622c8e7dc884dc1afb9af57f216f839d6634f5b94609603f778efd527c7c644ff42e946a78186c33f46371591f831e91c7e0602f9d1b2bc1d23e90c69b49ab100a12843c680c81e35d252;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h5ef7aed9f7e2907726baca7ba61e69c88f06ba1e1599d6a9434eaf452e933e70773cf70b4453039b191c4a7c4254496d3016183dfdd0eb7f1f9aca9a3920441c508d83989c975f76b6c34fe7ed91;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h13362fb817613dc080187902c4f66ef7476bbd57429ebd735862ba81c65e2a3f4b206e86db93c6396243e6904fd889f2ed4e6412272431167aedc9c2bec251eee3dbfd348a509157d96a9b5b012f4;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1bd44aa318959e32159c50abadcaf4091cb437d1b6453f45c0ae4b92f4b8a5845099d33c0c0fd9249153209db609a0a2607915148519a26c7a6f9bac91ba8a7fc6cbf2a38cd8748e6022a85fc587e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd3ab1e17e7f7e9340d2f22cd9a714cd39301790fe144d75d61e3a59dd0c1a3ec163eac147e51183f1dae1d551530dcf3203c06b3b8914c51ecec6afced6dbf12a9314025aaf3ba9d8a2289c6795e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb46d0b2bb0d24330541b5cd2bb94dc97a3cf4af9245ef523a96f78c51c614647665fd58e45d9a529bba72041882c64872a470244cf87146a5ee07332422ab55206635718e8ee0d15e068ea66d734;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10047a757f5d7af021ef9126dcd0ff3349db8a9ebb5329562b8b43b4442505434bbee7f868426895f0582b81539938982a17f483927b65a121b3cbaf1cf9d1fb4b606ec8ffbca94182fbba21d1f71;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h43e21e38a39c3ac3294b526f8806e0c1b47ad5a68c5d01f766a0a58aa1ab19032cee47123ea5e64c2d7a5efb76b5bd20c4dcc7221c2f6092ce1b3540a01ea01a02099fc31823e1c1d55dc284ed18;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h17b2a75bcb4b4d53f92da05ec271316cf0c5cf24239563e1e0ae519c54e65da90ef70572068aae48099398179744062cb7632c2d3da0fcc2b80a0f280e6aeea01281d529f595355da93847b2a919d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hfb5fc135186f30de93e3eb460f9925bffac8960822dbf32ae90803b3cc7b78cedb94826bc19d234d46e51d24ad2f07d8f9cf9159281fdd7254bfcfbc09e223bc76bbde82c6332fcee9c26461e945;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb5db542fe6c1af85b2124abe276877fae0997d78c75be508f8ba1c1a7e821150d8d9a09bac26cea585f809ee58833890fe2e6fb8b3d73b851c4b42f969bdc6c57d8013d7c0b343132965afde9b19;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e21193a7401871be5d6292c93a3685ddf4e9cdf5ae5edd80f07765e110b69fb4b12dbf30c84b61eb75dde08d744a5526a9a97eb5bc23582576ba0053659e8df313024cd2ab183b384045cf2d80ec;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h13f7edc3a9fd08e215c0925a8d8ed3f4b8174993d945eeb6eea42f77733742ee316c043604941db483167cb92ba18e5064594a5b0afaa09bc06873778c81d2f0b67749a00c1f4156aa10416fca133;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb6bc10594e604599407934296757b461e7af99e7a1fc1e1bafdd700aec57b85f41004de9ae8bac63c72f44d1b0907eaf736349cbfeb0cc6fb1c2d438516eca7ec1cd340fe1a6c6440a9fffec1b15;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h9dcbb76c6ff35f3a5f7f30b74da7a69b84965739453fcc5ba4b62f3041ca6a4b088393065a8ba7840445ef17678235e7ec9d4ccf2a840bea2a86795f541b4343648c5f122bd75f0942d2374081f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb609f56a17c0f2d75c74f325d018ca6e66e394f2dd3562ce67784f665fb7560270536c1e1abfe7ccb51821bc7dc5023825ab3d4bc5653317870fd8463999ae202ea825b91473fef08f49b2f55662;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h5dabcb3217591134447c1e34d177f68173644b6188e57e8be290cd7b4cbe1d3e989d0e4b3eaa05c605ab79ee986ddbf9831156b0f3bbf4889055c7cb756584603398a7e24f14b9e051b6bfe4984;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h4c923be0dcb3c952b01cf61ce86dc92ef71e98c16c3000091dd48578c839fcd78b335b4d722d405957c32919c027767288335cc4f39ea2e1662c320f105ba7302a91bcd3e26065cf5d8b46056bca;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1434f30c6766b0fc96107f1749831000151e16abb4aa49fa9d26f044d0f91002c33bbb72b38e7c0ce97c78b6f7e2f0c62267ee8497991280a603b302d19fd42a6f8fe81b0b2324ca53f61ff05492f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h9e01b3c8a5f9026a81c9ba9dbb62f0b5567150885378c2e42470aaa8de92263c443ac89c181d4984a7f1f3ab1f108e438c58faf5f4240b0cb0bfc0115dc002a297a5da84d4d183d4d026abadf7fe;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h11b72fcc5a6b7358829d05ecd9787ea2218a26cfa40de3008cc2ccb4b07c96b667fcb9a56ae7a2034ed38e8cf0612e0f50cbf3d669a23fae6aa5d5d644c30e0128fc3245d17f62b4a5ad11320b619;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h71fd218374de77813079c99f7ced1c6edb7cf9421b8ba8ec2be9884f0aa417eb019b12891342d9effe8eefe574417a811b4e5c9d63519ca12ba076ee05b52d98e8fd48b52773a03dac333fbe50a6;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hcae10ca3ba29392892a78c4c25de392a3a1a346f4fbe8822782028ccbb29da04cf09bb16a274b4efc59a5adba738cc88771c45df36ba261f87ae55e15ebbeb8d6f080a4161fe6de7e140babae43b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h189bd09d1052c6e075881cc8d0809814e655fcfc52078d17851cf78d17f9e18c9763eedd93e94249b953216ad81c141354411735c4f151f6de66816832ffe0fee18ffcbbe4e73691c5e3010b2b926;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ea3d2f6b019dc62d071a27443a3e55c0fe4acdeb4f54d7d4ee8f060c7c932f4db20011a104ef4fcc6b4d5bb2c2a25053a3e674d6fd64428138b2f76053ccc99bd610f91c256e69ce8517d31bbf9a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hfcaca9cfdc4e1ad551f120d6bbbd87998dad82fae194c3bc9968ce8444f8abbde40460593d9e38bdb68f3777634fd055ecba298d265a73535a87138a3b4f4661789a7b9a19bbaa8218048cf5f26d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h18e4c238e6f6185ab65951dbe0c4f873e6510e674c8ecdbcfca39c62be7a9960b4635c16f1d0410d6dd9014a88025f00359f434744e665b1f66e9a0658b7dd0687c682be64a865780c7cabaf913c8;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h128bc3699a5883383457185e4d8748da713820e1a5eeb02f9832fe26da1656c724b4a0ebce8c43ab15f5355a35cb6cdc8038ded227c19b8671217670ff8960831d187174f415a7bcad5c60a0e7b4e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h12ff7bc1bdf28140fa4b536d0e85247bc24c0332feaed8acd90971e518d8e5e38206b9a554093e5406915cf689966d8a3223c75be631b2b543e11cabf3478ad0728ab13b0a136c7fcea11f155a815;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e1cb3c8d2491fa1e2a3d57f834ea7d7df313923b0fb65732f001fee68bb1362f827da8b50743f3a327da1ac288158813e19911776d20ffd8dc5fcd22d9ebbcabecf7cefd4beff27be3a91ce57677;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h15f0affdad6a79f771591675efe1c6289186879fc73d3969a0daf765537255c669697af800294e072c43c62a8fb192c3b68ecc9c41e7733135e8acb7683113af5508db36a9f7cf726d8da7d1053e0;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h25f64da3f4673bc6eac774e459ea740df61de2ae827ea77941c561a5d47dffbb181fe94d0c3f62a297ffeae0d6a72f1e7dcc2dbad29476031c49e444d07dccb2f2a8b6af87cb329310b4161e1eb;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16f2c7aaaefc386a199b7d2bc1f480b01f974948acc51a71032d7dc4838c8e64afdbf5102d7ed666994ac6643e5960e5c38bb8b2a7e925b88ec36a58c9b86f81cbd6ee81fcb98058178f1aca29aa9;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h15c6addf45dca4f56fbe27c8c60265d699014773f1b3f7e702c931f494086b78c5d0c798d7ab9d2eb6d26c5a0b2f609d99cca9850995199986c54749cc7234f359bf2bbe6358eafca8dddba46c4b7;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h111c6dc6f653fc9ecf83f727e548be13a02cbd3685718152ddace4d9bf36625e6ee4a7b72c4a704040d44050ed0cd6bd16e9c7fe01e576ec7f98777a1817254bc9f3cc5bd23c4db10c3ea81c4d465;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h44dd11824935e1cfb01dccd8d36f478a477dd70ef894aabccc2d1956c61f808417f218cc13b00459d798cebbbb9ade54fcb7250741b1a0467080fa35234eac4bcef4471761a9766c9c6811edf883;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h9c39ffeba2450b7aa30f1100abb1aa666b87238bd577fc9d860d24354ef5d14df944ac945a5d3007324394734098b94a319314a7083b51b5203bb0b8f3ba94d4d04d61658732e845c09329528cc5;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1221c31d3358108e0d0b1466e0bbca9f0f9e25e049457f990e30b978442d8f08b766e40410a57f50e652199ffb210d33cc247d90b1c37a6a64ff093c4942f0f2865054f4e7ffba14a4e6606be8ebf;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f1b38dc7d124d857c1abebe1170dcb6028dddab4126155bb8c92eff088f4c8dff6a67393bae5c0f58cf171a81c0110f2e39dca8264d31c0d7f44eb79478c4008f0cc3a0f7b122fd1160676bf1999;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1dce4bc1cd407e5e4b425dd403a55e30f1ed2739071d26bd5aff82407aed6b910b39ccfeccda95ec6317e80d3618fe9dc52c8417715e98f329c5c99063a2ae17d7d2ab5844e3ea911bf6b8501158a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h68a0d1687334d0c2b1df02b321c5a3342d3650045d76335db5c2340f2c90b0dcf48357641a6c97adce2e358666936b90884f2836fbf4277cc601754538e8bdf1db50241f8bfbfcb5f1d0b792687a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f2baeca394c7cbe5d01814682dbf6b3374398c228becee3dd39cfc4bb8ee16dd644fc18675058778dc376386ee4a73829365270205fdf40224bccf1ff0f7591348381874f122e8c1660b805e5106;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb62e7c2eb82f3ad14657bd39290c51a9862ba8607131a2c1ee89ab3b61711d5ece422411688e292d74d81ff32229c51dd008b0b23cf682da5f44ae98270b74fcadea0eac127938a5233953a1122d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ddce03764d7f951a03c86be0747b328d0d113d39f86da29b28c12398c98fb48623dacdc216fe93e739332fbd6eea15efd349b1d61b8319a325a8009fce2ebdd84791971386f3a174bbbc4b36d7a9;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h11b66ffc75d7e33f5506f642da09cace6eadf89c78762b46e1ca2a0a4490c3c45df54acdc44f36ad89854fd4a09c24a05801c1e6303bcf1c8f6a3aec238071b731392a1480613a8a3871b926c42ea;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16f450269108e50fea6cb73490ede7c79a1a32ddc0be82088bce789c68138a24bef6bfc46a1b5e17d77ed70e66ab3f3822a91c0a7cd095a67a2f20559cfc9c1eff83b850e217b68fe677a89909718;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h69b27a78c8fefd2b7523e2471977046706de675ac464e7941e38bb41057cbe40fcc2a6b23e0b9a7ee9b60b1c80cf5dc5a3570ced925ce5074b2a3eed42ae932db78c73ad6b672f107825c98be40b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h97561fc44e64d77e7a609786406c72935a420c58f493b3eb48a83ce6307e6f8d24ec47bc4e1f16975d3940717f2d5bd46ada0f6655f7619d1a7134c53f056ae9606b5af5e8c3c7c9696f315e5701;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10132f0261340ecf640a7c58d88312c2fe1aa558a97da6517b799b8d428c02af97bc5c16c727a925ef641ae31f974c09d99b1d6525a73e515b4bcc6ec21a895f3c81cf42e09f1ec5467a3cf5246d0;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h145a0b73b8a1311e639fe9564bf3610be0d9eb1d8e629d96e04f9c511db4d4330d6038677255a007b04b5a9d0418ed39be448a47398a33ce79de42ef0feff8fdfddcfab2e1c19b0d212263e0ca97f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1197e5188a89f2523296c78b7025ee32d0882cf062ccf3db571ce61f5c8f31ed1db79b058acd3c296ef5f5d6d5f8cc090f6be62f816e6c1e52261191e96316985bde1baaac1c779f70ff9bf459ed8;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f86efb102946ac334f30dea745600cb49afdf4146e0c519eb15833ae5715884d77e3cfce636ad6b7653f3c7468f2aea2409c9a89ad9f944dcd67998c8759fb21c9efd81c0e59386050b53c32f930;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha436128375676634d61607c60cf52bf4704ff76561133cdb8a21a2dd336e0ee12f753739f091f2afc07131bbf81ef61987867a6e5eca49dccac41c183ea7bce13519a326df6e0f1e38286505eb4c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a1f1a6245ad5e54c137f153b10e7e1eb6f4112494f802391ab4caa4eee75eec04d7e35f7ec1e0865bd8384d14be632e72ad56170266c94a11901ec26920cf1b5a57700ddf16b5d25c04793fc965d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1751f2ac692435232493099754e754a3bad7de56d7de66be6e1dcebbdd9d994d5990f6b5fa57a59a90404e0b4c1191615a8aced1abb8c422b16f4612c4ca6473e3a9b81f8d9d0bb94e62596a1ebe1;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h6261d591f9d65ec07cd68fe61cc800d0f23c34a0ce16ab22e810ac00ba8c8502c100f670f462fa3df5eb9f65018e6f34b8e65c1417ff4d5c69fd283ae3acc9cd9dfa0ec0df87e4320bc9846d6735;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h6685beda7f994f7996e8ed158f0b165c62b08f6e56cec5b13f43ca42a4337a0764370862b7604166bef860339ee535e9cc35d2a4cff4f880e29bf6240116c9f3faa6bc5dc433d99da27ee6b82cc0;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb74c9cd880f1bc41a5efc6a43ddf14fc34c84fea01ad0434b58991ed513bbb9e42d2633cc74d5f51f833b82bca6fdd3fff3d6d2aaca0cb3e1664a17697b4c6fbaf8c95c2354415247adce45a1a48;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h193dcaae6d9052bf6532963bde9e35018569869f54cf0eb8629346bd6e09710037e3a23b7e96a0c4c8d5b8918419516c89efefca3e7304f87b8522ff013db0ad40d5ce7ccca030b725f13f6d549c5;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h2d4572fa255b4aad17c336a29a3555669b31e4cf8bae65d71964790f729f3f8567f5210eff5f5bb7df995d3af1f8beb1e9c74e95ffccf9b392c1243df1a91760efb8fac91c77c10a65a21448af30;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a2f67ca9c5fd9c97ee26e049d56bb98b7ac55d152a6744e2883696a6bd130244a41fdb9228d6e9f7cf32f8228d4b72146adb2fc3ea9f163e1482d2d74f2643e80521eeaddac696cc3952c7e132ba;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1eb699047c33b8e8c3d4d3fd2823e16610a5026f742f63fa44d001f5ea7e0eb9c924140d9b965b3cf41b7f8e65840c18360cd57097f7036a580db2d1eecb201ae28c3bb848766774eeef08eef961d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c92da404b6560a7199dc1867725975788fc029aad6ca9342ad1710dbbd76b71ff3970c84cfdbbdc1336435671469882917638c0aacf86fca77fb4f81585d721a2bcc6fe42c135918e9177e6bcc57;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h488f190be2c4f0fb15faee69b09112d2115c52f610db0fcee7a4e064b420da911d22ebf4c676fcd8e928655c3a90829b056000f4875aea9006ff9c271ec1246f0f379ff4fd5bef3e343677794a75;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h12dc929db7262ef93e24af513cb3f5fa5610b445c8ac80d297a883ce0e9eba436f783d0fd2a17daed8db3d8d0373a368ffcb4842b1862f29f1c57e9a9c0057f29881511c8e88d55dd2fefd0cf19ed;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h135e1101cbaf90454974145eb57ba5427505b7ac3290acda575ba13dd657c5d3c09d0522c970689c4ce85e987a6ad082b32981b4f46c36d5adcf3e790f06a9bcf4e82c9875db5940884f4c48b4ab3;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h5368edfeadd33889961a5690f6dc447b9289c5882df657de63c427c4e1f56005f2ea2245a801a6cb70c731b4d47d8b93f5850b91d4c0a8118129455cee21d9a5942935f45502d553eacbde3dcc82;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h8728a1c660be3251fb466aad39db9893b82fed5883d64e003137e24cf0ad2c191001525128c7bb6c2a2b38b1a47d8cb5f29a7e525f73dc231e5c6709a0e738b19aa2384a14b6286c7cb3932732cc;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1008a6c0e569e814154e613054b937a0520837bc59047bee73cfd9f91834ef0fc5b247eb240a993ef8671028713e597cd7ab1476267070ae31324ed6d9a6c6ed38abcdd1d8f36824ff4a4c4b1d411;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb799e6262084a0fe05cced864be87d815da36c20248675111acf38390c03e418261bc37758e8c05214e6db5a7fd320c3ee3f45061c1d2eddff2373dbba3a1a432045ae95534fbb95de7d3335c92a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf6f03177768556619446291c7da7528fa27fc6e9b940f405ebe233ac09cb1f74b6fa991c9ebd9c5601351b4d77756bf9dfd18402efc019ae7445f7b59bb012d9919a8bf4b1cfb3dc8d214478b697;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hcbb73f49d1b60ad19a3d0c61d1ce618da5a77080020e55692d6514e9e9e6c06a98c7ab8fd6b26fb2cba265031af1cf21737ac33a2d26e9f7ba4fb47f052bd06f55e1619999a3f514e8577b44a4cb;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h40bfacf399eefd0990d069467680f6095dc19e1a7734e2a7b48f96e88be43f7760b8fcbabb43056e873b175364be79547995c096f6b55343fa56cf23e2444de39add9a29b7a478288ca29354fa3c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h14c9cc66281204a77edc78240d7326aca547a3c7748a7869b2477c628c5b76ac53ef36830292b6d894bf395da4d3d82d7157e4dd04270a6012bec1031a95dd9f6238a76b487679145d932c59e1b87;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hcc2b87d81ce48b45ea30aae94e660a189090e5a37a08defb8fd0fdae471a6a58f2f792701eb41d51633b6445fd94e63a3ea32e490e4557bb860548f558bfd2101cae151ec8f860a10a5cfe4be90c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d75ab3e6e2621f2310b20c347b55aa4b06260c8381fbf90c821cf3d99f465323d72d6d0c2130baed6b141e0fbb4b8b0117bd2a6aff5eaae462dcba03251191e4185aa80b9dceba04acddf15ddfd3;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h165e06a65f48a5f61a66579219c20a26dda53d4bb94422e38fbc036551348ed7a1691ec76a08dbb9473a3ab11814d982d54516f4e46ce350f25dec152313188516800bc55fca961240ba4578d08a6;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e1f21e560cdb97d8daff7f20c2813d8e6c0f425223e1d3aaffd27fe514acd009e01e7938511b91912cd6a00d419e6ed958a56b0b448ed4951bdc736b5ca34f1dac0f1a951202f7e62d493466c7d9;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16c9f2e5de4b48337dfbaab26ca15cec6aca52d9be1d368ea18e70615ce7ed24c0c46c5c0cb58ef57448fd285a968023af0cbbb3698998569590ee9c283c828fba0395f9b561a425e2e797e9aa577;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hfd88439e40de49ca7bf3df33cffb3d58cdcfce3805490793ba18a74131133780575de7248ed86bf085ffbcd3cf3f17dce6c30a2d2b13524c92b6d266a72c9a82ccec97902a69e641001083e3daea;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b535ecf2c17d478e34227f4dd3ee513fc993a0b9a1977f2553a01b428523cbf70875330e93087cff46133a8f552c809645caaf52c6dd224a27080b129cb8e9b2654c363010da1805b56c14108b47;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h7b61251c7c52c31b2e7f7e8480e4dbe776e49c68490c3f7c8d7aeab308a96d3f3511e97a8b0b24d8bfc2db5913590e8eee0f2ae74913f3f6f612e8174c820ed482c657c98ca716fffa49c29c4f3e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he679b4fb6304fe687ea120c83b6b69e66521f2bc2e70e124dc9c0505a2e58033df35c2570ee8fd09c386e431dc175ef71de832919797ac63cda00278e005f7add0207af530a6dd7872b43fa2872d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hdee086d56f7049817e5070c8b1a8e91b2b3917f4bfe21c4cc4c215b6aad9d625fb9bb56f7cc674ed034f89e687d48829af062c7ce60e5b639bb3533d6d9938654293e5255398b23c7dac355fd33a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d46f793bab3626051799509d97bfce8aba36a083275788c4740940cea86ec908409f7f8550b6c8dfd14011402933db547915aeb1e6368b5c3cef0d21ef6b1fb3983bde84c278a054ece3390e4508;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h5b201f87981ea119e754af305e3dbac37e305e9590c73d4c00ead723d1de98aec02793547761245216a69e940719bce0b2c7dc5623b07ada60022cdf27f38d8e546d0a174328c99e0d1965e0c2ca;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h120d0057ec54195ea36b34a5b1de3dcef98b06c34200b6f49e01c0357283430b73de567307f50757e64248b7e57a23cdab4d4c2ad6e09c6807b6566e6c8006cf8fe7756257f4f409ff57b730c11ff;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d41af6b4f34cfc44392bd2b591386f25027c2f6d7a4dc8490e29d9f8146667a84c2a34c8ca41f03f06bd688701f6dabf2e2fa25d1b411762716ba713bcec0fcddb1e95d2b98ac53e7fb5a14179ea;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ecb9a231124550f0c5f4ea299c5d51a468929588bdfeee7ab63ff274f3d43a210d1366a8e270938f066dcfd1996fedf4e08970dfdf26316932b245ad2a55ddd14720a2df9b9a7b2cb3ac902d2cf9;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1edb6171f29edc404409016ade19fe7fa76b0419576869ce1ffaa9b7cfff633f93f69802f97cd8f6324f4c69ddcda26d1f202dc386dd692e77d89f836258b842fc863b080aa0101eca491fbe9258b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hfac078ab96350ed185ad1fa373b50d6c9e3f7fe83ab7aa861ffd69425abaf242fe30918461d82fab41a52c78fc5bf5d0f207bc3e6904192309a72703fdb7e135fc48432c912d280662aa783841f5;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h5e8bdabbd8449bf653dd7be27d67bc28d978ae7f6c0248c4669815feb8ed0abae064fdc5b3a7182363db6479fa28d20cb2e70db241ec43936c46927caa25ecf743582fea467fd4b0d1c3dd19efc2;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc39ff581c5cc6cccf419331b1c1a5d7bf80dec84c7e4ea9798869b86c64e31fb9d0a72b25448b89ada67fd209e536d346f83092c40ee097936cf9430319e9017adda97973230dc3f1dd0bd04e7db;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he1cecb1ef7557e6f5dcb871f3091567ac78d66986e7b854777412bfd85a3f98a4f95f8b53c2b6bc25dde8bb36390458addd554c842f551206a396d29b6b8d5002ac4fc7b351b5a37878bee1c640e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb9d7ee7d8ff186fea629609439cc30943ffd38ed8e42611ac2a1d74af463f82c55b12a8dc62158f302177ac780a05d1d18eceedbbcf9534899704b11e893c82d6b49d5db5ac2dd9fe7d9b30d0d6;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h28e8a72f80c7f2bf65b9182c2b6e2f749103cf6f6f7430153d3966acd92610e0b34bea4e9bb5bd120ffb63bbaf195ac7e88e072f2b963a026251959b26a27fb0bc8074a72fc55f96a0870e68bf43;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h164c5a09e7ea9ec2228cfd333dcb8bd6ad730779e6a6e7c32ab9811b75dda13fa695393d40daa18093e18974a472102d08be37acf3072a63b01ae52676e00ee91a0fd6432482b0873ebebeedd158b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1520253e620561e0851626124913e44950e63763781d9bef11e746abdac1d114740a7d09cafb50d590032411a8d490e5314e4fe24f5ff548f58f53105d4f0038c167d9440cf06a59330e1b4ac8e51;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h18410fc78ca4e36b67b316606f8d27b2ebac98d90ed6ec149015f76eff3a37a185bb20c8ba0dbc6da1e90f108a5fbe07eb9fb94461a2a2d16df20eeb6fee261c41cd8f0a08dd27d10027c72b69bdd;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1458039bc7118721d8f71abe41bd615812de1249aeaba812848d4fc0ebf16b1731fbb36a5900cace7c48f0c916e24c0d7cba056c7cd81dd8638db9bce64183fe8e6c29de41720b7bac3876dd7a6a4;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h150b8b51b1b07b59fcdaf5815fce49bc3ac75991c6c11322ac2172a1ab75f2b0c070ba74f97080375f8986c4dfcdf28369ca9b6abfdbea7432a1942840f4b05ae6aee2a19d211b45c47e6fbe5474a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h111be7b3a8d2e737e3fdef0d5da29c70c43a3aacd948a3faa855014e20188b7a9749c10a574188dd5acd98ca333cdb64ddc6f73451da0ef6b28d602caa7973844ba748e8f51af719ce10dae10a136;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h4d3daf33e02f065dd2d809de879628fc08e43a899253d617138c471f340ae93d0d98c4ddce999efbd5172da70412902f04168ac91ad0f879960e78687ad72a700680e25fdb280ee5d431b1c76131;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h39d1b4780f93919eb4598017e87e2fbe7d56187c13571e641e0007f333b08c608f0585e37fe3c84e57e0953baea78249197606556f4659326e8ab916d789fc8611c7d92600d7446aba14efa82476;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h19d2e056d1341b656c4aad7b7ac4848683d846bdf1708807df4fdd0713b468736ca6fad8237215f43e856e8fdeb70a4613f64ec5f7daeca1e197db3d90f8c7bc2bf6ec14ab8de200f09fc9bb5b039;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h4ce21fcab85f69c1535ad871517e6bb9c24a5bcb984bc3c332ac051b553555a733478de0ed56259de6836561a9a17037458757304e9051a7ba15c81f30610efa16aab3c36fd4b87838dada11e0cb;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h19d5aaf6078c58e593bb089041b706d921bf00d0a931368ee75e153166badce8844087866cb12d9b20941835665541d28f748810b0773f6c151221ea24a25710eb1bf69c2471320166bd30fba71eb;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he0abc0fe2e989d54b115fa3dadf7966dc7816e5cb1083502344eb9888b275ef4a78f5513c1b2b80813383f6bad1f89b6f4bc944d55839e48b2959a970c2ab4c2a70446caa676558436668c7d12c3;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h17af45a83fd0b823b3a29cab71fc0209bd1c3ef6f429b478504e16bafd547f655a1cd66cd18f32116b8a015c3cf87c38b00e29badbd73fb20c5a0f6cef646c80be99728288ea5d70fdb662038aadd;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he0fb7861ba63013d4bd9262e91428f94b95349a5775f188d42eeeecee4e8dc715efb09ea628fa5cf7dde68a458c1412f11d56fc623b48121ade01e3c1b86238085b1eb8c99850bcfe375fe95d042;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h11ea98de861e11a9fb30d7d8e5a84b1d2a8df05712740d312dbbeed72d8e42bd1f0628e7ad3a80c0ec70758784983ea9c55e4bc3d0721b92aa84ac3b870ea3fd60c4ec54e0333869cebd1d20c7114;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h18c663e325bf496a3e8873f1c6481eca5a1f89d6a20b936d463e96d1449a82ed7a7f37a1365ab3c59350101cd7bd14067e9571894675ebc0323f3e329b44309a1ed72c7ffe64135f25c4b8b3b78b1;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1010d25c64aa819dd3e542cf604794d5c0d758d955a49930b3f3f94ccb0f26e6a83cc3e74e3cd30854e62d61a28e977fd88a722998c6968d11f661b8795c03ce0ed5adcd0c34b4f8c94097ba09e8a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1396a287d32b67394e7e6fa46b4d7e4a69f0c985de6ca216c4f69959713aada2b5105a3b2b5d8e48561395e4a42b464ef60bc8e49f4d028e754092c4c607b4f6e2cce0b13c29935f85f6775e55ab2;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h19a6b06158b045649f4448f6383c38ffa7e37f6c7f4731e8b7f1c261431f01f68b0b0d019bb37b2d57ce43b4701a8e55f1a30f78c81e20cf03b373b27941cc288a743e7514091ca837859107cfa38;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h15ffe4407da6dccdd916fa158dd2ca72d2e3acbff8dad590ea24d9705b5a8e20ce9aa7155830578deb936ae4e53301a5b213feec549c1d0adac92492570e7e1aa50ba3ac82e1e21342f00e2411d6f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h199f78a6b942196f9c1ef98100754b6484592714be692dfb9f2286955bc8574985c7f173634ed93d72a314e28729e47f88bb58168022797526fa9b98a9f6ee3cf8adaecd6eac2213efd56afc2ce0;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e1addfb81ed2df0c5a49495e7860c85d07e63785cf1b6670bc1fd82162ebb7cd649bb64a91e972967a624593e8ba306a18468a2ae4a70cec623c4a9fe7760a80c8759252d7cb9c1fc3c64756a936;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h29a426b7294e1b338fc470ecdf760ea9491094ea694961dec9ac64e8ed5f96e315e8eb15d9e7602b23f74869a88323211af67c5d337c4b4295e978da99d0f5d4da5bed9993d8aeb92444d45c1ff2;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hbddf4b05846b06f44950c29077b21d0958720e85b9887d98b0988cb19b94d199b2eb44c95a5a80f807ab8fcad2696f28eb7e06e91c2471f815f59c26206c8a9d023eace43998d31be4955677ea73;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h5ebf6e9cab768b1a2d5b57e0d95ad080409aaafe1acb06c5952477a8a219bc3bb575e37384d6ffc7e6a6d94efa4144c366a1cfbd3c8d7b8e6d0f2d1facebba1c61be085e6095f27764671e3447ed;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1763f92f1f74bfec8596c4cdfbba0eebad27cebf85aed6714cfc78bc52e51b206938fae37a24e421f4802db453358fd3c41bff62bb2d7dfbf382c4ec8025b9d155c8170a5a62c580805f06e61b8c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha0afe2581125ebcd799370e9c9db67852e1ba929d32526f537e3762d0ad38a721b70e07dc2cc89bd291b6e9551b00d5295f3f12100b9f0bb8fa858b928b8320b073bad27ef49a226e1f41a7079df;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h85c69fd2c5252805dedf5b20764e85625768c5aa292e6fdd2a2099a8d4e2d6b6675d49062c53132eb80ea564b264faa69535138688cb30e920c32a3b48a395c2d229349e1dcbdac11ab7c2815568;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h281ca86dcf2942dea50b97f9c8d89c066902dce42723120d5ef7c02efe985076f19ac5e7e12c30e414d651351a1c25e07f6537ffd6ba25b10e512f97d22984fefa3a8cce0c5e17a2560a885870cc;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h17618d69e6b3e4d41bda794ece7614dd7b11923a7d7ff363d8fa7a4c2581093aa0061238bfc16ac3edba78df1d380df8572e51b065a8815ea63afa2faf0f37060758c694d1a3f2c6d9c9289acd509;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h609455d3780bebd10ac52a82fc3268c151b130cf3dbb73b7a46b31a63d48a5c3647ea82f7fa31a92b0bbcf1c60d50fc4474cd3d6678e50d161738d42f6f8998b4832a119250d9d60ca4222ed213;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1bfb54374f4021e45fab37c6d5793c853df7cc680904d048fa599abe0c57c33bd85f6fd6a98103ba2122a54caa44421bf456c3033eb2ee531b74d919400fd7e5adb1abf48cb9f147105f54325f465;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h18d22b80ba7621f607165a0684d0c0d36c18da7f394ee6644dc8cfc752510d21de659e98a21e580c6f7f23648db0b11f028f567b43d1065e0506f11c4ef7f601e94912d44f152285791ae3001972;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb84655a4a615e5b5bfbd3399776852c26ecd693d4d94172e933f48f3aad2a836dea404a5ff9022752ccf6603dd8f0c294b45c9a42a7aa99274998ab9aff4f101aab6fca17873e55579de1cff8c3d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h13772c565938845bb7f2f3e95e8dd8a3125b594f7141011d955fbc0484e6c65416909063f0fbe858142e6933cda6e646fca8500c39f10f7bd0ccc8786a7fe351f3a51457656e0de812a6236a3648b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h3f7b00cfb313d87fea297d190129a70c99441202f2c2028bfbeeb6ad51a733455d7df7138e15c92998002e567aeb9b7f99899f2dc996afb8c35e57da0af41f040bf880bdbb42f61259ba9fd4d4ac;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ab2dcdf1356fcb36039a3cf37efb2e05296df1c7521ddf6fd655cc22defa38365be44081d82f127a5b1b5ed3e347cabe59a9dcb1737839395834733fc8d7df476fef0768c8f3235afd11622f84f4;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h115793492387ca12738a26dbb2adb888a2f43e0b47a618b4d6ec1267872d0eb2feab0cf21fc5699789dfea592a21b961b50ca1eade8d6be5787d3bb3b873ba44ec696a89d683fdf3f4492446fa1e1;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h4d54644c5f9b884fd976891a6bbf8f722d211baa17720abd603b617baabe41207f13f0118b011eea7e01c01769c269b6dcf54842f838466f3ed56eabe7b0eaa4700f8d5c4fd3bcd2454056e52ed1;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hba8a98e8e9a4706c4ce98173f4491e21acba456482e668bf8f1d9bed8b41cbd63dde55c92a3502bd3c9a0c170ca507dd447a67d4d9901eaab4bad9f91d8bea97e5ed0446d8e15bb2115d4d907fdf;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h12b6b95aa53d3cf3747ec52ad12655da3a31638a86764a5ac45ad14766af9be3e09f4bf434be9f024375fd71435f77ca304fdfb067b60453c0c63997e3bfb60ee2199bbcb70973ab3e89f80b0f2f2;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h6d139aba7225c90374d1f52335994a460413c7105e83b88b043044d07478554a6277e509a30bcaeb00009b2640dde2a1aabd2493ef72beae78b4d6db8b0a87ee283913da3b3688488c4960e2cf8d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e815475ee640187d49486d2f3105f50aec411e492ece573594fd3fd713bde87cfc0ac024105d274031e5c72e1a8a45ddd02570f02ee4ce9e3980d206092df64e8fbdab1176e2cae0589eef5001a6;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h121bb8d4d82cc41802691a0b13f8d5e7bdbb5ff35da8c941e330e9889abd37deee4fcc88a2b2b66af7b4aa818caf721f187c27bf145cfb8c12bde73c0aae89c1e60e12bab681d7f3a4488ce5a83da;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h2b2c189928ebe12a71cc5963f520b380b6c6f919b4f292752bfdd137f97b7716d9b3e4f9ed2ec11d2117c4dca4da67cb378d41dff8f2736b69e72ec1e61ced474f724e80508d4c1c325e4be731da;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h159ce6035bb0c2b0693ec8d382c914da23e6d9c3435c29de22c16b7064452aae7de164695c692d34c79e49c7933a3bd065058c8a2bb4f52d9927782926246527306ad48f5c6b202390300b448f567;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c2d567c08bd73d32c67583dff3679bc519e75626432c8e711fcf80ab1c15d3a005f0c7c54e2b0424fb826cd3c8e32fb61b717357e491eaf2353f38c66948303c302a44bae12ef5e49fb1aafc79d3;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10c4c44eb3ec00c2f3a67c50fd12d9918c1ae4198ec297649cd7e56feb7f3c71305c4f9fa9f003217d7c917077110ed1b3bfaa26f1b6ae963a792c1c18c6bc47caf9dabe9deb26eb9297bcab297fe;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1910fc09d436d5a6135c9d17d40498936fb4dee53a4ddda1a836a2cb3c214f07987847bd0ea4217bf04c7d8c3af21570320ef6baf1f4a4d63658b00a84e9722dda6520ce0cec5ee144407fe9c54b4;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'haaa7d909b36d121443820dbf5541ebb90ee2836ebd220e5a19cb76a2e2ea543666c806278a6bfe99d05f71887b4fe6caf0c673ae8585f502fff0af325d348307f17b00725357be2128efe1fe4e8f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10a61a63f9fec46688bed6396edcb2d02e810cd33b023709f84378f960ac5cfbbcf33cd82a38fa2949ebf3f8bacbd63d44a42376afa5d11d8a7880eaa3438bf5b3ee2313e5b7dfc49f17f7abdf254;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h146905bad480827a32fb76dd077c9cbbc07ffcd6ba8b5ae2482f9e3f8ed5391a26f62f8195f5a6de3193dbd601a292a3b1aaffe073a40793464d1b4e54a7eb1d8d05689897214eacf9512f0b740be;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h20c6b07ded90ba283cb28962d68a2763a64e21510d8c70f898b03cfe31a0611b850a6cfaa1bb87c04bd4537513da21451dd30d56b51f8d43b0a63e80fe8312425aaa707a63847a44069b5cbd334a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he07dff6f9e7fff2e72f8a153687f2ee673d8c5dd473583014aea7ae01876f0cf5ae4ee1d0767a67b9977bee8961fa9a86ebd30221005a2f1c54d17d914a01b7723073b323f01c3a7ccdb0ed7e205;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d48f333cc65bd431f7d5a927986d536405273adf50883bfe34ba66d97e04c14b0d8e0072436eefec983fab13b405b3a6f38d10259c6cc2af8650831c4c0ec55caa95601ca5340e559f980601e5d7;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b1046e25320bff2a1b17f0acde915ed4d3200326d90856c9d39f387e2225892ac8a062532fc954a3ca284be9502802b61ec6a284416ec46ba9d538052a11f18cdf6593ffe4800596a88f12a23bb0;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h3b3d93cc750bbec7df7563963887e65096f31a58a05c156f580a52415b23caeae10681229c7fd7c3d0226f420ba7f0d5fa04fe64ddc06c37424cd03ea23173e4f19798e7eede26fe9387a7682429;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h18cb8b3864e9e870e3629c46f6f646ffaaaffaa0e6b2bef61202ffbf3182ee3318a5c894908ce6b6564a187313f2f66f15d3b8a5de1b2555460ae5030214342e0f01985c7e30ee499cc6ff1698fe0;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha64327cba4d9f8615edf1b50b7bc2fd4b2560d172d33802fcaddfd0edd93dfd1612a6fb3ffc312aa46a10a5249f7ef3629dacb858b49400e3ae8774a358b09ae15b2910bb160b67485e3db538bba;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h811a2dd99081e75dcfbf63105cc04b788fcc91f822ce1caf51adcf8a400878a575ef319ae998d2c489515ebeff574e7c5ec52b9b0a149b8d1d58b2aae9fce06eabb131674e10f2a403651b1b6d15;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h79ff76a2c246194ce46761b63434141724a24be0e42b026a5a894115226670cae6c776b26848abb2ee75e83083c8a1fb4834a01ae50b167029a913386f21516ef3d167b1078a02e89dc3d22e5720;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h7dcd6adfeca336dddcbe97b5dd7ef894a78b6f08e394c56482b731190a8a9091c33cafe43745011427e88d479516a05e8fe48e5c45dff4b0f32ab98a47a3f0779f18da500e9be3cc204916487a03;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a9e22acfb36d6a0473ac9ca094dff62e103446c06c61cc1c349e6f6a5ae192f936d2551731d1e9df0217619ea71b536ba2ac8a48d23b7fea3273e192b3ac6721bfacd70db39630289c7891b3dc8f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he14cd12f516b5c6ccd64c34a2ce960ffb59ba4ebce750eccef75dc1e9a216bf67896141b59f0483da929cbba68e6b3c2889ff4f86f666b17cd011aeb8ec04e55222af11f8f5b7a058124bd89bdd6;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h4420d5e25bf2fb47b00d8ded13e3441a4ce088663cfea33358de6590e3ced46a1ccef32fa9e195d0de4cc4e7f793d2e22e0187220d9c2c7f4554fcff14ac718c796b391208d3054d99e0f2a5bcdb;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hbed0be4d20b9b427014ddd8cff28260deb0239619512ad2908d35fe694e4b2a6b3255f21fb10aed7a9438a66163bac121ba0f622e7260d6bd0d3f8287990f9188f36edb4a37e2881a83a1323da15;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he72e98102f6caee353949a9c3ad6484b8b8d8b6727b3bac125922ba003c1277ddc0ae1a3ff4e15eb1898faa7a1d55acd5eff5a6662e001b38ac052aafae0c3fd0922ac2dd222cb3d9f5d18fb3c30;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ef72a3233b105d79f65d3c355a5dc6516bbbc5767b8e269de2bb36d3479c847f23f0f00eddc03187ccc4def8392043f9e7c6850777b1d26148e8701fe520e2884518b82f5f5523042be7bcb6cc94;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e132f65b4e6ea7ad13c0f352957a306c48b18bd69cf7a9bf452bdc0ec9192daa04570f1dc3144e9a9b0889b9c21f5945cf23dfc71d3902a746c481d15ce8d1eed9c76f28e4cd8da0aaf8e224383e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e5be01edaff9c7cdbc28b9c138736ffefd7a0887c6a469b6306699b16e8a66bc10e6e0f04624a12fb1789ad1f3bdfd6852d839e8c640dc2dc2298da96d93da4c81d5fe8ec97d3e431e3628181a9d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h145ff298802f3ff0637718a1b0201990d32b91a73df7bf503c77c34b4454a7e3f8845325761ab6c66d2279137fff4df57a3d4e8872490d1753ebdbaf33f32152c12d292870ef0528f68f4ac8bebe6;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hfc352cafe5f83b9dbf1e7db6822781f422dc2290033e5bc9c3163c46fb69e70f877b8ab180f7a6514f4a23946f41f16021461b9464288ccdacc250ff8710a53b85e3a335399a4c67bde3be3b667e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h65b1a9350e4935101758dd998ddd6ae5dae04d6b472e8ad511a669db2c8b72cf488de20632d5ce4de281d452ae80bda0d30a971591a2891ae773ae8dd5c2577747898a0b3a920c6aa6d3d10608e4;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h12562668a504af738740bcfd1fa4137ab62c8c84fa08aee135d9ccec27cde2b3a36b3c5a439036c3837bb0f9318631f8b8844e5558b86f183d20b5ba0b6f744ef1e528ccb13d96bef342ee56e0bf1;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e36b0f63878de587d2d1be02cfc73ce2a0b2ced598796574abfaf6ae6f2dec5a44b2a1e39438bc60cd8eb1a8edbbef6f80b9d448ae5f2ec073dd508dac4aca0f40ed09c0b5da82bcb030dc2a5da7;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1995f0b06052990e55c680637b23fe3d764ac5c61448d0f395c8a9dc45dfad6176b604b63fd628ade94c884391afff816c4be678f6ee494674457fcb96d5763b87669250ff6f245673cb78f1524eb;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h184af9fea5c79f83ce18648b89fb2faf4b36fe7ba64fabaeeac42d70e01ffb8fb2e14d3baa7fb09069478db4e65cd25fec4ae5d6b0a621bd49d32a129cf2e23e053de38107de7950a7f1e37ec11c9;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hcf1f2a53c9de6a5f7e67c6a46d9bf4a85920b562b0efef0691b81eb9b0d70015832776fb90995f94f5ddb7d0aacb111244c1f8e9598e7ea67562e34825aefc45c75c9b2e0bf20c02bada555dfb8b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h14359e5605a248f48b5a31989bf5b3e6a2411d7c3f714d0e5092de2485c4fee7981d5d0dab7470ba1d26b6439259d45c6264187e2743ca54064076ad2f24fcc47710bfe129e319769742a18adb1d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h17122a3e18daa545a9154f205ed07d013271d0cb9c278413749cb96fb26ae22c7a3311df953c431aea84df93d83ce5cef0e7ec6a3a07cb1805096521dea498004f05286bcd29a7cbc2da782c845ac;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf2a41f1f502e19ab71b677334de98084d01fc0d23ca14ed502e2539a1f650968c8d454befb7c79586324f1c42916ce8ee676607ac9fb39cfe2effea301954193df443abd51eacafacd84ba939353;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1fbe540591a74eb926ea7a81c486ef90ceae5d9d7cbc5284ade2f95cbc95b3849f9331c410162b5f4b5fa802bcb8b69718d652486153f26329ab0c92df85352813b958a396a350f3a0c4b61439d7e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd023210759f52fffa943dde0c486c6b5cfa791bfa440c6b40cb4008e72f6b0b53ccfd1b70d9e8fa81238bf2cd7af31088523dfaac98881551b5545cbcce962dde21f2f5ebce7fe716ce226ea0c09;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h39c1e44949ec75035ee20b136f4b74ef49e1a3160e15b8461f1e400b866010b4aab9f0cbbfff228ebc607462a4d467c1fd8dcaa73768fbe8912f741e77f530f1f40f77dfe6f721c191af26b5d894;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h4250681e1ae8d8df6902c9b306a175f83f444c103093a01832563e359b0118e5be72c385fbc8a16b46dcc8181108d3f7a9f7cb589366fa214dc737c45fa2401408c91b116ac739c0a33da8fb8098;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd5a2201fc0473ae3a0343698d4b6b88a89cd7dd42a677afdc213c657e9a21a4f259cc784105ed09b87f78eb598cd0946a0313c1a2c6c0f51fa8473d285f7cc1ad24cde42f0d94947487703a6d115;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f15b5bb6eb7a8b3d9c79ad119445daf80c1d0d5168a2af787cb95f0af6e1f6fac98e9127038664bd2d4b028bde2093c6513908202daadd4f4898c4d1785c4788993f14ed453c7ba7c73d61e82175;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1775bc31713884cfe773e09c267becffc8b09ee5cde786195c1181cf7ed413c04389a27bc9522ba5d5096078dd4f5602f5a55ceb0f5384a915838fe3e9ecbc1d8e8dbb1323f243e3563176391cebc;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h18edabf4b59cffe694874b3b96113e5b7e1bc0fc69be378f2d56fa8c884ecb15c58a81868de15c53e4942b3d2b20378c096f7233c11adeca2506198531113b02a619b9261d85406b23b3f077ef97b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h179b7c49c80028847deb52035e2e5c37bbe6cb11de49aca99ad11dd8265f64ea37a7a8ce66eb5d030a04760275959f1bed0f3d3dff774e2d7d2b6fbb90d6c797fe7a5408b30098eea6aa421faa88;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1003e58bd7a05e31e20bb948bbd18db2db02e9461e4031bf26b825acb891dba77a36fc15875c86ed3d3f799324804de69a65350acee6de8905c1aa7084cc96878e4c4bbd3f83fc29266410942d6e0;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h2d071b4915c22bf293f08dd19f656189d1fee4ec112f3ddfd95661efd5a5b13cdc6129e9b00f0ede812c1c0ec2f4454582ecbcd5d1261f7dcfd40ed9b5b1ac4171ac98e655724c63bf7fc689ecd5;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hefc12208972fb812c4cbc85a03b4abb2d7966149675b5e80ac0c576d5350abee746b00832623ce37702f9291240550a163b2b02d031a827813434e34c9cc955c34ec2e14ae9e10845040edad2079;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h8d6d1458436ca51ef253f7032cb12725e58b5ba2173e972d46b35f54018072c605e9bc1a4395d03816188284eadecadd99adb860d3592ce76a7f5e88a10a01d39cfaf9cc67d289563ced30c2860a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h11dc8a4d9b2690a58f656e37103a82ef73306f9ed776d1c94a8bbbc714f581095c8149944091f221a001141b0a0b9958ea15799cfec2734a49903235be8a63c4545dac6c35afb8980de1ede7972b5;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h18b597a97900ff04ae3dcac8b31bddb45569c89b4356451857d1c1bfe70b9f51b76b20de83378ec2d779358d7e629f6b5bde7c71910f174e56de654ca4fb7c9bca9f7889d8521080e57f3e587911a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1bc63fa9b6fab2c002a6ab35374e54a678fec48e56297f0e4a00bb78c4164c8b8b30745115e02b855ceb6db90a2e7e7604d34b4361793e6890f27ee0b272897330ff6dffb27c26644bc1b33115fef;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h2a0cbb0bf74861a1353d72afcd56c0afd8a01f0c416125a8e1cf5b4540af5435d82a7982724f1136fbbc8cccbc024721a400805862eb654008ae29b781daad5ced33dbf1ef6b750602f485447f3b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he4fdb20c149033ce16ca126a05c53b45382258219996b8ecf944f9a15923351b65be9f45b9a6259b333c2ef8f904e2a9d39df9115297dd3970fa44f92fb77b4b03e9e13e9835de7319aebc2dd24d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h11169cf305ad271515f72abf760c0d2bd9842584a4936455702dd0000e45e23c54fb6f8b88fe734897fde38293cb9e67a0b0ab32b75a6bc16b24bd03a4f53bd4af57a64341486e55237ea27fa7710;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h7cc6b2e6e018dc7886d9a70b316e9f3f8e5e949d48c4fb15d759556636fbbd4c34e506a886d138060c5deefa97b3226e3de5862c029ce28778e7e367e62154e4ef6998e91d522f5d9fc462b2de2b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h128fb6aae8e134841406401a8b2ba366a5481ae36fc304c4cebaad7d680426e8cc8c86c787bc0249166493d1145eb7f6bb045573f3c6870a9ec5dffcc4d7f235bb4eddd4360e9d6d68a26024995e4;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd5b259646818ec79f721583ef5726aea5fa4be688b5cf0b89d2a8a5850bfc9ebc485258611fa1d9fd6e50c5ba9b5ec8071dd86fef4829780de67f7a85ce12961f0c8cb55b14a6155153a068922dc;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h8a7101c30758eef29aaf5a796325a9139dd60ec59b9bf7385685eff3dd001169bc6ca3004d11e33d68ee3b832ca4d1dfa9d14631d6b8a0d96d7923b3f235ee5637270ca1ade45242c9abf31cea34;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b014301d5fb2bdc8bbe4de251a94a278eaa90b9aa5c3d01af5986f5be1438fa2645e7127ae336d09d2b62e728fc2a412f898ca92cc55441682873244a5052034fa87f37c9a586023679811ebf0a8;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h17a88630c1d008b5e449c7f625409086c62e8b93ae440fb5775ccd4ca1983f22763de6d20c842909885ebbf0667335190ba7467daf0824b957dea23ba04957cb57a1f7fdb4df66ba9eed827d667ff;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c0d3d75aa8a3d5e400fd19a71faa3787b945a90077e4a6ea37993c0a93e432ae859b85e9b6bf6686adc0c84f0232b5a9d488f0635fdc129aa96abc7579265f9dd146a92d5d43652ef012190f9196;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h192501e6afc4529562520e96bb36c44bb14cdf8d9e8c04bb160d000d883e1a49163979818ea6fe8f5e53f6788dd4f577b7c2e8d1086e8c2ec71b78d266478dd797ce5fc41662e53d1200c43c0c70f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h12cc0f1fd7b6be89387ae3eba87e32c81075012e76b70951609f242dbc68568b93c6d7abcbdd461c2fb0650f2a9413d67a6344a8201e726d475c5e294a9239398fd2ad64441f5ef01f4bcab16dffa;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a8a01cc2cebd10cb3365871c24095c5a36d3e0ed5ddcfd970b540d444d4455d97838ca8c9d148b942ecc921047b204d119a2eaafe323f9e4faaca97b46957cdae729f9f98e443dc862b49e1d2b5a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h11214d45b349d07b713fb4accf7e78f02ffafd14ea0af34f8be8b29ecede428c0e32b52c2e4247b5d6e80fdd3abfcbfb951f0221efe0fb3ee1b7e045f8995649a9902cce51490eaf74dd913f1daba;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h111c7e81eb1d9cebbf65d5abfab32cd3c2f61d532f046eb5d1a23408841e67f96bdc37256812a0d2c762e9b7fcf8e39df7e9909c1974953b00e3d11f33e5690b18eccb6b0c975e7f84ee712fd1455;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h170e845d31af0bb7a1bc9fa67fc8daa072b87c035ecfc305e79f24906cbf2fdbbab5ab7462a84e676fb2cac647b3a1cb0a01c65cceccef8f7293906d216511005bbef1c655d8c352a7f942d9f9def;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b7e2517de7bf98dfde4175f3eb28ec85a9535709c8694e68f9136bda91f9075e56d3255df825a030aa05ea4162216ec27caf9ea57ad092993ab795695801da4ece090e0e5819e50b71b2ea633028;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1338ac7606f93972d1e625feb77d432e2cb07c192eaa5a937f28d8dcdf5dd59ecae8182fbb807188119ff6a5a97b06f2be5326dfdcb8d5b234c470f506c13cf263267ffc4e3ce9a1805fa57ea1e35;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h2ce04dd9c4f0acbe2bad34faa28c519b59e7404fade1d30da84fd783b8716f21fa19a0b5505cb58f60b272ee3569602de0d026ed9001ac6a70e22a17ecdf4c9871d9cb3a9b84b843b669e1d07ec6;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h4e7459c5c1caae3bd58242362c5fd340053d26981e6d3f16121b76f62fdd511dd8627c6cd21579f6e82aa7ca801f0f17e624971d01b9fe6726525bbfa0f4f4dc06766a591e4470e113542e8648e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h133cdd06ac921925887570a0c8c92eb19ceb16f655033ff4a05140da54dc8d809fbca504387c82f1076f936829f7f07480c2807b4ec592f0b3d96980d30bc407384cb4c9005f1b05155f96e06cc52;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ca0ea3e4e38cc82d06991f11ba774f2ac358f49d6ee40334a1503a09b8ab64800427e4fd25131bf176f646143374630bba93f26a3b620e264a61080248018352451497256634e73a74d9ddd23dd;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he552bde3a4a932b5b049385106a05492f288b1fe053f5159eb44f46333f9b75f4baf3c331fe95c1710d5c7667ac74e0069578e6dc42c139d155297830cd096717432eac4714f02168151c03520b3;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf8d0684d674d12b8bba5a2aca88d9877c8e96451abefe12c92651f3e3a09f5bfed6450791717f73774f1919191eef3b7894a1b6ce9fac135a65d613f45fbe2bb5ba685ede658ad3af0e7d15a3770;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hea9932ec4ed60b64c36c5f7d3f3f502b809e01191d4fd68b10560983a00f579918f0e517d161256da989cfec01841db3bc617ae04c7d98089c8f84a172ab4c54f05e31b12a804a10a7921f85438d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h12bff86b43654306a493955d5dc5624345ab0eee14a92d79a8626fd0ba6176ad0671da2f7a1db8f9edbad4da1de4aa38665a31dfb387b99e38a1c803f1193400998b911f1f66e7eec4c74923a0a91;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h719cbc22d1956d286cc57aae7ba829dfecc1b15f3820198bf0a2c29fc9ac4bb5c08208a05aee47744c604f4414e2b978920a33bbba741a04079d671fc80ea0c86a581f41dcf7d6875664e5e1bc0d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hfe8787f45fe6825a63e9974d7de768bb90c094ddc0d366f24bf8250e44e0d314675f363ef9b5b0039eeb447a844cfd01e29722ef2d68fe9abd6afdaab3d40008fdcff96e6f89f94cbe34bd896dd8;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h146278c4d4522280994c9ca3dd49bc5b330994a8ec0c3befa57ada56499ed26217e5cb8838cd86eecad1211e9457346963b80fb2309357e81dccc9a6d1aa408e6d3ddaafec1e935f4e6f623f40807;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h70912815bea323523a346a8cb009b59cead2fe221dcc9081c088dc95b02b04057d90dc77e7441910eb664c7f5eaa500e9128ed0d00154ee9263dd8c8316c6920d8ab22c85cd42e441f97b659416d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h80de412e28fe5a460f0446cb6caf43ba3c90c165fb922f5f5c8b9c1e555d451e35cf82abefe064a59273b8d492d10bdf2dc9040d09b167ee3a20d55a5014c491079d1b8373aaf82e2724d8d0771f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h144c381a2d628b0db6c7bbf7c536ddf4bc77a8a8c2c1a7f1b8d1f16b0b047846f7d8bbf4f0fe41e03f5951be5ca21ad5e0918a18ea970fb02472709777a60a63bdeb727a459f8266c8b0b65fb48d4;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1bb418f7144114a2b7ab0fedc2b860455364637e9c60a97f7b434c04caae78e9ce97aa06d7b5cb4fb55c818b2e6d6fe0a0409ff9476dcfe19f58fe1b459d6987eef0e9c90ae85d274e338dca01201;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h216d0c7fbed554943a4bf543bb18bf7fb3a6e49cbb30712b6425c388a251d21679e95ca5c17de2d631bab94939c866eb06fead7ddf68c23ae41e68c0abc3523fe0c7d7b6906d80ef996e531de776;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h6653df02676c38f796e4b79207f1230737030258c5884102e8cdd65e2d0c6558ee68e165b35a3cffa5d6e01fefcbda631824da98db4b3e14a0f2fe5a59dc73c14b1dedff1442197d19db7820ba5e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h140e1556195970b1049ecd41fb59f06abcb42c26cf009a9e88bebcdeb8e69356cf687e26a38c497349830c3303ff094cf320d7fe21570ac445b8ea11c540f50d35c393e0c7fe4bfd926af0d13ee5e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd5b1e34f00dc2a0a72e64d59121c548a35d754a9c9837908a95c3e174f5bcc9f8286d77fbb88b2938bcb8333ebd437018444b76438f204ce3cad3b968126c62a360cd75accb5005c2e1a8f9f05ca;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a5866d66bd16dcfeeb9a2b981c3276dca9ea36a9dac130b35a04297b427fe1df18d35bd510c32cf26753fe74bdc36da86df45ecc3ce751d92c89aa3bbb2155c3a9ead071a636cef23a227e33052e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e78caa66b6758d2bc2e2b646b9bc7ebef4b855c488cd1bfd7eede1aa2460313551c0685ff87a6d92740ed1c757741d8221d6641c45fc4a8063e8a7531b1423189c6a224592c8111d9dee90b3e57d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h8bddd47df88e327814c698aa169d09ed295226426edc3a25dfb9d1e8c49bfef87c02210695902be91384bc94d0310094e509fb2c521b248f29dd1dd864b7a612a27edc64a18dc0e3aedf239189bc;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h5e23df1179e6c9081a491eca0c0d219abee72f50bf7f643325f3168d2f9acbf3166e71764450cc7978d5776c11617990c951caac0748da55175f2db3ea237c7c700f693fd7a350c1703e828e2b86;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b3490b55f0ccf06b0d8a406ce1a10e9f23253e8f8389c4e63b28bcdbfdf6ed580b73f055895682f4c2e3a67d38bc7047d421df277d5624d6f0aaedf1605035e2db1f0a9637f170c0d59d6ea05d98;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h534195b5f4794cbddfd00c304d3c9b0d1d690ce4eb0bc1e7db3ec236b87f4fc39513460ef706135944209b259ed43afbe0e186fc136b1c215ad9764a651d6e1ed9596e67215756acbd24d0103889;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b8a0eeb4953f5c8c8980b5f103cdb85f8a6c23a99ce2a840deff74551c5c7691fd6b8630b519085131eee1e2d97d5ba7f31e1afd9c76b2f727230180bb9532ec1179b3801108ecd259b6afdc5c13;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h5a23fba0f023652b938580ffb018793286a39681125205120dcb0c91114cbbe27a6938239e4eb668476bb3b47c6d52feeebac66c8d1aa3125d9d75b1ceb129a5d52750a704b247d826705c269f52;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h88e421785865499d3b993f392543fc088f644056cbc466352a3cc796b3e052be04aabc980bcf1b51441c6310cc0829b4e2625676fdff8f4ac335d54ad65faf6f6df1a9f3c1240b395e6d5cdb5b2;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h3f4a3da660921312bf9627144a253088b75d3a62b2ad02ec9d8ade3e4f60776686df2ad89c5a4bddebe1e5cbe44329f6be2f14b98e94bc38adb8066ad95f0930f84d6479ae5d1311c081c44c6734;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e87515b75e347cf9888bbd75a22b468adce53359f92af5be378edfc0ec7c59b6ae26c7c6cf7d6053e46456dd058efae654a2978895892a1983a86b25bfdeafec6d01b907b605e226f5780a6c2058;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e4a347ed392414b1af0196d46ec76bbd42f6d05bf2d07ad72daf2cc0cf763907d4b519e5b40c00fafc5c7a7905a0480888cf6a1809bab4171aeb32411ea5056ae5d7a6eadd42c1c6471bf336dd66;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h4e22655a9eff920c9ecab0608ac3b4f34c0dd099185d930369ade8fadb70a9236db42b666ab86bd6cbcc5eabd3783aa1a63f08baf1bae016ea8150d4bec1b00d75b64ccf725c4a0b60d18d317ee3;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ce755f0d4797003765df9c66987cb4316d2900b365dc6b19d0f65acf6ee877caa4da73e855c5d210a176c56b1dc9e7af4c874b1026e0df1dccb76e7f168d3c5528c45bfb24ea4a4605eeafa41bd0;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha716c39923a677dd3138585e8c30ea47f32b99b87205c34cf4a6756ab26cf82a19ee5ef17d5badfac5790b287adcb0758bc3193d9f4a1700a2459d9e2695ad2929b09165acf1841a498c053ccd24;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h12981d0174062341669af9b58778f890af7feccb8642aeee6c00b27cd467160738f769221b19e13b94952ec6cd52582268042acea8a49d22be7e673c3c610babc54486ab62d4a9e6082320a252f69;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h5574f472947f808a9f8a51b839154bebe5a5669956057f9ee3b5259148682f15d61550fed87c1a14d365981659defabda7f66b821bdd53d9bf7a571ffe53fc0ad8786844e2be32db422a6bef3084;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd7719efe72e27c476f26c6974743d43e5c703ff1f149b683b8d7781f956dc05b2d9bd5abe88eb44daacc607bfa6ccbebcb851c4243b0302a3214e98d890222822369e7cd08ffe28cff6c3a9b890b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16286b5b5b2e61e420d49e62400ad1bb2d3594add7989c7097776dbafd404355e1d44f590be85c56ec10cfef18fdb21454ecc20f338c9f69a8af8aae4aa81a88ce52a03c39147bfb8c3c81ada8e8c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h460fc876741167bc421d9e21a1e02b70933265d6d4fb29ed10a84f6f1c6a4e1308a70db711316d828e4c144b67c977bc1cbf723d1c4dc013b9c561f6c3d4fcdeba314c096240d8d83bbfc58f10a5;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h2ebef22fe91df1687378b39e8a3612377af995142419a3e5fe91c036d8dbea48931917e91b39cb348c2e7201694096c18a5110cbd74541a63d4404cb2138a900b433e5dd08edfbdb285d0a914089;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e41d2598e84c800fade2aa6d3e73d843ab965c7223cac54b585c81c2cf688db9069ddc355e542565d65eff9e1b4aec086ee7a03e99294729a1a830298ed975e5c2be876f2c23ecd038542b0a82f5;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h167e1c19ebe732ae5f0c285499208bea5f2fc083b45eeb305797562f0856eae6c4cbd45877e8567e504255f62b534382be2dddc92067e03524fd650d66b4b4bc113bd7ec1587184af242272f436d9;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hdb8a7a74560af20f1cf0582edb124897a280ba5cfb1f255686b405bf31b01c4c9aaa2f084214045e99158e8e04d59d391c39552c1d518f66134ef4f70b05339e8f818d45e4a9438206bd76a31c42;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h81819be63f55c31621854b212835d4dc75fbef7da6bfae67bd5cbe51a742022508d452c0985c584aabd172b7a55aa616437b309575648927cb08a7154bd5d6acf5ab5e914bc7d9c8bcd017b3b082;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h9172eeb17acd8512c26f335c4b236395cbfd9a9a1666471711af9c291341edf10ee4cf1eb463590a18398e9fa8f16049a4cb1b5e583fc33077afa7b38b375d3d964b24ce59ee2aa2cce7736eb539;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h7fe013914095dfbf604c6e6f4f6edc895e3cbd177158ccfe608c96675b3d9462b4248974c44e7d961dc77dd4e4a7bb2a0b412e40198ca8f72994254d96805c5706691a593681cf61101a0542efe8;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h19a9bc0a922745898992de48b1452b2adec4a4dbdb5f178f0f17db17c32ad077130428c587ade341c43e7a3c937cbbd0ded13ee906d09c71d5f311015ebd7a12d04eaa02ebe334c88197afba3c9b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h152b1c819f970de9811315a031e1dcb0384e016e585ffb04e427ffa7a17f0e2432cb8ed20c46be10396f1e7cf039f202bc72266405f2b9f58006d957daf653d49152a82874458fdbcfc9728c800;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a7f808180cce0d31b97ebe93fe28d697a2b7de3ef011f0588681cf5f8bbb95b738260143904ef33c288e125a769d3a4369459e387f7dce112420dc1444dae8ac003a9beedfba220507dd903728c1;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h109a83503fbede2bad5ab75d2a1e4e5f41b2250191540829e9907b01ce012c09e0c565525dce5361bb3922cc6e5373b660e8fc88dcb491f3947bbebf997b778d1f0d7462824426d08597dd782cf47;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h734ab4769a7faf1c8d6afaf105a4c8f71b53a26921a8a97910b0a906ec2c3a9be6cead17bfa541f80b5dae86417b2e6a79d56da5966f43c024067647a9bd2beb30b8c04cdf7d2b47df9129e4ac7d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f442c70c21f01aadde1b459ff3b52d6caba05b78f0f58bcb335bb5d95e8bd088dd5383557049f36bd28f4ce606bb00d9d1bc763bdf15cb57762dafefe85e4c0353d347126a247e01f141ea5b12e5;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ca628edc4f83bfd3cbcff9e07a0e5b782a490e4735bf3dab40c692cf119dd19e755064c65c038dc0becb3a8a2b38aaa80120da603981c0c5ca97b3cdc2cd851ae7ee9b708c7eba4cb472435ed76c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h78907179fa112df3b8c19acb026d1f00bdf96444289f2cd6868827b098bdc0f2b046343593c13ad1aad844214d1c6670b2e8391d3c16eb279ef5ef8a6d8405dd6cdc67a87c858cb072146c7e044d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h433f0462a9645500ff5e955ed2c606b13ddb4c61e266f18724198a227b4547761bab202620125685a01303212bd7627101a558ad545c4c070063ea86890a5a2315f2860f6231e45a6820ce6e9128;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha40e2ca979229de17ed5bae05a7438b645b73ee9fdd5400085e793af31c8973a4912c0f7073b3a3bb3f65d6c39b9b4d575f45c894aee085cab4c59e7f7ffaa8601dbee83001b0c33670c366e015e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he3027b116aacc8c87c23d28fc85f37ddb61f27215dee806cf2550077b5968bc94b7628920e7c1077fafc08dba704be6188b9e2fc22b026362441283ec1b49bd1e0066fed1fa1a9fe3862f1e551e6;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hdf6f6b7451102f0d21e20095fccf1f8e503c23a777441e6dd2234615ce372826ab561eb365b30bdb510f3f5641491d0bf34778773986d318ff2411201ea7850fab9df6bbaf08588f9eb0760e3669;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h81d25752c968b0014644a880e84b0d25f04f8c919ded0b678c3f62327f81dc3eb07f30a4c5cc9774168596e0934f62c72f2153571d3f61d77bdf64db577638f9bf30cb68b5b46030b23bd3f8170e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b2ff7f35b37f76fb9bef2afb01129dd8762308976890f5732bc7f7741fd5079078541f8493ab54efd61c6b4ef77546f9144bd09cfc1e724e2651b91da4b7b23c064282117b9ff1e336e3821e9875;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1223e8e82fb5429764fb0961fbcc13f378cd44acc2ead1aa857ea3326d91e0cb08c917fd03509e19337573c6701fdb8b5411c4a569d7530c5fde3b66d30a037809dcab8fcf2ca73efcc4154bf9cfe;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hdb93733b3fcad6ffc2168627a27f4b31f3e9ba0613afc45d719855859fb9b3daa96ee5c43f46ae3aead4464a788bbb31da7692f1b0b32c60c2bb4b08bdb272376e6433087ffec4f5f563ba0f0559;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h172fb6ca3d711a277d198b312c28759183d12c5c796cf025fe9697d63475e978214b32cece8693bb3913d167d850a8cf0dbdcd51afcc56d982903a8b1be87a2cb3f1a9373bd0bd4027500d1fb60f0;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1112ae28916f4abf69be4f8b8355ccb5ab97c7c021560d7a40ab41d01238b11c5075b500cad3e8e4e54c53129b342fc7178d9a4d588537a33582711e53edced5a3ca1084b597025f82729148ae4cf;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc454c4c1e98808062f38a7f0253e3b8bc7982a6cf36f162c4aec051b58db96b25718edad1956b1f361c23ea0f6e515583ec6f549b6eecd3b7143dfd2dee53bf2e807fce7a45da8701a8ebb1f678d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1aaebe6d52ffc5f0466e9394914bc6d21245ba3d74f3c1bd90458f240da61f3ee4b8106ac19c4c63d08f78ae06c7e484ee619c44250747d1ef605b27e98a7b2975ab96d8d2795e8e9eecd0e9976ae;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10fbf4ab458da7a105e9e7f215c05e6334fdad0e358d52e654fd5596ca52f6b3ec8d85ba8c98ec1218a3d5910b64cce72c115f51d0785f6ff4dd3fe5a2f4bbff34cee1eb7dc905681d82ed7f0a4e4;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1220e6760a90c5c7b6feb1d50292c7b735f2d8a1e4aa286ebcb5e05b042099491c10e268649b60b8b2429d8a550bd25c4d57c18632974b2dff89e0a184bd161767ece6997f4a319c2ebff0abeeede;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he0f8716ddcea7d3d6496a40e6bd003df2e6450893415ca90667778df1ad7ccce0fd93fcfab0823b718d4f23fa3c5e13f5be3e724d281388477c8b7fa6132ea328a685da404ffc159fd45f68fddb2;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he08c92b4a8ce2974610d9dcaabaca90a5ad97d3dcfba9adf3b523341d8f8b4ab53906212dbc67f0598439ef669a3d7da5921143319a311ad8ffd79e2792bed4ced3b362826395f891aa7545306ed;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb76ed4d1373d6a6c9b35c32bd09aaac49cb0d1080f59aa84b731959280591fcca5b21afa5b9526556b7f8ad075c0f641888ea846efa5da8ba47bba5fda0844a695ba656177dd843cf8cabacbacf5;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h9b1d9e41248470815964daf3b67b760a8b5b9740d3cee9ed15343a5d307f15bec7dfa8bf4d12ac902f4c0ea6a551cfca474e2f2645d6158d4b4d551155a10f2cdc763c9f66ec0faf26eed0027275;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h794bd11a7f5088c8b54413a03cbf3f86ccc93cbfd7d16a009193598f5672d44b4a6fdeb9bdde2bd3cd7cc0cdb3ce4f5fdec99c13e39f07bdc006cc046e09e163787e9e2666fbb8704cc27e05c3d4;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1cf63b5b1831687acb774f8610a591cf83d2793a2c6dff1d0f9194d988ae580c98ff74ec7ac478f732878da2c35a0c15cb225aaf665fd3ac0a8a48d59039bc334e15abbc979328248dd2d7243c483;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h134762d383274cb2cae130ece3695b676c37445cd0aaffd1f8bd4fe3ef4c632b911eb788952e423633ce9701580924dbe29a6da644a369368950b8d501ea000b0dea490715e2d4dafed59b167b7d6;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h168ba5476eea710d441bee20c75e1cd6b4eecf84d66ac646a17c7c03f1f975f9b773acef329e598755282f91575b2020900898c81e61223fa4dd0d76bdf07cc13df23bbbf8e3a00cd214beb151afd;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h2c735b7b0d394ee8f6efd6f9fc64a076ee8630ac8c3b59ec1956a3d1a2f32c0d9682a7aa33ec07fe29ff1ca0bc689057f5107ef4045eaf9b7caf1b1eb3d629b094ec2990904e6eb80a17c988b63c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha2f2c8aa96167fcb94454a4980898835acb6b9a9683b27269549837be505210b3e55352df11476fe497e639e6f36f5ec7aec10783fc9b0485a85f8fc9d77ebda3bcb07a0b9256cd853d80061fafd;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h180ab823f2d271555cbbf2f20212467b86ede3d62ce40cadd9e9271734764fe18d8bd571e55619d93fa26cf4e47a451c5f1c88e3658546af2090a3e1f6eb07482e760715d8ac64b657555bf37a667;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h11fb0b7864fd1a89db3748a4490f50c612bda38799cdb38b13882462821f4fbbdd97e482d52126ffadf50521d90508a7bc96884a6d257a387b3d885eb4368b2b23cb3115108fd19d63d01ce7e4c26;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h12e010b140dc76370deed659b959a79d7a203dc53a1931f2a35f4bc51b94d3b93700cc8c9c7fb4929fe01b3718011aa0ba05c2b7fbf7f5afb0e2a660c9da55cdb5abbac0b358fc3c248ebe6912a7f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h7efe16ec63f280b7a8a872f4ee1caea0adc7f4105bfb3e84d94e0888915a7a77a2301c96a16de28dae26a373af6d780d959a6389f8c4ae29fbfcd9011150b20e8dfb04c12b3f9695a742eba72d38;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hed784e79ea1763248627c96907490d76ef076990a5d95f314cc9d73dfafd5f9e3d5f9edd3bc95f1953e5ec323be98eaae0b3fb6ded59738c1640f8ba0808eebadf459d9a14f2dd987745b9b41a04;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16ab44ab16915c43c9abccfd8b996adbb4b8913a69ddf16df00ebb8a0ad2bf5c8390858b210d4f3ac773da4b5c9425ab3faed77a31d0d40785e6ee6918dfff94e3bdb1e92cc32672ee814509e97;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1741c5b3cae72706ff7c4d2c8c332b296da4fb9b75d8ad0e3ccd13ec78ebce8b3e20b88fa257f15050b27fcdc7f9d6ac7dc3a9387388fb0e17b9c2ebf01cf41785bba3504ec6b389cb49c9f4950cc;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h15431d7377041a99b1bbf7e52853eec872e207ee52342c8427671b8a992d12a68227ea35014522dd30f77ccbfaaed26b48b770d8fd23474e71cdedf0151ab32069d9bfc26ceba47a3d7474d667b7b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h9590d9d0b156fc6cf241519d12dbd2f64f4de80ceaeb97059e2842534389844a2ba65338b97a08eebe5281c7c7057b71787e71d52a86c00417fb6303840b9620686f9cfc44fda9dd109e61b13905;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ef7a9b5b1c654fdb523044016446aa4f0dc0e52a77fadf04543926f380e03f31b0377fedb7a39fa9f93aa4113e5b7a23f73542b9a93dded4558492a49bc0305de5ef9db2074de633b213cef17e6a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h64f6e918cf7937428e8caa391d4e071c171795d5f643d24f2f44a895d28d6f3fcd27a546e094f1adc7995c1c197e4e20969b741fae51748cd2d2760d186470c781b6536b96eeaacdb25c6b93c5ab;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h2ce686fa050218ce77c4fbb01c72dcd0ca5181370bab26b0104ecf4f9d822f60c34bfae2b5accb823ea86276f8cb5e1353a5a276b76141ba511e8246b10f6b855a545c2f13cd96d214565772f4f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h4f5a11a41eacd92df7142e872c77af639fa6af821534ea8267e479fe340ef9cdd10aa28ceb62cb643b1ec7a1ec025ab509b45dff641426cc96f1ee231bf88d0ecfe9e504b1810dc6f1e6dd2d8f11;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h14dc85984a30a72c778f1dbcf65a4b7e0d262b0511fd80c55334c2755903c6b30f2f130329dcf82f1849d72a1e1eee1f53e5820bf9234a59ef59210e35049227ed627b9c86c748c681f7e63f9ab7a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h467c42e757a00b49fb81d8db50dbbf36247a6b3e4a568f6778d018231e9e1acb74ebe2648be94955ab151a2e95b4c495fd6fd2bc1599cab1fafc380e9a71cb602beee194fbc0e3f1f93fa725974d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h8d4230f1c45f787747809c63d3d37a3ee84cc0dc139e1648609b55781c07b0ce94a15e3c95a205809da435bfe2abd4ac70ef3600ae27d8e5ab5a21f717e139d4a49c22980c72bdd2581a44d55b3a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd85063bb7eca4ff6d09b9023f80e61502801c590107a8c06cd41d548cadd809c680c3ad6b63b89344b408a5eed51d7e31179efb0ff2c27f75541f3596212cc6cf3e68e170bd54a9f9eeaf9648913;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h750e2dae8712b6d6c272e5ecd4b7b0f13a33bc83ea5cfcc1340e6d4b2c13815ecee05eff438c1fd5175dbf2253a8304ba3db1ccaae51035eb23685c6d4eee1f20aeaaacde8a496a2f9784eb3b8a6;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1df7ee18277820131544d100f28ac8d19b163dc5fa2b114d22a59f2f1c8f36737730157cf62e58a89fa5651291f23e3093ad7e4c50a9d5b07f65407e655d2b1b14780291fef803f0b02d85a2810e9;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h11a96019667191e40488fd0ce3a2ee4f84c6ce2a5cbf90894f7ad193189ad6f64be864fbb52a806710d54351a2c378c6b8cf69153de1856360ceeaeef57081b56ec2741bdfd247c909b393dc82e4e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h147ac6943fe54c2da231bbad7594ce55b797b9aa0752dfc9b5cc70642b559e6b2883f967b388b35dbac2e281e3a9107ee67ff02841c1f3175a6135e22da51f751bd8eb8b1fd80b07a9412768814f8;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc5a3cc89fe12955914bcfc85d863e29f47ff404b542227b8e9b856596dd9ba47cd0516a64c5c3991402254baabd4fd6027901ae89f67e78587ab61f27c6852afcb4d6982e1c0ae338f293a715fc1;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h150b16bd86d5446c22b83a3955b98f8dbe604797bc2e4cbf41cb721cef60e6dd4f9d0bffd4fa649aa7218e592b9533b33e73abec16592bf07d31bfbae2ea933c0b7d503da405e858085f151649a6f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf44b65a510b72fc4549a2aec82a616fce871a302d17df21255cb478c786a4404cfb88eeb7dfb8a40adc734c4ccb926d3854a7e01abb6e6ecbd4d223b3fc7ce126191fbc6819917375372770d4fe3;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc71f01e73907b30c1d18b99a71a6a6d0b73e55cd5fc37d612ef6fe93195ebe0d45d52518bad853978cdf27c5121abc48180554f06ec2660443a0b9a10de8219a26e15fee6301f8c86ad721cdd22e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f3b83096330a8283ef06192d4f2616309389b3ec807c244e51ecc0041524130ec991f400b42834e570367ed9145c5aa3708b4cebdb8cfbebfb6c66afec0263855ad419ed7ed67ebcbb87450ec738;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h896b890533fc18668e411118fad2e8f4b488b6c35904bc711f9ffd7adddecfa90e394f93a9c7ea9afc7f15ba5ff9e4ea5beb0fd18acf48c6d4866b611462f3736f4ebf290ab69de8be4e6009b86;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d9fa35f12abd727ca4962e324788b432f4c90597dc8c1469433d4c25b8ec4f4fa49778d3dc63ce40f72330c41ec13a847af442d31ebcb80b713231fd53242a1c87b846144fd90b5e2951cd986a45;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h416a62827318a3482081182d712b224748bc7ec5418761a052e950fed190cc76454729953d57f09187d22103cabbdbde2fa3e55ad33729f2cf2340ae86721742686f86ab03384a8fe2a6ff9ebf26;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h2bb3c4c9be7e71ddbd7626fb0243a4e9025cc7e4bad69a78007c179272271bca197b59cadbd47cb79f4b5a045f40b80506ae40c4e3a881f89985af6e864157a3a968d484dd7ce1cfeab23d424289;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h22fde90df2a11ca28fb41e05975626f9d54044948f44b483b5a88093a2fd8b0565b9c05e75ed12eeb60ef4edb53627f6b8d421dbaa8a77b6bb710d0dcda1eb3af0d2331e8b0104b8caba534c1a18;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h6c97c033f0e3f7df933e1e5c66ede77ad0dc8de941afa1fdd1ce23799070b0fae99fdbc7eed55a631cb5d49d2c050d7d4969b4745abb108f318a96071c7678f0badd85d282f72a46f49287ce9949;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd5c3481d0df5c272d2a4d79cdde59d11755f4f5ad27f913fb87eac5d4078970b9bbc2e3aaca203593c97a7647003484933c19e1c2ef60d646f3a08e4ecb7da216e91a9cd223a4fedd92f77a869ca;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h14e44e2c1f58aedf3a1e6e44c4d68280682035e1129bf7c5e04559867806b46203e600f7315dc88b1ec980d46872574172f5d0300ca156f7f28a2bbd84e6df5126800cf244ea355de6b78c3be66cf;
        #1
        $finish();
    end
endmodule
