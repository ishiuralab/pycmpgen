module shift_register(
        input wire clk,
        input wire src0_,
        input wire src1_,
        input wire src2_,
        input wire src3_,
        input wire src4_,
        input wire src5_,
        input wire src6_,
        input wire src7_,
        input wire src8_,
        input wire src9_,
        input wire src10_,
        input wire src11_,
        input wire src12_,
        input wire src13_,
        input wire src14_,
        input wire src15_,
        input wire src16_,
        input wire src17_,
        input wire src18_,
        input wire src19_,
        input wire src20_,
        input wire src21_,
        input wire src22_,
        input wire src23_,
        input wire src24_,
        input wire src25_,
        input wire src26_,
        input wire src27_,
        input wire src28_,
        input wire src29_,
        input wire src30_,
        input wire src31_,
        output wire [0:0] dst0,
        output wire [0:0] dst1,
        output wire [0:0] dst2,
        output wire [0:0] dst3,
        output wire [0:0] dst4,
        output wire [0:0] dst5,
        output wire [0:0] dst6,
        output wire [0:0] dst7,
        output wire [0:0] dst8,
        output wire [0:0] dst9,
        output wire [0:0] dst10,
        output wire [0:0] dst11,
        output wire [0:0] dst12,
        output wire [0:0] dst13,
        output wire [0:0] dst14,
        output wire [0:0] dst15,
        output wire [0:0] dst16,
        output wire [0:0] dst17,
        output wire [0:0] dst18,
        output wire [0:0] dst19,
        output wire [0:0] dst20,
        output wire [0:0] dst21,
        output wire [0:0] dst22,
        output wire [0:0] dst23,
        output wire [0:0] dst24,
        output wire [0:0] dst25,
        output wire [0:0] dst26,
        output wire [0:0] dst27,
        output wire [0:0] dst28,
        output wire [0:0] dst29,
        output wire [0:0] dst30,
        output wire [0:0] dst31,
        output wire [0:0] dst32,
        output wire [0:0] dst33,
        output wire [0:0] dst34,
        output wire [0:0] dst35,
        output wire [0:0] dst36,
        output wire [0:0] dst37,
        output wire [0:0] dst38,
        output wire [0:0] dst39,
        output wire [0:0] dst40);
    reg [511:0] src0;
    reg [511:0] src1;
    reg [511:0] src2;
    reg [511:0] src3;
    reg [511:0] src4;
    reg [511:0] src5;
    reg [511:0] src6;
    reg [511:0] src7;
    reg [511:0] src8;
    reg [511:0] src9;
    reg [511:0] src10;
    reg [511:0] src11;
    reg [511:0] src12;
    reg [511:0] src13;
    reg [511:0] src14;
    reg [511:0] src15;
    reg [511:0] src16;
    reg [511:0] src17;
    reg [511:0] src18;
    reg [511:0] src19;
    reg [511:0] src20;
    reg [511:0] src21;
    reg [511:0] src22;
    reg [511:0] src23;
    reg [511:0] src24;
    reg [511:0] src25;
    reg [511:0] src26;
    reg [511:0] src27;
    reg [511:0] src28;
    reg [511:0] src29;
    reg [511:0] src30;
    reg [511:0] src31;
    compressor2_1_512_32 compressor2_1_512_32(
            .src0(src0),
            .src1(src1),
            .src2(src2),
            .src3(src3),
            .src4(src4),
            .src5(src5),
            .src6(src6),
            .src7(src7),
            .src8(src8),
            .src9(src9),
            .src10(src10),
            .src11(src11),
            .src12(src12),
            .src13(src13),
            .src14(src14),
            .src15(src15),
            .src16(src16),
            .src17(src17),
            .src18(src18),
            .src19(src19),
            .src20(src20),
            .src21(src21),
            .src22(src22),
            .src23(src23),
            .src24(src24),
            .src25(src25),
            .src26(src26),
            .src27(src27),
            .src28(src28),
            .src29(src29),
            .src30(src30),
            .src31(src31),
            .dst0(dst0),
            .dst1(dst1),
            .dst2(dst2),
            .dst3(dst3),
            .dst4(dst4),
            .dst5(dst5),
            .dst6(dst6),
            .dst7(dst7),
            .dst8(dst8),
            .dst9(dst9),
            .dst10(dst10),
            .dst11(dst11),
            .dst12(dst12),
            .dst13(dst13),
            .dst14(dst14),
            .dst15(dst15),
            .dst16(dst16),
            .dst17(dst17),
            .dst18(dst18),
            .dst19(dst19),
            .dst20(dst20),
            .dst21(dst21),
            .dst22(dst22),
            .dst23(dst23),
            .dst24(dst24),
            .dst25(dst25),
            .dst26(dst26),
            .dst27(dst27),
            .dst28(dst28),
            .dst29(dst29),
            .dst30(dst30),
            .dst31(dst31),
            .dst32(dst32),
            .dst33(dst33),
            .dst34(dst34),
            .dst35(dst35),
            .dst36(dst36),
            .dst37(dst37),
            .dst38(dst38),
            .dst39(dst39),
            .dst40(dst40));
    initial begin
        src0 <= 512'h0;
        src1 <= 512'h0;
        src2 <= 512'h0;
        src3 <= 512'h0;
        src4 <= 512'h0;
        src5 <= 512'h0;
        src6 <= 512'h0;
        src7 <= 512'h0;
        src8 <= 512'h0;
        src9 <= 512'h0;
        src10 <= 512'h0;
        src11 <= 512'h0;
        src12 <= 512'h0;
        src13 <= 512'h0;
        src14 <= 512'h0;
        src15 <= 512'h0;
        src16 <= 512'h0;
        src17 <= 512'h0;
        src18 <= 512'h0;
        src19 <= 512'h0;
        src20 <= 512'h0;
        src21 <= 512'h0;
        src22 <= 512'h0;
        src23 <= 512'h0;
        src24 <= 512'h0;
        src25 <= 512'h0;
        src26 <= 512'h0;
        src27 <= 512'h0;
        src28 <= 512'h0;
        src29 <= 512'h0;
        src30 <= 512'h0;
        src31 <= 512'h0;
    end
    always @(posedge clk) begin
        src0 <= {src0, src0_};
        src1 <= {src1, src1_};
        src2 <= {src2, src2_};
        src3 <= {src3, src3_};
        src4 <= {src4, src4_};
        src5 <= {src5, src5_};
        src6 <= {src6, src6_};
        src7 <= {src7, src7_};
        src8 <= {src8, src8_};
        src9 <= {src9, src9_};
        src10 <= {src10, src10_};
        src11 <= {src11, src11_};
        src12 <= {src12, src12_};
        src13 <= {src13, src13_};
        src14 <= {src14, src14_};
        src15 <= {src15, src15_};
        src16 <= {src16, src16_};
        src17 <= {src17, src17_};
        src18 <= {src18, src18_};
        src19 <= {src19, src19_};
        src20 <= {src20, src20_};
        src21 <= {src21, src21_};
        src22 <= {src22, src22_};
        src23 <= {src23, src23_};
        src24 <= {src24, src24_};
        src25 <= {src25, src25_};
        src26 <= {src26, src26_};
        src27 <= {src27, src27_};
        src28 <= {src28, src28_};
        src29 <= {src29, src29_};
        src30 <= {src30, src30_};
        src31 <= {src31, src31_};
    end
endmodule
module compressor2_1_512_32(
    input [511:0]src0,
    input [511:0]src1,
    input [511:0]src2,
    input [511:0]src3,
    input [511:0]src4,
    input [511:0]src5,
    input [511:0]src6,
    input [511:0]src7,
    input [511:0]src8,
    input [511:0]src9,
    input [511:0]src10,
    input [511:0]src11,
    input [511:0]src12,
    input [511:0]src13,
    input [511:0]src14,
    input [511:0]src15,
    input [511:0]src16,
    input [511:0]src17,
    input [511:0]src18,
    input [511:0]src19,
    input [511:0]src20,
    input [511:0]src21,
    input [511:0]src22,
    input [511:0]src23,
    input [511:0]src24,
    input [511:0]src25,
    input [511:0]src26,
    input [511:0]src27,
    input [511:0]src28,
    input [511:0]src29,
    input [511:0]src30,
    input [511:0]src31,
    output dst0,
    output dst1,
    output dst2,
    output dst3,
    output dst4,
    output dst5,
    output dst6,
    output dst7,
    output dst8,
    output dst9,
    output dst10,
    output dst11,
    output dst12,
    output dst13,
    output dst14,
    output dst15,
    output dst16,
    output dst17,
    output dst18,
    output dst19,
    output dst20,
    output dst21,
    output dst22,
    output dst23,
    output dst24,
    output dst25,
    output dst26,
    output dst27,
    output dst28,
    output dst29,
    output dst30,
    output dst31,
    output dst32,
    output dst33,
    output dst34,
    output dst35,
    output dst36,
    output dst37,
    output dst38,
    output dst39,
    output dst40);

    wire [1:0] comp_out0;
    wire [1:0] comp_out1;
    wire [1:0] comp_out2;
    wire [1:0] comp_out3;
    wire [1:0] comp_out4;
    wire [1:0] comp_out5;
    wire [1:0] comp_out6;
    wire [1:0] comp_out7;
    wire [1:0] comp_out8;
    wire [1:0] comp_out9;
    wire [1:0] comp_out10;
    wire [1:0] comp_out11;
    wire [1:0] comp_out12;
    wire [1:0] comp_out13;
    wire [1:0] comp_out14;
    wire [1:0] comp_out15;
    wire [1:0] comp_out16;
    wire [1:0] comp_out17;
    wire [1:0] comp_out18;
    wire [1:0] comp_out19;
    wire [1:0] comp_out20;
    wire [1:0] comp_out21;
    wire [1:0] comp_out22;
    wire [1:0] comp_out23;
    wire [1:0] comp_out24;
    wire [1:0] comp_out25;
    wire [1:0] comp_out26;
    wire [1:0] comp_out27;
    wire [1:0] comp_out28;
    wire [1:0] comp_out29;
    wire [1:0] comp_out30;
    wire [1:0] comp_out31;
    wire [1:0] comp_out32;
    wire [1:0] comp_out33;
    wire [1:0] comp_out34;
    wire [1:0] comp_out35;
    wire [1:0] comp_out36;
    wire [1:0] comp_out37;
    wire [1:0] comp_out38;
    wire [1:0] comp_out39;
    wire [0:0] comp_out40;
    compressor compressor_inst(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .src31(src31),
        .dst0(comp_out0),
        .dst1(comp_out1),
        .dst2(comp_out2),
        .dst3(comp_out3),
        .dst4(comp_out4),
        .dst5(comp_out5),
        .dst6(comp_out6),
        .dst7(comp_out7),
        .dst8(comp_out8),
        .dst9(comp_out9),
        .dst10(comp_out10),
        .dst11(comp_out11),
        .dst12(comp_out12),
        .dst13(comp_out13),
        .dst14(comp_out14),
        .dst15(comp_out15),
        .dst16(comp_out16),
        .dst17(comp_out17),
        .dst18(comp_out18),
        .dst19(comp_out19),
        .dst20(comp_out20),
        .dst21(comp_out21),
        .dst22(comp_out22),
        .dst23(comp_out23),
        .dst24(comp_out24),
        .dst25(comp_out25),
        .dst26(comp_out26),
        .dst27(comp_out27),
        .dst28(comp_out28),
        .dst29(comp_out29),
        .dst30(comp_out30),
        .dst31(comp_out31),
        .dst32(comp_out32),
        .dst33(comp_out33),
        .dst34(comp_out34),
        .dst35(comp_out35),
        .dst36(comp_out36),
        .dst37(comp_out37),
        .dst38(comp_out38),
        .dst39(comp_out39),
        .dst40(comp_out40)
    );
    rowadder2_1_41 rowadder2_1inst(
        .src0({comp_out40[0], comp_out39[0], comp_out38[0], comp_out37[0], comp_out36[0], comp_out35[0], comp_out34[0], comp_out33[0], comp_out32[0], comp_out31[0], comp_out30[0], comp_out29[0], comp_out28[0], comp_out27[0], comp_out26[0], comp_out25[0], comp_out24[0], comp_out23[0], comp_out22[0], comp_out21[0], comp_out20[0], comp_out19[0], comp_out18[0], comp_out17[0], comp_out16[0], comp_out15[0], comp_out14[0], comp_out13[0], comp_out12[0], comp_out11[0], comp_out10[0], comp_out9[0], comp_out8[0], comp_out7[0], comp_out6[0], comp_out5[0], comp_out4[0], comp_out3[0], comp_out2[0], comp_out1[0], comp_out0[0]}),
        .src1({1'h0, comp_out39[1], comp_out38[1], comp_out37[1], comp_out36[1], comp_out35[1], comp_out34[1], comp_out33[1], comp_out32[1], comp_out31[1], comp_out30[1], comp_out29[1], comp_out28[1], comp_out27[1], comp_out26[1], comp_out25[1], comp_out24[1], comp_out23[1], comp_out22[1], comp_out21[1], comp_out20[1], comp_out19[1], comp_out18[1], comp_out17[1], comp_out16[1], comp_out15[1], comp_out14[1], comp_out13[1], comp_out12[1], comp_out11[1], comp_out10[1], comp_out9[1], comp_out8[1], comp_out7[1], comp_out6[1], comp_out5[1], comp_out4[1], comp_out3[1], comp_out2[1], comp_out1[1], comp_out0[1]}),
        .dst0({dst40, dst39, dst38, dst37, dst36, dst35, dst34, dst33, dst32, dst31, dst30, dst29, dst28, dst27, dst26, dst25, dst24, dst23, dst22, dst21, dst20, dst19, dst18, dst17, dst16, dst15, dst14, dst13, dst12, dst11, dst10, dst9, dst8, dst7, dst6, dst5, dst4, dst3, dst2, dst1, dst0})
    );
endmodule
module compressor (
      input wire [511:0] src0,
      input wire [511:0] src1,
      input wire [511:0] src2,
      input wire [511:0] src3,
      input wire [511:0] src4,
      input wire [511:0] src5,
      input wire [511:0] src6,
      input wire [511:0] src7,
      input wire [511:0] src8,
      input wire [511:0] src9,
      input wire [511:0] src10,
      input wire [511:0] src11,
      input wire [511:0] src12,
      input wire [511:0] src13,
      input wire [511:0] src14,
      input wire [511:0] src15,
      input wire [511:0] src16,
      input wire [511:0] src17,
      input wire [511:0] src18,
      input wire [511:0] src19,
      input wire [511:0] src20,
      input wire [511:0] src21,
      input wire [511:0] src22,
      input wire [511:0] src23,
      input wire [511:0] src24,
      input wire [511:0] src25,
      input wire [511:0] src26,
      input wire [511:0] src27,
      input wire [511:0] src28,
      input wire [511:0] src29,
      input wire [511:0] src30,
      input wire [511:0] src31,
      output wire [1:0] dst0,
      output wire [1:0] dst1,
      output wire [1:0] dst2,
      output wire [1:0] dst3,
      output wire [1:0] dst4,
      output wire [1:0] dst5,
      output wire [1:0] dst6,
      output wire [1:0] dst7,
      output wire [1:0] dst8,
      output wire [1:0] dst9,
      output wire [1:0] dst10,
      output wire [1:0] dst11,
      output wire [1:0] dst12,
      output wire [1:0] dst13,
      output wire [1:0] dst14,
      output wire [1:0] dst15,
      output wire [1:0] dst16,
      output wire [1:0] dst17,
      output wire [1:0] dst18,
      output wire [1:0] dst19,
      output wire [1:0] dst20,
      output wire [1:0] dst21,
      output wire [1:0] dst22,
      output wire [1:0] dst23,
      output wire [1:0] dst24,
      output wire [1:0] dst25,
      output wire [1:0] dst26,
      output wire [1:0] dst27,
      output wire [1:0] dst28,
      output wire [1:0] dst29,
      output wire [1:0] dst30,
      output wire [1:0] dst31,
      output wire [1:0] dst32,
      output wire [1:0] dst33,
      output wire [1:0] dst34,
      output wire [1:0] dst35,
      output wire [1:0] dst36,
      output wire [1:0] dst37,
      output wire [1:0] dst38,
      output wire [1:0] dst39,
      output wire [0:0] dst40);

   wire [511:0] stage0_0;
   wire [511:0] stage0_1;
   wire [511:0] stage0_2;
   wire [511:0] stage0_3;
   wire [511:0] stage0_4;
   wire [511:0] stage0_5;
   wire [511:0] stage0_6;
   wire [511:0] stage0_7;
   wire [511:0] stage0_8;
   wire [511:0] stage0_9;
   wire [511:0] stage0_10;
   wire [511:0] stage0_11;
   wire [511:0] stage0_12;
   wire [511:0] stage0_13;
   wire [511:0] stage0_14;
   wire [511:0] stage0_15;
   wire [511:0] stage0_16;
   wire [511:0] stage0_17;
   wire [511:0] stage0_18;
   wire [511:0] stage0_19;
   wire [511:0] stage0_20;
   wire [511:0] stage0_21;
   wire [511:0] stage0_22;
   wire [511:0] stage0_23;
   wire [511:0] stage0_24;
   wire [511:0] stage0_25;
   wire [511:0] stage0_26;
   wire [511:0] stage0_27;
   wire [511:0] stage0_28;
   wire [511:0] stage0_29;
   wire [511:0] stage0_30;
   wire [511:0] stage0_31;
   wire [110:0] stage1_0;
   wire [198:0] stage1_1;
   wire [187:0] stage1_2;
   wire [276:0] stage1_3;
   wire [244:0] stage1_4;
   wire [205:0] stage1_5;
   wire [242:0] stage1_6;
   wire [185:0] stage1_7;
   wire [348:0] stage1_8;
   wire [211:0] stage1_9;
   wire [181:0] stage1_10;
   wire [205:0] stage1_11;
   wire [221:0] stage1_12;
   wire [231:0] stage1_13;
   wire [231:0] stage1_14;
   wire [236:0] stage1_15;
   wire [213:0] stage1_16;
   wire [223:0] stage1_17;
   wire [202:0] stage1_18;
   wire [262:0] stage1_19;
   wire [213:0] stage1_20;
   wire [269:0] stage1_21;
   wire [273:0] stage1_22;
   wire [165:0] stage1_23;
   wire [220:0] stage1_24;
   wire [273:0] stage1_25;
   wire [190:0] stage1_26;
   wire [199:0] stage1_27;
   wire [247:0] stage1_28;
   wire [242:0] stage1_29;
   wire [206:0] stage1_30;
   wire [242:0] stage1_31;
   wire [149:0] stage1_32;
   wire [70:0] stage1_33;
   wire [62:0] stage2_0;
   wire [55:0] stage2_1;
   wire [94:0] stage2_2;
   wire [76:0] stage2_3;
   wire [118:0] stage2_4;
   wire [93:0] stage2_5;
   wire [95:0] stage2_6;
   wire [108:0] stage2_7;
   wire [97:0] stage2_8;
   wire [107:0] stage2_9;
   wire [94:0] stage2_10;
   wire [115:0] stage2_11;
   wire [101:0] stage2_12;
   wire [123:0] stage2_13;
   wire [69:0] stage2_14;
   wire [97:0] stage2_15;
   wire [124:0] stage2_16;
   wire [127:0] stage2_17;
   wire [72:0] stage2_18;
   wire [97:0] stage2_19;
   wire [109:0] stage2_20;
   wire [124:0] stage2_21;
   wire [94:0] stage2_22;
   wire [122:0] stage2_23;
   wire [89:0] stage2_24;
   wire [102:0] stage2_25;
   wire [99:0] stage2_26;
   wire [84:0] stage2_27;
   wire [170:0] stage2_28;
   wire [142:0] stage2_29;
   wire [91:0] stage2_30;
   wire [101:0] stage2_31;
   wire [73:0] stage2_32;
   wire [59:0] stage2_33;
   wire [34:0] stage2_34;
   wire [11:0] stage2_35;
   wire [10:0] stage3_0;
   wire [25:0] stage3_1;
   wire [35:0] stage3_2;
   wire [27:0] stage3_3;
   wire [46:0] stage3_4;
   wire [58:0] stage3_5;
   wire [37:0] stage3_6;
   wire [46:0] stage3_7;
   wire [92:0] stage3_8;
   wire [49:0] stage3_9;
   wire [37:0] stage3_10;
   wire [54:0] stage3_11;
   wire [46:0] stage3_12;
   wire [36:0] stage3_13;
   wire [55:0] stage3_14;
   wire [70:0] stage3_15;
   wire [66:0] stage3_16;
   wire [76:0] stage3_17;
   wire [34:0] stage3_18;
   wire [69:0] stage3_19;
   wire [29:0] stage3_20;
   wire [62:0] stage3_21;
   wire [50:0] stage3_22;
   wire [45:0] stage3_23;
   wire [60:0] stage3_24;
   wire [48:0] stage3_25;
   wire [50:0] stage3_26;
   wire [54:0] stage3_27;
   wire [73:0] stage3_28;
   wire [57:0] stage3_29;
   wire [70:0] stage3_30;
   wire [57:0] stage3_31;
   wire [57:0] stage3_32;
   wire [26:0] stage3_33;
   wire [26:0] stage3_34;
   wire [12:0] stage3_35;
   wire [5:0] stage3_36;
   wire [1:0] stage3_37;
   wire [10:0] stage4_0;
   wire [15:0] stage4_1;
   wire [12:0] stage4_2;
   wire [22:0] stage4_3;
   wire [23:0] stage4_4;
   wire [45:0] stage4_5;
   wire [22:0] stage4_6;
   wire [14:0] stage4_7;
   wire [28:0] stage4_8;
   wire [41:0] stage4_9;
   wire [17:0] stage4_10;
   wire [42:0] stage4_11;
   wire [23:0] stage4_12;
   wire [18:0] stage4_13;
   wire [34:0] stage4_14;
   wire [38:0] stage4_15;
   wire [19:0] stage4_16;
   wire [42:0] stage4_17;
   wire [28:0] stage4_18;
   wire [31:0] stage4_19;
   wire [18:0] stage4_20;
   wire [18:0] stage4_21;
   wire [30:0] stage4_22;
   wire [37:0] stage4_23;
   wire [29:0] stage4_24;
   wire [18:0] stage4_25;
   wire [22:0] stage4_26;
   wire [26:0] stage4_27;
   wire [24:0] stage4_28;
   wire [25:0] stage4_29;
   wire [26:0] stage4_30;
   wire [30:0] stage4_31;
   wire [42:0] stage4_32;
   wire [18:0] stage4_33;
   wire [12:0] stage4_34;
   wire [14:0] stage4_35;
   wire [10:0] stage4_36;
   wire [2:0] stage4_37;
   wire [10:0] stage5_0;
   wire [10:0] stage5_1;
   wire [9:0] stage5_2;
   wire [5:0] stage5_3;
   wire [9:0] stage5_4;
   wire [10:0] stage5_5;
   wire [12:0] stage5_6;
   wire [19:0] stage5_7;
   wire [9:0] stage5_8;
   wire [10:0] stage5_9;
   wire [12:0] stage5_10;
   wire [15:0] stage5_11;
   wire [10:0] stage5_12;
   wire [14:0] stage5_13;
   wire [9:0] stage5_14;
   wire [12:0] stage5_15;
   wire [14:0] stage5_16;
   wire [14:0] stage5_17;
   wire [16:0] stage5_18;
   wire [23:0] stage5_19;
   wire [13:0] stage5_20;
   wire [8:0] stage5_21;
   wire [16:0] stage5_22;
   wire [9:0] stage5_23;
   wire [13:0] stage5_24;
   wire [11:0] stage5_25;
   wire [13:0] stage5_26;
   wire [13:0] stage5_27;
   wire [6:0] stage5_28;
   wire [12:0] stage5_29;
   wire [16:0] stage5_30;
   wire [12:0] stage5_31;
   wire [25:0] stage5_32;
   wire [10:0] stage5_33;
   wire [9:0] stage5_34;
   wire [7:0] stage5_35;
   wire [3:0] stage5_36;
   wire [6:0] stage5_37;
   wire [1:0] stage5_38;
   wire [6:0] stage6_0;
   wire [4:0] stage6_1;
   wire [5:0] stage6_2;
   wire [5:0] stage6_3;
   wire [5:0] stage6_4;
   wire [4:0] stage6_5;
   wire [3:0] stage6_6;
   wire [5:0] stage6_7;
   wire [5:0] stage6_8;
   wire [5:0] stage6_9;
   wire [3:0] stage6_10;
   wire [7:0] stage6_11;
   wire [6:0] stage6_12;
   wire [8:0] stage6_13;
   wire [5:0] stage6_14;
   wire [3:0] stage6_15;
   wire [5:0] stage6_16;
   wire [9:0] stage6_17;
   wire [5:0] stage6_18;
   wire [14:0] stage6_19;
   wire [5:0] stage6_20;
   wire [12:0] stage6_21;
   wire [7:0] stage6_22;
   wire [3:0] stage6_23;
   wire [5:0] stage6_24;
   wire [5:0] stage6_25;
   wire [4:0] stage6_26;
   wire [7:0] stage6_27;
   wire [4:0] stage6_28;
   wire [3:0] stage6_29;
   wire [5:0] stage6_30;
   wire [7:0] stage6_31;
   wire [5:0] stage6_32;
   wire [5:0] stage6_33;
   wire [9:0] stage6_34;
   wire [5:0] stage6_35;
   wire [2:0] stage6_36;
   wire [1:0] stage6_37;
   wire [1:0] stage6_38;
   wire [1:0] stage6_39;
   wire [0:0] stage6_40;
   wire [6:0] stage7_0;
   wire [0:0] stage7_1;
   wire [6:0] stage7_2;
   wire [0:0] stage7_3;
   wire [6:0] stage7_4;
   wire [1:0] stage7_5;
   wire [3:0] stage7_6;
   wire [1:0] stage7_7;
   wire [6:0] stage7_8;
   wire [0:0] stage7_9;
   wire [4:0] stage7_10;
   wire [2:0] stage7_11;
   wire [3:0] stage7_12;
   wire [1:0] stage7_13;
   wire [6:0] stage7_14;
   wire [5:0] stage7_15;
   wire [1:0] stage7_16;
   wire [3:0] stage7_17;
   wire [1:0] stage7_18;
   wire [4:0] stage7_19;
   wire [5:0] stage7_20;
   wire [2:0] stage7_21;
   wire [5:0] stage7_22;
   wire [6:0] stage7_23;
   wire [0:0] stage7_24;
   wire [1:0] stage7_25;
   wire [2:0] stage7_26;
   wire [2:0] stage7_27;
   wire [6:0] stage7_28;
   wire [4:0] stage7_29;
   wire [0:0] stage7_30;
   wire [8:0] stage7_31;
   wire [0:0] stage7_32;
   wire [1:0] stage7_33;
   wire [6:0] stage7_34;
   wire [1:0] stage7_35;
   wire [1:0] stage7_36;
   wire [3:0] stage7_37;
   wire [2:0] stage7_38;
   wire [1:0] stage7_39;
   wire [0:0] stage7_40;
   wire [1:0] stage8_0;
   wire [1:0] stage8_1;
   wire [1:0] stage8_2;
   wire [1:0] stage8_3;
   wire [1:0] stage8_4;
   wire [1:0] stage8_5;
   wire [1:0] stage8_6;
   wire [1:0] stage8_7;
   wire [1:0] stage8_8;
   wire [1:0] stage8_9;
   wire [1:0] stage8_10;
   wire [1:0] stage8_11;
   wire [1:0] stage8_12;
   wire [1:0] stage8_13;
   wire [1:0] stage8_14;
   wire [1:0] stage8_15;
   wire [1:0] stage8_16;
   wire [1:0] stage8_17;
   wire [1:0] stage8_18;
   wire [1:0] stage8_19;
   wire [1:0] stage8_20;
   wire [1:0] stage8_21;
   wire [1:0] stage8_22;
   wire [1:0] stage8_23;
   wire [1:0] stage8_24;
   wire [1:0] stage8_25;
   wire [1:0] stage8_26;
   wire [1:0] stage8_27;
   wire [1:0] stage8_28;
   wire [1:0] stage8_29;
   wire [1:0] stage8_30;
   wire [1:0] stage8_31;
   wire [1:0] stage8_32;
   wire [1:0] stage8_33;
   wire [1:0] stage8_34;
   wire [1:0] stage8_35;
   wire [1:0] stage8_36;
   wire [1:0] stage8_37;
   wire [1:0] stage8_38;
   wire [1:0] stage8_39;
   wire [0:0] stage8_40;

   assign stage0_0 = src0;
   assign stage0_1 = src1;
   assign stage0_2 = src2;
   assign stage0_3 = src3;
   assign stage0_4 = src4;
   assign stage0_5 = src5;
   assign stage0_6 = src6;
   assign stage0_7 = src7;
   assign stage0_8 = src8;
   assign stage0_9 = src9;
   assign stage0_10 = src10;
   assign stage0_11 = src11;
   assign stage0_12 = src12;
   assign stage0_13 = src13;
   assign stage0_14 = src14;
   assign stage0_15 = src15;
   assign stage0_16 = src16;
   assign stage0_17 = src17;
   assign stage0_18 = src18;
   assign stage0_19 = src19;
   assign stage0_20 = src20;
   assign stage0_21 = src21;
   assign stage0_22 = src22;
   assign stage0_23 = src23;
   assign stage0_24 = src24;
   assign stage0_25 = src25;
   assign stage0_26 = src26;
   assign stage0_27 = src27;
   assign stage0_28 = src28;
   assign stage0_29 = src29;
   assign stage0_30 = src30;
   assign stage0_31 = src31;
   assign dst0 = stage8_0;
   assign dst1 = stage8_1;
   assign dst2 = stage8_2;
   assign dst3 = stage8_3;
   assign dst4 = stage8_4;
   assign dst5 = stage8_5;
   assign dst6 = stage8_6;
   assign dst7 = stage8_7;
   assign dst8 = stage8_8;
   assign dst9 = stage8_9;
   assign dst10 = stage8_10;
   assign dst11 = stage8_11;
   assign dst12 = stage8_12;
   assign dst13 = stage8_13;
   assign dst14 = stage8_14;
   assign dst15 = stage8_15;
   assign dst16 = stage8_16;
   assign dst17 = stage8_17;
   assign dst18 = stage8_18;
   assign dst19 = stage8_19;
   assign dst20 = stage8_20;
   assign dst21 = stage8_21;
   assign dst22 = stage8_22;
   assign dst23 = stage8_23;
   assign dst24 = stage8_24;
   assign dst25 = stage8_25;
   assign dst26 = stage8_26;
   assign dst27 = stage8_27;
   assign dst28 = stage8_28;
   assign dst29 = stage8_29;
   assign dst30 = stage8_30;
   assign dst31 = stage8_31;
   assign dst32 = stage8_32;
   assign dst33 = stage8_33;
   assign dst34 = stage8_34;
   assign dst35 = stage8_35;
   assign dst36 = stage8_36;
   assign dst37 = stage8_37;
   assign dst38 = stage8_38;
   assign dst39 = stage8_39;
   assign dst40 = stage8_40;

   gpc2135_5 gpc0 (
      {stage0_0[0], stage0_0[1], stage0_0[2], stage0_0[3], stage0_0[4]},
      {stage0_1[0], stage0_1[1], stage0_1[2]},
      {stage0_2[0]},
      {stage0_3[0], stage0_3[1]},
      {stage1_4[0],stage1_3[0],stage1_2[0],stage1_1[0],stage1_0[0]}
   );
   gpc2135_5 gpc1 (
      {stage0_0[5], stage0_0[6], stage0_0[7], stage0_0[8], stage0_0[9]},
      {stage0_1[3], stage0_1[4], stage0_1[5]},
      {stage0_2[1]},
      {stage0_3[2], stage0_3[3]},
      {stage1_4[1],stage1_3[1],stage1_2[1],stage1_1[1],stage1_0[1]}
   );
   gpc2135_5 gpc2 (
      {stage0_0[10], stage0_0[11], stage0_0[12], stage0_0[13], stage0_0[14]},
      {stage0_1[6], stage0_1[7], stage0_1[8]},
      {stage0_2[2]},
      {stage0_3[4], stage0_3[5]},
      {stage1_4[2],stage1_3[2],stage1_2[2],stage1_1[2],stage1_0[2]}
   );
   gpc2135_5 gpc3 (
      {stage0_0[15], stage0_0[16], stage0_0[17], stage0_0[18], stage0_0[19]},
      {stage0_1[9], stage0_1[10], stage0_1[11]},
      {stage0_2[3]},
      {stage0_3[6], stage0_3[7]},
      {stage1_4[3],stage1_3[3],stage1_2[3],stage1_1[3],stage1_0[3]}
   );
   gpc2135_5 gpc4 (
      {stage0_0[20], stage0_0[21], stage0_0[22], stage0_0[23], stage0_0[24]},
      {stage0_1[12], stage0_1[13], stage0_1[14]},
      {stage0_2[4]},
      {stage0_3[8], stage0_3[9]},
      {stage1_4[4],stage1_3[4],stage1_2[4],stage1_1[4],stage1_0[4]}
   );
   gpc2135_5 gpc5 (
      {stage0_0[25], stage0_0[26], stage0_0[27], stage0_0[28], stage0_0[29]},
      {stage0_1[15], stage0_1[16], stage0_1[17]},
      {stage0_2[5]},
      {stage0_3[10], stage0_3[11]},
      {stage1_4[5],stage1_3[5],stage1_2[5],stage1_1[5],stage1_0[5]}
   );
   gpc2135_5 gpc6 (
      {stage0_0[30], stage0_0[31], stage0_0[32], stage0_0[33], stage0_0[34]},
      {stage0_1[18], stage0_1[19], stage0_1[20]},
      {stage0_2[6]},
      {stage0_3[12], stage0_3[13]},
      {stage1_4[6],stage1_3[6],stage1_2[6],stage1_1[6],stage1_0[6]}
   );
   gpc2135_5 gpc7 (
      {stage0_0[35], stage0_0[36], stage0_0[37], stage0_0[38], stage0_0[39]},
      {stage0_1[21], stage0_1[22], stage0_1[23]},
      {stage0_2[7]},
      {stage0_3[14], stage0_3[15]},
      {stage1_4[7],stage1_3[7],stage1_2[7],stage1_1[7],stage1_0[7]}
   );
   gpc2135_5 gpc8 (
      {stage0_0[40], stage0_0[41], stage0_0[42], stage0_0[43], stage0_0[44]},
      {stage0_1[24], stage0_1[25], stage0_1[26]},
      {stage0_2[8]},
      {stage0_3[16], stage0_3[17]},
      {stage1_4[8],stage1_3[8],stage1_2[8],stage1_1[8],stage1_0[8]}
   );
   gpc2135_5 gpc9 (
      {stage0_0[45], stage0_0[46], stage0_0[47], stage0_0[48], stage0_0[49]},
      {stage0_1[27], stage0_1[28], stage0_1[29]},
      {stage0_2[9]},
      {stage0_3[18], stage0_3[19]},
      {stage1_4[9],stage1_3[9],stage1_2[9],stage1_1[9],stage1_0[9]}
   );
   gpc2135_5 gpc10 (
      {stage0_0[50], stage0_0[51], stage0_0[52], stage0_0[53], stage0_0[54]},
      {stage0_1[30], stage0_1[31], stage0_1[32]},
      {stage0_2[10]},
      {stage0_3[20], stage0_3[21]},
      {stage1_4[10],stage1_3[10],stage1_2[10],stage1_1[10],stage1_0[10]}
   );
   gpc1163_5 gpc11 (
      {stage0_0[55], stage0_0[56], stage0_0[57]},
      {stage0_1[33], stage0_1[34], stage0_1[35], stage0_1[36], stage0_1[37], stage0_1[38]},
      {stage0_2[11]},
      {stage0_3[22]},
      {stage1_4[11],stage1_3[11],stage1_2[11],stage1_1[11],stage1_0[11]}
   );
   gpc1163_5 gpc12 (
      {stage0_0[58], stage0_0[59], stage0_0[60]},
      {stage0_1[39], stage0_1[40], stage0_1[41], stage0_1[42], stage0_1[43], stage0_1[44]},
      {stage0_2[12]},
      {stage0_3[23]},
      {stage1_4[12],stage1_3[12],stage1_2[12],stage1_1[12],stage1_0[12]}
   );
   gpc1163_5 gpc13 (
      {stage0_0[61], stage0_0[62], stage0_0[63]},
      {stage0_1[45], stage0_1[46], stage0_1[47], stage0_1[48], stage0_1[49], stage0_1[50]},
      {stage0_2[13]},
      {stage0_3[24]},
      {stage1_4[13],stage1_3[13],stage1_2[13],stage1_1[13],stage1_0[13]}
   );
   gpc1163_5 gpc14 (
      {stage0_0[64], stage0_0[65], stage0_0[66]},
      {stage0_1[51], stage0_1[52], stage0_1[53], stage0_1[54], stage0_1[55], stage0_1[56]},
      {stage0_2[14]},
      {stage0_3[25]},
      {stage1_4[14],stage1_3[14],stage1_2[14],stage1_1[14],stage1_0[14]}
   );
   gpc1163_5 gpc15 (
      {stage0_0[67], stage0_0[68], stage0_0[69]},
      {stage0_1[57], stage0_1[58], stage0_1[59], stage0_1[60], stage0_1[61], stage0_1[62]},
      {stage0_2[15]},
      {stage0_3[26]},
      {stage1_4[15],stage1_3[15],stage1_2[15],stage1_1[15],stage1_0[15]}
   );
   gpc1163_5 gpc16 (
      {stage0_0[70], stage0_0[71], stage0_0[72]},
      {stage0_1[63], stage0_1[64], stage0_1[65], stage0_1[66], stage0_1[67], stage0_1[68]},
      {stage0_2[16]},
      {stage0_3[27]},
      {stage1_4[16],stage1_3[16],stage1_2[16],stage1_1[16],stage1_0[16]}
   );
   gpc1163_5 gpc17 (
      {stage0_0[73], stage0_0[74], stage0_0[75]},
      {stage0_1[69], stage0_1[70], stage0_1[71], stage0_1[72], stage0_1[73], stage0_1[74]},
      {stage0_2[17]},
      {stage0_3[28]},
      {stage1_4[17],stage1_3[17],stage1_2[17],stage1_1[17],stage1_0[17]}
   );
   gpc1163_5 gpc18 (
      {stage0_0[76], stage0_0[77], stage0_0[78]},
      {stage0_1[75], stage0_1[76], stage0_1[77], stage0_1[78], stage0_1[79], stage0_1[80]},
      {stage0_2[18]},
      {stage0_3[29]},
      {stage1_4[18],stage1_3[18],stage1_2[18],stage1_1[18],stage1_0[18]}
   );
   gpc1163_5 gpc19 (
      {stage0_0[79], stage0_0[80], stage0_0[81]},
      {stage0_1[81], stage0_1[82], stage0_1[83], stage0_1[84], stage0_1[85], stage0_1[86]},
      {stage0_2[19]},
      {stage0_3[30]},
      {stage1_4[19],stage1_3[19],stage1_2[19],stage1_1[19],stage1_0[19]}
   );
   gpc1163_5 gpc20 (
      {stage0_0[82], stage0_0[83], stage0_0[84]},
      {stage0_1[87], stage0_1[88], stage0_1[89], stage0_1[90], stage0_1[91], stage0_1[92]},
      {stage0_2[20]},
      {stage0_3[31]},
      {stage1_4[20],stage1_3[20],stage1_2[20],stage1_1[20],stage1_0[20]}
   );
   gpc1163_5 gpc21 (
      {stage0_0[85], stage0_0[86], stage0_0[87]},
      {stage0_1[93], stage0_1[94], stage0_1[95], stage0_1[96], stage0_1[97], stage0_1[98]},
      {stage0_2[21]},
      {stage0_3[32]},
      {stage1_4[21],stage1_3[21],stage1_2[21],stage1_1[21],stage1_0[21]}
   );
   gpc1163_5 gpc22 (
      {stage0_0[88], stage0_0[89], stage0_0[90]},
      {stage0_1[99], stage0_1[100], stage0_1[101], stage0_1[102], stage0_1[103], stage0_1[104]},
      {stage0_2[22]},
      {stage0_3[33]},
      {stage1_4[22],stage1_3[22],stage1_2[22],stage1_1[22],stage1_0[22]}
   );
   gpc1163_5 gpc23 (
      {stage0_0[91], stage0_0[92], stage0_0[93]},
      {stage0_1[105], stage0_1[106], stage0_1[107], stage0_1[108], stage0_1[109], stage0_1[110]},
      {stage0_2[23]},
      {stage0_3[34]},
      {stage1_4[23],stage1_3[23],stage1_2[23],stage1_1[23],stage1_0[23]}
   );
   gpc1163_5 gpc24 (
      {stage0_0[94], stage0_0[95], stage0_0[96]},
      {stage0_1[111], stage0_1[112], stage0_1[113], stage0_1[114], stage0_1[115], stage0_1[116]},
      {stage0_2[24]},
      {stage0_3[35]},
      {stage1_4[24],stage1_3[24],stage1_2[24],stage1_1[24],stage1_0[24]}
   );
   gpc1163_5 gpc25 (
      {stage0_0[97], stage0_0[98], stage0_0[99]},
      {stage0_1[117], stage0_1[118], stage0_1[119], stage0_1[120], stage0_1[121], stage0_1[122]},
      {stage0_2[25]},
      {stage0_3[36]},
      {stage1_4[25],stage1_3[25],stage1_2[25],stage1_1[25],stage1_0[25]}
   );
   gpc1163_5 gpc26 (
      {stage0_0[100], stage0_0[101], stage0_0[102]},
      {stage0_1[123], stage0_1[124], stage0_1[125], stage0_1[126], stage0_1[127], stage0_1[128]},
      {stage0_2[26]},
      {stage0_3[37]},
      {stage1_4[26],stage1_3[26],stage1_2[26],stage1_1[26],stage1_0[26]}
   );
   gpc1163_5 gpc27 (
      {stage0_0[103], stage0_0[104], stage0_0[105]},
      {stage0_1[129], stage0_1[130], stage0_1[131], stage0_1[132], stage0_1[133], stage0_1[134]},
      {stage0_2[27]},
      {stage0_3[38]},
      {stage1_4[27],stage1_3[27],stage1_2[27],stage1_1[27],stage1_0[27]}
   );
   gpc1163_5 gpc28 (
      {stage0_0[106], stage0_0[107], stage0_0[108]},
      {stage0_1[135], stage0_1[136], stage0_1[137], stage0_1[138], stage0_1[139], stage0_1[140]},
      {stage0_2[28]},
      {stage0_3[39]},
      {stage1_4[28],stage1_3[28],stage1_2[28],stage1_1[28],stage1_0[28]}
   );
   gpc1163_5 gpc29 (
      {stage0_0[109], stage0_0[110], stage0_0[111]},
      {stage0_1[141], stage0_1[142], stage0_1[143], stage0_1[144], stage0_1[145], stage0_1[146]},
      {stage0_2[29]},
      {stage0_3[40]},
      {stage1_4[29],stage1_3[29],stage1_2[29],stage1_1[29],stage1_0[29]}
   );
   gpc1163_5 gpc30 (
      {stage0_0[112], stage0_0[113], stage0_0[114]},
      {stage0_1[147], stage0_1[148], stage0_1[149], stage0_1[150], stage0_1[151], stage0_1[152]},
      {stage0_2[30]},
      {stage0_3[41]},
      {stage1_4[30],stage1_3[30],stage1_2[30],stage1_1[30],stage1_0[30]}
   );
   gpc1163_5 gpc31 (
      {stage0_0[115], stage0_0[116], stage0_0[117]},
      {stage0_1[153], stage0_1[154], stage0_1[155], stage0_1[156], stage0_1[157], stage0_1[158]},
      {stage0_2[31]},
      {stage0_3[42]},
      {stage1_4[31],stage1_3[31],stage1_2[31],stage1_1[31],stage1_0[31]}
   );
   gpc1163_5 gpc32 (
      {stage0_0[118], stage0_0[119], stage0_0[120]},
      {stage0_1[159], stage0_1[160], stage0_1[161], stage0_1[162], stage0_1[163], stage0_1[164]},
      {stage0_2[32]},
      {stage0_3[43]},
      {stage1_4[32],stage1_3[32],stage1_2[32],stage1_1[32],stage1_0[32]}
   );
   gpc1163_5 gpc33 (
      {stage0_0[121], stage0_0[122], stage0_0[123]},
      {stage0_1[165], stage0_1[166], stage0_1[167], stage0_1[168], stage0_1[169], stage0_1[170]},
      {stage0_2[33]},
      {stage0_3[44]},
      {stage1_4[33],stage1_3[33],stage1_2[33],stage1_1[33],stage1_0[33]}
   );
   gpc1163_5 gpc34 (
      {stage0_0[124], stage0_0[125], stage0_0[126]},
      {stage0_1[171], stage0_1[172], stage0_1[173], stage0_1[174], stage0_1[175], stage0_1[176]},
      {stage0_2[34]},
      {stage0_3[45]},
      {stage1_4[34],stage1_3[34],stage1_2[34],stage1_1[34],stage1_0[34]}
   );
   gpc1163_5 gpc35 (
      {stage0_0[127], stage0_0[128], stage0_0[129]},
      {stage0_1[177], stage0_1[178], stage0_1[179], stage0_1[180], stage0_1[181], stage0_1[182]},
      {stage0_2[35]},
      {stage0_3[46]},
      {stage1_4[35],stage1_3[35],stage1_2[35],stage1_1[35],stage1_0[35]}
   );
   gpc1163_5 gpc36 (
      {stage0_0[130], stage0_0[131], stage0_0[132]},
      {stage0_1[183], stage0_1[184], stage0_1[185], stage0_1[186], stage0_1[187], stage0_1[188]},
      {stage0_2[36]},
      {stage0_3[47]},
      {stage1_4[36],stage1_3[36],stage1_2[36],stage1_1[36],stage1_0[36]}
   );
   gpc1163_5 gpc37 (
      {stage0_0[133], stage0_0[134], stage0_0[135]},
      {stage0_1[189], stage0_1[190], stage0_1[191], stage0_1[192], stage0_1[193], stage0_1[194]},
      {stage0_2[37]},
      {stage0_3[48]},
      {stage1_4[37],stage1_3[37],stage1_2[37],stage1_1[37],stage1_0[37]}
   );
   gpc1163_5 gpc38 (
      {stage0_0[136], stage0_0[137], stage0_0[138]},
      {stage0_1[195], stage0_1[196], stage0_1[197], stage0_1[198], stage0_1[199], stage0_1[200]},
      {stage0_2[38]},
      {stage0_3[49]},
      {stage1_4[38],stage1_3[38],stage1_2[38],stage1_1[38],stage1_0[38]}
   );
   gpc1163_5 gpc39 (
      {stage0_0[139], stage0_0[140], stage0_0[141]},
      {stage0_1[201], stage0_1[202], stage0_1[203], stage0_1[204], stage0_1[205], stage0_1[206]},
      {stage0_2[39]},
      {stage0_3[50]},
      {stage1_4[39],stage1_3[39],stage1_2[39],stage1_1[39],stage1_0[39]}
   );
   gpc1163_5 gpc40 (
      {stage0_0[142], stage0_0[143], stage0_0[144]},
      {stage0_1[207], stage0_1[208], stage0_1[209], stage0_1[210], stage0_1[211], stage0_1[212]},
      {stage0_2[40]},
      {stage0_3[51]},
      {stage1_4[40],stage1_3[40],stage1_2[40],stage1_1[40],stage1_0[40]}
   );
   gpc1163_5 gpc41 (
      {stage0_0[145], stage0_0[146], stage0_0[147]},
      {stage0_1[213], stage0_1[214], stage0_1[215], stage0_1[216], stage0_1[217], stage0_1[218]},
      {stage0_2[41]},
      {stage0_3[52]},
      {stage1_4[41],stage1_3[41],stage1_2[41],stage1_1[41],stage1_0[41]}
   );
   gpc606_5 gpc42 (
      {stage0_0[148], stage0_0[149], stage0_0[150], stage0_0[151], stage0_0[152], stage0_0[153]},
      {stage0_2[42], stage0_2[43], stage0_2[44], stage0_2[45], stage0_2[46], stage0_2[47]},
      {stage1_4[42],stage1_3[42],stage1_2[42],stage1_1[42],stage1_0[42]}
   );
   gpc606_5 gpc43 (
      {stage0_0[154], stage0_0[155], stage0_0[156], stage0_0[157], stage0_0[158], stage0_0[159]},
      {stage0_2[48], stage0_2[49], stage0_2[50], stage0_2[51], stage0_2[52], stage0_2[53]},
      {stage1_4[43],stage1_3[43],stage1_2[43],stage1_1[43],stage1_0[43]}
   );
   gpc606_5 gpc44 (
      {stage0_0[160], stage0_0[161], stage0_0[162], stage0_0[163], stage0_0[164], stage0_0[165]},
      {stage0_2[54], stage0_2[55], stage0_2[56], stage0_2[57], stage0_2[58], stage0_2[59]},
      {stage1_4[44],stage1_3[44],stage1_2[44],stage1_1[44],stage1_0[44]}
   );
   gpc606_5 gpc45 (
      {stage0_0[166], stage0_0[167], stage0_0[168], stage0_0[169], stage0_0[170], stage0_0[171]},
      {stage0_2[60], stage0_2[61], stage0_2[62], stage0_2[63], stage0_2[64], stage0_2[65]},
      {stage1_4[45],stage1_3[45],stage1_2[45],stage1_1[45],stage1_0[45]}
   );
   gpc606_5 gpc46 (
      {stage0_0[172], stage0_0[173], stage0_0[174], stage0_0[175], stage0_0[176], stage0_0[177]},
      {stage0_2[66], stage0_2[67], stage0_2[68], stage0_2[69], stage0_2[70], stage0_2[71]},
      {stage1_4[46],stage1_3[46],stage1_2[46],stage1_1[46],stage1_0[46]}
   );
   gpc606_5 gpc47 (
      {stage0_0[178], stage0_0[179], stage0_0[180], stage0_0[181], stage0_0[182], stage0_0[183]},
      {stage0_2[72], stage0_2[73], stage0_2[74], stage0_2[75], stage0_2[76], stage0_2[77]},
      {stage1_4[47],stage1_3[47],stage1_2[47],stage1_1[47],stage1_0[47]}
   );
   gpc606_5 gpc48 (
      {stage0_0[184], stage0_0[185], stage0_0[186], stage0_0[187], stage0_0[188], stage0_0[189]},
      {stage0_2[78], stage0_2[79], stage0_2[80], stage0_2[81], stage0_2[82], stage0_2[83]},
      {stage1_4[48],stage1_3[48],stage1_2[48],stage1_1[48],stage1_0[48]}
   );
   gpc606_5 gpc49 (
      {stage0_0[190], stage0_0[191], stage0_0[192], stage0_0[193], stage0_0[194], stage0_0[195]},
      {stage0_2[84], stage0_2[85], stage0_2[86], stage0_2[87], stage0_2[88], stage0_2[89]},
      {stage1_4[49],stage1_3[49],stage1_2[49],stage1_1[49],stage1_0[49]}
   );
   gpc606_5 gpc50 (
      {stage0_0[196], stage0_0[197], stage0_0[198], stage0_0[199], stage0_0[200], stage0_0[201]},
      {stage0_2[90], stage0_2[91], stage0_2[92], stage0_2[93], stage0_2[94], stage0_2[95]},
      {stage1_4[50],stage1_3[50],stage1_2[50],stage1_1[50],stage1_0[50]}
   );
   gpc606_5 gpc51 (
      {stage0_0[202], stage0_0[203], stage0_0[204], stage0_0[205], stage0_0[206], stage0_0[207]},
      {stage0_2[96], stage0_2[97], stage0_2[98], stage0_2[99], stage0_2[100], stage0_2[101]},
      {stage1_4[51],stage1_3[51],stage1_2[51],stage1_1[51],stage1_0[51]}
   );
   gpc606_5 gpc52 (
      {stage0_0[208], stage0_0[209], stage0_0[210], stage0_0[211], stage0_0[212], stage0_0[213]},
      {stage0_2[102], stage0_2[103], stage0_2[104], stage0_2[105], stage0_2[106], stage0_2[107]},
      {stage1_4[52],stage1_3[52],stage1_2[52],stage1_1[52],stage1_0[52]}
   );
   gpc606_5 gpc53 (
      {stage0_0[214], stage0_0[215], stage0_0[216], stage0_0[217], stage0_0[218], stage0_0[219]},
      {stage0_2[108], stage0_2[109], stage0_2[110], stage0_2[111], stage0_2[112], stage0_2[113]},
      {stage1_4[53],stage1_3[53],stage1_2[53],stage1_1[53],stage1_0[53]}
   );
   gpc606_5 gpc54 (
      {stage0_0[220], stage0_0[221], stage0_0[222], stage0_0[223], stage0_0[224], stage0_0[225]},
      {stage0_2[114], stage0_2[115], stage0_2[116], stage0_2[117], stage0_2[118], stage0_2[119]},
      {stage1_4[54],stage1_3[54],stage1_2[54],stage1_1[54],stage1_0[54]}
   );
   gpc606_5 gpc55 (
      {stage0_0[226], stage0_0[227], stage0_0[228], stage0_0[229], stage0_0[230], stage0_0[231]},
      {stage0_2[120], stage0_2[121], stage0_2[122], stage0_2[123], stage0_2[124], stage0_2[125]},
      {stage1_4[55],stage1_3[55],stage1_2[55],stage1_1[55],stage1_0[55]}
   );
   gpc606_5 gpc56 (
      {stage0_0[232], stage0_0[233], stage0_0[234], stage0_0[235], stage0_0[236], stage0_0[237]},
      {stage0_2[126], stage0_2[127], stage0_2[128], stage0_2[129], stage0_2[130], stage0_2[131]},
      {stage1_4[56],stage1_3[56],stage1_2[56],stage1_1[56],stage1_0[56]}
   );
   gpc606_5 gpc57 (
      {stage0_0[238], stage0_0[239], stage0_0[240], stage0_0[241], stage0_0[242], stage0_0[243]},
      {stage0_2[132], stage0_2[133], stage0_2[134], stage0_2[135], stage0_2[136], stage0_2[137]},
      {stage1_4[57],stage1_3[57],stage1_2[57],stage1_1[57],stage1_0[57]}
   );
   gpc606_5 gpc58 (
      {stage0_0[244], stage0_0[245], stage0_0[246], stage0_0[247], stage0_0[248], stage0_0[249]},
      {stage0_2[138], stage0_2[139], stage0_2[140], stage0_2[141], stage0_2[142], stage0_2[143]},
      {stage1_4[58],stage1_3[58],stage1_2[58],stage1_1[58],stage1_0[58]}
   );
   gpc606_5 gpc59 (
      {stage0_0[250], stage0_0[251], stage0_0[252], stage0_0[253], stage0_0[254], stage0_0[255]},
      {stage0_2[144], stage0_2[145], stage0_2[146], stage0_2[147], stage0_2[148], stage0_2[149]},
      {stage1_4[59],stage1_3[59],stage1_2[59],stage1_1[59],stage1_0[59]}
   );
   gpc606_5 gpc60 (
      {stage0_0[256], stage0_0[257], stage0_0[258], stage0_0[259], stage0_0[260], stage0_0[261]},
      {stage0_2[150], stage0_2[151], stage0_2[152], stage0_2[153], stage0_2[154], stage0_2[155]},
      {stage1_4[60],stage1_3[60],stage1_2[60],stage1_1[60],stage1_0[60]}
   );
   gpc606_5 gpc61 (
      {stage0_0[262], stage0_0[263], stage0_0[264], stage0_0[265], stage0_0[266], stage0_0[267]},
      {stage0_2[156], stage0_2[157], stage0_2[158], stage0_2[159], stage0_2[160], stage0_2[161]},
      {stage1_4[61],stage1_3[61],stage1_2[61],stage1_1[61],stage1_0[61]}
   );
   gpc606_5 gpc62 (
      {stage0_0[268], stage0_0[269], stage0_0[270], stage0_0[271], stage0_0[272], stage0_0[273]},
      {stage0_2[162], stage0_2[163], stage0_2[164], stage0_2[165], stage0_2[166], stage0_2[167]},
      {stage1_4[62],stage1_3[62],stage1_2[62],stage1_1[62],stage1_0[62]}
   );
   gpc606_5 gpc63 (
      {stage0_0[274], stage0_0[275], stage0_0[276], stage0_0[277], stage0_0[278], stage0_0[279]},
      {stage0_2[168], stage0_2[169], stage0_2[170], stage0_2[171], stage0_2[172], stage0_2[173]},
      {stage1_4[63],stage1_3[63],stage1_2[63],stage1_1[63],stage1_0[63]}
   );
   gpc606_5 gpc64 (
      {stage0_0[280], stage0_0[281], stage0_0[282], stage0_0[283], stage0_0[284], stage0_0[285]},
      {stage0_2[174], stage0_2[175], stage0_2[176], stage0_2[177], stage0_2[178], stage0_2[179]},
      {stage1_4[64],stage1_3[64],stage1_2[64],stage1_1[64],stage1_0[64]}
   );
   gpc606_5 gpc65 (
      {stage0_0[286], stage0_0[287], stage0_0[288], stage0_0[289], stage0_0[290], stage0_0[291]},
      {stage0_2[180], stage0_2[181], stage0_2[182], stage0_2[183], stage0_2[184], stage0_2[185]},
      {stage1_4[65],stage1_3[65],stage1_2[65],stage1_1[65],stage1_0[65]}
   );
   gpc606_5 gpc66 (
      {stage0_0[292], stage0_0[293], stage0_0[294], stage0_0[295], stage0_0[296], stage0_0[297]},
      {stage0_2[186], stage0_2[187], stage0_2[188], stage0_2[189], stage0_2[190], stage0_2[191]},
      {stage1_4[66],stage1_3[66],stage1_2[66],stage1_1[66],stage1_0[66]}
   );
   gpc606_5 gpc67 (
      {stage0_0[298], stage0_0[299], stage0_0[300], stage0_0[301], stage0_0[302], stage0_0[303]},
      {stage0_2[192], stage0_2[193], stage0_2[194], stage0_2[195], stage0_2[196], stage0_2[197]},
      {stage1_4[67],stage1_3[67],stage1_2[67],stage1_1[67],stage1_0[67]}
   );
   gpc606_5 gpc68 (
      {stage0_0[304], stage0_0[305], stage0_0[306], stage0_0[307], stage0_0[308], stage0_0[309]},
      {stage0_2[198], stage0_2[199], stage0_2[200], stage0_2[201], stage0_2[202], stage0_2[203]},
      {stage1_4[68],stage1_3[68],stage1_2[68],stage1_1[68],stage1_0[68]}
   );
   gpc606_5 gpc69 (
      {stage0_0[310], stage0_0[311], stage0_0[312], stage0_0[313], stage0_0[314], stage0_0[315]},
      {stage0_2[204], stage0_2[205], stage0_2[206], stage0_2[207], stage0_2[208], stage0_2[209]},
      {stage1_4[69],stage1_3[69],stage1_2[69],stage1_1[69],stage1_0[69]}
   );
   gpc606_5 gpc70 (
      {stage0_0[316], stage0_0[317], stage0_0[318], stage0_0[319], stage0_0[320], stage0_0[321]},
      {stage0_2[210], stage0_2[211], stage0_2[212], stage0_2[213], stage0_2[214], stage0_2[215]},
      {stage1_4[70],stage1_3[70],stage1_2[70],stage1_1[70],stage1_0[70]}
   );
   gpc606_5 gpc71 (
      {stage0_0[322], stage0_0[323], stage0_0[324], stage0_0[325], stage0_0[326], stage0_0[327]},
      {stage0_2[216], stage0_2[217], stage0_2[218], stage0_2[219], stage0_2[220], stage0_2[221]},
      {stage1_4[71],stage1_3[71],stage1_2[71],stage1_1[71],stage1_0[71]}
   );
   gpc606_5 gpc72 (
      {stage0_0[328], stage0_0[329], stage0_0[330], stage0_0[331], stage0_0[332], stage0_0[333]},
      {stage0_2[222], stage0_2[223], stage0_2[224], stage0_2[225], stage0_2[226], stage0_2[227]},
      {stage1_4[72],stage1_3[72],stage1_2[72],stage1_1[72],stage1_0[72]}
   );
   gpc606_5 gpc73 (
      {stage0_0[334], stage0_0[335], stage0_0[336], stage0_0[337], stage0_0[338], stage0_0[339]},
      {stage0_2[228], stage0_2[229], stage0_2[230], stage0_2[231], stage0_2[232], stage0_2[233]},
      {stage1_4[73],stage1_3[73],stage1_2[73],stage1_1[73],stage1_0[73]}
   );
   gpc606_5 gpc74 (
      {stage0_0[340], stage0_0[341], stage0_0[342], stage0_0[343], stage0_0[344], stage0_0[345]},
      {stage0_2[234], stage0_2[235], stage0_2[236], stage0_2[237], stage0_2[238], stage0_2[239]},
      {stage1_4[74],stage1_3[74],stage1_2[74],stage1_1[74],stage1_0[74]}
   );
   gpc606_5 gpc75 (
      {stage0_0[346], stage0_0[347], stage0_0[348], stage0_0[349], stage0_0[350], stage0_0[351]},
      {stage0_2[240], stage0_2[241], stage0_2[242], stage0_2[243], stage0_2[244], stage0_2[245]},
      {stage1_4[75],stage1_3[75],stage1_2[75],stage1_1[75],stage1_0[75]}
   );
   gpc606_5 gpc76 (
      {stage0_0[352], stage0_0[353], stage0_0[354], stage0_0[355], stage0_0[356], stage0_0[357]},
      {stage0_2[246], stage0_2[247], stage0_2[248], stage0_2[249], stage0_2[250], stage0_2[251]},
      {stage1_4[76],stage1_3[76],stage1_2[76],stage1_1[76],stage1_0[76]}
   );
   gpc606_5 gpc77 (
      {stage0_0[358], stage0_0[359], stage0_0[360], stage0_0[361], stage0_0[362], stage0_0[363]},
      {stage0_2[252], stage0_2[253], stage0_2[254], stage0_2[255], stage0_2[256], stage0_2[257]},
      {stage1_4[77],stage1_3[77],stage1_2[77],stage1_1[77],stage1_0[77]}
   );
   gpc606_5 gpc78 (
      {stage0_0[364], stage0_0[365], stage0_0[366], stage0_0[367], stage0_0[368], stage0_0[369]},
      {stage0_2[258], stage0_2[259], stage0_2[260], stage0_2[261], stage0_2[262], stage0_2[263]},
      {stage1_4[78],stage1_3[78],stage1_2[78],stage1_1[78],stage1_0[78]}
   );
   gpc606_5 gpc79 (
      {stage0_0[370], stage0_0[371], stage0_0[372], stage0_0[373], stage0_0[374], stage0_0[375]},
      {stage0_2[264], stage0_2[265], stage0_2[266], stage0_2[267], stage0_2[268], stage0_2[269]},
      {stage1_4[79],stage1_3[79],stage1_2[79],stage1_1[79],stage1_0[79]}
   );
   gpc606_5 gpc80 (
      {stage0_0[376], stage0_0[377], stage0_0[378], stage0_0[379], stage0_0[380], stage0_0[381]},
      {stage0_2[270], stage0_2[271], stage0_2[272], stage0_2[273], stage0_2[274], stage0_2[275]},
      {stage1_4[80],stage1_3[80],stage1_2[80],stage1_1[80],stage1_0[80]}
   );
   gpc606_5 gpc81 (
      {stage0_0[382], stage0_0[383], stage0_0[384], stage0_0[385], stage0_0[386], stage0_0[387]},
      {stage0_2[276], stage0_2[277], stage0_2[278], stage0_2[279], stage0_2[280], stage0_2[281]},
      {stage1_4[81],stage1_3[81],stage1_2[81],stage1_1[81],stage1_0[81]}
   );
   gpc606_5 gpc82 (
      {stage0_0[388], stage0_0[389], stage0_0[390], stage0_0[391], stage0_0[392], stage0_0[393]},
      {stage0_2[282], stage0_2[283], stage0_2[284], stage0_2[285], stage0_2[286], stage0_2[287]},
      {stage1_4[82],stage1_3[82],stage1_2[82],stage1_1[82],stage1_0[82]}
   );
   gpc606_5 gpc83 (
      {stage0_0[394], stage0_0[395], stage0_0[396], stage0_0[397], stage0_0[398], stage0_0[399]},
      {stage0_2[288], stage0_2[289], stage0_2[290], stage0_2[291], stage0_2[292], stage0_2[293]},
      {stage1_4[83],stage1_3[83],stage1_2[83],stage1_1[83],stage1_0[83]}
   );
   gpc606_5 gpc84 (
      {stage0_0[400], stage0_0[401], stage0_0[402], stage0_0[403], stage0_0[404], stage0_0[405]},
      {stage0_2[294], stage0_2[295], stage0_2[296], stage0_2[297], stage0_2[298], stage0_2[299]},
      {stage1_4[84],stage1_3[84],stage1_2[84],stage1_1[84],stage1_0[84]}
   );
   gpc606_5 gpc85 (
      {stage0_0[406], stage0_0[407], stage0_0[408], stage0_0[409], stage0_0[410], stage0_0[411]},
      {stage0_2[300], stage0_2[301], stage0_2[302], stage0_2[303], stage0_2[304], stage0_2[305]},
      {stage1_4[85],stage1_3[85],stage1_2[85],stage1_1[85],stage1_0[85]}
   );
   gpc606_5 gpc86 (
      {stage0_0[412], stage0_0[413], stage0_0[414], stage0_0[415], stage0_0[416], stage0_0[417]},
      {stage0_2[306], stage0_2[307], stage0_2[308], stage0_2[309], stage0_2[310], stage0_2[311]},
      {stage1_4[86],stage1_3[86],stage1_2[86],stage1_1[86],stage1_0[86]}
   );
   gpc606_5 gpc87 (
      {stage0_0[418], stage0_0[419], stage0_0[420], stage0_0[421], stage0_0[422], stage0_0[423]},
      {stage0_2[312], stage0_2[313], stage0_2[314], stage0_2[315], stage0_2[316], stage0_2[317]},
      {stage1_4[87],stage1_3[87],stage1_2[87],stage1_1[87],stage1_0[87]}
   );
   gpc606_5 gpc88 (
      {stage0_0[424], stage0_0[425], stage0_0[426], stage0_0[427], stage0_0[428], stage0_0[429]},
      {stage0_2[318], stage0_2[319], stage0_2[320], stage0_2[321], stage0_2[322], stage0_2[323]},
      {stage1_4[88],stage1_3[88],stage1_2[88],stage1_1[88],stage1_0[88]}
   );
   gpc606_5 gpc89 (
      {stage0_0[430], stage0_0[431], stage0_0[432], stage0_0[433], stage0_0[434], stage0_0[435]},
      {stage0_2[324], stage0_2[325], stage0_2[326], stage0_2[327], stage0_2[328], stage0_2[329]},
      {stage1_4[89],stage1_3[89],stage1_2[89],stage1_1[89],stage1_0[89]}
   );
   gpc606_5 gpc90 (
      {stage0_0[436], stage0_0[437], stage0_0[438], stage0_0[439], stage0_0[440], stage0_0[441]},
      {stage0_2[330], stage0_2[331], stage0_2[332], stage0_2[333], stage0_2[334], stage0_2[335]},
      {stage1_4[90],stage1_3[90],stage1_2[90],stage1_1[90],stage1_0[90]}
   );
   gpc606_5 gpc91 (
      {stage0_0[442], stage0_0[443], stage0_0[444], stage0_0[445], stage0_0[446], stage0_0[447]},
      {stage0_2[336], stage0_2[337], stage0_2[338], stage0_2[339], stage0_2[340], stage0_2[341]},
      {stage1_4[91],stage1_3[91],stage1_2[91],stage1_1[91],stage1_0[91]}
   );
   gpc606_5 gpc92 (
      {stage0_0[448], stage0_0[449], stage0_0[450], stage0_0[451], stage0_0[452], stage0_0[453]},
      {stage0_2[342], stage0_2[343], stage0_2[344], stage0_2[345], stage0_2[346], stage0_2[347]},
      {stage1_4[92],stage1_3[92],stage1_2[92],stage1_1[92],stage1_0[92]}
   );
   gpc606_5 gpc93 (
      {stage0_0[454], stage0_0[455], stage0_0[456], stage0_0[457], stage0_0[458], stage0_0[459]},
      {stage0_2[348], stage0_2[349], stage0_2[350], stage0_2[351], stage0_2[352], stage0_2[353]},
      {stage1_4[93],stage1_3[93],stage1_2[93],stage1_1[93],stage1_0[93]}
   );
   gpc606_5 gpc94 (
      {stage0_0[460], stage0_0[461], stage0_0[462], stage0_0[463], stage0_0[464], stage0_0[465]},
      {stage0_2[354], stage0_2[355], stage0_2[356], stage0_2[357], stage0_2[358], stage0_2[359]},
      {stage1_4[94],stage1_3[94],stage1_2[94],stage1_1[94],stage1_0[94]}
   );
   gpc606_5 gpc95 (
      {stage0_0[466], stage0_0[467], stage0_0[468], stage0_0[469], stage0_0[470], stage0_0[471]},
      {stage0_2[360], stage0_2[361], stage0_2[362], stage0_2[363], stage0_2[364], stage0_2[365]},
      {stage1_4[95],stage1_3[95],stage1_2[95],stage1_1[95],stage1_0[95]}
   );
   gpc606_5 gpc96 (
      {stage0_0[472], stage0_0[473], stage0_0[474], stage0_0[475], stage0_0[476], stage0_0[477]},
      {stage0_2[366], stage0_2[367], stage0_2[368], stage0_2[369], stage0_2[370], stage0_2[371]},
      {stage1_4[96],stage1_3[96],stage1_2[96],stage1_1[96],stage1_0[96]}
   );
   gpc606_5 gpc97 (
      {stage0_0[478], stage0_0[479], stage0_0[480], stage0_0[481], stage0_0[482], stage0_0[483]},
      {stage0_2[372], stage0_2[373], stage0_2[374], stage0_2[375], stage0_2[376], stage0_2[377]},
      {stage1_4[97],stage1_3[97],stage1_2[97],stage1_1[97],stage1_0[97]}
   );
   gpc606_5 gpc98 (
      {stage0_0[484], stage0_0[485], stage0_0[486], stage0_0[487], stage0_0[488], stage0_0[489]},
      {stage0_2[378], stage0_2[379], stage0_2[380], stage0_2[381], stage0_2[382], stage0_2[383]},
      {stage1_4[98],stage1_3[98],stage1_2[98],stage1_1[98],stage1_0[98]}
   );
   gpc606_5 gpc99 (
      {stage0_0[490], stage0_0[491], stage0_0[492], stage0_0[493], stage0_0[494], stage0_0[495]},
      {stage0_2[384], stage0_2[385], stage0_2[386], stage0_2[387], stage0_2[388], stage0_2[389]},
      {stage1_4[99],stage1_3[99],stage1_2[99],stage1_1[99],stage1_0[99]}
   );
   gpc606_5 gpc100 (
      {stage0_0[496], stage0_0[497], stage0_0[498], stage0_0[499], stage0_0[500], stage0_0[501]},
      {stage0_2[390], stage0_2[391], stage0_2[392], stage0_2[393], stage0_2[394], stage0_2[395]},
      {stage1_4[100],stage1_3[100],stage1_2[100],stage1_1[100],stage1_0[100]}
   );
   gpc606_5 gpc101 (
      {stage0_1[219], stage0_1[220], stage0_1[221], stage0_1[222], stage0_1[223], stage0_1[224]},
      {stage0_3[53], stage0_3[54], stage0_3[55], stage0_3[56], stage0_3[57], stage0_3[58]},
      {stage1_5[0],stage1_4[101],stage1_3[101],stage1_2[101],stage1_1[101]}
   );
   gpc606_5 gpc102 (
      {stage0_1[225], stage0_1[226], stage0_1[227], stage0_1[228], stage0_1[229], stage0_1[230]},
      {stage0_3[59], stage0_3[60], stage0_3[61], stage0_3[62], stage0_3[63], stage0_3[64]},
      {stage1_5[1],stage1_4[102],stage1_3[102],stage1_2[102],stage1_1[102]}
   );
   gpc606_5 gpc103 (
      {stage0_1[231], stage0_1[232], stage0_1[233], stage0_1[234], stage0_1[235], stage0_1[236]},
      {stage0_3[65], stage0_3[66], stage0_3[67], stage0_3[68], stage0_3[69], stage0_3[70]},
      {stage1_5[2],stage1_4[103],stage1_3[103],stage1_2[103],stage1_1[103]}
   );
   gpc606_5 gpc104 (
      {stage0_1[237], stage0_1[238], stage0_1[239], stage0_1[240], stage0_1[241], stage0_1[242]},
      {stage0_3[71], stage0_3[72], stage0_3[73], stage0_3[74], stage0_3[75], stage0_3[76]},
      {stage1_5[3],stage1_4[104],stage1_3[104],stage1_2[104],stage1_1[104]}
   );
   gpc606_5 gpc105 (
      {stage0_1[243], stage0_1[244], stage0_1[245], stage0_1[246], stage0_1[247], stage0_1[248]},
      {stage0_3[77], stage0_3[78], stage0_3[79], stage0_3[80], stage0_3[81], stage0_3[82]},
      {stage1_5[4],stage1_4[105],stage1_3[105],stage1_2[105],stage1_1[105]}
   );
   gpc606_5 gpc106 (
      {stage0_1[249], stage0_1[250], stage0_1[251], stage0_1[252], stage0_1[253], stage0_1[254]},
      {stage0_3[83], stage0_3[84], stage0_3[85], stage0_3[86], stage0_3[87], stage0_3[88]},
      {stage1_5[5],stage1_4[106],stage1_3[106],stage1_2[106],stage1_1[106]}
   );
   gpc606_5 gpc107 (
      {stage0_1[255], stage0_1[256], stage0_1[257], stage0_1[258], stage0_1[259], stage0_1[260]},
      {stage0_3[89], stage0_3[90], stage0_3[91], stage0_3[92], stage0_3[93], stage0_3[94]},
      {stage1_5[6],stage1_4[107],stage1_3[107],stage1_2[107],stage1_1[107]}
   );
   gpc606_5 gpc108 (
      {stage0_1[261], stage0_1[262], stage0_1[263], stage0_1[264], stage0_1[265], stage0_1[266]},
      {stage0_3[95], stage0_3[96], stage0_3[97], stage0_3[98], stage0_3[99], stage0_3[100]},
      {stage1_5[7],stage1_4[108],stage1_3[108],stage1_2[108],stage1_1[108]}
   );
   gpc606_5 gpc109 (
      {stage0_1[267], stage0_1[268], stage0_1[269], stage0_1[270], stage0_1[271], stage0_1[272]},
      {stage0_3[101], stage0_3[102], stage0_3[103], stage0_3[104], stage0_3[105], stage0_3[106]},
      {stage1_5[8],stage1_4[109],stage1_3[109],stage1_2[109],stage1_1[109]}
   );
   gpc606_5 gpc110 (
      {stage0_1[273], stage0_1[274], stage0_1[275], stage0_1[276], stage0_1[277], stage0_1[278]},
      {stage0_3[107], stage0_3[108], stage0_3[109], stage0_3[110], stage0_3[111], stage0_3[112]},
      {stage1_5[9],stage1_4[110],stage1_3[110],stage1_2[110],stage1_1[110]}
   );
   gpc606_5 gpc111 (
      {stage0_1[279], stage0_1[280], stage0_1[281], stage0_1[282], stage0_1[283], stage0_1[284]},
      {stage0_3[113], stage0_3[114], stage0_3[115], stage0_3[116], stage0_3[117], stage0_3[118]},
      {stage1_5[10],stage1_4[111],stage1_3[111],stage1_2[111],stage1_1[111]}
   );
   gpc606_5 gpc112 (
      {stage0_1[285], stage0_1[286], stage0_1[287], stage0_1[288], stage0_1[289], stage0_1[290]},
      {stage0_3[119], stage0_3[120], stage0_3[121], stage0_3[122], stage0_3[123], stage0_3[124]},
      {stage1_5[11],stage1_4[112],stage1_3[112],stage1_2[112],stage1_1[112]}
   );
   gpc606_5 gpc113 (
      {stage0_1[291], stage0_1[292], stage0_1[293], stage0_1[294], stage0_1[295], stage0_1[296]},
      {stage0_3[125], stage0_3[126], stage0_3[127], stage0_3[128], stage0_3[129], stage0_3[130]},
      {stage1_5[12],stage1_4[113],stage1_3[113],stage1_2[113],stage1_1[113]}
   );
   gpc606_5 gpc114 (
      {stage0_1[297], stage0_1[298], stage0_1[299], stage0_1[300], stage0_1[301], stage0_1[302]},
      {stage0_3[131], stage0_3[132], stage0_3[133], stage0_3[134], stage0_3[135], stage0_3[136]},
      {stage1_5[13],stage1_4[114],stage1_3[114],stage1_2[114],stage1_1[114]}
   );
   gpc606_5 gpc115 (
      {stage0_1[303], stage0_1[304], stage0_1[305], stage0_1[306], stage0_1[307], stage0_1[308]},
      {stage0_3[137], stage0_3[138], stage0_3[139], stage0_3[140], stage0_3[141], stage0_3[142]},
      {stage1_5[14],stage1_4[115],stage1_3[115],stage1_2[115],stage1_1[115]}
   );
   gpc606_5 gpc116 (
      {stage0_1[309], stage0_1[310], stage0_1[311], stage0_1[312], stage0_1[313], stage0_1[314]},
      {stage0_3[143], stage0_3[144], stage0_3[145], stage0_3[146], stage0_3[147], stage0_3[148]},
      {stage1_5[15],stage1_4[116],stage1_3[116],stage1_2[116],stage1_1[116]}
   );
   gpc606_5 gpc117 (
      {stage0_1[315], stage0_1[316], stage0_1[317], stage0_1[318], stage0_1[319], stage0_1[320]},
      {stage0_3[149], stage0_3[150], stage0_3[151], stage0_3[152], stage0_3[153], stage0_3[154]},
      {stage1_5[16],stage1_4[117],stage1_3[117],stage1_2[117],stage1_1[117]}
   );
   gpc606_5 gpc118 (
      {stage0_1[321], stage0_1[322], stage0_1[323], stage0_1[324], stage0_1[325], stage0_1[326]},
      {stage0_3[155], stage0_3[156], stage0_3[157], stage0_3[158], stage0_3[159], stage0_3[160]},
      {stage1_5[17],stage1_4[118],stage1_3[118],stage1_2[118],stage1_1[118]}
   );
   gpc606_5 gpc119 (
      {stage0_1[327], stage0_1[328], stage0_1[329], stage0_1[330], stage0_1[331], stage0_1[332]},
      {stage0_3[161], stage0_3[162], stage0_3[163], stage0_3[164], stage0_3[165], stage0_3[166]},
      {stage1_5[18],stage1_4[119],stage1_3[119],stage1_2[119],stage1_1[119]}
   );
   gpc606_5 gpc120 (
      {stage0_1[333], stage0_1[334], stage0_1[335], stage0_1[336], stage0_1[337], stage0_1[338]},
      {stage0_3[167], stage0_3[168], stage0_3[169], stage0_3[170], stage0_3[171], stage0_3[172]},
      {stage1_5[19],stage1_4[120],stage1_3[120],stage1_2[120],stage1_1[120]}
   );
   gpc606_5 gpc121 (
      {stage0_1[339], stage0_1[340], stage0_1[341], stage0_1[342], stage0_1[343], stage0_1[344]},
      {stage0_3[173], stage0_3[174], stage0_3[175], stage0_3[176], stage0_3[177], stage0_3[178]},
      {stage1_5[20],stage1_4[121],stage1_3[121],stage1_2[121],stage1_1[121]}
   );
   gpc606_5 gpc122 (
      {stage0_1[345], stage0_1[346], stage0_1[347], stage0_1[348], stage0_1[349], stage0_1[350]},
      {stage0_3[179], stage0_3[180], stage0_3[181], stage0_3[182], stage0_3[183], stage0_3[184]},
      {stage1_5[21],stage1_4[122],stage1_3[122],stage1_2[122],stage1_1[122]}
   );
   gpc606_5 gpc123 (
      {stage0_1[351], stage0_1[352], stage0_1[353], stage0_1[354], stage0_1[355], stage0_1[356]},
      {stage0_3[185], stage0_3[186], stage0_3[187], stage0_3[188], stage0_3[189], stage0_3[190]},
      {stage1_5[22],stage1_4[123],stage1_3[123],stage1_2[123],stage1_1[123]}
   );
   gpc606_5 gpc124 (
      {stage0_1[357], stage0_1[358], stage0_1[359], stage0_1[360], stage0_1[361], stage0_1[362]},
      {stage0_3[191], stage0_3[192], stage0_3[193], stage0_3[194], stage0_3[195], stage0_3[196]},
      {stage1_5[23],stage1_4[124],stage1_3[124],stage1_2[124],stage1_1[124]}
   );
   gpc606_5 gpc125 (
      {stage0_1[363], stage0_1[364], stage0_1[365], stage0_1[366], stage0_1[367], stage0_1[368]},
      {stage0_3[197], stage0_3[198], stage0_3[199], stage0_3[200], stage0_3[201], stage0_3[202]},
      {stage1_5[24],stage1_4[125],stage1_3[125],stage1_2[125],stage1_1[125]}
   );
   gpc606_5 gpc126 (
      {stage0_1[369], stage0_1[370], stage0_1[371], stage0_1[372], stage0_1[373], stage0_1[374]},
      {stage0_3[203], stage0_3[204], stage0_3[205], stage0_3[206], stage0_3[207], stage0_3[208]},
      {stage1_5[25],stage1_4[126],stage1_3[126],stage1_2[126],stage1_1[126]}
   );
   gpc606_5 gpc127 (
      {stage0_1[375], stage0_1[376], stage0_1[377], stage0_1[378], stage0_1[379], stage0_1[380]},
      {stage0_3[209], stage0_3[210], stage0_3[211], stage0_3[212], stage0_3[213], stage0_3[214]},
      {stage1_5[26],stage1_4[127],stage1_3[127],stage1_2[127],stage1_1[127]}
   );
   gpc606_5 gpc128 (
      {stage0_1[381], stage0_1[382], stage0_1[383], stage0_1[384], stage0_1[385], stage0_1[386]},
      {stage0_3[215], stage0_3[216], stage0_3[217], stage0_3[218], stage0_3[219], stage0_3[220]},
      {stage1_5[27],stage1_4[128],stage1_3[128],stage1_2[128],stage1_1[128]}
   );
   gpc606_5 gpc129 (
      {stage0_1[387], stage0_1[388], stage0_1[389], stage0_1[390], stage0_1[391], stage0_1[392]},
      {stage0_3[221], stage0_3[222], stage0_3[223], stage0_3[224], stage0_3[225], stage0_3[226]},
      {stage1_5[28],stage1_4[129],stage1_3[129],stage1_2[129],stage1_1[129]}
   );
   gpc606_5 gpc130 (
      {stage0_1[393], stage0_1[394], stage0_1[395], stage0_1[396], stage0_1[397], stage0_1[398]},
      {stage0_3[227], stage0_3[228], stage0_3[229], stage0_3[230], stage0_3[231], stage0_3[232]},
      {stage1_5[29],stage1_4[130],stage1_3[130],stage1_2[130],stage1_1[130]}
   );
   gpc606_5 gpc131 (
      {stage0_1[399], stage0_1[400], stage0_1[401], stage0_1[402], stage0_1[403], stage0_1[404]},
      {stage0_3[233], stage0_3[234], stage0_3[235], stage0_3[236], stage0_3[237], stage0_3[238]},
      {stage1_5[30],stage1_4[131],stage1_3[131],stage1_2[131],stage1_1[131]}
   );
   gpc606_5 gpc132 (
      {stage0_1[405], stage0_1[406], stage0_1[407], stage0_1[408], stage0_1[409], stage0_1[410]},
      {stage0_3[239], stage0_3[240], stage0_3[241], stage0_3[242], stage0_3[243], stage0_3[244]},
      {stage1_5[31],stage1_4[132],stage1_3[132],stage1_2[132],stage1_1[132]}
   );
   gpc606_5 gpc133 (
      {stage0_1[411], stage0_1[412], stage0_1[413], stage0_1[414], stage0_1[415], stage0_1[416]},
      {stage0_3[245], stage0_3[246], stage0_3[247], stage0_3[248], stage0_3[249], stage0_3[250]},
      {stage1_5[32],stage1_4[133],stage1_3[133],stage1_2[133],stage1_1[133]}
   );
   gpc606_5 gpc134 (
      {stage0_1[417], stage0_1[418], stage0_1[419], stage0_1[420], stage0_1[421], stage0_1[422]},
      {stage0_3[251], stage0_3[252], stage0_3[253], stage0_3[254], stage0_3[255], stage0_3[256]},
      {stage1_5[33],stage1_4[134],stage1_3[134],stage1_2[134],stage1_1[134]}
   );
   gpc606_5 gpc135 (
      {stage0_1[423], stage0_1[424], stage0_1[425], stage0_1[426], stage0_1[427], stage0_1[428]},
      {stage0_3[257], stage0_3[258], stage0_3[259], stage0_3[260], stage0_3[261], stage0_3[262]},
      {stage1_5[34],stage1_4[135],stage1_3[135],stage1_2[135],stage1_1[135]}
   );
   gpc606_5 gpc136 (
      {stage0_1[429], stage0_1[430], stage0_1[431], stage0_1[432], stage0_1[433], stage0_1[434]},
      {stage0_3[263], stage0_3[264], stage0_3[265], stage0_3[266], stage0_3[267], stage0_3[268]},
      {stage1_5[35],stage1_4[136],stage1_3[136],stage1_2[136],stage1_1[136]}
   );
   gpc606_5 gpc137 (
      {stage0_1[435], stage0_1[436], stage0_1[437], stage0_1[438], stage0_1[439], stage0_1[440]},
      {stage0_3[269], stage0_3[270], stage0_3[271], stage0_3[272], stage0_3[273], stage0_3[274]},
      {stage1_5[36],stage1_4[137],stage1_3[137],stage1_2[137],stage1_1[137]}
   );
   gpc606_5 gpc138 (
      {stage0_1[441], stage0_1[442], stage0_1[443], stage0_1[444], stage0_1[445], stage0_1[446]},
      {stage0_3[275], stage0_3[276], stage0_3[277], stage0_3[278], stage0_3[279], stage0_3[280]},
      {stage1_5[37],stage1_4[138],stage1_3[138],stage1_2[138],stage1_1[138]}
   );
   gpc606_5 gpc139 (
      {stage0_1[447], stage0_1[448], stage0_1[449], stage0_1[450], stage0_1[451], stage0_1[452]},
      {stage0_3[281], stage0_3[282], stage0_3[283], stage0_3[284], stage0_3[285], stage0_3[286]},
      {stage1_5[38],stage1_4[139],stage1_3[139],stage1_2[139],stage1_1[139]}
   );
   gpc615_5 gpc140 (
      {stage0_2[396], stage0_2[397], stage0_2[398], stage0_2[399], stage0_2[400]},
      {stage0_3[287]},
      {stage0_4[0], stage0_4[1], stage0_4[2], stage0_4[3], stage0_4[4], stage0_4[5]},
      {stage1_6[0],stage1_5[39],stage1_4[140],stage1_3[140],stage1_2[140]}
   );
   gpc615_5 gpc141 (
      {stage0_2[401], stage0_2[402], stage0_2[403], stage0_2[404], stage0_2[405]},
      {stage0_3[288]},
      {stage0_4[6], stage0_4[7], stage0_4[8], stage0_4[9], stage0_4[10], stage0_4[11]},
      {stage1_6[1],stage1_5[40],stage1_4[141],stage1_3[141],stage1_2[141]}
   );
   gpc615_5 gpc142 (
      {stage0_2[406], stage0_2[407], stage0_2[408], stage0_2[409], stage0_2[410]},
      {stage0_3[289]},
      {stage0_4[12], stage0_4[13], stage0_4[14], stage0_4[15], stage0_4[16], stage0_4[17]},
      {stage1_6[2],stage1_5[41],stage1_4[142],stage1_3[142],stage1_2[142]}
   );
   gpc615_5 gpc143 (
      {stage0_2[411], stage0_2[412], stage0_2[413], stage0_2[414], stage0_2[415]},
      {stage0_3[290]},
      {stage0_4[18], stage0_4[19], stage0_4[20], stage0_4[21], stage0_4[22], stage0_4[23]},
      {stage1_6[3],stage1_5[42],stage1_4[143],stage1_3[143],stage1_2[143]}
   );
   gpc615_5 gpc144 (
      {stage0_2[416], stage0_2[417], stage0_2[418], stage0_2[419], stage0_2[420]},
      {stage0_3[291]},
      {stage0_4[24], stage0_4[25], stage0_4[26], stage0_4[27], stage0_4[28], stage0_4[29]},
      {stage1_6[4],stage1_5[43],stage1_4[144],stage1_3[144],stage1_2[144]}
   );
   gpc615_5 gpc145 (
      {stage0_2[421], stage0_2[422], stage0_2[423], stage0_2[424], stage0_2[425]},
      {stage0_3[292]},
      {stage0_4[30], stage0_4[31], stage0_4[32], stage0_4[33], stage0_4[34], stage0_4[35]},
      {stage1_6[5],stage1_5[44],stage1_4[145],stage1_3[145],stage1_2[145]}
   );
   gpc615_5 gpc146 (
      {stage0_2[426], stage0_2[427], stage0_2[428], stage0_2[429], stage0_2[430]},
      {stage0_3[293]},
      {stage0_4[36], stage0_4[37], stage0_4[38], stage0_4[39], stage0_4[40], stage0_4[41]},
      {stage1_6[6],stage1_5[45],stage1_4[146],stage1_3[146],stage1_2[146]}
   );
   gpc615_5 gpc147 (
      {stage0_2[431], stage0_2[432], stage0_2[433], stage0_2[434], stage0_2[435]},
      {stage0_3[294]},
      {stage0_4[42], stage0_4[43], stage0_4[44], stage0_4[45], stage0_4[46], stage0_4[47]},
      {stage1_6[7],stage1_5[46],stage1_4[147],stage1_3[147],stage1_2[147]}
   );
   gpc615_5 gpc148 (
      {stage0_2[436], stage0_2[437], stage0_2[438], stage0_2[439], stage0_2[440]},
      {stage0_3[295]},
      {stage0_4[48], stage0_4[49], stage0_4[50], stage0_4[51], stage0_4[52], stage0_4[53]},
      {stage1_6[8],stage1_5[47],stage1_4[148],stage1_3[148],stage1_2[148]}
   );
   gpc615_5 gpc149 (
      {stage0_2[441], stage0_2[442], stage0_2[443], stage0_2[444], stage0_2[445]},
      {stage0_3[296]},
      {stage0_4[54], stage0_4[55], stage0_4[56], stage0_4[57], stage0_4[58], stage0_4[59]},
      {stage1_6[9],stage1_5[48],stage1_4[149],stage1_3[149],stage1_2[149]}
   );
   gpc615_5 gpc150 (
      {stage0_2[446], stage0_2[447], stage0_2[448], stage0_2[449], stage0_2[450]},
      {stage0_3[297]},
      {stage0_4[60], stage0_4[61], stage0_4[62], stage0_4[63], stage0_4[64], stage0_4[65]},
      {stage1_6[10],stage1_5[49],stage1_4[150],stage1_3[150],stage1_2[150]}
   );
   gpc615_5 gpc151 (
      {stage0_2[451], stage0_2[452], stage0_2[453], stage0_2[454], stage0_2[455]},
      {stage0_3[298]},
      {stage0_4[66], stage0_4[67], stage0_4[68], stage0_4[69], stage0_4[70], stage0_4[71]},
      {stage1_6[11],stage1_5[50],stage1_4[151],stage1_3[151],stage1_2[151]}
   );
   gpc615_5 gpc152 (
      {stage0_2[456], stage0_2[457], stage0_2[458], stage0_2[459], stage0_2[460]},
      {stage0_3[299]},
      {stage0_4[72], stage0_4[73], stage0_4[74], stage0_4[75], stage0_4[76], stage0_4[77]},
      {stage1_6[12],stage1_5[51],stage1_4[152],stage1_3[152],stage1_2[152]}
   );
   gpc615_5 gpc153 (
      {stage0_2[461], stage0_2[462], stage0_2[463], stage0_2[464], stage0_2[465]},
      {stage0_3[300]},
      {stage0_4[78], stage0_4[79], stage0_4[80], stage0_4[81], stage0_4[82], stage0_4[83]},
      {stage1_6[13],stage1_5[52],stage1_4[153],stage1_3[153],stage1_2[153]}
   );
   gpc615_5 gpc154 (
      {stage0_2[466], stage0_2[467], stage0_2[468], stage0_2[469], stage0_2[470]},
      {stage0_3[301]},
      {stage0_4[84], stage0_4[85], stage0_4[86], stage0_4[87], stage0_4[88], stage0_4[89]},
      {stage1_6[14],stage1_5[53],stage1_4[154],stage1_3[154],stage1_2[154]}
   );
   gpc615_5 gpc155 (
      {stage0_2[471], stage0_2[472], stage0_2[473], stage0_2[474], stage0_2[475]},
      {stage0_3[302]},
      {stage0_4[90], stage0_4[91], stage0_4[92], stage0_4[93], stage0_4[94], stage0_4[95]},
      {stage1_6[15],stage1_5[54],stage1_4[155],stage1_3[155],stage1_2[155]}
   );
   gpc615_5 gpc156 (
      {stage0_2[476], stage0_2[477], stage0_2[478], stage0_2[479], stage0_2[480]},
      {stage0_3[303]},
      {stage0_4[96], stage0_4[97], stage0_4[98], stage0_4[99], stage0_4[100], stage0_4[101]},
      {stage1_6[16],stage1_5[55],stage1_4[156],stage1_3[156],stage1_2[156]}
   );
   gpc615_5 gpc157 (
      {stage0_3[304], stage0_3[305], stage0_3[306], stage0_3[307], stage0_3[308]},
      {stage0_4[102]},
      {stage0_5[0], stage0_5[1], stage0_5[2], stage0_5[3], stage0_5[4], stage0_5[5]},
      {stage1_7[0],stage1_6[17],stage1_5[56],stage1_4[157],stage1_3[157]}
   );
   gpc615_5 gpc158 (
      {stage0_3[309], stage0_3[310], stage0_3[311], stage0_3[312], stage0_3[313]},
      {stage0_4[103]},
      {stage0_5[6], stage0_5[7], stage0_5[8], stage0_5[9], stage0_5[10], stage0_5[11]},
      {stage1_7[1],stage1_6[18],stage1_5[57],stage1_4[158],stage1_3[158]}
   );
   gpc615_5 gpc159 (
      {stage0_3[314], stage0_3[315], stage0_3[316], stage0_3[317], stage0_3[318]},
      {stage0_4[104]},
      {stage0_5[12], stage0_5[13], stage0_5[14], stage0_5[15], stage0_5[16], stage0_5[17]},
      {stage1_7[2],stage1_6[19],stage1_5[58],stage1_4[159],stage1_3[159]}
   );
   gpc615_5 gpc160 (
      {stage0_3[319], stage0_3[320], stage0_3[321], stage0_3[322], stage0_3[323]},
      {stage0_4[105]},
      {stage0_5[18], stage0_5[19], stage0_5[20], stage0_5[21], stage0_5[22], stage0_5[23]},
      {stage1_7[3],stage1_6[20],stage1_5[59],stage1_4[160],stage1_3[160]}
   );
   gpc615_5 gpc161 (
      {stage0_3[324], stage0_3[325], stage0_3[326], stage0_3[327], stage0_3[328]},
      {stage0_4[106]},
      {stage0_5[24], stage0_5[25], stage0_5[26], stage0_5[27], stage0_5[28], stage0_5[29]},
      {stage1_7[4],stage1_6[21],stage1_5[60],stage1_4[161],stage1_3[161]}
   );
   gpc615_5 gpc162 (
      {stage0_3[329], stage0_3[330], stage0_3[331], stage0_3[332], stage0_3[333]},
      {stage0_4[107]},
      {stage0_5[30], stage0_5[31], stage0_5[32], stage0_5[33], stage0_5[34], stage0_5[35]},
      {stage1_7[5],stage1_6[22],stage1_5[61],stage1_4[162],stage1_3[162]}
   );
   gpc615_5 gpc163 (
      {stage0_3[334], stage0_3[335], stage0_3[336], stage0_3[337], stage0_3[338]},
      {stage0_4[108]},
      {stage0_5[36], stage0_5[37], stage0_5[38], stage0_5[39], stage0_5[40], stage0_5[41]},
      {stage1_7[6],stage1_6[23],stage1_5[62],stage1_4[163],stage1_3[163]}
   );
   gpc615_5 gpc164 (
      {stage0_3[339], stage0_3[340], stage0_3[341], stage0_3[342], stage0_3[343]},
      {stage0_4[109]},
      {stage0_5[42], stage0_5[43], stage0_5[44], stage0_5[45], stage0_5[46], stage0_5[47]},
      {stage1_7[7],stage1_6[24],stage1_5[63],stage1_4[164],stage1_3[164]}
   );
   gpc615_5 gpc165 (
      {stage0_3[344], stage0_3[345], stage0_3[346], stage0_3[347], stage0_3[348]},
      {stage0_4[110]},
      {stage0_5[48], stage0_5[49], stage0_5[50], stage0_5[51], stage0_5[52], stage0_5[53]},
      {stage1_7[8],stage1_6[25],stage1_5[64],stage1_4[165],stage1_3[165]}
   );
   gpc615_5 gpc166 (
      {stage0_3[349], stage0_3[350], stage0_3[351], stage0_3[352], stage0_3[353]},
      {stage0_4[111]},
      {stage0_5[54], stage0_5[55], stage0_5[56], stage0_5[57], stage0_5[58], stage0_5[59]},
      {stage1_7[9],stage1_6[26],stage1_5[65],stage1_4[166],stage1_3[166]}
   );
   gpc615_5 gpc167 (
      {stage0_3[354], stage0_3[355], stage0_3[356], stage0_3[357], stage0_3[358]},
      {stage0_4[112]},
      {stage0_5[60], stage0_5[61], stage0_5[62], stage0_5[63], stage0_5[64], stage0_5[65]},
      {stage1_7[10],stage1_6[27],stage1_5[66],stage1_4[167],stage1_3[167]}
   );
   gpc615_5 gpc168 (
      {stage0_3[359], stage0_3[360], stage0_3[361], stage0_3[362], stage0_3[363]},
      {stage0_4[113]},
      {stage0_5[66], stage0_5[67], stage0_5[68], stage0_5[69], stage0_5[70], stage0_5[71]},
      {stage1_7[11],stage1_6[28],stage1_5[67],stage1_4[168],stage1_3[168]}
   );
   gpc615_5 gpc169 (
      {stage0_3[364], stage0_3[365], stage0_3[366], stage0_3[367], stage0_3[368]},
      {stage0_4[114]},
      {stage0_5[72], stage0_5[73], stage0_5[74], stage0_5[75], stage0_5[76], stage0_5[77]},
      {stage1_7[12],stage1_6[29],stage1_5[68],stage1_4[169],stage1_3[169]}
   );
   gpc615_5 gpc170 (
      {stage0_3[369], stage0_3[370], stage0_3[371], stage0_3[372], stage0_3[373]},
      {stage0_4[115]},
      {stage0_5[78], stage0_5[79], stage0_5[80], stage0_5[81], stage0_5[82], stage0_5[83]},
      {stage1_7[13],stage1_6[30],stage1_5[69],stage1_4[170],stage1_3[170]}
   );
   gpc615_5 gpc171 (
      {stage0_3[374], stage0_3[375], stage0_3[376], stage0_3[377], stage0_3[378]},
      {stage0_4[116]},
      {stage0_5[84], stage0_5[85], stage0_5[86], stage0_5[87], stage0_5[88], stage0_5[89]},
      {stage1_7[14],stage1_6[31],stage1_5[70],stage1_4[171],stage1_3[171]}
   );
   gpc615_5 gpc172 (
      {stage0_3[379], stage0_3[380], stage0_3[381], stage0_3[382], stage0_3[383]},
      {stage0_4[117]},
      {stage0_5[90], stage0_5[91], stage0_5[92], stage0_5[93], stage0_5[94], stage0_5[95]},
      {stage1_7[15],stage1_6[32],stage1_5[71],stage1_4[172],stage1_3[172]}
   );
   gpc615_5 gpc173 (
      {stage0_3[384], stage0_3[385], stage0_3[386], stage0_3[387], stage0_3[388]},
      {stage0_4[118]},
      {stage0_5[96], stage0_5[97], stage0_5[98], stage0_5[99], stage0_5[100], stage0_5[101]},
      {stage1_7[16],stage1_6[33],stage1_5[72],stage1_4[173],stage1_3[173]}
   );
   gpc615_5 gpc174 (
      {stage0_3[389], stage0_3[390], stage0_3[391], stage0_3[392], stage0_3[393]},
      {stage0_4[119]},
      {stage0_5[102], stage0_5[103], stage0_5[104], stage0_5[105], stage0_5[106], stage0_5[107]},
      {stage1_7[17],stage1_6[34],stage1_5[73],stage1_4[174],stage1_3[174]}
   );
   gpc615_5 gpc175 (
      {stage0_3[394], stage0_3[395], stage0_3[396], stage0_3[397], stage0_3[398]},
      {stage0_4[120]},
      {stage0_5[108], stage0_5[109], stage0_5[110], stage0_5[111], stage0_5[112], stage0_5[113]},
      {stage1_7[18],stage1_6[35],stage1_5[74],stage1_4[175],stage1_3[175]}
   );
   gpc615_5 gpc176 (
      {stage0_3[399], stage0_3[400], stage0_3[401], stage0_3[402], stage0_3[403]},
      {stage0_4[121]},
      {stage0_5[114], stage0_5[115], stage0_5[116], stage0_5[117], stage0_5[118], stage0_5[119]},
      {stage1_7[19],stage1_6[36],stage1_5[75],stage1_4[176],stage1_3[176]}
   );
   gpc615_5 gpc177 (
      {stage0_3[404], stage0_3[405], stage0_3[406], stage0_3[407], stage0_3[408]},
      {stage0_4[122]},
      {stage0_5[120], stage0_5[121], stage0_5[122], stage0_5[123], stage0_5[124], stage0_5[125]},
      {stage1_7[20],stage1_6[37],stage1_5[76],stage1_4[177],stage1_3[177]}
   );
   gpc615_5 gpc178 (
      {stage0_3[409], stage0_3[410], stage0_3[411], stage0_3[412], stage0_3[413]},
      {stage0_4[123]},
      {stage0_5[126], stage0_5[127], stage0_5[128], stage0_5[129], stage0_5[130], stage0_5[131]},
      {stage1_7[21],stage1_6[38],stage1_5[77],stage1_4[178],stage1_3[178]}
   );
   gpc606_5 gpc179 (
      {stage0_4[124], stage0_4[125], stage0_4[126], stage0_4[127], stage0_4[128], stage0_4[129]},
      {stage0_6[0], stage0_6[1], stage0_6[2], stage0_6[3], stage0_6[4], stage0_6[5]},
      {stage1_8[0],stage1_7[22],stage1_6[39],stage1_5[78],stage1_4[179]}
   );
   gpc606_5 gpc180 (
      {stage0_4[130], stage0_4[131], stage0_4[132], stage0_4[133], stage0_4[134], stage0_4[135]},
      {stage0_6[6], stage0_6[7], stage0_6[8], stage0_6[9], stage0_6[10], stage0_6[11]},
      {stage1_8[1],stage1_7[23],stage1_6[40],stage1_5[79],stage1_4[180]}
   );
   gpc606_5 gpc181 (
      {stage0_4[136], stage0_4[137], stage0_4[138], stage0_4[139], stage0_4[140], stage0_4[141]},
      {stage0_6[12], stage0_6[13], stage0_6[14], stage0_6[15], stage0_6[16], stage0_6[17]},
      {stage1_8[2],stage1_7[24],stage1_6[41],stage1_5[80],stage1_4[181]}
   );
   gpc606_5 gpc182 (
      {stage0_4[142], stage0_4[143], stage0_4[144], stage0_4[145], stage0_4[146], stage0_4[147]},
      {stage0_6[18], stage0_6[19], stage0_6[20], stage0_6[21], stage0_6[22], stage0_6[23]},
      {stage1_8[3],stage1_7[25],stage1_6[42],stage1_5[81],stage1_4[182]}
   );
   gpc606_5 gpc183 (
      {stage0_4[148], stage0_4[149], stage0_4[150], stage0_4[151], stage0_4[152], stage0_4[153]},
      {stage0_6[24], stage0_6[25], stage0_6[26], stage0_6[27], stage0_6[28], stage0_6[29]},
      {stage1_8[4],stage1_7[26],stage1_6[43],stage1_5[82],stage1_4[183]}
   );
   gpc606_5 gpc184 (
      {stage0_4[154], stage0_4[155], stage0_4[156], stage0_4[157], stage0_4[158], stage0_4[159]},
      {stage0_6[30], stage0_6[31], stage0_6[32], stage0_6[33], stage0_6[34], stage0_6[35]},
      {stage1_8[5],stage1_7[27],stage1_6[44],stage1_5[83],stage1_4[184]}
   );
   gpc606_5 gpc185 (
      {stage0_4[160], stage0_4[161], stage0_4[162], stage0_4[163], stage0_4[164], stage0_4[165]},
      {stage0_6[36], stage0_6[37], stage0_6[38], stage0_6[39], stage0_6[40], stage0_6[41]},
      {stage1_8[6],stage1_7[28],stage1_6[45],stage1_5[84],stage1_4[185]}
   );
   gpc606_5 gpc186 (
      {stage0_4[166], stage0_4[167], stage0_4[168], stage0_4[169], stage0_4[170], stage0_4[171]},
      {stage0_6[42], stage0_6[43], stage0_6[44], stage0_6[45], stage0_6[46], stage0_6[47]},
      {stage1_8[7],stage1_7[29],stage1_6[46],stage1_5[85],stage1_4[186]}
   );
   gpc606_5 gpc187 (
      {stage0_4[172], stage0_4[173], stage0_4[174], stage0_4[175], stage0_4[176], stage0_4[177]},
      {stage0_6[48], stage0_6[49], stage0_6[50], stage0_6[51], stage0_6[52], stage0_6[53]},
      {stage1_8[8],stage1_7[30],stage1_6[47],stage1_5[86],stage1_4[187]}
   );
   gpc606_5 gpc188 (
      {stage0_4[178], stage0_4[179], stage0_4[180], stage0_4[181], stage0_4[182], stage0_4[183]},
      {stage0_6[54], stage0_6[55], stage0_6[56], stage0_6[57], stage0_6[58], stage0_6[59]},
      {stage1_8[9],stage1_7[31],stage1_6[48],stage1_5[87],stage1_4[188]}
   );
   gpc606_5 gpc189 (
      {stage0_4[184], stage0_4[185], stage0_4[186], stage0_4[187], stage0_4[188], stage0_4[189]},
      {stage0_6[60], stage0_6[61], stage0_6[62], stage0_6[63], stage0_6[64], stage0_6[65]},
      {stage1_8[10],stage1_7[32],stage1_6[49],stage1_5[88],stage1_4[189]}
   );
   gpc606_5 gpc190 (
      {stage0_4[190], stage0_4[191], stage0_4[192], stage0_4[193], stage0_4[194], stage0_4[195]},
      {stage0_6[66], stage0_6[67], stage0_6[68], stage0_6[69], stage0_6[70], stage0_6[71]},
      {stage1_8[11],stage1_7[33],stage1_6[50],stage1_5[89],stage1_4[190]}
   );
   gpc606_5 gpc191 (
      {stage0_4[196], stage0_4[197], stage0_4[198], stage0_4[199], stage0_4[200], stage0_4[201]},
      {stage0_6[72], stage0_6[73], stage0_6[74], stage0_6[75], stage0_6[76], stage0_6[77]},
      {stage1_8[12],stage1_7[34],stage1_6[51],stage1_5[90],stage1_4[191]}
   );
   gpc606_5 gpc192 (
      {stage0_4[202], stage0_4[203], stage0_4[204], stage0_4[205], stage0_4[206], stage0_4[207]},
      {stage0_6[78], stage0_6[79], stage0_6[80], stage0_6[81], stage0_6[82], stage0_6[83]},
      {stage1_8[13],stage1_7[35],stage1_6[52],stage1_5[91],stage1_4[192]}
   );
   gpc606_5 gpc193 (
      {stage0_4[208], stage0_4[209], stage0_4[210], stage0_4[211], stage0_4[212], stage0_4[213]},
      {stage0_6[84], stage0_6[85], stage0_6[86], stage0_6[87], stage0_6[88], stage0_6[89]},
      {stage1_8[14],stage1_7[36],stage1_6[53],stage1_5[92],stage1_4[193]}
   );
   gpc606_5 gpc194 (
      {stage0_4[214], stage0_4[215], stage0_4[216], stage0_4[217], stage0_4[218], stage0_4[219]},
      {stage0_6[90], stage0_6[91], stage0_6[92], stage0_6[93], stage0_6[94], stage0_6[95]},
      {stage1_8[15],stage1_7[37],stage1_6[54],stage1_5[93],stage1_4[194]}
   );
   gpc606_5 gpc195 (
      {stage0_4[220], stage0_4[221], stage0_4[222], stage0_4[223], stage0_4[224], stage0_4[225]},
      {stage0_6[96], stage0_6[97], stage0_6[98], stage0_6[99], stage0_6[100], stage0_6[101]},
      {stage1_8[16],stage1_7[38],stage1_6[55],stage1_5[94],stage1_4[195]}
   );
   gpc606_5 gpc196 (
      {stage0_4[226], stage0_4[227], stage0_4[228], stage0_4[229], stage0_4[230], stage0_4[231]},
      {stage0_6[102], stage0_6[103], stage0_6[104], stage0_6[105], stage0_6[106], stage0_6[107]},
      {stage1_8[17],stage1_7[39],stage1_6[56],stage1_5[95],stage1_4[196]}
   );
   gpc606_5 gpc197 (
      {stage0_4[232], stage0_4[233], stage0_4[234], stage0_4[235], stage0_4[236], stage0_4[237]},
      {stage0_6[108], stage0_6[109], stage0_6[110], stage0_6[111], stage0_6[112], stage0_6[113]},
      {stage1_8[18],stage1_7[40],stage1_6[57],stage1_5[96],stage1_4[197]}
   );
   gpc606_5 gpc198 (
      {stage0_4[238], stage0_4[239], stage0_4[240], stage0_4[241], stage0_4[242], stage0_4[243]},
      {stage0_6[114], stage0_6[115], stage0_6[116], stage0_6[117], stage0_6[118], stage0_6[119]},
      {stage1_8[19],stage1_7[41],stage1_6[58],stage1_5[97],stage1_4[198]}
   );
   gpc606_5 gpc199 (
      {stage0_4[244], stage0_4[245], stage0_4[246], stage0_4[247], stage0_4[248], stage0_4[249]},
      {stage0_6[120], stage0_6[121], stage0_6[122], stage0_6[123], stage0_6[124], stage0_6[125]},
      {stage1_8[20],stage1_7[42],stage1_6[59],stage1_5[98],stage1_4[199]}
   );
   gpc606_5 gpc200 (
      {stage0_4[250], stage0_4[251], stage0_4[252], stage0_4[253], stage0_4[254], stage0_4[255]},
      {stage0_6[126], stage0_6[127], stage0_6[128], stage0_6[129], stage0_6[130], stage0_6[131]},
      {stage1_8[21],stage1_7[43],stage1_6[60],stage1_5[99],stage1_4[200]}
   );
   gpc606_5 gpc201 (
      {stage0_4[256], stage0_4[257], stage0_4[258], stage0_4[259], stage0_4[260], stage0_4[261]},
      {stage0_6[132], stage0_6[133], stage0_6[134], stage0_6[135], stage0_6[136], stage0_6[137]},
      {stage1_8[22],stage1_7[44],stage1_6[61],stage1_5[100],stage1_4[201]}
   );
   gpc606_5 gpc202 (
      {stage0_4[262], stage0_4[263], stage0_4[264], stage0_4[265], stage0_4[266], stage0_4[267]},
      {stage0_6[138], stage0_6[139], stage0_6[140], stage0_6[141], stage0_6[142], stage0_6[143]},
      {stage1_8[23],stage1_7[45],stage1_6[62],stage1_5[101],stage1_4[202]}
   );
   gpc606_5 gpc203 (
      {stage0_4[268], stage0_4[269], stage0_4[270], stage0_4[271], stage0_4[272], stage0_4[273]},
      {stage0_6[144], stage0_6[145], stage0_6[146], stage0_6[147], stage0_6[148], stage0_6[149]},
      {stage1_8[24],stage1_7[46],stage1_6[63],stage1_5[102],stage1_4[203]}
   );
   gpc606_5 gpc204 (
      {stage0_4[274], stage0_4[275], stage0_4[276], stage0_4[277], stage0_4[278], stage0_4[279]},
      {stage0_6[150], stage0_6[151], stage0_6[152], stage0_6[153], stage0_6[154], stage0_6[155]},
      {stage1_8[25],stage1_7[47],stage1_6[64],stage1_5[103],stage1_4[204]}
   );
   gpc606_5 gpc205 (
      {stage0_4[280], stage0_4[281], stage0_4[282], stage0_4[283], stage0_4[284], stage0_4[285]},
      {stage0_6[156], stage0_6[157], stage0_6[158], stage0_6[159], stage0_6[160], stage0_6[161]},
      {stage1_8[26],stage1_7[48],stage1_6[65],stage1_5[104],stage1_4[205]}
   );
   gpc606_5 gpc206 (
      {stage0_4[286], stage0_4[287], stage0_4[288], stage0_4[289], stage0_4[290], stage0_4[291]},
      {stage0_6[162], stage0_6[163], stage0_6[164], stage0_6[165], stage0_6[166], stage0_6[167]},
      {stage1_8[27],stage1_7[49],stage1_6[66],stage1_5[105],stage1_4[206]}
   );
   gpc606_5 gpc207 (
      {stage0_4[292], stage0_4[293], stage0_4[294], stage0_4[295], stage0_4[296], stage0_4[297]},
      {stage0_6[168], stage0_6[169], stage0_6[170], stage0_6[171], stage0_6[172], stage0_6[173]},
      {stage1_8[28],stage1_7[50],stage1_6[67],stage1_5[106],stage1_4[207]}
   );
   gpc606_5 gpc208 (
      {stage0_4[298], stage0_4[299], stage0_4[300], stage0_4[301], stage0_4[302], stage0_4[303]},
      {stage0_6[174], stage0_6[175], stage0_6[176], stage0_6[177], stage0_6[178], stage0_6[179]},
      {stage1_8[29],stage1_7[51],stage1_6[68],stage1_5[107],stage1_4[208]}
   );
   gpc606_5 gpc209 (
      {stage0_4[304], stage0_4[305], stage0_4[306], stage0_4[307], stage0_4[308], stage0_4[309]},
      {stage0_6[180], stage0_6[181], stage0_6[182], stage0_6[183], stage0_6[184], stage0_6[185]},
      {stage1_8[30],stage1_7[52],stage1_6[69],stage1_5[108],stage1_4[209]}
   );
   gpc606_5 gpc210 (
      {stage0_4[310], stage0_4[311], stage0_4[312], stage0_4[313], stage0_4[314], stage0_4[315]},
      {stage0_6[186], stage0_6[187], stage0_6[188], stage0_6[189], stage0_6[190], stage0_6[191]},
      {stage1_8[31],stage1_7[53],stage1_6[70],stage1_5[109],stage1_4[210]}
   );
   gpc606_5 gpc211 (
      {stage0_4[316], stage0_4[317], stage0_4[318], stage0_4[319], stage0_4[320], stage0_4[321]},
      {stage0_6[192], stage0_6[193], stage0_6[194], stage0_6[195], stage0_6[196], stage0_6[197]},
      {stage1_8[32],stage1_7[54],stage1_6[71],stage1_5[110],stage1_4[211]}
   );
   gpc606_5 gpc212 (
      {stage0_4[322], stage0_4[323], stage0_4[324], stage0_4[325], stage0_4[326], stage0_4[327]},
      {stage0_6[198], stage0_6[199], stage0_6[200], stage0_6[201], stage0_6[202], stage0_6[203]},
      {stage1_8[33],stage1_7[55],stage1_6[72],stage1_5[111],stage1_4[212]}
   );
   gpc606_5 gpc213 (
      {stage0_4[328], stage0_4[329], stage0_4[330], stage0_4[331], stage0_4[332], stage0_4[333]},
      {stage0_6[204], stage0_6[205], stage0_6[206], stage0_6[207], stage0_6[208], stage0_6[209]},
      {stage1_8[34],stage1_7[56],stage1_6[73],stage1_5[112],stage1_4[213]}
   );
   gpc606_5 gpc214 (
      {stage0_4[334], stage0_4[335], stage0_4[336], stage0_4[337], stage0_4[338], stage0_4[339]},
      {stage0_6[210], stage0_6[211], stage0_6[212], stage0_6[213], stage0_6[214], stage0_6[215]},
      {stage1_8[35],stage1_7[57],stage1_6[74],stage1_5[113],stage1_4[214]}
   );
   gpc606_5 gpc215 (
      {stage0_4[340], stage0_4[341], stage0_4[342], stage0_4[343], stage0_4[344], stage0_4[345]},
      {stage0_6[216], stage0_6[217], stage0_6[218], stage0_6[219], stage0_6[220], stage0_6[221]},
      {stage1_8[36],stage1_7[58],stage1_6[75],stage1_5[114],stage1_4[215]}
   );
   gpc606_5 gpc216 (
      {stage0_4[346], stage0_4[347], stage0_4[348], stage0_4[349], stage0_4[350], stage0_4[351]},
      {stage0_6[222], stage0_6[223], stage0_6[224], stage0_6[225], stage0_6[226], stage0_6[227]},
      {stage1_8[37],stage1_7[59],stage1_6[76],stage1_5[115],stage1_4[216]}
   );
   gpc606_5 gpc217 (
      {stage0_4[352], stage0_4[353], stage0_4[354], stage0_4[355], stage0_4[356], stage0_4[357]},
      {stage0_6[228], stage0_6[229], stage0_6[230], stage0_6[231], stage0_6[232], stage0_6[233]},
      {stage1_8[38],stage1_7[60],stage1_6[77],stage1_5[116],stage1_4[217]}
   );
   gpc606_5 gpc218 (
      {stage0_4[358], stage0_4[359], stage0_4[360], stage0_4[361], stage0_4[362], stage0_4[363]},
      {stage0_6[234], stage0_6[235], stage0_6[236], stage0_6[237], stage0_6[238], stage0_6[239]},
      {stage1_8[39],stage1_7[61],stage1_6[78],stage1_5[117],stage1_4[218]}
   );
   gpc606_5 gpc219 (
      {stage0_4[364], stage0_4[365], stage0_4[366], stage0_4[367], stage0_4[368], stage0_4[369]},
      {stage0_6[240], stage0_6[241], stage0_6[242], stage0_6[243], stage0_6[244], stage0_6[245]},
      {stage1_8[40],stage1_7[62],stage1_6[79],stage1_5[118],stage1_4[219]}
   );
   gpc606_5 gpc220 (
      {stage0_4[370], stage0_4[371], stage0_4[372], stage0_4[373], stage0_4[374], stage0_4[375]},
      {stage0_6[246], stage0_6[247], stage0_6[248], stage0_6[249], stage0_6[250], stage0_6[251]},
      {stage1_8[41],stage1_7[63],stage1_6[80],stage1_5[119],stage1_4[220]}
   );
   gpc606_5 gpc221 (
      {stage0_4[376], stage0_4[377], stage0_4[378], stage0_4[379], stage0_4[380], stage0_4[381]},
      {stage0_6[252], stage0_6[253], stage0_6[254], stage0_6[255], stage0_6[256], stage0_6[257]},
      {stage1_8[42],stage1_7[64],stage1_6[81],stage1_5[120],stage1_4[221]}
   );
   gpc606_5 gpc222 (
      {stage0_4[382], stage0_4[383], stage0_4[384], stage0_4[385], stage0_4[386], stage0_4[387]},
      {stage0_6[258], stage0_6[259], stage0_6[260], stage0_6[261], stage0_6[262], stage0_6[263]},
      {stage1_8[43],stage1_7[65],stage1_6[82],stage1_5[121],stage1_4[222]}
   );
   gpc606_5 gpc223 (
      {stage0_4[388], stage0_4[389], stage0_4[390], stage0_4[391], stage0_4[392], stage0_4[393]},
      {stage0_6[264], stage0_6[265], stage0_6[266], stage0_6[267], stage0_6[268], stage0_6[269]},
      {stage1_8[44],stage1_7[66],stage1_6[83],stage1_5[122],stage1_4[223]}
   );
   gpc606_5 gpc224 (
      {stage0_4[394], stage0_4[395], stage0_4[396], stage0_4[397], stage0_4[398], stage0_4[399]},
      {stage0_6[270], stage0_6[271], stage0_6[272], stage0_6[273], stage0_6[274], stage0_6[275]},
      {stage1_8[45],stage1_7[67],stage1_6[84],stage1_5[123],stage1_4[224]}
   );
   gpc606_5 gpc225 (
      {stage0_4[400], stage0_4[401], stage0_4[402], stage0_4[403], stage0_4[404], stage0_4[405]},
      {stage0_6[276], stage0_6[277], stage0_6[278], stage0_6[279], stage0_6[280], stage0_6[281]},
      {stage1_8[46],stage1_7[68],stage1_6[85],stage1_5[124],stage1_4[225]}
   );
   gpc606_5 gpc226 (
      {stage0_4[406], stage0_4[407], stage0_4[408], stage0_4[409], stage0_4[410], stage0_4[411]},
      {stage0_6[282], stage0_6[283], stage0_6[284], stage0_6[285], stage0_6[286], stage0_6[287]},
      {stage1_8[47],stage1_7[69],stage1_6[86],stage1_5[125],stage1_4[226]}
   );
   gpc606_5 gpc227 (
      {stage0_4[412], stage0_4[413], stage0_4[414], stage0_4[415], stage0_4[416], stage0_4[417]},
      {stage0_6[288], stage0_6[289], stage0_6[290], stage0_6[291], stage0_6[292], stage0_6[293]},
      {stage1_8[48],stage1_7[70],stage1_6[87],stage1_5[126],stage1_4[227]}
   );
   gpc606_5 gpc228 (
      {stage0_4[418], stage0_4[419], stage0_4[420], stage0_4[421], stage0_4[422], stage0_4[423]},
      {stage0_6[294], stage0_6[295], stage0_6[296], stage0_6[297], stage0_6[298], stage0_6[299]},
      {stage1_8[49],stage1_7[71],stage1_6[88],stage1_5[127],stage1_4[228]}
   );
   gpc606_5 gpc229 (
      {stage0_4[424], stage0_4[425], stage0_4[426], stage0_4[427], stage0_4[428], stage0_4[429]},
      {stage0_6[300], stage0_6[301], stage0_6[302], stage0_6[303], stage0_6[304], stage0_6[305]},
      {stage1_8[50],stage1_7[72],stage1_6[89],stage1_5[128],stage1_4[229]}
   );
   gpc606_5 gpc230 (
      {stage0_4[430], stage0_4[431], stage0_4[432], stage0_4[433], stage0_4[434], stage0_4[435]},
      {stage0_6[306], stage0_6[307], stage0_6[308], stage0_6[309], stage0_6[310], stage0_6[311]},
      {stage1_8[51],stage1_7[73],stage1_6[90],stage1_5[129],stage1_4[230]}
   );
   gpc606_5 gpc231 (
      {stage0_4[436], stage0_4[437], stage0_4[438], stage0_4[439], stage0_4[440], stage0_4[441]},
      {stage0_6[312], stage0_6[313], stage0_6[314], stage0_6[315], stage0_6[316], stage0_6[317]},
      {stage1_8[52],stage1_7[74],stage1_6[91],stage1_5[130],stage1_4[231]}
   );
   gpc606_5 gpc232 (
      {stage0_4[442], stage0_4[443], stage0_4[444], stage0_4[445], stage0_4[446], stage0_4[447]},
      {stage0_6[318], stage0_6[319], stage0_6[320], stage0_6[321], stage0_6[322], stage0_6[323]},
      {stage1_8[53],stage1_7[75],stage1_6[92],stage1_5[131],stage1_4[232]}
   );
   gpc606_5 gpc233 (
      {stage0_4[448], stage0_4[449], stage0_4[450], stage0_4[451], stage0_4[452], stage0_4[453]},
      {stage0_6[324], stage0_6[325], stage0_6[326], stage0_6[327], stage0_6[328], stage0_6[329]},
      {stage1_8[54],stage1_7[76],stage1_6[93],stage1_5[132],stage1_4[233]}
   );
   gpc606_5 gpc234 (
      {stage0_4[454], stage0_4[455], stage0_4[456], stage0_4[457], stage0_4[458], stage0_4[459]},
      {stage0_6[330], stage0_6[331], stage0_6[332], stage0_6[333], stage0_6[334], stage0_6[335]},
      {stage1_8[55],stage1_7[77],stage1_6[94],stage1_5[133],stage1_4[234]}
   );
   gpc606_5 gpc235 (
      {stage0_4[460], stage0_4[461], stage0_4[462], stage0_4[463], stage0_4[464], stage0_4[465]},
      {stage0_6[336], stage0_6[337], stage0_6[338], stage0_6[339], stage0_6[340], stage0_6[341]},
      {stage1_8[56],stage1_7[78],stage1_6[95],stage1_5[134],stage1_4[235]}
   );
   gpc606_5 gpc236 (
      {stage0_4[466], stage0_4[467], stage0_4[468], stage0_4[469], stage0_4[470], stage0_4[471]},
      {stage0_6[342], stage0_6[343], stage0_6[344], stage0_6[345], stage0_6[346], stage0_6[347]},
      {stage1_8[57],stage1_7[79],stage1_6[96],stage1_5[135],stage1_4[236]}
   );
   gpc615_5 gpc237 (
      {stage0_4[472], stage0_4[473], stage0_4[474], stage0_4[475], stage0_4[476]},
      {stage0_5[132]},
      {stage0_6[348], stage0_6[349], stage0_6[350], stage0_6[351], stage0_6[352], stage0_6[353]},
      {stage1_8[58],stage1_7[80],stage1_6[97],stage1_5[136],stage1_4[237]}
   );
   gpc615_5 gpc238 (
      {stage0_4[477], stage0_4[478], stage0_4[479], stage0_4[480], stage0_4[481]},
      {stage0_5[133]},
      {stage0_6[354], stage0_6[355], stage0_6[356], stage0_6[357], stage0_6[358], stage0_6[359]},
      {stage1_8[59],stage1_7[81],stage1_6[98],stage1_5[137],stage1_4[238]}
   );
   gpc615_5 gpc239 (
      {stage0_4[482], stage0_4[483], stage0_4[484], stage0_4[485], stage0_4[486]},
      {stage0_5[134]},
      {stage0_6[360], stage0_6[361], stage0_6[362], stage0_6[363], stage0_6[364], stage0_6[365]},
      {stage1_8[60],stage1_7[82],stage1_6[99],stage1_5[138],stage1_4[239]}
   );
   gpc615_5 gpc240 (
      {stage0_4[487], stage0_4[488], stage0_4[489], stage0_4[490], stage0_4[491]},
      {stage0_5[135]},
      {stage0_6[366], stage0_6[367], stage0_6[368], stage0_6[369], stage0_6[370], stage0_6[371]},
      {stage1_8[61],stage1_7[83],stage1_6[100],stage1_5[139],stage1_4[240]}
   );
   gpc615_5 gpc241 (
      {stage0_4[492], stage0_4[493], stage0_4[494], stage0_4[495], stage0_4[496]},
      {stage0_5[136]},
      {stage0_6[372], stage0_6[373], stage0_6[374], stage0_6[375], stage0_6[376], stage0_6[377]},
      {stage1_8[62],stage1_7[84],stage1_6[101],stage1_5[140],stage1_4[241]}
   );
   gpc615_5 gpc242 (
      {stage0_4[497], stage0_4[498], stage0_4[499], stage0_4[500], stage0_4[501]},
      {stage0_5[137]},
      {stage0_6[378], stage0_6[379], stage0_6[380], stage0_6[381], stage0_6[382], stage0_6[383]},
      {stage1_8[63],stage1_7[85],stage1_6[102],stage1_5[141],stage1_4[242]}
   );
   gpc615_5 gpc243 (
      {stage0_4[502], stage0_4[503], stage0_4[504], stage0_4[505], stage0_4[506]},
      {stage0_5[138]},
      {stage0_6[384], stage0_6[385], stage0_6[386], stage0_6[387], stage0_6[388], stage0_6[389]},
      {stage1_8[64],stage1_7[86],stage1_6[103],stage1_5[142],stage1_4[243]}
   );
   gpc615_5 gpc244 (
      {stage0_4[507], stage0_4[508], stage0_4[509], stage0_4[510], stage0_4[511]},
      {stage0_5[139]},
      {stage0_6[390], stage0_6[391], stage0_6[392], stage0_6[393], stage0_6[394], stage0_6[395]},
      {stage1_8[65],stage1_7[87],stage1_6[104],stage1_5[143],stage1_4[244]}
   );
   gpc606_5 gpc245 (
      {stage0_5[140], stage0_5[141], stage0_5[142], stage0_5[143], stage0_5[144], stage0_5[145]},
      {stage0_7[0], stage0_7[1], stage0_7[2], stage0_7[3], stage0_7[4], stage0_7[5]},
      {stage1_9[0],stage1_8[66],stage1_7[88],stage1_6[105],stage1_5[144]}
   );
   gpc606_5 gpc246 (
      {stage0_5[146], stage0_5[147], stage0_5[148], stage0_5[149], stage0_5[150], stage0_5[151]},
      {stage0_7[6], stage0_7[7], stage0_7[8], stage0_7[9], stage0_7[10], stage0_7[11]},
      {stage1_9[1],stage1_8[67],stage1_7[89],stage1_6[106],stage1_5[145]}
   );
   gpc606_5 gpc247 (
      {stage0_5[152], stage0_5[153], stage0_5[154], stage0_5[155], stage0_5[156], stage0_5[157]},
      {stage0_7[12], stage0_7[13], stage0_7[14], stage0_7[15], stage0_7[16], stage0_7[17]},
      {stage1_9[2],stage1_8[68],stage1_7[90],stage1_6[107],stage1_5[146]}
   );
   gpc606_5 gpc248 (
      {stage0_5[158], stage0_5[159], stage0_5[160], stage0_5[161], stage0_5[162], stage0_5[163]},
      {stage0_7[18], stage0_7[19], stage0_7[20], stage0_7[21], stage0_7[22], stage0_7[23]},
      {stage1_9[3],stage1_8[69],stage1_7[91],stage1_6[108],stage1_5[147]}
   );
   gpc606_5 gpc249 (
      {stage0_5[164], stage0_5[165], stage0_5[166], stage0_5[167], stage0_5[168], stage0_5[169]},
      {stage0_7[24], stage0_7[25], stage0_7[26], stage0_7[27], stage0_7[28], stage0_7[29]},
      {stage1_9[4],stage1_8[70],stage1_7[92],stage1_6[109],stage1_5[148]}
   );
   gpc606_5 gpc250 (
      {stage0_5[170], stage0_5[171], stage0_5[172], stage0_5[173], stage0_5[174], stage0_5[175]},
      {stage0_7[30], stage0_7[31], stage0_7[32], stage0_7[33], stage0_7[34], stage0_7[35]},
      {stage1_9[5],stage1_8[71],stage1_7[93],stage1_6[110],stage1_5[149]}
   );
   gpc606_5 gpc251 (
      {stage0_5[176], stage0_5[177], stage0_5[178], stage0_5[179], stage0_5[180], stage0_5[181]},
      {stage0_7[36], stage0_7[37], stage0_7[38], stage0_7[39], stage0_7[40], stage0_7[41]},
      {stage1_9[6],stage1_8[72],stage1_7[94],stage1_6[111],stage1_5[150]}
   );
   gpc606_5 gpc252 (
      {stage0_5[182], stage0_5[183], stage0_5[184], stage0_5[185], stage0_5[186], stage0_5[187]},
      {stage0_7[42], stage0_7[43], stage0_7[44], stage0_7[45], stage0_7[46], stage0_7[47]},
      {stage1_9[7],stage1_8[73],stage1_7[95],stage1_6[112],stage1_5[151]}
   );
   gpc606_5 gpc253 (
      {stage0_5[188], stage0_5[189], stage0_5[190], stage0_5[191], stage0_5[192], stage0_5[193]},
      {stage0_7[48], stage0_7[49], stage0_7[50], stage0_7[51], stage0_7[52], stage0_7[53]},
      {stage1_9[8],stage1_8[74],stage1_7[96],stage1_6[113],stage1_5[152]}
   );
   gpc606_5 gpc254 (
      {stage0_5[194], stage0_5[195], stage0_5[196], stage0_5[197], stage0_5[198], stage0_5[199]},
      {stage0_7[54], stage0_7[55], stage0_7[56], stage0_7[57], stage0_7[58], stage0_7[59]},
      {stage1_9[9],stage1_8[75],stage1_7[97],stage1_6[114],stage1_5[153]}
   );
   gpc606_5 gpc255 (
      {stage0_5[200], stage0_5[201], stage0_5[202], stage0_5[203], stage0_5[204], stage0_5[205]},
      {stage0_7[60], stage0_7[61], stage0_7[62], stage0_7[63], stage0_7[64], stage0_7[65]},
      {stage1_9[10],stage1_8[76],stage1_7[98],stage1_6[115],stage1_5[154]}
   );
   gpc606_5 gpc256 (
      {stage0_5[206], stage0_5[207], stage0_5[208], stage0_5[209], stage0_5[210], stage0_5[211]},
      {stage0_7[66], stage0_7[67], stage0_7[68], stage0_7[69], stage0_7[70], stage0_7[71]},
      {stage1_9[11],stage1_8[77],stage1_7[99],stage1_6[116],stage1_5[155]}
   );
   gpc606_5 gpc257 (
      {stage0_5[212], stage0_5[213], stage0_5[214], stage0_5[215], stage0_5[216], stage0_5[217]},
      {stage0_7[72], stage0_7[73], stage0_7[74], stage0_7[75], stage0_7[76], stage0_7[77]},
      {stage1_9[12],stage1_8[78],stage1_7[100],stage1_6[117],stage1_5[156]}
   );
   gpc606_5 gpc258 (
      {stage0_5[218], stage0_5[219], stage0_5[220], stage0_5[221], stage0_5[222], stage0_5[223]},
      {stage0_7[78], stage0_7[79], stage0_7[80], stage0_7[81], stage0_7[82], stage0_7[83]},
      {stage1_9[13],stage1_8[79],stage1_7[101],stage1_6[118],stage1_5[157]}
   );
   gpc606_5 gpc259 (
      {stage0_5[224], stage0_5[225], stage0_5[226], stage0_5[227], stage0_5[228], stage0_5[229]},
      {stage0_7[84], stage0_7[85], stage0_7[86], stage0_7[87], stage0_7[88], stage0_7[89]},
      {stage1_9[14],stage1_8[80],stage1_7[102],stage1_6[119],stage1_5[158]}
   );
   gpc606_5 gpc260 (
      {stage0_5[230], stage0_5[231], stage0_5[232], stage0_5[233], stage0_5[234], stage0_5[235]},
      {stage0_7[90], stage0_7[91], stage0_7[92], stage0_7[93], stage0_7[94], stage0_7[95]},
      {stage1_9[15],stage1_8[81],stage1_7[103],stage1_6[120],stage1_5[159]}
   );
   gpc606_5 gpc261 (
      {stage0_5[236], stage0_5[237], stage0_5[238], stage0_5[239], stage0_5[240], stage0_5[241]},
      {stage0_7[96], stage0_7[97], stage0_7[98], stage0_7[99], stage0_7[100], stage0_7[101]},
      {stage1_9[16],stage1_8[82],stage1_7[104],stage1_6[121],stage1_5[160]}
   );
   gpc606_5 gpc262 (
      {stage0_5[242], stage0_5[243], stage0_5[244], stage0_5[245], stage0_5[246], stage0_5[247]},
      {stage0_7[102], stage0_7[103], stage0_7[104], stage0_7[105], stage0_7[106], stage0_7[107]},
      {stage1_9[17],stage1_8[83],stage1_7[105],stage1_6[122],stage1_5[161]}
   );
   gpc606_5 gpc263 (
      {stage0_5[248], stage0_5[249], stage0_5[250], stage0_5[251], stage0_5[252], stage0_5[253]},
      {stage0_7[108], stage0_7[109], stage0_7[110], stage0_7[111], stage0_7[112], stage0_7[113]},
      {stage1_9[18],stage1_8[84],stage1_7[106],stage1_6[123],stage1_5[162]}
   );
   gpc606_5 gpc264 (
      {stage0_5[254], stage0_5[255], stage0_5[256], stage0_5[257], stage0_5[258], stage0_5[259]},
      {stage0_7[114], stage0_7[115], stage0_7[116], stage0_7[117], stage0_7[118], stage0_7[119]},
      {stage1_9[19],stage1_8[85],stage1_7[107],stage1_6[124],stage1_5[163]}
   );
   gpc606_5 gpc265 (
      {stage0_5[260], stage0_5[261], stage0_5[262], stage0_5[263], stage0_5[264], stage0_5[265]},
      {stage0_7[120], stage0_7[121], stage0_7[122], stage0_7[123], stage0_7[124], stage0_7[125]},
      {stage1_9[20],stage1_8[86],stage1_7[108],stage1_6[125],stage1_5[164]}
   );
   gpc606_5 gpc266 (
      {stage0_5[266], stage0_5[267], stage0_5[268], stage0_5[269], stage0_5[270], stage0_5[271]},
      {stage0_7[126], stage0_7[127], stage0_7[128], stage0_7[129], stage0_7[130], stage0_7[131]},
      {stage1_9[21],stage1_8[87],stage1_7[109],stage1_6[126],stage1_5[165]}
   );
   gpc606_5 gpc267 (
      {stage0_5[272], stage0_5[273], stage0_5[274], stage0_5[275], stage0_5[276], stage0_5[277]},
      {stage0_7[132], stage0_7[133], stage0_7[134], stage0_7[135], stage0_7[136], stage0_7[137]},
      {stage1_9[22],stage1_8[88],stage1_7[110],stage1_6[127],stage1_5[166]}
   );
   gpc606_5 gpc268 (
      {stage0_5[278], stage0_5[279], stage0_5[280], stage0_5[281], stage0_5[282], stage0_5[283]},
      {stage0_7[138], stage0_7[139], stage0_7[140], stage0_7[141], stage0_7[142], stage0_7[143]},
      {stage1_9[23],stage1_8[89],stage1_7[111],stage1_6[128],stage1_5[167]}
   );
   gpc606_5 gpc269 (
      {stage0_5[284], stage0_5[285], stage0_5[286], stage0_5[287], stage0_5[288], stage0_5[289]},
      {stage0_7[144], stage0_7[145], stage0_7[146], stage0_7[147], stage0_7[148], stage0_7[149]},
      {stage1_9[24],stage1_8[90],stage1_7[112],stage1_6[129],stage1_5[168]}
   );
   gpc606_5 gpc270 (
      {stage0_5[290], stage0_5[291], stage0_5[292], stage0_5[293], stage0_5[294], stage0_5[295]},
      {stage0_7[150], stage0_7[151], stage0_7[152], stage0_7[153], stage0_7[154], stage0_7[155]},
      {stage1_9[25],stage1_8[91],stage1_7[113],stage1_6[130],stage1_5[169]}
   );
   gpc606_5 gpc271 (
      {stage0_5[296], stage0_5[297], stage0_5[298], stage0_5[299], stage0_5[300], stage0_5[301]},
      {stage0_7[156], stage0_7[157], stage0_7[158], stage0_7[159], stage0_7[160], stage0_7[161]},
      {stage1_9[26],stage1_8[92],stage1_7[114],stage1_6[131],stage1_5[170]}
   );
   gpc606_5 gpc272 (
      {stage0_5[302], stage0_5[303], stage0_5[304], stage0_5[305], stage0_5[306], stage0_5[307]},
      {stage0_7[162], stage0_7[163], stage0_7[164], stage0_7[165], stage0_7[166], stage0_7[167]},
      {stage1_9[27],stage1_8[93],stage1_7[115],stage1_6[132],stage1_5[171]}
   );
   gpc606_5 gpc273 (
      {stage0_5[308], stage0_5[309], stage0_5[310], stage0_5[311], stage0_5[312], stage0_5[313]},
      {stage0_7[168], stage0_7[169], stage0_7[170], stage0_7[171], stage0_7[172], stage0_7[173]},
      {stage1_9[28],stage1_8[94],stage1_7[116],stage1_6[133],stage1_5[172]}
   );
   gpc606_5 gpc274 (
      {stage0_5[314], stage0_5[315], stage0_5[316], stage0_5[317], stage0_5[318], stage0_5[319]},
      {stage0_7[174], stage0_7[175], stage0_7[176], stage0_7[177], stage0_7[178], stage0_7[179]},
      {stage1_9[29],stage1_8[95],stage1_7[117],stage1_6[134],stage1_5[173]}
   );
   gpc606_5 gpc275 (
      {stage0_5[320], stage0_5[321], stage0_5[322], stage0_5[323], stage0_5[324], stage0_5[325]},
      {stage0_7[180], stage0_7[181], stage0_7[182], stage0_7[183], stage0_7[184], stage0_7[185]},
      {stage1_9[30],stage1_8[96],stage1_7[118],stage1_6[135],stage1_5[174]}
   );
   gpc606_5 gpc276 (
      {stage0_5[326], stage0_5[327], stage0_5[328], stage0_5[329], stage0_5[330], stage0_5[331]},
      {stage0_7[186], stage0_7[187], stage0_7[188], stage0_7[189], stage0_7[190], stage0_7[191]},
      {stage1_9[31],stage1_8[97],stage1_7[119],stage1_6[136],stage1_5[175]}
   );
   gpc606_5 gpc277 (
      {stage0_5[332], stage0_5[333], stage0_5[334], stage0_5[335], stage0_5[336], stage0_5[337]},
      {stage0_7[192], stage0_7[193], stage0_7[194], stage0_7[195], stage0_7[196], stage0_7[197]},
      {stage1_9[32],stage1_8[98],stage1_7[120],stage1_6[137],stage1_5[176]}
   );
   gpc606_5 gpc278 (
      {stage0_5[338], stage0_5[339], stage0_5[340], stage0_5[341], stage0_5[342], stage0_5[343]},
      {stage0_7[198], stage0_7[199], stage0_7[200], stage0_7[201], stage0_7[202], stage0_7[203]},
      {stage1_9[33],stage1_8[99],stage1_7[121],stage1_6[138],stage1_5[177]}
   );
   gpc606_5 gpc279 (
      {stage0_5[344], stage0_5[345], stage0_5[346], stage0_5[347], stage0_5[348], stage0_5[349]},
      {stage0_7[204], stage0_7[205], stage0_7[206], stage0_7[207], stage0_7[208], stage0_7[209]},
      {stage1_9[34],stage1_8[100],stage1_7[122],stage1_6[139],stage1_5[178]}
   );
   gpc606_5 gpc280 (
      {stage0_5[350], stage0_5[351], stage0_5[352], stage0_5[353], stage0_5[354], stage0_5[355]},
      {stage0_7[210], stage0_7[211], stage0_7[212], stage0_7[213], stage0_7[214], stage0_7[215]},
      {stage1_9[35],stage1_8[101],stage1_7[123],stage1_6[140],stage1_5[179]}
   );
   gpc606_5 gpc281 (
      {stage0_5[356], stage0_5[357], stage0_5[358], stage0_5[359], stage0_5[360], stage0_5[361]},
      {stage0_7[216], stage0_7[217], stage0_7[218], stage0_7[219], stage0_7[220], stage0_7[221]},
      {stage1_9[36],stage1_8[102],stage1_7[124],stage1_6[141],stage1_5[180]}
   );
   gpc606_5 gpc282 (
      {stage0_5[362], stage0_5[363], stage0_5[364], stage0_5[365], stage0_5[366], stage0_5[367]},
      {stage0_7[222], stage0_7[223], stage0_7[224], stage0_7[225], stage0_7[226], stage0_7[227]},
      {stage1_9[37],stage1_8[103],stage1_7[125],stage1_6[142],stage1_5[181]}
   );
   gpc606_5 gpc283 (
      {stage0_5[368], stage0_5[369], stage0_5[370], stage0_5[371], stage0_5[372], stage0_5[373]},
      {stage0_7[228], stage0_7[229], stage0_7[230], stage0_7[231], stage0_7[232], stage0_7[233]},
      {stage1_9[38],stage1_8[104],stage1_7[126],stage1_6[143],stage1_5[182]}
   );
   gpc606_5 gpc284 (
      {stage0_5[374], stage0_5[375], stage0_5[376], stage0_5[377], stage0_5[378], stage0_5[379]},
      {stage0_7[234], stage0_7[235], stage0_7[236], stage0_7[237], stage0_7[238], stage0_7[239]},
      {stage1_9[39],stage1_8[105],stage1_7[127],stage1_6[144],stage1_5[183]}
   );
   gpc606_5 gpc285 (
      {stage0_5[380], stage0_5[381], stage0_5[382], stage0_5[383], stage0_5[384], stage0_5[385]},
      {stage0_7[240], stage0_7[241], stage0_7[242], stage0_7[243], stage0_7[244], stage0_7[245]},
      {stage1_9[40],stage1_8[106],stage1_7[128],stage1_6[145],stage1_5[184]}
   );
   gpc606_5 gpc286 (
      {stage0_5[386], stage0_5[387], stage0_5[388], stage0_5[389], stage0_5[390], stage0_5[391]},
      {stage0_7[246], stage0_7[247], stage0_7[248], stage0_7[249], stage0_7[250], stage0_7[251]},
      {stage1_9[41],stage1_8[107],stage1_7[129],stage1_6[146],stage1_5[185]}
   );
   gpc606_5 gpc287 (
      {stage0_5[392], stage0_5[393], stage0_5[394], stage0_5[395], stage0_5[396], stage0_5[397]},
      {stage0_7[252], stage0_7[253], stage0_7[254], stage0_7[255], stage0_7[256], stage0_7[257]},
      {stage1_9[42],stage1_8[108],stage1_7[130],stage1_6[147],stage1_5[186]}
   );
   gpc606_5 gpc288 (
      {stage0_5[398], stage0_5[399], stage0_5[400], stage0_5[401], stage0_5[402], stage0_5[403]},
      {stage0_7[258], stage0_7[259], stage0_7[260], stage0_7[261], stage0_7[262], stage0_7[263]},
      {stage1_9[43],stage1_8[109],stage1_7[131],stage1_6[148],stage1_5[187]}
   );
   gpc606_5 gpc289 (
      {stage0_5[404], stage0_5[405], stage0_5[406], stage0_5[407], stage0_5[408], stage0_5[409]},
      {stage0_7[264], stage0_7[265], stage0_7[266], stage0_7[267], stage0_7[268], stage0_7[269]},
      {stage1_9[44],stage1_8[110],stage1_7[132],stage1_6[149],stage1_5[188]}
   );
   gpc606_5 gpc290 (
      {stage0_5[410], stage0_5[411], stage0_5[412], stage0_5[413], stage0_5[414], stage0_5[415]},
      {stage0_7[270], stage0_7[271], stage0_7[272], stage0_7[273], stage0_7[274], stage0_7[275]},
      {stage1_9[45],stage1_8[111],stage1_7[133],stage1_6[150],stage1_5[189]}
   );
   gpc606_5 gpc291 (
      {stage0_5[416], stage0_5[417], stage0_5[418], stage0_5[419], stage0_5[420], stage0_5[421]},
      {stage0_7[276], stage0_7[277], stage0_7[278], stage0_7[279], stage0_7[280], stage0_7[281]},
      {stage1_9[46],stage1_8[112],stage1_7[134],stage1_6[151],stage1_5[190]}
   );
   gpc606_5 gpc292 (
      {stage0_5[422], stage0_5[423], stage0_5[424], stage0_5[425], stage0_5[426], stage0_5[427]},
      {stage0_7[282], stage0_7[283], stage0_7[284], stage0_7[285], stage0_7[286], stage0_7[287]},
      {stage1_9[47],stage1_8[113],stage1_7[135],stage1_6[152],stage1_5[191]}
   );
   gpc606_5 gpc293 (
      {stage0_5[428], stage0_5[429], stage0_5[430], stage0_5[431], stage0_5[432], stage0_5[433]},
      {stage0_7[288], stage0_7[289], stage0_7[290], stage0_7[291], stage0_7[292], stage0_7[293]},
      {stage1_9[48],stage1_8[114],stage1_7[136],stage1_6[153],stage1_5[192]}
   );
   gpc606_5 gpc294 (
      {stage0_5[434], stage0_5[435], stage0_5[436], stage0_5[437], stage0_5[438], stage0_5[439]},
      {stage0_7[294], stage0_7[295], stage0_7[296], stage0_7[297], stage0_7[298], stage0_7[299]},
      {stage1_9[49],stage1_8[115],stage1_7[137],stage1_6[154],stage1_5[193]}
   );
   gpc606_5 gpc295 (
      {stage0_5[440], stage0_5[441], stage0_5[442], stage0_5[443], stage0_5[444], stage0_5[445]},
      {stage0_7[300], stage0_7[301], stage0_7[302], stage0_7[303], stage0_7[304], stage0_7[305]},
      {stage1_9[50],stage1_8[116],stage1_7[138],stage1_6[155],stage1_5[194]}
   );
   gpc606_5 gpc296 (
      {stage0_5[446], stage0_5[447], stage0_5[448], stage0_5[449], stage0_5[450], stage0_5[451]},
      {stage0_7[306], stage0_7[307], stage0_7[308], stage0_7[309], stage0_7[310], stage0_7[311]},
      {stage1_9[51],stage1_8[117],stage1_7[139],stage1_6[156],stage1_5[195]}
   );
   gpc606_5 gpc297 (
      {stage0_5[452], stage0_5[453], stage0_5[454], stage0_5[455], stage0_5[456], stage0_5[457]},
      {stage0_7[312], stage0_7[313], stage0_7[314], stage0_7[315], stage0_7[316], stage0_7[317]},
      {stage1_9[52],stage1_8[118],stage1_7[140],stage1_6[157],stage1_5[196]}
   );
   gpc606_5 gpc298 (
      {stage0_5[458], stage0_5[459], stage0_5[460], stage0_5[461], stage0_5[462], stage0_5[463]},
      {stage0_7[318], stage0_7[319], stage0_7[320], stage0_7[321], stage0_7[322], stage0_7[323]},
      {stage1_9[53],stage1_8[119],stage1_7[141],stage1_6[158],stage1_5[197]}
   );
   gpc606_5 gpc299 (
      {stage0_5[464], stage0_5[465], stage0_5[466], stage0_5[467], stage0_5[468], stage0_5[469]},
      {stage0_7[324], stage0_7[325], stage0_7[326], stage0_7[327], stage0_7[328], stage0_7[329]},
      {stage1_9[54],stage1_8[120],stage1_7[142],stage1_6[159],stage1_5[198]}
   );
   gpc606_5 gpc300 (
      {stage0_5[470], stage0_5[471], stage0_5[472], stage0_5[473], stage0_5[474], stage0_5[475]},
      {stage0_7[330], stage0_7[331], stage0_7[332], stage0_7[333], stage0_7[334], stage0_7[335]},
      {stage1_9[55],stage1_8[121],stage1_7[143],stage1_6[160],stage1_5[199]}
   );
   gpc606_5 gpc301 (
      {stage0_5[476], stage0_5[477], stage0_5[478], stage0_5[479], stage0_5[480], stage0_5[481]},
      {stage0_7[336], stage0_7[337], stage0_7[338], stage0_7[339], stage0_7[340], stage0_7[341]},
      {stage1_9[56],stage1_8[122],stage1_7[144],stage1_6[161],stage1_5[200]}
   );
   gpc606_5 gpc302 (
      {stage0_5[482], stage0_5[483], stage0_5[484], stage0_5[485], stage0_5[486], stage0_5[487]},
      {stage0_7[342], stage0_7[343], stage0_7[344], stage0_7[345], stage0_7[346], stage0_7[347]},
      {stage1_9[57],stage1_8[123],stage1_7[145],stage1_6[162],stage1_5[201]}
   );
   gpc606_5 gpc303 (
      {stage0_5[488], stage0_5[489], stage0_5[490], stage0_5[491], stage0_5[492], stage0_5[493]},
      {stage0_7[348], stage0_7[349], stage0_7[350], stage0_7[351], stage0_7[352], stage0_7[353]},
      {stage1_9[58],stage1_8[124],stage1_7[146],stage1_6[163],stage1_5[202]}
   );
   gpc606_5 gpc304 (
      {stage0_5[494], stage0_5[495], stage0_5[496], stage0_5[497], stage0_5[498], stage0_5[499]},
      {stage0_7[354], stage0_7[355], stage0_7[356], stage0_7[357], stage0_7[358], stage0_7[359]},
      {stage1_9[59],stage1_8[125],stage1_7[147],stage1_6[164],stage1_5[203]}
   );
   gpc606_5 gpc305 (
      {stage0_5[500], stage0_5[501], stage0_5[502], stage0_5[503], stage0_5[504], stage0_5[505]},
      {stage0_7[360], stage0_7[361], stage0_7[362], stage0_7[363], stage0_7[364], stage0_7[365]},
      {stage1_9[60],stage1_8[126],stage1_7[148],stage1_6[165],stage1_5[204]}
   );
   gpc606_5 gpc306 (
      {stage0_5[506], stage0_5[507], stage0_5[508], stage0_5[509], stage0_5[510], stage0_5[511]},
      {stage0_7[366], stage0_7[367], stage0_7[368], stage0_7[369], stage0_7[370], stage0_7[371]},
      {stage1_9[61],stage1_8[127],stage1_7[149],stage1_6[166],stage1_5[205]}
   );
   gpc615_5 gpc307 (
      {stage0_6[396], stage0_6[397], stage0_6[398], stage0_6[399], stage0_6[400]},
      {stage0_7[372]},
      {stage0_8[0], stage0_8[1], stage0_8[2], stage0_8[3], stage0_8[4], stage0_8[5]},
      {stage1_10[0],stage1_9[62],stage1_8[128],stage1_7[150],stage1_6[167]}
   );
   gpc615_5 gpc308 (
      {stage0_6[401], stage0_6[402], stage0_6[403], stage0_6[404], stage0_6[405]},
      {stage0_7[373]},
      {stage0_8[6], stage0_8[7], stage0_8[8], stage0_8[9], stage0_8[10], stage0_8[11]},
      {stage1_10[1],stage1_9[63],stage1_8[129],stage1_7[151],stage1_6[168]}
   );
   gpc615_5 gpc309 (
      {stage0_6[406], stage0_6[407], stage0_6[408], stage0_6[409], stage0_6[410]},
      {stage0_7[374]},
      {stage0_8[12], stage0_8[13], stage0_8[14], stage0_8[15], stage0_8[16], stage0_8[17]},
      {stage1_10[2],stage1_9[64],stage1_8[130],stage1_7[152],stage1_6[169]}
   );
   gpc615_5 gpc310 (
      {stage0_6[411], stage0_6[412], stage0_6[413], stage0_6[414], stage0_6[415]},
      {stage0_7[375]},
      {stage0_8[18], stage0_8[19], stage0_8[20], stage0_8[21], stage0_8[22], stage0_8[23]},
      {stage1_10[3],stage1_9[65],stage1_8[131],stage1_7[153],stage1_6[170]}
   );
   gpc615_5 gpc311 (
      {stage0_6[416], stage0_6[417], stage0_6[418], stage0_6[419], stage0_6[420]},
      {stage0_7[376]},
      {stage0_8[24], stage0_8[25], stage0_8[26], stage0_8[27], stage0_8[28], stage0_8[29]},
      {stage1_10[4],stage1_9[66],stage1_8[132],stage1_7[154],stage1_6[171]}
   );
   gpc615_5 gpc312 (
      {stage0_6[421], stage0_6[422], stage0_6[423], stage0_6[424], stage0_6[425]},
      {stage0_7[377]},
      {stage0_8[30], stage0_8[31], stage0_8[32], stage0_8[33], stage0_8[34], stage0_8[35]},
      {stage1_10[5],stage1_9[67],stage1_8[133],stage1_7[155],stage1_6[172]}
   );
   gpc615_5 gpc313 (
      {stage0_6[426], stage0_6[427], stage0_6[428], stage0_6[429], stage0_6[430]},
      {stage0_7[378]},
      {stage0_8[36], stage0_8[37], stage0_8[38], stage0_8[39], stage0_8[40], stage0_8[41]},
      {stage1_10[6],stage1_9[68],stage1_8[134],stage1_7[156],stage1_6[173]}
   );
   gpc615_5 gpc314 (
      {stage0_6[431], stage0_6[432], stage0_6[433], stage0_6[434], stage0_6[435]},
      {stage0_7[379]},
      {stage0_8[42], stage0_8[43], stage0_8[44], stage0_8[45], stage0_8[46], stage0_8[47]},
      {stage1_10[7],stage1_9[69],stage1_8[135],stage1_7[157],stage1_6[174]}
   );
   gpc615_5 gpc315 (
      {stage0_6[436], stage0_6[437], stage0_6[438], stage0_6[439], stage0_6[440]},
      {stage0_7[380]},
      {stage0_8[48], stage0_8[49], stage0_8[50], stage0_8[51], stage0_8[52], stage0_8[53]},
      {stage1_10[8],stage1_9[70],stage1_8[136],stage1_7[158],stage1_6[175]}
   );
   gpc615_5 gpc316 (
      {stage0_6[441], stage0_6[442], stage0_6[443], stage0_6[444], stage0_6[445]},
      {stage0_7[381]},
      {stage0_8[54], stage0_8[55], stage0_8[56], stage0_8[57], stage0_8[58], stage0_8[59]},
      {stage1_10[9],stage1_9[71],stage1_8[137],stage1_7[159],stage1_6[176]}
   );
   gpc615_5 gpc317 (
      {stage0_7[382], stage0_7[383], stage0_7[384], stage0_7[385], stage0_7[386]},
      {stage0_8[60]},
      {stage0_9[0], stage0_9[1], stage0_9[2], stage0_9[3], stage0_9[4], stage0_9[5]},
      {stage1_11[0],stage1_10[10],stage1_9[72],stage1_8[138],stage1_7[160]}
   );
   gpc615_5 gpc318 (
      {stage0_7[387], stage0_7[388], stage0_7[389], stage0_7[390], stage0_7[391]},
      {stage0_8[61]},
      {stage0_9[6], stage0_9[7], stage0_9[8], stage0_9[9], stage0_9[10], stage0_9[11]},
      {stage1_11[1],stage1_10[11],stage1_9[73],stage1_8[139],stage1_7[161]}
   );
   gpc615_5 gpc319 (
      {stage0_7[392], stage0_7[393], stage0_7[394], stage0_7[395], stage0_7[396]},
      {stage0_8[62]},
      {stage0_9[12], stage0_9[13], stage0_9[14], stage0_9[15], stage0_9[16], stage0_9[17]},
      {stage1_11[2],stage1_10[12],stage1_9[74],stage1_8[140],stage1_7[162]}
   );
   gpc615_5 gpc320 (
      {stage0_7[397], stage0_7[398], stage0_7[399], stage0_7[400], stage0_7[401]},
      {stage0_8[63]},
      {stage0_9[18], stage0_9[19], stage0_9[20], stage0_9[21], stage0_9[22], stage0_9[23]},
      {stage1_11[3],stage1_10[13],stage1_9[75],stage1_8[141],stage1_7[163]}
   );
   gpc615_5 gpc321 (
      {stage0_7[402], stage0_7[403], stage0_7[404], stage0_7[405], stage0_7[406]},
      {stage0_8[64]},
      {stage0_9[24], stage0_9[25], stage0_9[26], stage0_9[27], stage0_9[28], stage0_9[29]},
      {stage1_11[4],stage1_10[14],stage1_9[76],stage1_8[142],stage1_7[164]}
   );
   gpc615_5 gpc322 (
      {stage0_7[407], stage0_7[408], stage0_7[409], stage0_7[410], stage0_7[411]},
      {stage0_8[65]},
      {stage0_9[30], stage0_9[31], stage0_9[32], stage0_9[33], stage0_9[34], stage0_9[35]},
      {stage1_11[5],stage1_10[15],stage1_9[77],stage1_8[143],stage1_7[165]}
   );
   gpc615_5 gpc323 (
      {stage0_7[412], stage0_7[413], stage0_7[414], stage0_7[415], stage0_7[416]},
      {stage0_8[66]},
      {stage0_9[36], stage0_9[37], stage0_9[38], stage0_9[39], stage0_9[40], stage0_9[41]},
      {stage1_11[6],stage1_10[16],stage1_9[78],stage1_8[144],stage1_7[166]}
   );
   gpc615_5 gpc324 (
      {stage0_7[417], stage0_7[418], stage0_7[419], stage0_7[420], stage0_7[421]},
      {stage0_8[67]},
      {stage0_9[42], stage0_9[43], stage0_9[44], stage0_9[45], stage0_9[46], stage0_9[47]},
      {stage1_11[7],stage1_10[17],stage1_9[79],stage1_8[145],stage1_7[167]}
   );
   gpc615_5 gpc325 (
      {stage0_7[422], stage0_7[423], stage0_7[424], stage0_7[425], stage0_7[426]},
      {stage0_8[68]},
      {stage0_9[48], stage0_9[49], stage0_9[50], stage0_9[51], stage0_9[52], stage0_9[53]},
      {stage1_11[8],stage1_10[18],stage1_9[80],stage1_8[146],stage1_7[168]}
   );
   gpc615_5 gpc326 (
      {stage0_7[427], stage0_7[428], stage0_7[429], stage0_7[430], stage0_7[431]},
      {stage0_8[69]},
      {stage0_9[54], stage0_9[55], stage0_9[56], stage0_9[57], stage0_9[58], stage0_9[59]},
      {stage1_11[9],stage1_10[19],stage1_9[81],stage1_8[147],stage1_7[169]}
   );
   gpc615_5 gpc327 (
      {stage0_7[432], stage0_7[433], stage0_7[434], stage0_7[435], stage0_7[436]},
      {stage0_8[70]},
      {stage0_9[60], stage0_9[61], stage0_9[62], stage0_9[63], stage0_9[64], stage0_9[65]},
      {stage1_11[10],stage1_10[20],stage1_9[82],stage1_8[148],stage1_7[170]}
   );
   gpc615_5 gpc328 (
      {stage0_7[437], stage0_7[438], stage0_7[439], stage0_7[440], stage0_7[441]},
      {stage0_8[71]},
      {stage0_9[66], stage0_9[67], stage0_9[68], stage0_9[69], stage0_9[70], stage0_9[71]},
      {stage1_11[11],stage1_10[21],stage1_9[83],stage1_8[149],stage1_7[171]}
   );
   gpc615_5 gpc329 (
      {stage0_7[442], stage0_7[443], stage0_7[444], stage0_7[445], stage0_7[446]},
      {stage0_8[72]},
      {stage0_9[72], stage0_9[73], stage0_9[74], stage0_9[75], stage0_9[76], stage0_9[77]},
      {stage1_11[12],stage1_10[22],stage1_9[84],stage1_8[150],stage1_7[172]}
   );
   gpc615_5 gpc330 (
      {stage0_7[447], stage0_7[448], stage0_7[449], stage0_7[450], stage0_7[451]},
      {stage0_8[73]},
      {stage0_9[78], stage0_9[79], stage0_9[80], stage0_9[81], stage0_9[82], stage0_9[83]},
      {stage1_11[13],stage1_10[23],stage1_9[85],stage1_8[151],stage1_7[173]}
   );
   gpc615_5 gpc331 (
      {stage0_7[452], stage0_7[453], stage0_7[454], stage0_7[455], stage0_7[456]},
      {stage0_8[74]},
      {stage0_9[84], stage0_9[85], stage0_9[86], stage0_9[87], stage0_9[88], stage0_9[89]},
      {stage1_11[14],stage1_10[24],stage1_9[86],stage1_8[152],stage1_7[174]}
   );
   gpc615_5 gpc332 (
      {stage0_7[457], stage0_7[458], stage0_7[459], stage0_7[460], stage0_7[461]},
      {stage0_8[75]},
      {stage0_9[90], stage0_9[91], stage0_9[92], stage0_9[93], stage0_9[94], stage0_9[95]},
      {stage1_11[15],stage1_10[25],stage1_9[87],stage1_8[153],stage1_7[175]}
   );
   gpc615_5 gpc333 (
      {stage0_7[462], stage0_7[463], stage0_7[464], stage0_7[465], stage0_7[466]},
      {stage0_8[76]},
      {stage0_9[96], stage0_9[97], stage0_9[98], stage0_9[99], stage0_9[100], stage0_9[101]},
      {stage1_11[16],stage1_10[26],stage1_9[88],stage1_8[154],stage1_7[176]}
   );
   gpc615_5 gpc334 (
      {stage0_7[467], stage0_7[468], stage0_7[469], stage0_7[470], stage0_7[471]},
      {stage0_8[77]},
      {stage0_9[102], stage0_9[103], stage0_9[104], stage0_9[105], stage0_9[106], stage0_9[107]},
      {stage1_11[17],stage1_10[27],stage1_9[89],stage1_8[155],stage1_7[177]}
   );
   gpc615_5 gpc335 (
      {stage0_7[472], stage0_7[473], stage0_7[474], stage0_7[475], stage0_7[476]},
      {stage0_8[78]},
      {stage0_9[108], stage0_9[109], stage0_9[110], stage0_9[111], stage0_9[112], stage0_9[113]},
      {stage1_11[18],stage1_10[28],stage1_9[90],stage1_8[156],stage1_7[178]}
   );
   gpc615_5 gpc336 (
      {stage0_7[477], stage0_7[478], stage0_7[479], stage0_7[480], stage0_7[481]},
      {stage0_8[79]},
      {stage0_9[114], stage0_9[115], stage0_9[116], stage0_9[117], stage0_9[118], stage0_9[119]},
      {stage1_11[19],stage1_10[29],stage1_9[91],stage1_8[157],stage1_7[179]}
   );
   gpc615_5 gpc337 (
      {stage0_7[482], stage0_7[483], stage0_7[484], stage0_7[485], stage0_7[486]},
      {stage0_8[80]},
      {stage0_9[120], stage0_9[121], stage0_9[122], stage0_9[123], stage0_9[124], stage0_9[125]},
      {stage1_11[20],stage1_10[30],stage1_9[92],stage1_8[158],stage1_7[180]}
   );
   gpc615_5 gpc338 (
      {stage0_7[487], stage0_7[488], stage0_7[489], stage0_7[490], stage0_7[491]},
      {stage0_8[81]},
      {stage0_9[126], stage0_9[127], stage0_9[128], stage0_9[129], stage0_9[130], stage0_9[131]},
      {stage1_11[21],stage1_10[31],stage1_9[93],stage1_8[159],stage1_7[181]}
   );
   gpc615_5 gpc339 (
      {stage0_7[492], stage0_7[493], stage0_7[494], stage0_7[495], stage0_7[496]},
      {stage0_8[82]},
      {stage0_9[132], stage0_9[133], stage0_9[134], stage0_9[135], stage0_9[136], stage0_9[137]},
      {stage1_11[22],stage1_10[32],stage1_9[94],stage1_8[160],stage1_7[182]}
   );
   gpc615_5 gpc340 (
      {stage0_7[497], stage0_7[498], stage0_7[499], stage0_7[500], stage0_7[501]},
      {stage0_8[83]},
      {stage0_9[138], stage0_9[139], stage0_9[140], stage0_9[141], stage0_9[142], stage0_9[143]},
      {stage1_11[23],stage1_10[33],stage1_9[95],stage1_8[161],stage1_7[183]}
   );
   gpc615_5 gpc341 (
      {stage0_7[502], stage0_7[503], stage0_7[504], stage0_7[505], stage0_7[506]},
      {stage0_8[84]},
      {stage0_9[144], stage0_9[145], stage0_9[146], stage0_9[147], stage0_9[148], stage0_9[149]},
      {stage1_11[24],stage1_10[34],stage1_9[96],stage1_8[162],stage1_7[184]}
   );
   gpc615_5 gpc342 (
      {stage0_7[507], stage0_7[508], stage0_7[509], stage0_7[510], stage0_7[511]},
      {stage0_8[85]},
      {stage0_9[150], stage0_9[151], stage0_9[152], stage0_9[153], stage0_9[154], stage0_9[155]},
      {stage1_11[25],stage1_10[35],stage1_9[97],stage1_8[163],stage1_7[185]}
   );
   gpc606_5 gpc343 (
      {stage0_8[86], stage0_8[87], stage0_8[88], stage0_8[89], stage0_8[90], stage0_8[91]},
      {stage0_10[0], stage0_10[1], stage0_10[2], stage0_10[3], stage0_10[4], stage0_10[5]},
      {stage1_12[0],stage1_11[26],stage1_10[36],stage1_9[98],stage1_8[164]}
   );
   gpc606_5 gpc344 (
      {stage0_8[92], stage0_8[93], stage0_8[94], stage0_8[95], stage0_8[96], stage0_8[97]},
      {stage0_10[6], stage0_10[7], stage0_10[8], stage0_10[9], stage0_10[10], stage0_10[11]},
      {stage1_12[1],stage1_11[27],stage1_10[37],stage1_9[99],stage1_8[165]}
   );
   gpc606_5 gpc345 (
      {stage0_8[98], stage0_8[99], stage0_8[100], stage0_8[101], stage0_8[102], stage0_8[103]},
      {stage0_10[12], stage0_10[13], stage0_10[14], stage0_10[15], stage0_10[16], stage0_10[17]},
      {stage1_12[2],stage1_11[28],stage1_10[38],stage1_9[100],stage1_8[166]}
   );
   gpc606_5 gpc346 (
      {stage0_8[104], stage0_8[105], stage0_8[106], stage0_8[107], stage0_8[108], stage0_8[109]},
      {stage0_10[18], stage0_10[19], stage0_10[20], stage0_10[21], stage0_10[22], stage0_10[23]},
      {stage1_12[3],stage1_11[29],stage1_10[39],stage1_9[101],stage1_8[167]}
   );
   gpc606_5 gpc347 (
      {stage0_8[110], stage0_8[111], stage0_8[112], stage0_8[113], stage0_8[114], stage0_8[115]},
      {stage0_10[24], stage0_10[25], stage0_10[26], stage0_10[27], stage0_10[28], stage0_10[29]},
      {stage1_12[4],stage1_11[30],stage1_10[40],stage1_9[102],stage1_8[168]}
   );
   gpc606_5 gpc348 (
      {stage0_8[116], stage0_8[117], stage0_8[118], stage0_8[119], stage0_8[120], stage0_8[121]},
      {stage0_10[30], stage0_10[31], stage0_10[32], stage0_10[33], stage0_10[34], stage0_10[35]},
      {stage1_12[5],stage1_11[31],stage1_10[41],stage1_9[103],stage1_8[169]}
   );
   gpc606_5 gpc349 (
      {stage0_8[122], stage0_8[123], stage0_8[124], stage0_8[125], stage0_8[126], stage0_8[127]},
      {stage0_10[36], stage0_10[37], stage0_10[38], stage0_10[39], stage0_10[40], stage0_10[41]},
      {stage1_12[6],stage1_11[32],stage1_10[42],stage1_9[104],stage1_8[170]}
   );
   gpc606_5 gpc350 (
      {stage0_8[128], stage0_8[129], stage0_8[130], stage0_8[131], stage0_8[132], stage0_8[133]},
      {stage0_10[42], stage0_10[43], stage0_10[44], stage0_10[45], stage0_10[46], stage0_10[47]},
      {stage1_12[7],stage1_11[33],stage1_10[43],stage1_9[105],stage1_8[171]}
   );
   gpc606_5 gpc351 (
      {stage0_8[134], stage0_8[135], stage0_8[136], stage0_8[137], stage0_8[138], stage0_8[139]},
      {stage0_10[48], stage0_10[49], stage0_10[50], stage0_10[51], stage0_10[52], stage0_10[53]},
      {stage1_12[8],stage1_11[34],stage1_10[44],stage1_9[106],stage1_8[172]}
   );
   gpc606_5 gpc352 (
      {stage0_8[140], stage0_8[141], stage0_8[142], stage0_8[143], stage0_8[144], stage0_8[145]},
      {stage0_10[54], stage0_10[55], stage0_10[56], stage0_10[57], stage0_10[58], stage0_10[59]},
      {stage1_12[9],stage1_11[35],stage1_10[45],stage1_9[107],stage1_8[173]}
   );
   gpc606_5 gpc353 (
      {stage0_8[146], stage0_8[147], stage0_8[148], stage0_8[149], stage0_8[150], stage0_8[151]},
      {stage0_10[60], stage0_10[61], stage0_10[62], stage0_10[63], stage0_10[64], stage0_10[65]},
      {stage1_12[10],stage1_11[36],stage1_10[46],stage1_9[108],stage1_8[174]}
   );
   gpc606_5 gpc354 (
      {stage0_8[152], stage0_8[153], stage0_8[154], stage0_8[155], stage0_8[156], stage0_8[157]},
      {stage0_10[66], stage0_10[67], stage0_10[68], stage0_10[69], stage0_10[70], stage0_10[71]},
      {stage1_12[11],stage1_11[37],stage1_10[47],stage1_9[109],stage1_8[175]}
   );
   gpc606_5 gpc355 (
      {stage0_8[158], stage0_8[159], stage0_8[160], stage0_8[161], stage0_8[162], stage0_8[163]},
      {stage0_10[72], stage0_10[73], stage0_10[74], stage0_10[75], stage0_10[76], stage0_10[77]},
      {stage1_12[12],stage1_11[38],stage1_10[48],stage1_9[110],stage1_8[176]}
   );
   gpc606_5 gpc356 (
      {stage0_8[164], stage0_8[165], stage0_8[166], stage0_8[167], stage0_8[168], stage0_8[169]},
      {stage0_10[78], stage0_10[79], stage0_10[80], stage0_10[81], stage0_10[82], stage0_10[83]},
      {stage1_12[13],stage1_11[39],stage1_10[49],stage1_9[111],stage1_8[177]}
   );
   gpc606_5 gpc357 (
      {stage0_8[170], stage0_8[171], stage0_8[172], stage0_8[173], stage0_8[174], stage0_8[175]},
      {stage0_10[84], stage0_10[85], stage0_10[86], stage0_10[87], stage0_10[88], stage0_10[89]},
      {stage1_12[14],stage1_11[40],stage1_10[50],stage1_9[112],stage1_8[178]}
   );
   gpc606_5 gpc358 (
      {stage0_8[176], stage0_8[177], stage0_8[178], stage0_8[179], stage0_8[180], stage0_8[181]},
      {stage0_10[90], stage0_10[91], stage0_10[92], stage0_10[93], stage0_10[94], stage0_10[95]},
      {stage1_12[15],stage1_11[41],stage1_10[51],stage1_9[113],stage1_8[179]}
   );
   gpc606_5 gpc359 (
      {stage0_8[182], stage0_8[183], stage0_8[184], stage0_8[185], stage0_8[186], stage0_8[187]},
      {stage0_10[96], stage0_10[97], stage0_10[98], stage0_10[99], stage0_10[100], stage0_10[101]},
      {stage1_12[16],stage1_11[42],stage1_10[52],stage1_9[114],stage1_8[180]}
   );
   gpc606_5 gpc360 (
      {stage0_8[188], stage0_8[189], stage0_8[190], stage0_8[191], stage0_8[192], stage0_8[193]},
      {stage0_10[102], stage0_10[103], stage0_10[104], stage0_10[105], stage0_10[106], stage0_10[107]},
      {stage1_12[17],stage1_11[43],stage1_10[53],stage1_9[115],stage1_8[181]}
   );
   gpc606_5 gpc361 (
      {stage0_8[194], stage0_8[195], stage0_8[196], stage0_8[197], stage0_8[198], stage0_8[199]},
      {stage0_10[108], stage0_10[109], stage0_10[110], stage0_10[111], stage0_10[112], stage0_10[113]},
      {stage1_12[18],stage1_11[44],stage1_10[54],stage1_9[116],stage1_8[182]}
   );
   gpc606_5 gpc362 (
      {stage0_8[200], stage0_8[201], stage0_8[202], stage0_8[203], stage0_8[204], stage0_8[205]},
      {stage0_10[114], stage0_10[115], stage0_10[116], stage0_10[117], stage0_10[118], stage0_10[119]},
      {stage1_12[19],stage1_11[45],stage1_10[55],stage1_9[117],stage1_8[183]}
   );
   gpc606_5 gpc363 (
      {stage0_8[206], stage0_8[207], stage0_8[208], stage0_8[209], stage0_8[210], stage0_8[211]},
      {stage0_10[120], stage0_10[121], stage0_10[122], stage0_10[123], stage0_10[124], stage0_10[125]},
      {stage1_12[20],stage1_11[46],stage1_10[56],stage1_9[118],stage1_8[184]}
   );
   gpc606_5 gpc364 (
      {stage0_8[212], stage0_8[213], stage0_8[214], stage0_8[215], stage0_8[216], stage0_8[217]},
      {stage0_10[126], stage0_10[127], stage0_10[128], stage0_10[129], stage0_10[130], stage0_10[131]},
      {stage1_12[21],stage1_11[47],stage1_10[57],stage1_9[119],stage1_8[185]}
   );
   gpc606_5 gpc365 (
      {stage0_8[218], stage0_8[219], stage0_8[220], stage0_8[221], stage0_8[222], stage0_8[223]},
      {stage0_10[132], stage0_10[133], stage0_10[134], stage0_10[135], stage0_10[136], stage0_10[137]},
      {stage1_12[22],stage1_11[48],stage1_10[58],stage1_9[120],stage1_8[186]}
   );
   gpc606_5 gpc366 (
      {stage0_8[224], stage0_8[225], stage0_8[226], stage0_8[227], stage0_8[228], stage0_8[229]},
      {stage0_10[138], stage0_10[139], stage0_10[140], stage0_10[141], stage0_10[142], stage0_10[143]},
      {stage1_12[23],stage1_11[49],stage1_10[59],stage1_9[121],stage1_8[187]}
   );
   gpc606_5 gpc367 (
      {stage0_8[230], stage0_8[231], stage0_8[232], stage0_8[233], stage0_8[234], stage0_8[235]},
      {stage0_10[144], stage0_10[145], stage0_10[146], stage0_10[147], stage0_10[148], stage0_10[149]},
      {stage1_12[24],stage1_11[50],stage1_10[60],stage1_9[122],stage1_8[188]}
   );
   gpc606_5 gpc368 (
      {stage0_8[236], stage0_8[237], stage0_8[238], stage0_8[239], stage0_8[240], stage0_8[241]},
      {stage0_10[150], stage0_10[151], stage0_10[152], stage0_10[153], stage0_10[154], stage0_10[155]},
      {stage1_12[25],stage1_11[51],stage1_10[61],stage1_9[123],stage1_8[189]}
   );
   gpc606_5 gpc369 (
      {stage0_8[242], stage0_8[243], stage0_8[244], stage0_8[245], stage0_8[246], stage0_8[247]},
      {stage0_10[156], stage0_10[157], stage0_10[158], stage0_10[159], stage0_10[160], stage0_10[161]},
      {stage1_12[26],stage1_11[52],stage1_10[62],stage1_9[124],stage1_8[190]}
   );
   gpc606_5 gpc370 (
      {stage0_8[248], stage0_8[249], stage0_8[250], stage0_8[251], stage0_8[252], stage0_8[253]},
      {stage0_10[162], stage0_10[163], stage0_10[164], stage0_10[165], stage0_10[166], stage0_10[167]},
      {stage1_12[27],stage1_11[53],stage1_10[63],stage1_9[125],stage1_8[191]}
   );
   gpc606_5 gpc371 (
      {stage0_8[254], stage0_8[255], stage0_8[256], stage0_8[257], stage0_8[258], stage0_8[259]},
      {stage0_10[168], stage0_10[169], stage0_10[170], stage0_10[171], stage0_10[172], stage0_10[173]},
      {stage1_12[28],stage1_11[54],stage1_10[64],stage1_9[126],stage1_8[192]}
   );
   gpc606_5 gpc372 (
      {stage0_8[260], stage0_8[261], stage0_8[262], stage0_8[263], stage0_8[264], stage0_8[265]},
      {stage0_10[174], stage0_10[175], stage0_10[176], stage0_10[177], stage0_10[178], stage0_10[179]},
      {stage1_12[29],stage1_11[55],stage1_10[65],stage1_9[127],stage1_8[193]}
   );
   gpc606_5 gpc373 (
      {stage0_8[266], stage0_8[267], stage0_8[268], stage0_8[269], stage0_8[270], stage0_8[271]},
      {stage0_10[180], stage0_10[181], stage0_10[182], stage0_10[183], stage0_10[184], stage0_10[185]},
      {stage1_12[30],stage1_11[56],stage1_10[66],stage1_9[128],stage1_8[194]}
   );
   gpc606_5 gpc374 (
      {stage0_8[272], stage0_8[273], stage0_8[274], stage0_8[275], stage0_8[276], stage0_8[277]},
      {stage0_10[186], stage0_10[187], stage0_10[188], stage0_10[189], stage0_10[190], stage0_10[191]},
      {stage1_12[31],stage1_11[57],stage1_10[67],stage1_9[129],stage1_8[195]}
   );
   gpc606_5 gpc375 (
      {stage0_8[278], stage0_8[279], stage0_8[280], stage0_8[281], stage0_8[282], stage0_8[283]},
      {stage0_10[192], stage0_10[193], stage0_10[194], stage0_10[195], stage0_10[196], stage0_10[197]},
      {stage1_12[32],stage1_11[58],stage1_10[68],stage1_9[130],stage1_8[196]}
   );
   gpc606_5 gpc376 (
      {stage0_8[284], stage0_8[285], stage0_8[286], stage0_8[287], stage0_8[288], stage0_8[289]},
      {stage0_10[198], stage0_10[199], stage0_10[200], stage0_10[201], stage0_10[202], stage0_10[203]},
      {stage1_12[33],stage1_11[59],stage1_10[69],stage1_9[131],stage1_8[197]}
   );
   gpc606_5 gpc377 (
      {stage0_8[290], stage0_8[291], stage0_8[292], stage0_8[293], stage0_8[294], stage0_8[295]},
      {stage0_10[204], stage0_10[205], stage0_10[206], stage0_10[207], stage0_10[208], stage0_10[209]},
      {stage1_12[34],stage1_11[60],stage1_10[70],stage1_9[132],stage1_8[198]}
   );
   gpc606_5 gpc378 (
      {stage0_8[296], stage0_8[297], stage0_8[298], stage0_8[299], stage0_8[300], stage0_8[301]},
      {stage0_10[210], stage0_10[211], stage0_10[212], stage0_10[213], stage0_10[214], stage0_10[215]},
      {stage1_12[35],stage1_11[61],stage1_10[71],stage1_9[133],stage1_8[199]}
   );
   gpc606_5 gpc379 (
      {stage0_8[302], stage0_8[303], stage0_8[304], stage0_8[305], stage0_8[306], stage0_8[307]},
      {stage0_10[216], stage0_10[217], stage0_10[218], stage0_10[219], stage0_10[220], stage0_10[221]},
      {stage1_12[36],stage1_11[62],stage1_10[72],stage1_9[134],stage1_8[200]}
   );
   gpc606_5 gpc380 (
      {stage0_8[308], stage0_8[309], stage0_8[310], stage0_8[311], stage0_8[312], stage0_8[313]},
      {stage0_10[222], stage0_10[223], stage0_10[224], stage0_10[225], stage0_10[226], stage0_10[227]},
      {stage1_12[37],stage1_11[63],stage1_10[73],stage1_9[135],stage1_8[201]}
   );
   gpc606_5 gpc381 (
      {stage0_8[314], stage0_8[315], stage0_8[316], stage0_8[317], stage0_8[318], stage0_8[319]},
      {stage0_10[228], stage0_10[229], stage0_10[230], stage0_10[231], stage0_10[232], stage0_10[233]},
      {stage1_12[38],stage1_11[64],stage1_10[74],stage1_9[136],stage1_8[202]}
   );
   gpc606_5 gpc382 (
      {stage0_8[320], stage0_8[321], stage0_8[322], stage0_8[323], stage0_8[324], stage0_8[325]},
      {stage0_10[234], stage0_10[235], stage0_10[236], stage0_10[237], stage0_10[238], stage0_10[239]},
      {stage1_12[39],stage1_11[65],stage1_10[75],stage1_9[137],stage1_8[203]}
   );
   gpc606_5 gpc383 (
      {stage0_8[326], stage0_8[327], stage0_8[328], stage0_8[329], stage0_8[330], stage0_8[331]},
      {stage0_10[240], stage0_10[241], stage0_10[242], stage0_10[243], stage0_10[244], stage0_10[245]},
      {stage1_12[40],stage1_11[66],stage1_10[76],stage1_9[138],stage1_8[204]}
   );
   gpc615_5 gpc384 (
      {stage0_8[332], stage0_8[333], stage0_8[334], stage0_8[335], stage0_8[336]},
      {stage0_9[156]},
      {stage0_10[246], stage0_10[247], stage0_10[248], stage0_10[249], stage0_10[250], stage0_10[251]},
      {stage1_12[41],stage1_11[67],stage1_10[77],stage1_9[139],stage1_8[205]}
   );
   gpc615_5 gpc385 (
      {stage0_8[337], stage0_8[338], stage0_8[339], stage0_8[340], stage0_8[341]},
      {stage0_9[157]},
      {stage0_10[252], stage0_10[253], stage0_10[254], stage0_10[255], stage0_10[256], stage0_10[257]},
      {stage1_12[42],stage1_11[68],stage1_10[78],stage1_9[140],stage1_8[206]}
   );
   gpc615_5 gpc386 (
      {stage0_8[342], stage0_8[343], stage0_8[344], stage0_8[345], stage0_8[346]},
      {stage0_9[158]},
      {stage0_10[258], stage0_10[259], stage0_10[260], stage0_10[261], stage0_10[262], stage0_10[263]},
      {stage1_12[43],stage1_11[69],stage1_10[79],stage1_9[141],stage1_8[207]}
   );
   gpc615_5 gpc387 (
      {stage0_8[347], stage0_8[348], stage0_8[349], stage0_8[350], stage0_8[351]},
      {stage0_9[159]},
      {stage0_10[264], stage0_10[265], stage0_10[266], stage0_10[267], stage0_10[268], stage0_10[269]},
      {stage1_12[44],stage1_11[70],stage1_10[80],stage1_9[142],stage1_8[208]}
   );
   gpc615_5 gpc388 (
      {stage0_8[352], stage0_8[353], stage0_8[354], stage0_8[355], stage0_8[356]},
      {stage0_9[160]},
      {stage0_10[270], stage0_10[271], stage0_10[272], stage0_10[273], stage0_10[274], stage0_10[275]},
      {stage1_12[45],stage1_11[71],stage1_10[81],stage1_9[143],stage1_8[209]}
   );
   gpc615_5 gpc389 (
      {stage0_8[357], stage0_8[358], stage0_8[359], stage0_8[360], stage0_8[361]},
      {stage0_9[161]},
      {stage0_10[276], stage0_10[277], stage0_10[278], stage0_10[279], stage0_10[280], stage0_10[281]},
      {stage1_12[46],stage1_11[72],stage1_10[82],stage1_9[144],stage1_8[210]}
   );
   gpc615_5 gpc390 (
      {stage0_8[362], stage0_8[363], stage0_8[364], stage0_8[365], stage0_8[366]},
      {stage0_9[162]},
      {stage0_10[282], stage0_10[283], stage0_10[284], stage0_10[285], stage0_10[286], stage0_10[287]},
      {stage1_12[47],stage1_11[73],stage1_10[83],stage1_9[145],stage1_8[211]}
   );
   gpc615_5 gpc391 (
      {stage0_8[367], stage0_8[368], stage0_8[369], stage0_8[370], stage0_8[371]},
      {stage0_9[163]},
      {stage0_10[288], stage0_10[289], stage0_10[290], stage0_10[291], stage0_10[292], stage0_10[293]},
      {stage1_12[48],stage1_11[74],stage1_10[84],stage1_9[146],stage1_8[212]}
   );
   gpc615_5 gpc392 (
      {stage0_8[372], stage0_8[373], stage0_8[374], stage0_8[375], stage0_8[376]},
      {stage0_9[164]},
      {stage0_10[294], stage0_10[295], stage0_10[296], stage0_10[297], stage0_10[298], stage0_10[299]},
      {stage1_12[49],stage1_11[75],stage1_10[85],stage1_9[147],stage1_8[213]}
   );
   gpc606_5 gpc393 (
      {stage0_9[165], stage0_9[166], stage0_9[167], stage0_9[168], stage0_9[169], stage0_9[170]},
      {stage0_11[0], stage0_11[1], stage0_11[2], stage0_11[3], stage0_11[4], stage0_11[5]},
      {stage1_13[0],stage1_12[50],stage1_11[76],stage1_10[86],stage1_9[148]}
   );
   gpc606_5 gpc394 (
      {stage0_9[171], stage0_9[172], stage0_9[173], stage0_9[174], stage0_9[175], stage0_9[176]},
      {stage0_11[6], stage0_11[7], stage0_11[8], stage0_11[9], stage0_11[10], stage0_11[11]},
      {stage1_13[1],stage1_12[51],stage1_11[77],stage1_10[87],stage1_9[149]}
   );
   gpc606_5 gpc395 (
      {stage0_9[177], stage0_9[178], stage0_9[179], stage0_9[180], stage0_9[181], stage0_9[182]},
      {stage0_11[12], stage0_11[13], stage0_11[14], stage0_11[15], stage0_11[16], stage0_11[17]},
      {stage1_13[2],stage1_12[52],stage1_11[78],stage1_10[88],stage1_9[150]}
   );
   gpc606_5 gpc396 (
      {stage0_9[183], stage0_9[184], stage0_9[185], stage0_9[186], stage0_9[187], stage0_9[188]},
      {stage0_11[18], stage0_11[19], stage0_11[20], stage0_11[21], stage0_11[22], stage0_11[23]},
      {stage1_13[3],stage1_12[53],stage1_11[79],stage1_10[89],stage1_9[151]}
   );
   gpc606_5 gpc397 (
      {stage0_9[189], stage0_9[190], stage0_9[191], stage0_9[192], stage0_9[193], stage0_9[194]},
      {stage0_11[24], stage0_11[25], stage0_11[26], stage0_11[27], stage0_11[28], stage0_11[29]},
      {stage1_13[4],stage1_12[54],stage1_11[80],stage1_10[90],stage1_9[152]}
   );
   gpc606_5 gpc398 (
      {stage0_9[195], stage0_9[196], stage0_9[197], stage0_9[198], stage0_9[199], stage0_9[200]},
      {stage0_11[30], stage0_11[31], stage0_11[32], stage0_11[33], stage0_11[34], stage0_11[35]},
      {stage1_13[5],stage1_12[55],stage1_11[81],stage1_10[91],stage1_9[153]}
   );
   gpc606_5 gpc399 (
      {stage0_9[201], stage0_9[202], stage0_9[203], stage0_9[204], stage0_9[205], stage0_9[206]},
      {stage0_11[36], stage0_11[37], stage0_11[38], stage0_11[39], stage0_11[40], stage0_11[41]},
      {stage1_13[6],stage1_12[56],stage1_11[82],stage1_10[92],stage1_9[154]}
   );
   gpc606_5 gpc400 (
      {stage0_9[207], stage0_9[208], stage0_9[209], stage0_9[210], stage0_9[211], stage0_9[212]},
      {stage0_11[42], stage0_11[43], stage0_11[44], stage0_11[45], stage0_11[46], stage0_11[47]},
      {stage1_13[7],stage1_12[57],stage1_11[83],stage1_10[93],stage1_9[155]}
   );
   gpc606_5 gpc401 (
      {stage0_9[213], stage0_9[214], stage0_9[215], stage0_9[216], stage0_9[217], stage0_9[218]},
      {stage0_11[48], stage0_11[49], stage0_11[50], stage0_11[51], stage0_11[52], stage0_11[53]},
      {stage1_13[8],stage1_12[58],stage1_11[84],stage1_10[94],stage1_9[156]}
   );
   gpc606_5 gpc402 (
      {stage0_9[219], stage0_9[220], stage0_9[221], stage0_9[222], stage0_9[223], stage0_9[224]},
      {stage0_11[54], stage0_11[55], stage0_11[56], stage0_11[57], stage0_11[58], stage0_11[59]},
      {stage1_13[9],stage1_12[59],stage1_11[85],stage1_10[95],stage1_9[157]}
   );
   gpc606_5 gpc403 (
      {stage0_9[225], stage0_9[226], stage0_9[227], stage0_9[228], stage0_9[229], stage0_9[230]},
      {stage0_11[60], stage0_11[61], stage0_11[62], stage0_11[63], stage0_11[64], stage0_11[65]},
      {stage1_13[10],stage1_12[60],stage1_11[86],stage1_10[96],stage1_9[158]}
   );
   gpc606_5 gpc404 (
      {stage0_9[231], stage0_9[232], stage0_9[233], stage0_9[234], stage0_9[235], stage0_9[236]},
      {stage0_11[66], stage0_11[67], stage0_11[68], stage0_11[69], stage0_11[70], stage0_11[71]},
      {stage1_13[11],stage1_12[61],stage1_11[87],stage1_10[97],stage1_9[159]}
   );
   gpc606_5 gpc405 (
      {stage0_9[237], stage0_9[238], stage0_9[239], stage0_9[240], stage0_9[241], stage0_9[242]},
      {stage0_11[72], stage0_11[73], stage0_11[74], stage0_11[75], stage0_11[76], stage0_11[77]},
      {stage1_13[12],stage1_12[62],stage1_11[88],stage1_10[98],stage1_9[160]}
   );
   gpc606_5 gpc406 (
      {stage0_9[243], stage0_9[244], stage0_9[245], stage0_9[246], stage0_9[247], stage0_9[248]},
      {stage0_11[78], stage0_11[79], stage0_11[80], stage0_11[81], stage0_11[82], stage0_11[83]},
      {stage1_13[13],stage1_12[63],stage1_11[89],stage1_10[99],stage1_9[161]}
   );
   gpc606_5 gpc407 (
      {stage0_9[249], stage0_9[250], stage0_9[251], stage0_9[252], stage0_9[253], stage0_9[254]},
      {stage0_11[84], stage0_11[85], stage0_11[86], stage0_11[87], stage0_11[88], stage0_11[89]},
      {stage1_13[14],stage1_12[64],stage1_11[90],stage1_10[100],stage1_9[162]}
   );
   gpc606_5 gpc408 (
      {stage0_9[255], stage0_9[256], stage0_9[257], stage0_9[258], stage0_9[259], stage0_9[260]},
      {stage0_11[90], stage0_11[91], stage0_11[92], stage0_11[93], stage0_11[94], stage0_11[95]},
      {stage1_13[15],stage1_12[65],stage1_11[91],stage1_10[101],stage1_9[163]}
   );
   gpc606_5 gpc409 (
      {stage0_9[261], stage0_9[262], stage0_9[263], stage0_9[264], stage0_9[265], stage0_9[266]},
      {stage0_11[96], stage0_11[97], stage0_11[98], stage0_11[99], stage0_11[100], stage0_11[101]},
      {stage1_13[16],stage1_12[66],stage1_11[92],stage1_10[102],stage1_9[164]}
   );
   gpc606_5 gpc410 (
      {stage0_9[267], stage0_9[268], stage0_9[269], stage0_9[270], stage0_9[271], stage0_9[272]},
      {stage0_11[102], stage0_11[103], stage0_11[104], stage0_11[105], stage0_11[106], stage0_11[107]},
      {stage1_13[17],stage1_12[67],stage1_11[93],stage1_10[103],stage1_9[165]}
   );
   gpc606_5 gpc411 (
      {stage0_9[273], stage0_9[274], stage0_9[275], stage0_9[276], stage0_9[277], stage0_9[278]},
      {stage0_11[108], stage0_11[109], stage0_11[110], stage0_11[111], stage0_11[112], stage0_11[113]},
      {stage1_13[18],stage1_12[68],stage1_11[94],stage1_10[104],stage1_9[166]}
   );
   gpc606_5 gpc412 (
      {stage0_9[279], stage0_9[280], stage0_9[281], stage0_9[282], stage0_9[283], stage0_9[284]},
      {stage0_11[114], stage0_11[115], stage0_11[116], stage0_11[117], stage0_11[118], stage0_11[119]},
      {stage1_13[19],stage1_12[69],stage1_11[95],stage1_10[105],stage1_9[167]}
   );
   gpc606_5 gpc413 (
      {stage0_9[285], stage0_9[286], stage0_9[287], stage0_9[288], stage0_9[289], stage0_9[290]},
      {stage0_11[120], stage0_11[121], stage0_11[122], stage0_11[123], stage0_11[124], stage0_11[125]},
      {stage1_13[20],stage1_12[70],stage1_11[96],stage1_10[106],stage1_9[168]}
   );
   gpc606_5 gpc414 (
      {stage0_9[291], stage0_9[292], stage0_9[293], stage0_9[294], stage0_9[295], stage0_9[296]},
      {stage0_11[126], stage0_11[127], stage0_11[128], stage0_11[129], stage0_11[130], stage0_11[131]},
      {stage1_13[21],stage1_12[71],stage1_11[97],stage1_10[107],stage1_9[169]}
   );
   gpc606_5 gpc415 (
      {stage0_9[297], stage0_9[298], stage0_9[299], stage0_9[300], stage0_9[301], stage0_9[302]},
      {stage0_11[132], stage0_11[133], stage0_11[134], stage0_11[135], stage0_11[136], stage0_11[137]},
      {stage1_13[22],stage1_12[72],stage1_11[98],stage1_10[108],stage1_9[170]}
   );
   gpc606_5 gpc416 (
      {stage0_9[303], stage0_9[304], stage0_9[305], stage0_9[306], stage0_9[307], stage0_9[308]},
      {stage0_11[138], stage0_11[139], stage0_11[140], stage0_11[141], stage0_11[142], stage0_11[143]},
      {stage1_13[23],stage1_12[73],stage1_11[99],stage1_10[109],stage1_9[171]}
   );
   gpc606_5 gpc417 (
      {stage0_9[309], stage0_9[310], stage0_9[311], stage0_9[312], stage0_9[313], stage0_9[314]},
      {stage0_11[144], stage0_11[145], stage0_11[146], stage0_11[147], stage0_11[148], stage0_11[149]},
      {stage1_13[24],stage1_12[74],stage1_11[100],stage1_10[110],stage1_9[172]}
   );
   gpc606_5 gpc418 (
      {stage0_9[315], stage0_9[316], stage0_9[317], stage0_9[318], stage0_9[319], stage0_9[320]},
      {stage0_11[150], stage0_11[151], stage0_11[152], stage0_11[153], stage0_11[154], stage0_11[155]},
      {stage1_13[25],stage1_12[75],stage1_11[101],stage1_10[111],stage1_9[173]}
   );
   gpc606_5 gpc419 (
      {stage0_9[321], stage0_9[322], stage0_9[323], stage0_9[324], stage0_9[325], stage0_9[326]},
      {stage0_11[156], stage0_11[157], stage0_11[158], stage0_11[159], stage0_11[160], stage0_11[161]},
      {stage1_13[26],stage1_12[76],stage1_11[102],stage1_10[112],stage1_9[174]}
   );
   gpc606_5 gpc420 (
      {stage0_9[327], stage0_9[328], stage0_9[329], stage0_9[330], stage0_9[331], stage0_9[332]},
      {stage0_11[162], stage0_11[163], stage0_11[164], stage0_11[165], stage0_11[166], stage0_11[167]},
      {stage1_13[27],stage1_12[77],stage1_11[103],stage1_10[113],stage1_9[175]}
   );
   gpc606_5 gpc421 (
      {stage0_9[333], stage0_9[334], stage0_9[335], stage0_9[336], stage0_9[337], stage0_9[338]},
      {stage0_11[168], stage0_11[169], stage0_11[170], stage0_11[171], stage0_11[172], stage0_11[173]},
      {stage1_13[28],stage1_12[78],stage1_11[104],stage1_10[114],stage1_9[176]}
   );
   gpc606_5 gpc422 (
      {stage0_9[339], stage0_9[340], stage0_9[341], stage0_9[342], stage0_9[343], stage0_9[344]},
      {stage0_11[174], stage0_11[175], stage0_11[176], stage0_11[177], stage0_11[178], stage0_11[179]},
      {stage1_13[29],stage1_12[79],stage1_11[105],stage1_10[115],stage1_9[177]}
   );
   gpc606_5 gpc423 (
      {stage0_9[345], stage0_9[346], stage0_9[347], stage0_9[348], stage0_9[349], stage0_9[350]},
      {stage0_11[180], stage0_11[181], stage0_11[182], stage0_11[183], stage0_11[184], stage0_11[185]},
      {stage1_13[30],stage1_12[80],stage1_11[106],stage1_10[116],stage1_9[178]}
   );
   gpc606_5 gpc424 (
      {stage0_9[351], stage0_9[352], stage0_9[353], stage0_9[354], stage0_9[355], stage0_9[356]},
      {stage0_11[186], stage0_11[187], stage0_11[188], stage0_11[189], stage0_11[190], stage0_11[191]},
      {stage1_13[31],stage1_12[81],stage1_11[107],stage1_10[117],stage1_9[179]}
   );
   gpc606_5 gpc425 (
      {stage0_9[357], stage0_9[358], stage0_9[359], stage0_9[360], stage0_9[361], stage0_9[362]},
      {stage0_11[192], stage0_11[193], stage0_11[194], stage0_11[195], stage0_11[196], stage0_11[197]},
      {stage1_13[32],stage1_12[82],stage1_11[108],stage1_10[118],stage1_9[180]}
   );
   gpc606_5 gpc426 (
      {stage0_9[363], stage0_9[364], stage0_9[365], stage0_9[366], stage0_9[367], stage0_9[368]},
      {stage0_11[198], stage0_11[199], stage0_11[200], stage0_11[201], stage0_11[202], stage0_11[203]},
      {stage1_13[33],stage1_12[83],stage1_11[109],stage1_10[119],stage1_9[181]}
   );
   gpc606_5 gpc427 (
      {stage0_9[369], stage0_9[370], stage0_9[371], stage0_9[372], stage0_9[373], stage0_9[374]},
      {stage0_11[204], stage0_11[205], stage0_11[206], stage0_11[207], stage0_11[208], stage0_11[209]},
      {stage1_13[34],stage1_12[84],stage1_11[110],stage1_10[120],stage1_9[182]}
   );
   gpc606_5 gpc428 (
      {stage0_9[375], stage0_9[376], stage0_9[377], stage0_9[378], stage0_9[379], stage0_9[380]},
      {stage0_11[210], stage0_11[211], stage0_11[212], stage0_11[213], stage0_11[214], stage0_11[215]},
      {stage1_13[35],stage1_12[85],stage1_11[111],stage1_10[121],stage1_9[183]}
   );
   gpc606_5 gpc429 (
      {stage0_9[381], stage0_9[382], stage0_9[383], stage0_9[384], stage0_9[385], stage0_9[386]},
      {stage0_11[216], stage0_11[217], stage0_11[218], stage0_11[219], stage0_11[220], stage0_11[221]},
      {stage1_13[36],stage1_12[86],stage1_11[112],stage1_10[122],stage1_9[184]}
   );
   gpc606_5 gpc430 (
      {stage0_9[387], stage0_9[388], stage0_9[389], stage0_9[390], stage0_9[391], stage0_9[392]},
      {stage0_11[222], stage0_11[223], stage0_11[224], stage0_11[225], stage0_11[226], stage0_11[227]},
      {stage1_13[37],stage1_12[87],stage1_11[113],stage1_10[123],stage1_9[185]}
   );
   gpc606_5 gpc431 (
      {stage0_9[393], stage0_9[394], stage0_9[395], stage0_9[396], stage0_9[397], stage0_9[398]},
      {stage0_11[228], stage0_11[229], stage0_11[230], stage0_11[231], stage0_11[232], stage0_11[233]},
      {stage1_13[38],stage1_12[88],stage1_11[114],stage1_10[124],stage1_9[186]}
   );
   gpc615_5 gpc432 (
      {stage0_9[399], stage0_9[400], stage0_9[401], stage0_9[402], stage0_9[403]},
      {stage0_10[300]},
      {stage0_11[234], stage0_11[235], stage0_11[236], stage0_11[237], stage0_11[238], stage0_11[239]},
      {stage1_13[39],stage1_12[89],stage1_11[115],stage1_10[125],stage1_9[187]}
   );
   gpc615_5 gpc433 (
      {stage0_9[404], stage0_9[405], stage0_9[406], stage0_9[407], stage0_9[408]},
      {stage0_10[301]},
      {stage0_11[240], stage0_11[241], stage0_11[242], stage0_11[243], stage0_11[244], stage0_11[245]},
      {stage1_13[40],stage1_12[90],stage1_11[116],stage1_10[126],stage1_9[188]}
   );
   gpc615_5 gpc434 (
      {stage0_9[409], stage0_9[410], stage0_9[411], stage0_9[412], stage0_9[413]},
      {stage0_10[302]},
      {stage0_11[246], stage0_11[247], stage0_11[248], stage0_11[249], stage0_11[250], stage0_11[251]},
      {stage1_13[41],stage1_12[91],stage1_11[117],stage1_10[127],stage1_9[189]}
   );
   gpc615_5 gpc435 (
      {stage0_9[414], stage0_9[415], stage0_9[416], stage0_9[417], stage0_9[418]},
      {stage0_10[303]},
      {stage0_11[252], stage0_11[253], stage0_11[254], stage0_11[255], stage0_11[256], stage0_11[257]},
      {stage1_13[42],stage1_12[92],stage1_11[118],stage1_10[128],stage1_9[190]}
   );
   gpc615_5 gpc436 (
      {stage0_9[419], stage0_9[420], stage0_9[421], stage0_9[422], stage0_9[423]},
      {stage0_10[304]},
      {stage0_11[258], stage0_11[259], stage0_11[260], stage0_11[261], stage0_11[262], stage0_11[263]},
      {stage1_13[43],stage1_12[93],stage1_11[119],stage1_10[129],stage1_9[191]}
   );
   gpc615_5 gpc437 (
      {stage0_9[424], stage0_9[425], stage0_9[426], stage0_9[427], stage0_9[428]},
      {stage0_10[305]},
      {stage0_11[264], stage0_11[265], stage0_11[266], stage0_11[267], stage0_11[268], stage0_11[269]},
      {stage1_13[44],stage1_12[94],stage1_11[120],stage1_10[130],stage1_9[192]}
   );
   gpc615_5 gpc438 (
      {stage0_9[429], stage0_9[430], stage0_9[431], stage0_9[432], stage0_9[433]},
      {stage0_10[306]},
      {stage0_11[270], stage0_11[271], stage0_11[272], stage0_11[273], stage0_11[274], stage0_11[275]},
      {stage1_13[45],stage1_12[95],stage1_11[121],stage1_10[131],stage1_9[193]}
   );
   gpc615_5 gpc439 (
      {stage0_9[434], stage0_9[435], stage0_9[436], stage0_9[437], stage0_9[438]},
      {stage0_10[307]},
      {stage0_11[276], stage0_11[277], stage0_11[278], stage0_11[279], stage0_11[280], stage0_11[281]},
      {stage1_13[46],stage1_12[96],stage1_11[122],stage1_10[132],stage1_9[194]}
   );
   gpc615_5 gpc440 (
      {stage0_9[439], stage0_9[440], stage0_9[441], stage0_9[442], stage0_9[443]},
      {stage0_10[308]},
      {stage0_11[282], stage0_11[283], stage0_11[284], stage0_11[285], stage0_11[286], stage0_11[287]},
      {stage1_13[47],stage1_12[97],stage1_11[123],stage1_10[133],stage1_9[195]}
   );
   gpc615_5 gpc441 (
      {stage0_9[444], stage0_9[445], stage0_9[446], stage0_9[447], stage0_9[448]},
      {stage0_10[309]},
      {stage0_11[288], stage0_11[289], stage0_11[290], stage0_11[291], stage0_11[292], stage0_11[293]},
      {stage1_13[48],stage1_12[98],stage1_11[124],stage1_10[134],stage1_9[196]}
   );
   gpc615_5 gpc442 (
      {stage0_9[449], stage0_9[450], stage0_9[451], stage0_9[452], stage0_9[453]},
      {stage0_10[310]},
      {stage0_11[294], stage0_11[295], stage0_11[296], stage0_11[297], stage0_11[298], stage0_11[299]},
      {stage1_13[49],stage1_12[99],stage1_11[125],stage1_10[135],stage1_9[197]}
   );
   gpc615_5 gpc443 (
      {stage0_9[454], stage0_9[455], stage0_9[456], stage0_9[457], stage0_9[458]},
      {stage0_10[311]},
      {stage0_11[300], stage0_11[301], stage0_11[302], stage0_11[303], stage0_11[304], stage0_11[305]},
      {stage1_13[50],stage1_12[100],stage1_11[126],stage1_10[136],stage1_9[198]}
   );
   gpc615_5 gpc444 (
      {stage0_9[459], stage0_9[460], stage0_9[461], stage0_9[462], stage0_9[463]},
      {stage0_10[312]},
      {stage0_11[306], stage0_11[307], stage0_11[308], stage0_11[309], stage0_11[310], stage0_11[311]},
      {stage1_13[51],stage1_12[101],stage1_11[127],stage1_10[137],stage1_9[199]}
   );
   gpc615_5 gpc445 (
      {stage0_9[464], stage0_9[465], stage0_9[466], stage0_9[467], stage0_9[468]},
      {stage0_10[313]},
      {stage0_11[312], stage0_11[313], stage0_11[314], stage0_11[315], stage0_11[316], stage0_11[317]},
      {stage1_13[52],stage1_12[102],stage1_11[128],stage1_10[138],stage1_9[200]}
   );
   gpc615_5 gpc446 (
      {stage0_9[469], stage0_9[470], stage0_9[471], stage0_9[472], stage0_9[473]},
      {stage0_10[314]},
      {stage0_11[318], stage0_11[319], stage0_11[320], stage0_11[321], stage0_11[322], stage0_11[323]},
      {stage1_13[53],stage1_12[103],stage1_11[129],stage1_10[139],stage1_9[201]}
   );
   gpc615_5 gpc447 (
      {stage0_9[474], stage0_9[475], stage0_9[476], stage0_9[477], stage0_9[478]},
      {stage0_10[315]},
      {stage0_11[324], stage0_11[325], stage0_11[326], stage0_11[327], stage0_11[328], stage0_11[329]},
      {stage1_13[54],stage1_12[104],stage1_11[130],stage1_10[140],stage1_9[202]}
   );
   gpc615_5 gpc448 (
      {stage0_9[479], stage0_9[480], stage0_9[481], stage0_9[482], stage0_9[483]},
      {stage0_10[316]},
      {stage0_11[330], stage0_11[331], stage0_11[332], stage0_11[333], stage0_11[334], stage0_11[335]},
      {stage1_13[55],stage1_12[105],stage1_11[131],stage1_10[141],stage1_9[203]}
   );
   gpc615_5 gpc449 (
      {stage0_9[484], stage0_9[485], stage0_9[486], stage0_9[487], stage0_9[488]},
      {stage0_10[317]},
      {stage0_11[336], stage0_11[337], stage0_11[338], stage0_11[339], stage0_11[340], stage0_11[341]},
      {stage1_13[56],stage1_12[106],stage1_11[132],stage1_10[142],stage1_9[204]}
   );
   gpc615_5 gpc450 (
      {stage0_9[489], stage0_9[490], stage0_9[491], stage0_9[492], stage0_9[493]},
      {stage0_10[318]},
      {stage0_11[342], stage0_11[343], stage0_11[344], stage0_11[345], stage0_11[346], stage0_11[347]},
      {stage1_13[57],stage1_12[107],stage1_11[133],stage1_10[143],stage1_9[205]}
   );
   gpc615_5 gpc451 (
      {stage0_9[494], stage0_9[495], stage0_9[496], stage0_9[497], stage0_9[498]},
      {stage0_10[319]},
      {stage0_11[348], stage0_11[349], stage0_11[350], stage0_11[351], stage0_11[352], stage0_11[353]},
      {stage1_13[58],stage1_12[108],stage1_11[134],stage1_10[144],stage1_9[206]}
   );
   gpc615_5 gpc452 (
      {stage0_9[499], stage0_9[500], stage0_9[501], stage0_9[502], stage0_9[503]},
      {stage0_10[320]},
      {stage0_11[354], stage0_11[355], stage0_11[356], stage0_11[357], stage0_11[358], stage0_11[359]},
      {stage1_13[59],stage1_12[109],stage1_11[135],stage1_10[145],stage1_9[207]}
   );
   gpc615_5 gpc453 (
      {stage0_9[504], stage0_9[505], stage0_9[506], stage0_9[507], stage0_9[508]},
      {stage0_10[321]},
      {stage0_11[360], stage0_11[361], stage0_11[362], stage0_11[363], stage0_11[364], stage0_11[365]},
      {stage1_13[60],stage1_12[110],stage1_11[136],stage1_10[146],stage1_9[208]}
   );
   gpc606_5 gpc454 (
      {stage0_10[322], stage0_10[323], stage0_10[324], stage0_10[325], stage0_10[326], stage0_10[327]},
      {stage0_12[0], stage0_12[1], stage0_12[2], stage0_12[3], stage0_12[4], stage0_12[5]},
      {stage1_14[0],stage1_13[61],stage1_12[111],stage1_11[137],stage1_10[147]}
   );
   gpc606_5 gpc455 (
      {stage0_10[328], stage0_10[329], stage0_10[330], stage0_10[331], stage0_10[332], stage0_10[333]},
      {stage0_12[6], stage0_12[7], stage0_12[8], stage0_12[9], stage0_12[10], stage0_12[11]},
      {stage1_14[1],stage1_13[62],stage1_12[112],stage1_11[138],stage1_10[148]}
   );
   gpc606_5 gpc456 (
      {stage0_10[334], stage0_10[335], stage0_10[336], stage0_10[337], stage0_10[338], stage0_10[339]},
      {stage0_12[12], stage0_12[13], stage0_12[14], stage0_12[15], stage0_12[16], stage0_12[17]},
      {stage1_14[2],stage1_13[63],stage1_12[113],stage1_11[139],stage1_10[149]}
   );
   gpc606_5 gpc457 (
      {stage0_10[340], stage0_10[341], stage0_10[342], stage0_10[343], stage0_10[344], stage0_10[345]},
      {stage0_12[18], stage0_12[19], stage0_12[20], stage0_12[21], stage0_12[22], stage0_12[23]},
      {stage1_14[3],stage1_13[64],stage1_12[114],stage1_11[140],stage1_10[150]}
   );
   gpc606_5 gpc458 (
      {stage0_10[346], stage0_10[347], stage0_10[348], stage0_10[349], stage0_10[350], stage0_10[351]},
      {stage0_12[24], stage0_12[25], stage0_12[26], stage0_12[27], stage0_12[28], stage0_12[29]},
      {stage1_14[4],stage1_13[65],stage1_12[115],stage1_11[141],stage1_10[151]}
   );
   gpc606_5 gpc459 (
      {stage0_10[352], stage0_10[353], stage0_10[354], stage0_10[355], stage0_10[356], stage0_10[357]},
      {stage0_12[30], stage0_12[31], stage0_12[32], stage0_12[33], stage0_12[34], stage0_12[35]},
      {stage1_14[5],stage1_13[66],stage1_12[116],stage1_11[142],stage1_10[152]}
   );
   gpc606_5 gpc460 (
      {stage0_10[358], stage0_10[359], stage0_10[360], stage0_10[361], stage0_10[362], stage0_10[363]},
      {stage0_12[36], stage0_12[37], stage0_12[38], stage0_12[39], stage0_12[40], stage0_12[41]},
      {stage1_14[6],stage1_13[67],stage1_12[117],stage1_11[143],stage1_10[153]}
   );
   gpc606_5 gpc461 (
      {stage0_10[364], stage0_10[365], stage0_10[366], stage0_10[367], stage0_10[368], stage0_10[369]},
      {stage0_12[42], stage0_12[43], stage0_12[44], stage0_12[45], stage0_12[46], stage0_12[47]},
      {stage1_14[7],stage1_13[68],stage1_12[118],stage1_11[144],stage1_10[154]}
   );
   gpc606_5 gpc462 (
      {stage0_10[370], stage0_10[371], stage0_10[372], stage0_10[373], stage0_10[374], stage0_10[375]},
      {stage0_12[48], stage0_12[49], stage0_12[50], stage0_12[51], stage0_12[52], stage0_12[53]},
      {stage1_14[8],stage1_13[69],stage1_12[119],stage1_11[145],stage1_10[155]}
   );
   gpc606_5 gpc463 (
      {stage0_10[376], stage0_10[377], stage0_10[378], stage0_10[379], stage0_10[380], stage0_10[381]},
      {stage0_12[54], stage0_12[55], stage0_12[56], stage0_12[57], stage0_12[58], stage0_12[59]},
      {stage1_14[9],stage1_13[70],stage1_12[120],stage1_11[146],stage1_10[156]}
   );
   gpc606_5 gpc464 (
      {stage0_10[382], stage0_10[383], stage0_10[384], stage0_10[385], stage0_10[386], stage0_10[387]},
      {stage0_12[60], stage0_12[61], stage0_12[62], stage0_12[63], stage0_12[64], stage0_12[65]},
      {stage1_14[10],stage1_13[71],stage1_12[121],stage1_11[147],stage1_10[157]}
   );
   gpc606_5 gpc465 (
      {stage0_10[388], stage0_10[389], stage0_10[390], stage0_10[391], stage0_10[392], stage0_10[393]},
      {stage0_12[66], stage0_12[67], stage0_12[68], stage0_12[69], stage0_12[70], stage0_12[71]},
      {stage1_14[11],stage1_13[72],stage1_12[122],stage1_11[148],stage1_10[158]}
   );
   gpc606_5 gpc466 (
      {stage0_10[394], stage0_10[395], stage0_10[396], stage0_10[397], stage0_10[398], stage0_10[399]},
      {stage0_12[72], stage0_12[73], stage0_12[74], stage0_12[75], stage0_12[76], stage0_12[77]},
      {stage1_14[12],stage1_13[73],stage1_12[123],stage1_11[149],stage1_10[159]}
   );
   gpc606_5 gpc467 (
      {stage0_10[400], stage0_10[401], stage0_10[402], stage0_10[403], stage0_10[404], stage0_10[405]},
      {stage0_12[78], stage0_12[79], stage0_12[80], stage0_12[81], stage0_12[82], stage0_12[83]},
      {stage1_14[13],stage1_13[74],stage1_12[124],stage1_11[150],stage1_10[160]}
   );
   gpc606_5 gpc468 (
      {stage0_10[406], stage0_10[407], stage0_10[408], stage0_10[409], stage0_10[410], stage0_10[411]},
      {stage0_12[84], stage0_12[85], stage0_12[86], stage0_12[87], stage0_12[88], stage0_12[89]},
      {stage1_14[14],stage1_13[75],stage1_12[125],stage1_11[151],stage1_10[161]}
   );
   gpc615_5 gpc469 (
      {stage0_10[412], stage0_10[413], stage0_10[414], stage0_10[415], stage0_10[416]},
      {stage0_11[366]},
      {stage0_12[90], stage0_12[91], stage0_12[92], stage0_12[93], stage0_12[94], stage0_12[95]},
      {stage1_14[15],stage1_13[76],stage1_12[126],stage1_11[152],stage1_10[162]}
   );
   gpc615_5 gpc470 (
      {stage0_10[417], stage0_10[418], stage0_10[419], stage0_10[420], stage0_10[421]},
      {stage0_11[367]},
      {stage0_12[96], stage0_12[97], stage0_12[98], stage0_12[99], stage0_12[100], stage0_12[101]},
      {stage1_14[16],stage1_13[77],stage1_12[127],stage1_11[153],stage1_10[163]}
   );
   gpc615_5 gpc471 (
      {stage0_10[422], stage0_10[423], stage0_10[424], stage0_10[425], stage0_10[426]},
      {stage0_11[368]},
      {stage0_12[102], stage0_12[103], stage0_12[104], stage0_12[105], stage0_12[106], stage0_12[107]},
      {stage1_14[17],stage1_13[78],stage1_12[128],stage1_11[154],stage1_10[164]}
   );
   gpc615_5 gpc472 (
      {stage0_10[427], stage0_10[428], stage0_10[429], stage0_10[430], stage0_10[431]},
      {stage0_11[369]},
      {stage0_12[108], stage0_12[109], stage0_12[110], stage0_12[111], stage0_12[112], stage0_12[113]},
      {stage1_14[18],stage1_13[79],stage1_12[129],stage1_11[155],stage1_10[165]}
   );
   gpc615_5 gpc473 (
      {stage0_10[432], stage0_10[433], stage0_10[434], stage0_10[435], stage0_10[436]},
      {stage0_11[370]},
      {stage0_12[114], stage0_12[115], stage0_12[116], stage0_12[117], stage0_12[118], stage0_12[119]},
      {stage1_14[19],stage1_13[80],stage1_12[130],stage1_11[156],stage1_10[166]}
   );
   gpc615_5 gpc474 (
      {stage0_10[437], stage0_10[438], stage0_10[439], stage0_10[440], stage0_10[441]},
      {stage0_11[371]},
      {stage0_12[120], stage0_12[121], stage0_12[122], stage0_12[123], stage0_12[124], stage0_12[125]},
      {stage1_14[20],stage1_13[81],stage1_12[131],stage1_11[157],stage1_10[167]}
   );
   gpc615_5 gpc475 (
      {stage0_10[442], stage0_10[443], stage0_10[444], stage0_10[445], stage0_10[446]},
      {stage0_11[372]},
      {stage0_12[126], stage0_12[127], stage0_12[128], stage0_12[129], stage0_12[130], stage0_12[131]},
      {stage1_14[21],stage1_13[82],stage1_12[132],stage1_11[158],stage1_10[168]}
   );
   gpc615_5 gpc476 (
      {stage0_10[447], stage0_10[448], stage0_10[449], stage0_10[450], stage0_10[451]},
      {stage0_11[373]},
      {stage0_12[132], stage0_12[133], stage0_12[134], stage0_12[135], stage0_12[136], stage0_12[137]},
      {stage1_14[22],stage1_13[83],stage1_12[133],stage1_11[159],stage1_10[169]}
   );
   gpc615_5 gpc477 (
      {stage0_10[452], stage0_10[453], stage0_10[454], stage0_10[455], stage0_10[456]},
      {stage0_11[374]},
      {stage0_12[138], stage0_12[139], stage0_12[140], stage0_12[141], stage0_12[142], stage0_12[143]},
      {stage1_14[23],stage1_13[84],stage1_12[134],stage1_11[160],stage1_10[170]}
   );
   gpc615_5 gpc478 (
      {stage0_10[457], stage0_10[458], stage0_10[459], stage0_10[460], stage0_10[461]},
      {stage0_11[375]},
      {stage0_12[144], stage0_12[145], stage0_12[146], stage0_12[147], stage0_12[148], stage0_12[149]},
      {stage1_14[24],stage1_13[85],stage1_12[135],stage1_11[161],stage1_10[171]}
   );
   gpc615_5 gpc479 (
      {stage0_10[462], stage0_10[463], stage0_10[464], stage0_10[465], stage0_10[466]},
      {stage0_11[376]},
      {stage0_12[150], stage0_12[151], stage0_12[152], stage0_12[153], stage0_12[154], stage0_12[155]},
      {stage1_14[25],stage1_13[86],stage1_12[136],stage1_11[162],stage1_10[172]}
   );
   gpc615_5 gpc480 (
      {stage0_10[467], stage0_10[468], stage0_10[469], stage0_10[470], stage0_10[471]},
      {stage0_11[377]},
      {stage0_12[156], stage0_12[157], stage0_12[158], stage0_12[159], stage0_12[160], stage0_12[161]},
      {stage1_14[26],stage1_13[87],stage1_12[137],stage1_11[163],stage1_10[173]}
   );
   gpc615_5 gpc481 (
      {stage0_10[472], stage0_10[473], stage0_10[474], stage0_10[475], stage0_10[476]},
      {stage0_11[378]},
      {stage0_12[162], stage0_12[163], stage0_12[164], stage0_12[165], stage0_12[166], stage0_12[167]},
      {stage1_14[27],stage1_13[88],stage1_12[138],stage1_11[164],stage1_10[174]}
   );
   gpc615_5 gpc482 (
      {stage0_10[477], stage0_10[478], stage0_10[479], stage0_10[480], stage0_10[481]},
      {stage0_11[379]},
      {stage0_12[168], stage0_12[169], stage0_12[170], stage0_12[171], stage0_12[172], stage0_12[173]},
      {stage1_14[28],stage1_13[89],stage1_12[139],stage1_11[165],stage1_10[175]}
   );
   gpc615_5 gpc483 (
      {stage0_10[482], stage0_10[483], stage0_10[484], stage0_10[485], stage0_10[486]},
      {stage0_11[380]},
      {stage0_12[174], stage0_12[175], stage0_12[176], stage0_12[177], stage0_12[178], stage0_12[179]},
      {stage1_14[29],stage1_13[90],stage1_12[140],stage1_11[166],stage1_10[176]}
   );
   gpc615_5 gpc484 (
      {stage0_10[487], stage0_10[488], stage0_10[489], stage0_10[490], stage0_10[491]},
      {stage0_11[381]},
      {stage0_12[180], stage0_12[181], stage0_12[182], stage0_12[183], stage0_12[184], stage0_12[185]},
      {stage1_14[30],stage1_13[91],stage1_12[141],stage1_11[167],stage1_10[177]}
   );
   gpc615_5 gpc485 (
      {stage0_10[492], stage0_10[493], stage0_10[494], stage0_10[495], stage0_10[496]},
      {stage0_11[382]},
      {stage0_12[186], stage0_12[187], stage0_12[188], stage0_12[189], stage0_12[190], stage0_12[191]},
      {stage1_14[31],stage1_13[92],stage1_12[142],stage1_11[168],stage1_10[178]}
   );
   gpc615_5 gpc486 (
      {stage0_10[497], stage0_10[498], stage0_10[499], stage0_10[500], stage0_10[501]},
      {stage0_11[383]},
      {stage0_12[192], stage0_12[193], stage0_12[194], stage0_12[195], stage0_12[196], stage0_12[197]},
      {stage1_14[32],stage1_13[93],stage1_12[143],stage1_11[169],stage1_10[179]}
   );
   gpc615_5 gpc487 (
      {stage0_10[502], stage0_10[503], stage0_10[504], stage0_10[505], stage0_10[506]},
      {stage0_11[384]},
      {stage0_12[198], stage0_12[199], stage0_12[200], stage0_12[201], stage0_12[202], stage0_12[203]},
      {stage1_14[33],stage1_13[94],stage1_12[144],stage1_11[170],stage1_10[180]}
   );
   gpc615_5 gpc488 (
      {stage0_10[507], stage0_10[508], stage0_10[509], stage0_10[510], stage0_10[511]},
      {stage0_11[385]},
      {stage0_12[204], stage0_12[205], stage0_12[206], stage0_12[207], stage0_12[208], stage0_12[209]},
      {stage1_14[34],stage1_13[95],stage1_12[145],stage1_11[171],stage1_10[181]}
   );
   gpc615_5 gpc489 (
      {stage0_11[386], stage0_11[387], stage0_11[388], stage0_11[389], stage0_11[390]},
      {stage0_12[210]},
      {stage0_13[0], stage0_13[1], stage0_13[2], stage0_13[3], stage0_13[4], stage0_13[5]},
      {stage1_15[0],stage1_14[35],stage1_13[96],stage1_12[146],stage1_11[172]}
   );
   gpc615_5 gpc490 (
      {stage0_11[391], stage0_11[392], stage0_11[393], stage0_11[394], stage0_11[395]},
      {stage0_12[211]},
      {stage0_13[6], stage0_13[7], stage0_13[8], stage0_13[9], stage0_13[10], stage0_13[11]},
      {stage1_15[1],stage1_14[36],stage1_13[97],stage1_12[147],stage1_11[173]}
   );
   gpc615_5 gpc491 (
      {stage0_11[396], stage0_11[397], stage0_11[398], stage0_11[399], stage0_11[400]},
      {stage0_12[212]},
      {stage0_13[12], stage0_13[13], stage0_13[14], stage0_13[15], stage0_13[16], stage0_13[17]},
      {stage1_15[2],stage1_14[37],stage1_13[98],stage1_12[148],stage1_11[174]}
   );
   gpc615_5 gpc492 (
      {stage0_11[401], stage0_11[402], stage0_11[403], stage0_11[404], stage0_11[405]},
      {stage0_12[213]},
      {stage0_13[18], stage0_13[19], stage0_13[20], stage0_13[21], stage0_13[22], stage0_13[23]},
      {stage1_15[3],stage1_14[38],stage1_13[99],stage1_12[149],stage1_11[175]}
   );
   gpc615_5 gpc493 (
      {stage0_11[406], stage0_11[407], stage0_11[408], stage0_11[409], stage0_11[410]},
      {stage0_12[214]},
      {stage0_13[24], stage0_13[25], stage0_13[26], stage0_13[27], stage0_13[28], stage0_13[29]},
      {stage1_15[4],stage1_14[39],stage1_13[100],stage1_12[150],stage1_11[176]}
   );
   gpc615_5 gpc494 (
      {stage0_11[411], stage0_11[412], stage0_11[413], stage0_11[414], stage0_11[415]},
      {stage0_12[215]},
      {stage0_13[30], stage0_13[31], stage0_13[32], stage0_13[33], stage0_13[34], stage0_13[35]},
      {stage1_15[5],stage1_14[40],stage1_13[101],stage1_12[151],stage1_11[177]}
   );
   gpc615_5 gpc495 (
      {stage0_11[416], stage0_11[417], stage0_11[418], stage0_11[419], stage0_11[420]},
      {stage0_12[216]},
      {stage0_13[36], stage0_13[37], stage0_13[38], stage0_13[39], stage0_13[40], stage0_13[41]},
      {stage1_15[6],stage1_14[41],stage1_13[102],stage1_12[152],stage1_11[178]}
   );
   gpc615_5 gpc496 (
      {stage0_11[421], stage0_11[422], stage0_11[423], stage0_11[424], stage0_11[425]},
      {stage0_12[217]},
      {stage0_13[42], stage0_13[43], stage0_13[44], stage0_13[45], stage0_13[46], stage0_13[47]},
      {stage1_15[7],stage1_14[42],stage1_13[103],stage1_12[153],stage1_11[179]}
   );
   gpc615_5 gpc497 (
      {stage0_11[426], stage0_11[427], stage0_11[428], stage0_11[429], stage0_11[430]},
      {stage0_12[218]},
      {stage0_13[48], stage0_13[49], stage0_13[50], stage0_13[51], stage0_13[52], stage0_13[53]},
      {stage1_15[8],stage1_14[43],stage1_13[104],stage1_12[154],stage1_11[180]}
   );
   gpc615_5 gpc498 (
      {stage0_11[431], stage0_11[432], stage0_11[433], stage0_11[434], stage0_11[435]},
      {stage0_12[219]},
      {stage0_13[54], stage0_13[55], stage0_13[56], stage0_13[57], stage0_13[58], stage0_13[59]},
      {stage1_15[9],stage1_14[44],stage1_13[105],stage1_12[155],stage1_11[181]}
   );
   gpc615_5 gpc499 (
      {stage0_11[436], stage0_11[437], stage0_11[438], stage0_11[439], stage0_11[440]},
      {stage0_12[220]},
      {stage0_13[60], stage0_13[61], stage0_13[62], stage0_13[63], stage0_13[64], stage0_13[65]},
      {stage1_15[10],stage1_14[45],stage1_13[106],stage1_12[156],stage1_11[182]}
   );
   gpc615_5 gpc500 (
      {stage0_11[441], stage0_11[442], stage0_11[443], stage0_11[444], stage0_11[445]},
      {stage0_12[221]},
      {stage0_13[66], stage0_13[67], stage0_13[68], stage0_13[69], stage0_13[70], stage0_13[71]},
      {stage1_15[11],stage1_14[46],stage1_13[107],stage1_12[157],stage1_11[183]}
   );
   gpc615_5 gpc501 (
      {stage0_11[446], stage0_11[447], stage0_11[448], stage0_11[449], stage0_11[450]},
      {stage0_12[222]},
      {stage0_13[72], stage0_13[73], stage0_13[74], stage0_13[75], stage0_13[76], stage0_13[77]},
      {stage1_15[12],stage1_14[47],stage1_13[108],stage1_12[158],stage1_11[184]}
   );
   gpc615_5 gpc502 (
      {stage0_11[451], stage0_11[452], stage0_11[453], stage0_11[454], stage0_11[455]},
      {stage0_12[223]},
      {stage0_13[78], stage0_13[79], stage0_13[80], stage0_13[81], stage0_13[82], stage0_13[83]},
      {stage1_15[13],stage1_14[48],stage1_13[109],stage1_12[159],stage1_11[185]}
   );
   gpc615_5 gpc503 (
      {stage0_11[456], stage0_11[457], stage0_11[458], stage0_11[459], stage0_11[460]},
      {stage0_12[224]},
      {stage0_13[84], stage0_13[85], stage0_13[86], stage0_13[87], stage0_13[88], stage0_13[89]},
      {stage1_15[14],stage1_14[49],stage1_13[110],stage1_12[160],stage1_11[186]}
   );
   gpc615_5 gpc504 (
      {stage0_11[461], stage0_11[462], stage0_11[463], stage0_11[464], stage0_11[465]},
      {stage0_12[225]},
      {stage0_13[90], stage0_13[91], stage0_13[92], stage0_13[93], stage0_13[94], stage0_13[95]},
      {stage1_15[15],stage1_14[50],stage1_13[111],stage1_12[161],stage1_11[187]}
   );
   gpc615_5 gpc505 (
      {stage0_11[466], stage0_11[467], stage0_11[468], stage0_11[469], stage0_11[470]},
      {stage0_12[226]},
      {stage0_13[96], stage0_13[97], stage0_13[98], stage0_13[99], stage0_13[100], stage0_13[101]},
      {stage1_15[16],stage1_14[51],stage1_13[112],stage1_12[162],stage1_11[188]}
   );
   gpc615_5 gpc506 (
      {stage0_11[471], stage0_11[472], stage0_11[473], stage0_11[474], stage0_11[475]},
      {stage0_12[227]},
      {stage0_13[102], stage0_13[103], stage0_13[104], stage0_13[105], stage0_13[106], stage0_13[107]},
      {stage1_15[17],stage1_14[52],stage1_13[113],stage1_12[163],stage1_11[189]}
   );
   gpc615_5 gpc507 (
      {stage0_11[476], stage0_11[477], stage0_11[478], stage0_11[479], stage0_11[480]},
      {stage0_12[228]},
      {stage0_13[108], stage0_13[109], stage0_13[110], stage0_13[111], stage0_13[112], stage0_13[113]},
      {stage1_15[18],stage1_14[53],stage1_13[114],stage1_12[164],stage1_11[190]}
   );
   gpc615_5 gpc508 (
      {stage0_11[481], stage0_11[482], stage0_11[483], stage0_11[484], stage0_11[485]},
      {stage0_12[229]},
      {stage0_13[114], stage0_13[115], stage0_13[116], stage0_13[117], stage0_13[118], stage0_13[119]},
      {stage1_15[19],stage1_14[54],stage1_13[115],stage1_12[165],stage1_11[191]}
   );
   gpc615_5 gpc509 (
      {stage0_11[486], stage0_11[487], stage0_11[488], stage0_11[489], stage0_11[490]},
      {stage0_12[230]},
      {stage0_13[120], stage0_13[121], stage0_13[122], stage0_13[123], stage0_13[124], stage0_13[125]},
      {stage1_15[20],stage1_14[55],stage1_13[116],stage1_12[166],stage1_11[192]}
   );
   gpc615_5 gpc510 (
      {stage0_11[491], stage0_11[492], stage0_11[493], stage0_11[494], stage0_11[495]},
      {stage0_12[231]},
      {stage0_13[126], stage0_13[127], stage0_13[128], stage0_13[129], stage0_13[130], stage0_13[131]},
      {stage1_15[21],stage1_14[56],stage1_13[117],stage1_12[167],stage1_11[193]}
   );
   gpc615_5 gpc511 (
      {stage0_11[496], stage0_11[497], stage0_11[498], stage0_11[499], stage0_11[500]},
      {stage0_12[232]},
      {stage0_13[132], stage0_13[133], stage0_13[134], stage0_13[135], stage0_13[136], stage0_13[137]},
      {stage1_15[22],stage1_14[57],stage1_13[118],stage1_12[168],stage1_11[194]}
   );
   gpc606_5 gpc512 (
      {stage0_12[233], stage0_12[234], stage0_12[235], stage0_12[236], stage0_12[237], stage0_12[238]},
      {stage0_14[0], stage0_14[1], stage0_14[2], stage0_14[3], stage0_14[4], stage0_14[5]},
      {stage1_16[0],stage1_15[23],stage1_14[58],stage1_13[119],stage1_12[169]}
   );
   gpc606_5 gpc513 (
      {stage0_12[239], stage0_12[240], stage0_12[241], stage0_12[242], stage0_12[243], stage0_12[244]},
      {stage0_14[6], stage0_14[7], stage0_14[8], stage0_14[9], stage0_14[10], stage0_14[11]},
      {stage1_16[1],stage1_15[24],stage1_14[59],stage1_13[120],stage1_12[170]}
   );
   gpc606_5 gpc514 (
      {stage0_12[245], stage0_12[246], stage0_12[247], stage0_12[248], stage0_12[249], stage0_12[250]},
      {stage0_14[12], stage0_14[13], stage0_14[14], stage0_14[15], stage0_14[16], stage0_14[17]},
      {stage1_16[2],stage1_15[25],stage1_14[60],stage1_13[121],stage1_12[171]}
   );
   gpc606_5 gpc515 (
      {stage0_12[251], stage0_12[252], stage0_12[253], stage0_12[254], stage0_12[255], stage0_12[256]},
      {stage0_14[18], stage0_14[19], stage0_14[20], stage0_14[21], stage0_14[22], stage0_14[23]},
      {stage1_16[3],stage1_15[26],stage1_14[61],stage1_13[122],stage1_12[172]}
   );
   gpc606_5 gpc516 (
      {stage0_12[257], stage0_12[258], stage0_12[259], stage0_12[260], stage0_12[261], stage0_12[262]},
      {stage0_14[24], stage0_14[25], stage0_14[26], stage0_14[27], stage0_14[28], stage0_14[29]},
      {stage1_16[4],stage1_15[27],stage1_14[62],stage1_13[123],stage1_12[173]}
   );
   gpc606_5 gpc517 (
      {stage0_12[263], stage0_12[264], stage0_12[265], stage0_12[266], stage0_12[267], stage0_12[268]},
      {stage0_14[30], stage0_14[31], stage0_14[32], stage0_14[33], stage0_14[34], stage0_14[35]},
      {stage1_16[5],stage1_15[28],stage1_14[63],stage1_13[124],stage1_12[174]}
   );
   gpc606_5 gpc518 (
      {stage0_12[269], stage0_12[270], stage0_12[271], stage0_12[272], stage0_12[273], stage0_12[274]},
      {stage0_14[36], stage0_14[37], stage0_14[38], stage0_14[39], stage0_14[40], stage0_14[41]},
      {stage1_16[6],stage1_15[29],stage1_14[64],stage1_13[125],stage1_12[175]}
   );
   gpc606_5 gpc519 (
      {stage0_12[275], stage0_12[276], stage0_12[277], stage0_12[278], stage0_12[279], stage0_12[280]},
      {stage0_14[42], stage0_14[43], stage0_14[44], stage0_14[45], stage0_14[46], stage0_14[47]},
      {stage1_16[7],stage1_15[30],stage1_14[65],stage1_13[126],stage1_12[176]}
   );
   gpc606_5 gpc520 (
      {stage0_12[281], stage0_12[282], stage0_12[283], stage0_12[284], stage0_12[285], stage0_12[286]},
      {stage0_14[48], stage0_14[49], stage0_14[50], stage0_14[51], stage0_14[52], stage0_14[53]},
      {stage1_16[8],stage1_15[31],stage1_14[66],stage1_13[127],stage1_12[177]}
   );
   gpc606_5 gpc521 (
      {stage0_12[287], stage0_12[288], stage0_12[289], stage0_12[290], stage0_12[291], stage0_12[292]},
      {stage0_14[54], stage0_14[55], stage0_14[56], stage0_14[57], stage0_14[58], stage0_14[59]},
      {stage1_16[9],stage1_15[32],stage1_14[67],stage1_13[128],stage1_12[178]}
   );
   gpc606_5 gpc522 (
      {stage0_12[293], stage0_12[294], stage0_12[295], stage0_12[296], stage0_12[297], stage0_12[298]},
      {stage0_14[60], stage0_14[61], stage0_14[62], stage0_14[63], stage0_14[64], stage0_14[65]},
      {stage1_16[10],stage1_15[33],stage1_14[68],stage1_13[129],stage1_12[179]}
   );
   gpc606_5 gpc523 (
      {stage0_12[299], stage0_12[300], stage0_12[301], stage0_12[302], stage0_12[303], stage0_12[304]},
      {stage0_14[66], stage0_14[67], stage0_14[68], stage0_14[69], stage0_14[70], stage0_14[71]},
      {stage1_16[11],stage1_15[34],stage1_14[69],stage1_13[130],stage1_12[180]}
   );
   gpc606_5 gpc524 (
      {stage0_12[305], stage0_12[306], stage0_12[307], stage0_12[308], stage0_12[309], stage0_12[310]},
      {stage0_14[72], stage0_14[73], stage0_14[74], stage0_14[75], stage0_14[76], stage0_14[77]},
      {stage1_16[12],stage1_15[35],stage1_14[70],stage1_13[131],stage1_12[181]}
   );
   gpc606_5 gpc525 (
      {stage0_12[311], stage0_12[312], stage0_12[313], stage0_12[314], stage0_12[315], stage0_12[316]},
      {stage0_14[78], stage0_14[79], stage0_14[80], stage0_14[81], stage0_14[82], stage0_14[83]},
      {stage1_16[13],stage1_15[36],stage1_14[71],stage1_13[132],stage1_12[182]}
   );
   gpc615_5 gpc526 (
      {stage0_12[317], stage0_12[318], stage0_12[319], stage0_12[320], stage0_12[321]},
      {stage0_13[138]},
      {stage0_14[84], stage0_14[85], stage0_14[86], stage0_14[87], stage0_14[88], stage0_14[89]},
      {stage1_16[14],stage1_15[37],stage1_14[72],stage1_13[133],stage1_12[183]}
   );
   gpc615_5 gpc527 (
      {stage0_12[322], stage0_12[323], stage0_12[324], stage0_12[325], stage0_12[326]},
      {stage0_13[139]},
      {stage0_14[90], stage0_14[91], stage0_14[92], stage0_14[93], stage0_14[94], stage0_14[95]},
      {stage1_16[15],stage1_15[38],stage1_14[73],stage1_13[134],stage1_12[184]}
   );
   gpc615_5 gpc528 (
      {stage0_12[327], stage0_12[328], stage0_12[329], stage0_12[330], stage0_12[331]},
      {stage0_13[140]},
      {stage0_14[96], stage0_14[97], stage0_14[98], stage0_14[99], stage0_14[100], stage0_14[101]},
      {stage1_16[16],stage1_15[39],stage1_14[74],stage1_13[135],stage1_12[185]}
   );
   gpc615_5 gpc529 (
      {stage0_12[332], stage0_12[333], stage0_12[334], stage0_12[335], stage0_12[336]},
      {stage0_13[141]},
      {stage0_14[102], stage0_14[103], stage0_14[104], stage0_14[105], stage0_14[106], stage0_14[107]},
      {stage1_16[17],stage1_15[40],stage1_14[75],stage1_13[136],stage1_12[186]}
   );
   gpc615_5 gpc530 (
      {stage0_12[337], stage0_12[338], stage0_12[339], stage0_12[340], stage0_12[341]},
      {stage0_13[142]},
      {stage0_14[108], stage0_14[109], stage0_14[110], stage0_14[111], stage0_14[112], stage0_14[113]},
      {stage1_16[18],stage1_15[41],stage1_14[76],stage1_13[137],stage1_12[187]}
   );
   gpc615_5 gpc531 (
      {stage0_12[342], stage0_12[343], stage0_12[344], stage0_12[345], stage0_12[346]},
      {stage0_13[143]},
      {stage0_14[114], stage0_14[115], stage0_14[116], stage0_14[117], stage0_14[118], stage0_14[119]},
      {stage1_16[19],stage1_15[42],stage1_14[77],stage1_13[138],stage1_12[188]}
   );
   gpc615_5 gpc532 (
      {stage0_12[347], stage0_12[348], stage0_12[349], stage0_12[350], stage0_12[351]},
      {stage0_13[144]},
      {stage0_14[120], stage0_14[121], stage0_14[122], stage0_14[123], stage0_14[124], stage0_14[125]},
      {stage1_16[20],stage1_15[43],stage1_14[78],stage1_13[139],stage1_12[189]}
   );
   gpc615_5 gpc533 (
      {stage0_12[352], stage0_12[353], stage0_12[354], stage0_12[355], stage0_12[356]},
      {stage0_13[145]},
      {stage0_14[126], stage0_14[127], stage0_14[128], stage0_14[129], stage0_14[130], stage0_14[131]},
      {stage1_16[21],stage1_15[44],stage1_14[79],stage1_13[140],stage1_12[190]}
   );
   gpc615_5 gpc534 (
      {stage0_12[357], stage0_12[358], stage0_12[359], stage0_12[360], stage0_12[361]},
      {stage0_13[146]},
      {stage0_14[132], stage0_14[133], stage0_14[134], stage0_14[135], stage0_14[136], stage0_14[137]},
      {stage1_16[22],stage1_15[45],stage1_14[80],stage1_13[141],stage1_12[191]}
   );
   gpc615_5 gpc535 (
      {stage0_12[362], stage0_12[363], stage0_12[364], stage0_12[365], stage0_12[366]},
      {stage0_13[147]},
      {stage0_14[138], stage0_14[139], stage0_14[140], stage0_14[141], stage0_14[142], stage0_14[143]},
      {stage1_16[23],stage1_15[46],stage1_14[81],stage1_13[142],stage1_12[192]}
   );
   gpc615_5 gpc536 (
      {stage0_12[367], stage0_12[368], stage0_12[369], stage0_12[370], stage0_12[371]},
      {stage0_13[148]},
      {stage0_14[144], stage0_14[145], stage0_14[146], stage0_14[147], stage0_14[148], stage0_14[149]},
      {stage1_16[24],stage1_15[47],stage1_14[82],stage1_13[143],stage1_12[193]}
   );
   gpc615_5 gpc537 (
      {stage0_12[372], stage0_12[373], stage0_12[374], stage0_12[375], stage0_12[376]},
      {stage0_13[149]},
      {stage0_14[150], stage0_14[151], stage0_14[152], stage0_14[153], stage0_14[154], stage0_14[155]},
      {stage1_16[25],stage1_15[48],stage1_14[83],stage1_13[144],stage1_12[194]}
   );
   gpc615_5 gpc538 (
      {stage0_12[377], stage0_12[378], stage0_12[379], stage0_12[380], stage0_12[381]},
      {stage0_13[150]},
      {stage0_14[156], stage0_14[157], stage0_14[158], stage0_14[159], stage0_14[160], stage0_14[161]},
      {stage1_16[26],stage1_15[49],stage1_14[84],stage1_13[145],stage1_12[195]}
   );
   gpc615_5 gpc539 (
      {stage0_12[382], stage0_12[383], stage0_12[384], stage0_12[385], stage0_12[386]},
      {stage0_13[151]},
      {stage0_14[162], stage0_14[163], stage0_14[164], stage0_14[165], stage0_14[166], stage0_14[167]},
      {stage1_16[27],stage1_15[50],stage1_14[85],stage1_13[146],stage1_12[196]}
   );
   gpc615_5 gpc540 (
      {stage0_12[387], stage0_12[388], stage0_12[389], stage0_12[390], stage0_12[391]},
      {stage0_13[152]},
      {stage0_14[168], stage0_14[169], stage0_14[170], stage0_14[171], stage0_14[172], stage0_14[173]},
      {stage1_16[28],stage1_15[51],stage1_14[86],stage1_13[147],stage1_12[197]}
   );
   gpc615_5 gpc541 (
      {stage0_12[392], stage0_12[393], stage0_12[394], stage0_12[395], stage0_12[396]},
      {stage0_13[153]},
      {stage0_14[174], stage0_14[175], stage0_14[176], stage0_14[177], stage0_14[178], stage0_14[179]},
      {stage1_16[29],stage1_15[52],stage1_14[87],stage1_13[148],stage1_12[198]}
   );
   gpc615_5 gpc542 (
      {stage0_12[397], stage0_12[398], stage0_12[399], stage0_12[400], stage0_12[401]},
      {stage0_13[154]},
      {stage0_14[180], stage0_14[181], stage0_14[182], stage0_14[183], stage0_14[184], stage0_14[185]},
      {stage1_16[30],stage1_15[53],stage1_14[88],stage1_13[149],stage1_12[199]}
   );
   gpc615_5 gpc543 (
      {stage0_12[402], stage0_12[403], stage0_12[404], stage0_12[405], stage0_12[406]},
      {stage0_13[155]},
      {stage0_14[186], stage0_14[187], stage0_14[188], stage0_14[189], stage0_14[190], stage0_14[191]},
      {stage1_16[31],stage1_15[54],stage1_14[89],stage1_13[150],stage1_12[200]}
   );
   gpc615_5 gpc544 (
      {stage0_12[407], stage0_12[408], stage0_12[409], stage0_12[410], stage0_12[411]},
      {stage0_13[156]},
      {stage0_14[192], stage0_14[193], stage0_14[194], stage0_14[195], stage0_14[196], stage0_14[197]},
      {stage1_16[32],stage1_15[55],stage1_14[90],stage1_13[151],stage1_12[201]}
   );
   gpc615_5 gpc545 (
      {stage0_12[412], stage0_12[413], stage0_12[414], stage0_12[415], stage0_12[416]},
      {stage0_13[157]},
      {stage0_14[198], stage0_14[199], stage0_14[200], stage0_14[201], stage0_14[202], stage0_14[203]},
      {stage1_16[33],stage1_15[56],stage1_14[91],stage1_13[152],stage1_12[202]}
   );
   gpc615_5 gpc546 (
      {stage0_12[417], stage0_12[418], stage0_12[419], stage0_12[420], stage0_12[421]},
      {stage0_13[158]},
      {stage0_14[204], stage0_14[205], stage0_14[206], stage0_14[207], stage0_14[208], stage0_14[209]},
      {stage1_16[34],stage1_15[57],stage1_14[92],stage1_13[153],stage1_12[203]}
   );
   gpc615_5 gpc547 (
      {stage0_12[422], stage0_12[423], stage0_12[424], stage0_12[425], stage0_12[426]},
      {stage0_13[159]},
      {stage0_14[210], stage0_14[211], stage0_14[212], stage0_14[213], stage0_14[214], stage0_14[215]},
      {stage1_16[35],stage1_15[58],stage1_14[93],stage1_13[154],stage1_12[204]}
   );
   gpc615_5 gpc548 (
      {stage0_12[427], stage0_12[428], stage0_12[429], stage0_12[430], stage0_12[431]},
      {stage0_13[160]},
      {stage0_14[216], stage0_14[217], stage0_14[218], stage0_14[219], stage0_14[220], stage0_14[221]},
      {stage1_16[36],stage1_15[59],stage1_14[94],stage1_13[155],stage1_12[205]}
   );
   gpc615_5 gpc549 (
      {stage0_12[432], stage0_12[433], stage0_12[434], stage0_12[435], stage0_12[436]},
      {stage0_13[161]},
      {stage0_14[222], stage0_14[223], stage0_14[224], stage0_14[225], stage0_14[226], stage0_14[227]},
      {stage1_16[37],stage1_15[60],stage1_14[95],stage1_13[156],stage1_12[206]}
   );
   gpc615_5 gpc550 (
      {stage0_12[437], stage0_12[438], stage0_12[439], stage0_12[440], stage0_12[441]},
      {stage0_13[162]},
      {stage0_14[228], stage0_14[229], stage0_14[230], stage0_14[231], stage0_14[232], stage0_14[233]},
      {stage1_16[38],stage1_15[61],stage1_14[96],stage1_13[157],stage1_12[207]}
   );
   gpc615_5 gpc551 (
      {stage0_12[442], stage0_12[443], stage0_12[444], stage0_12[445], stage0_12[446]},
      {stage0_13[163]},
      {stage0_14[234], stage0_14[235], stage0_14[236], stage0_14[237], stage0_14[238], stage0_14[239]},
      {stage1_16[39],stage1_15[62],stage1_14[97],stage1_13[158],stage1_12[208]}
   );
   gpc615_5 gpc552 (
      {stage0_12[447], stage0_12[448], stage0_12[449], stage0_12[450], stage0_12[451]},
      {stage0_13[164]},
      {stage0_14[240], stage0_14[241], stage0_14[242], stage0_14[243], stage0_14[244], stage0_14[245]},
      {stage1_16[40],stage1_15[63],stage1_14[98],stage1_13[159],stage1_12[209]}
   );
   gpc615_5 gpc553 (
      {stage0_12[452], stage0_12[453], stage0_12[454], stage0_12[455], stage0_12[456]},
      {stage0_13[165]},
      {stage0_14[246], stage0_14[247], stage0_14[248], stage0_14[249], stage0_14[250], stage0_14[251]},
      {stage1_16[41],stage1_15[64],stage1_14[99],stage1_13[160],stage1_12[210]}
   );
   gpc615_5 gpc554 (
      {stage0_12[457], stage0_12[458], stage0_12[459], stage0_12[460], stage0_12[461]},
      {stage0_13[166]},
      {stage0_14[252], stage0_14[253], stage0_14[254], stage0_14[255], stage0_14[256], stage0_14[257]},
      {stage1_16[42],stage1_15[65],stage1_14[100],stage1_13[161],stage1_12[211]}
   );
   gpc615_5 gpc555 (
      {stage0_12[462], stage0_12[463], stage0_12[464], stage0_12[465], stage0_12[466]},
      {stage0_13[167]},
      {stage0_14[258], stage0_14[259], stage0_14[260], stage0_14[261], stage0_14[262], stage0_14[263]},
      {stage1_16[43],stage1_15[66],stage1_14[101],stage1_13[162],stage1_12[212]}
   );
   gpc615_5 gpc556 (
      {stage0_12[467], stage0_12[468], stage0_12[469], stage0_12[470], stage0_12[471]},
      {stage0_13[168]},
      {stage0_14[264], stage0_14[265], stage0_14[266], stage0_14[267], stage0_14[268], stage0_14[269]},
      {stage1_16[44],stage1_15[67],stage1_14[102],stage1_13[163],stage1_12[213]}
   );
   gpc615_5 gpc557 (
      {stage0_12[472], stage0_12[473], stage0_12[474], stage0_12[475], stage0_12[476]},
      {stage0_13[169]},
      {stage0_14[270], stage0_14[271], stage0_14[272], stage0_14[273], stage0_14[274], stage0_14[275]},
      {stage1_16[45],stage1_15[68],stage1_14[103],stage1_13[164],stage1_12[214]}
   );
   gpc615_5 gpc558 (
      {stage0_12[477], stage0_12[478], stage0_12[479], stage0_12[480], stage0_12[481]},
      {stage0_13[170]},
      {stage0_14[276], stage0_14[277], stage0_14[278], stage0_14[279], stage0_14[280], stage0_14[281]},
      {stage1_16[46],stage1_15[69],stage1_14[104],stage1_13[165],stage1_12[215]}
   );
   gpc615_5 gpc559 (
      {stage0_12[482], stage0_12[483], stage0_12[484], stage0_12[485], stage0_12[486]},
      {stage0_13[171]},
      {stage0_14[282], stage0_14[283], stage0_14[284], stage0_14[285], stage0_14[286], stage0_14[287]},
      {stage1_16[47],stage1_15[70],stage1_14[105],stage1_13[166],stage1_12[216]}
   );
   gpc615_5 gpc560 (
      {stage0_12[487], stage0_12[488], stage0_12[489], stage0_12[490], stage0_12[491]},
      {stage0_13[172]},
      {stage0_14[288], stage0_14[289], stage0_14[290], stage0_14[291], stage0_14[292], stage0_14[293]},
      {stage1_16[48],stage1_15[71],stage1_14[106],stage1_13[167],stage1_12[217]}
   );
   gpc615_5 gpc561 (
      {stage0_12[492], stage0_12[493], stage0_12[494], stage0_12[495], stage0_12[496]},
      {stage0_13[173]},
      {stage0_14[294], stage0_14[295], stage0_14[296], stage0_14[297], stage0_14[298], stage0_14[299]},
      {stage1_16[49],stage1_15[72],stage1_14[107],stage1_13[168],stage1_12[218]}
   );
   gpc615_5 gpc562 (
      {stage0_12[497], stage0_12[498], stage0_12[499], stage0_12[500], stage0_12[501]},
      {stage0_13[174]},
      {stage0_14[300], stage0_14[301], stage0_14[302], stage0_14[303], stage0_14[304], stage0_14[305]},
      {stage1_16[50],stage1_15[73],stage1_14[108],stage1_13[169],stage1_12[219]}
   );
   gpc615_5 gpc563 (
      {stage0_12[502], stage0_12[503], stage0_12[504], stage0_12[505], stage0_12[506]},
      {stage0_13[175]},
      {stage0_14[306], stage0_14[307], stage0_14[308], stage0_14[309], stage0_14[310], stage0_14[311]},
      {stage1_16[51],stage1_15[74],stage1_14[109],stage1_13[170],stage1_12[220]}
   );
   gpc615_5 gpc564 (
      {stage0_12[507], stage0_12[508], stage0_12[509], stage0_12[510], stage0_12[511]},
      {stage0_13[176]},
      {stage0_14[312], stage0_14[313], stage0_14[314], stage0_14[315], stage0_14[316], stage0_14[317]},
      {stage1_16[52],stage1_15[75],stage1_14[110],stage1_13[171],stage1_12[221]}
   );
   gpc606_5 gpc565 (
      {stage0_13[177], stage0_13[178], stage0_13[179], stage0_13[180], stage0_13[181], stage0_13[182]},
      {stage0_15[0], stage0_15[1], stage0_15[2], stage0_15[3], stage0_15[4], stage0_15[5]},
      {stage1_17[0],stage1_16[53],stage1_15[76],stage1_14[111],stage1_13[172]}
   );
   gpc606_5 gpc566 (
      {stage0_13[183], stage0_13[184], stage0_13[185], stage0_13[186], stage0_13[187], stage0_13[188]},
      {stage0_15[6], stage0_15[7], stage0_15[8], stage0_15[9], stage0_15[10], stage0_15[11]},
      {stage1_17[1],stage1_16[54],stage1_15[77],stage1_14[112],stage1_13[173]}
   );
   gpc606_5 gpc567 (
      {stage0_13[189], stage0_13[190], stage0_13[191], stage0_13[192], stage0_13[193], stage0_13[194]},
      {stage0_15[12], stage0_15[13], stage0_15[14], stage0_15[15], stage0_15[16], stage0_15[17]},
      {stage1_17[2],stage1_16[55],stage1_15[78],stage1_14[113],stage1_13[174]}
   );
   gpc606_5 gpc568 (
      {stage0_13[195], stage0_13[196], stage0_13[197], stage0_13[198], stage0_13[199], stage0_13[200]},
      {stage0_15[18], stage0_15[19], stage0_15[20], stage0_15[21], stage0_15[22], stage0_15[23]},
      {stage1_17[3],stage1_16[56],stage1_15[79],stage1_14[114],stage1_13[175]}
   );
   gpc606_5 gpc569 (
      {stage0_13[201], stage0_13[202], stage0_13[203], stage0_13[204], stage0_13[205], stage0_13[206]},
      {stage0_15[24], stage0_15[25], stage0_15[26], stage0_15[27], stage0_15[28], stage0_15[29]},
      {stage1_17[4],stage1_16[57],stage1_15[80],stage1_14[115],stage1_13[176]}
   );
   gpc606_5 gpc570 (
      {stage0_13[207], stage0_13[208], stage0_13[209], stage0_13[210], stage0_13[211], stage0_13[212]},
      {stage0_15[30], stage0_15[31], stage0_15[32], stage0_15[33], stage0_15[34], stage0_15[35]},
      {stage1_17[5],stage1_16[58],stage1_15[81],stage1_14[116],stage1_13[177]}
   );
   gpc606_5 gpc571 (
      {stage0_13[213], stage0_13[214], stage0_13[215], stage0_13[216], stage0_13[217], stage0_13[218]},
      {stage0_15[36], stage0_15[37], stage0_15[38], stage0_15[39], stage0_15[40], stage0_15[41]},
      {stage1_17[6],stage1_16[59],stage1_15[82],stage1_14[117],stage1_13[178]}
   );
   gpc606_5 gpc572 (
      {stage0_13[219], stage0_13[220], stage0_13[221], stage0_13[222], stage0_13[223], stage0_13[224]},
      {stage0_15[42], stage0_15[43], stage0_15[44], stage0_15[45], stage0_15[46], stage0_15[47]},
      {stage1_17[7],stage1_16[60],stage1_15[83],stage1_14[118],stage1_13[179]}
   );
   gpc606_5 gpc573 (
      {stage0_13[225], stage0_13[226], stage0_13[227], stage0_13[228], stage0_13[229], stage0_13[230]},
      {stage0_15[48], stage0_15[49], stage0_15[50], stage0_15[51], stage0_15[52], stage0_15[53]},
      {stage1_17[8],stage1_16[61],stage1_15[84],stage1_14[119],stage1_13[180]}
   );
   gpc606_5 gpc574 (
      {stage0_13[231], stage0_13[232], stage0_13[233], stage0_13[234], stage0_13[235], stage0_13[236]},
      {stage0_15[54], stage0_15[55], stage0_15[56], stage0_15[57], stage0_15[58], stage0_15[59]},
      {stage1_17[9],stage1_16[62],stage1_15[85],stage1_14[120],stage1_13[181]}
   );
   gpc606_5 gpc575 (
      {stage0_13[237], stage0_13[238], stage0_13[239], stage0_13[240], stage0_13[241], stage0_13[242]},
      {stage0_15[60], stage0_15[61], stage0_15[62], stage0_15[63], stage0_15[64], stage0_15[65]},
      {stage1_17[10],stage1_16[63],stage1_15[86],stage1_14[121],stage1_13[182]}
   );
   gpc606_5 gpc576 (
      {stage0_13[243], stage0_13[244], stage0_13[245], stage0_13[246], stage0_13[247], stage0_13[248]},
      {stage0_15[66], stage0_15[67], stage0_15[68], stage0_15[69], stage0_15[70], stage0_15[71]},
      {stage1_17[11],stage1_16[64],stage1_15[87],stage1_14[122],stage1_13[183]}
   );
   gpc606_5 gpc577 (
      {stage0_13[249], stage0_13[250], stage0_13[251], stage0_13[252], stage0_13[253], stage0_13[254]},
      {stage0_15[72], stage0_15[73], stage0_15[74], stage0_15[75], stage0_15[76], stage0_15[77]},
      {stage1_17[12],stage1_16[65],stage1_15[88],stage1_14[123],stage1_13[184]}
   );
   gpc606_5 gpc578 (
      {stage0_13[255], stage0_13[256], stage0_13[257], stage0_13[258], stage0_13[259], stage0_13[260]},
      {stage0_15[78], stage0_15[79], stage0_15[80], stage0_15[81], stage0_15[82], stage0_15[83]},
      {stage1_17[13],stage1_16[66],stage1_15[89],stage1_14[124],stage1_13[185]}
   );
   gpc606_5 gpc579 (
      {stage0_13[261], stage0_13[262], stage0_13[263], stage0_13[264], stage0_13[265], stage0_13[266]},
      {stage0_15[84], stage0_15[85], stage0_15[86], stage0_15[87], stage0_15[88], stage0_15[89]},
      {stage1_17[14],stage1_16[67],stage1_15[90],stage1_14[125],stage1_13[186]}
   );
   gpc606_5 gpc580 (
      {stage0_13[267], stage0_13[268], stage0_13[269], stage0_13[270], stage0_13[271], stage0_13[272]},
      {stage0_15[90], stage0_15[91], stage0_15[92], stage0_15[93], stage0_15[94], stage0_15[95]},
      {stage1_17[15],stage1_16[68],stage1_15[91],stage1_14[126],stage1_13[187]}
   );
   gpc606_5 gpc581 (
      {stage0_13[273], stage0_13[274], stage0_13[275], stage0_13[276], stage0_13[277], stage0_13[278]},
      {stage0_15[96], stage0_15[97], stage0_15[98], stage0_15[99], stage0_15[100], stage0_15[101]},
      {stage1_17[16],stage1_16[69],stage1_15[92],stage1_14[127],stage1_13[188]}
   );
   gpc606_5 gpc582 (
      {stage0_13[279], stage0_13[280], stage0_13[281], stage0_13[282], stage0_13[283], stage0_13[284]},
      {stage0_15[102], stage0_15[103], stage0_15[104], stage0_15[105], stage0_15[106], stage0_15[107]},
      {stage1_17[17],stage1_16[70],stage1_15[93],stage1_14[128],stage1_13[189]}
   );
   gpc606_5 gpc583 (
      {stage0_13[285], stage0_13[286], stage0_13[287], stage0_13[288], stage0_13[289], stage0_13[290]},
      {stage0_15[108], stage0_15[109], stage0_15[110], stage0_15[111], stage0_15[112], stage0_15[113]},
      {stage1_17[18],stage1_16[71],stage1_15[94],stage1_14[129],stage1_13[190]}
   );
   gpc606_5 gpc584 (
      {stage0_13[291], stage0_13[292], stage0_13[293], stage0_13[294], stage0_13[295], stage0_13[296]},
      {stage0_15[114], stage0_15[115], stage0_15[116], stage0_15[117], stage0_15[118], stage0_15[119]},
      {stage1_17[19],stage1_16[72],stage1_15[95],stage1_14[130],stage1_13[191]}
   );
   gpc606_5 gpc585 (
      {stage0_13[297], stage0_13[298], stage0_13[299], stage0_13[300], stage0_13[301], stage0_13[302]},
      {stage0_15[120], stage0_15[121], stage0_15[122], stage0_15[123], stage0_15[124], stage0_15[125]},
      {stage1_17[20],stage1_16[73],stage1_15[96],stage1_14[131],stage1_13[192]}
   );
   gpc606_5 gpc586 (
      {stage0_13[303], stage0_13[304], stage0_13[305], stage0_13[306], stage0_13[307], stage0_13[308]},
      {stage0_15[126], stage0_15[127], stage0_15[128], stage0_15[129], stage0_15[130], stage0_15[131]},
      {stage1_17[21],stage1_16[74],stage1_15[97],stage1_14[132],stage1_13[193]}
   );
   gpc606_5 gpc587 (
      {stage0_13[309], stage0_13[310], stage0_13[311], stage0_13[312], stage0_13[313], stage0_13[314]},
      {stage0_15[132], stage0_15[133], stage0_15[134], stage0_15[135], stage0_15[136], stage0_15[137]},
      {stage1_17[22],stage1_16[75],stage1_15[98],stage1_14[133],stage1_13[194]}
   );
   gpc606_5 gpc588 (
      {stage0_13[315], stage0_13[316], stage0_13[317], stage0_13[318], stage0_13[319], stage0_13[320]},
      {stage0_15[138], stage0_15[139], stage0_15[140], stage0_15[141], stage0_15[142], stage0_15[143]},
      {stage1_17[23],stage1_16[76],stage1_15[99],stage1_14[134],stage1_13[195]}
   );
   gpc606_5 gpc589 (
      {stage0_13[321], stage0_13[322], stage0_13[323], stage0_13[324], stage0_13[325], stage0_13[326]},
      {stage0_15[144], stage0_15[145], stage0_15[146], stage0_15[147], stage0_15[148], stage0_15[149]},
      {stage1_17[24],stage1_16[77],stage1_15[100],stage1_14[135],stage1_13[196]}
   );
   gpc606_5 gpc590 (
      {stage0_13[327], stage0_13[328], stage0_13[329], stage0_13[330], stage0_13[331], stage0_13[332]},
      {stage0_15[150], stage0_15[151], stage0_15[152], stage0_15[153], stage0_15[154], stage0_15[155]},
      {stage1_17[25],stage1_16[78],stage1_15[101],stage1_14[136],stage1_13[197]}
   );
   gpc606_5 gpc591 (
      {stage0_13[333], stage0_13[334], stage0_13[335], stage0_13[336], stage0_13[337], stage0_13[338]},
      {stage0_15[156], stage0_15[157], stage0_15[158], stage0_15[159], stage0_15[160], stage0_15[161]},
      {stage1_17[26],stage1_16[79],stage1_15[102],stage1_14[137],stage1_13[198]}
   );
   gpc606_5 gpc592 (
      {stage0_13[339], stage0_13[340], stage0_13[341], stage0_13[342], stage0_13[343], stage0_13[344]},
      {stage0_15[162], stage0_15[163], stage0_15[164], stage0_15[165], stage0_15[166], stage0_15[167]},
      {stage1_17[27],stage1_16[80],stage1_15[103],stage1_14[138],stage1_13[199]}
   );
   gpc606_5 gpc593 (
      {stage0_13[345], stage0_13[346], stage0_13[347], stage0_13[348], stage0_13[349], stage0_13[350]},
      {stage0_15[168], stage0_15[169], stage0_15[170], stage0_15[171], stage0_15[172], stage0_15[173]},
      {stage1_17[28],stage1_16[81],stage1_15[104],stage1_14[139],stage1_13[200]}
   );
   gpc606_5 gpc594 (
      {stage0_13[351], stage0_13[352], stage0_13[353], stage0_13[354], stage0_13[355], stage0_13[356]},
      {stage0_15[174], stage0_15[175], stage0_15[176], stage0_15[177], stage0_15[178], stage0_15[179]},
      {stage1_17[29],stage1_16[82],stage1_15[105],stage1_14[140],stage1_13[201]}
   );
   gpc606_5 gpc595 (
      {stage0_13[357], stage0_13[358], stage0_13[359], stage0_13[360], stage0_13[361], stage0_13[362]},
      {stage0_15[180], stage0_15[181], stage0_15[182], stage0_15[183], stage0_15[184], stage0_15[185]},
      {stage1_17[30],stage1_16[83],stage1_15[106],stage1_14[141],stage1_13[202]}
   );
   gpc606_5 gpc596 (
      {stage0_13[363], stage0_13[364], stage0_13[365], stage0_13[366], stage0_13[367], stage0_13[368]},
      {stage0_15[186], stage0_15[187], stage0_15[188], stage0_15[189], stage0_15[190], stage0_15[191]},
      {stage1_17[31],stage1_16[84],stage1_15[107],stage1_14[142],stage1_13[203]}
   );
   gpc606_5 gpc597 (
      {stage0_13[369], stage0_13[370], stage0_13[371], stage0_13[372], stage0_13[373], stage0_13[374]},
      {stage0_15[192], stage0_15[193], stage0_15[194], stage0_15[195], stage0_15[196], stage0_15[197]},
      {stage1_17[32],stage1_16[85],stage1_15[108],stage1_14[143],stage1_13[204]}
   );
   gpc606_5 gpc598 (
      {stage0_13[375], stage0_13[376], stage0_13[377], stage0_13[378], stage0_13[379], stage0_13[380]},
      {stage0_15[198], stage0_15[199], stage0_15[200], stage0_15[201], stage0_15[202], stage0_15[203]},
      {stage1_17[33],stage1_16[86],stage1_15[109],stage1_14[144],stage1_13[205]}
   );
   gpc606_5 gpc599 (
      {stage0_13[381], stage0_13[382], stage0_13[383], stage0_13[384], stage0_13[385], stage0_13[386]},
      {stage0_15[204], stage0_15[205], stage0_15[206], stage0_15[207], stage0_15[208], stage0_15[209]},
      {stage1_17[34],stage1_16[87],stage1_15[110],stage1_14[145],stage1_13[206]}
   );
   gpc606_5 gpc600 (
      {stage0_13[387], stage0_13[388], stage0_13[389], stage0_13[390], stage0_13[391], stage0_13[392]},
      {stage0_15[210], stage0_15[211], stage0_15[212], stage0_15[213], stage0_15[214], stage0_15[215]},
      {stage1_17[35],stage1_16[88],stage1_15[111],stage1_14[146],stage1_13[207]}
   );
   gpc606_5 gpc601 (
      {stage0_13[393], stage0_13[394], stage0_13[395], stage0_13[396], stage0_13[397], stage0_13[398]},
      {stage0_15[216], stage0_15[217], stage0_15[218], stage0_15[219], stage0_15[220], stage0_15[221]},
      {stage1_17[36],stage1_16[89],stage1_15[112],stage1_14[147],stage1_13[208]}
   );
   gpc606_5 gpc602 (
      {stage0_13[399], stage0_13[400], stage0_13[401], stage0_13[402], stage0_13[403], stage0_13[404]},
      {stage0_15[222], stage0_15[223], stage0_15[224], stage0_15[225], stage0_15[226], stage0_15[227]},
      {stage1_17[37],stage1_16[90],stage1_15[113],stage1_14[148],stage1_13[209]}
   );
   gpc606_5 gpc603 (
      {stage0_13[405], stage0_13[406], stage0_13[407], stage0_13[408], stage0_13[409], stage0_13[410]},
      {stage0_15[228], stage0_15[229], stage0_15[230], stage0_15[231], stage0_15[232], stage0_15[233]},
      {stage1_17[38],stage1_16[91],stage1_15[114],stage1_14[149],stage1_13[210]}
   );
   gpc606_5 gpc604 (
      {stage0_13[411], stage0_13[412], stage0_13[413], stage0_13[414], stage0_13[415], stage0_13[416]},
      {stage0_15[234], stage0_15[235], stage0_15[236], stage0_15[237], stage0_15[238], stage0_15[239]},
      {stage1_17[39],stage1_16[92],stage1_15[115],stage1_14[150],stage1_13[211]}
   );
   gpc606_5 gpc605 (
      {stage0_13[417], stage0_13[418], stage0_13[419], stage0_13[420], stage0_13[421], stage0_13[422]},
      {stage0_15[240], stage0_15[241], stage0_15[242], stage0_15[243], stage0_15[244], stage0_15[245]},
      {stage1_17[40],stage1_16[93],stage1_15[116],stage1_14[151],stage1_13[212]}
   );
   gpc606_5 gpc606 (
      {stage0_13[423], stage0_13[424], stage0_13[425], stage0_13[426], stage0_13[427], stage0_13[428]},
      {stage0_15[246], stage0_15[247], stage0_15[248], stage0_15[249], stage0_15[250], stage0_15[251]},
      {stage1_17[41],stage1_16[94],stage1_15[117],stage1_14[152],stage1_13[213]}
   );
   gpc606_5 gpc607 (
      {stage0_13[429], stage0_13[430], stage0_13[431], stage0_13[432], stage0_13[433], stage0_13[434]},
      {stage0_15[252], stage0_15[253], stage0_15[254], stage0_15[255], stage0_15[256], stage0_15[257]},
      {stage1_17[42],stage1_16[95],stage1_15[118],stage1_14[153],stage1_13[214]}
   );
   gpc606_5 gpc608 (
      {stage0_13[435], stage0_13[436], stage0_13[437], stage0_13[438], stage0_13[439], stage0_13[440]},
      {stage0_15[258], stage0_15[259], stage0_15[260], stage0_15[261], stage0_15[262], stage0_15[263]},
      {stage1_17[43],stage1_16[96],stage1_15[119],stage1_14[154],stage1_13[215]}
   );
   gpc606_5 gpc609 (
      {stage0_13[441], stage0_13[442], stage0_13[443], stage0_13[444], stage0_13[445], stage0_13[446]},
      {stage0_15[264], stage0_15[265], stage0_15[266], stage0_15[267], stage0_15[268], stage0_15[269]},
      {stage1_17[44],stage1_16[97],stage1_15[120],stage1_14[155],stage1_13[216]}
   );
   gpc606_5 gpc610 (
      {stage0_13[447], stage0_13[448], stage0_13[449], stage0_13[450], stage0_13[451], stage0_13[452]},
      {stage0_15[270], stage0_15[271], stage0_15[272], stage0_15[273], stage0_15[274], stage0_15[275]},
      {stage1_17[45],stage1_16[98],stage1_15[121],stage1_14[156],stage1_13[217]}
   );
   gpc606_5 gpc611 (
      {stage0_13[453], stage0_13[454], stage0_13[455], stage0_13[456], stage0_13[457], stage0_13[458]},
      {stage0_15[276], stage0_15[277], stage0_15[278], stage0_15[279], stage0_15[280], stage0_15[281]},
      {stage1_17[46],stage1_16[99],stage1_15[122],stage1_14[157],stage1_13[218]}
   );
   gpc606_5 gpc612 (
      {stage0_13[459], stage0_13[460], stage0_13[461], stage0_13[462], stage0_13[463], stage0_13[464]},
      {stage0_15[282], stage0_15[283], stage0_15[284], stage0_15[285], stage0_15[286], stage0_15[287]},
      {stage1_17[47],stage1_16[100],stage1_15[123],stage1_14[158],stage1_13[219]}
   );
   gpc606_5 gpc613 (
      {stage0_13[465], stage0_13[466], stage0_13[467], stage0_13[468], stage0_13[469], stage0_13[470]},
      {stage0_15[288], stage0_15[289], stage0_15[290], stage0_15[291], stage0_15[292], stage0_15[293]},
      {stage1_17[48],stage1_16[101],stage1_15[124],stage1_14[159],stage1_13[220]}
   );
   gpc606_5 gpc614 (
      {stage0_13[471], stage0_13[472], stage0_13[473], stage0_13[474], stage0_13[475], stage0_13[476]},
      {stage0_15[294], stage0_15[295], stage0_15[296], stage0_15[297], stage0_15[298], stage0_15[299]},
      {stage1_17[49],stage1_16[102],stage1_15[125],stage1_14[160],stage1_13[221]}
   );
   gpc606_5 gpc615 (
      {stage0_13[477], stage0_13[478], stage0_13[479], stage0_13[480], stage0_13[481], stage0_13[482]},
      {stage0_15[300], stage0_15[301], stage0_15[302], stage0_15[303], stage0_15[304], stage0_15[305]},
      {stage1_17[50],stage1_16[103],stage1_15[126],stage1_14[161],stage1_13[222]}
   );
   gpc606_5 gpc616 (
      {stage0_13[483], stage0_13[484], stage0_13[485], stage0_13[486], stage0_13[487], stage0_13[488]},
      {stage0_15[306], stage0_15[307], stage0_15[308], stage0_15[309], stage0_15[310], stage0_15[311]},
      {stage1_17[51],stage1_16[104],stage1_15[127],stage1_14[162],stage1_13[223]}
   );
   gpc606_5 gpc617 (
      {stage0_13[489], stage0_13[490], stage0_13[491], stage0_13[492], stage0_13[493], stage0_13[494]},
      {stage0_15[312], stage0_15[313], stage0_15[314], stage0_15[315], stage0_15[316], stage0_15[317]},
      {stage1_17[52],stage1_16[105],stage1_15[128],stage1_14[163],stage1_13[224]}
   );
   gpc606_5 gpc618 (
      {stage0_13[495], stage0_13[496], stage0_13[497], stage0_13[498], stage0_13[499], stage0_13[500]},
      {stage0_15[318], stage0_15[319], stage0_15[320], stage0_15[321], stage0_15[322], stage0_15[323]},
      {stage1_17[53],stage1_16[106],stage1_15[129],stage1_14[164],stage1_13[225]}
   );
   gpc606_5 gpc619 (
      {stage0_13[501], stage0_13[502], stage0_13[503], stage0_13[504], stage0_13[505], stage0_13[506]},
      {stage0_15[324], stage0_15[325], stage0_15[326], stage0_15[327], stage0_15[328], stage0_15[329]},
      {stage1_17[54],stage1_16[107],stage1_15[130],stage1_14[165],stage1_13[226]}
   );
   gpc606_5 gpc620 (
      {stage0_14[318], stage0_14[319], stage0_14[320], stage0_14[321], stage0_14[322], stage0_14[323]},
      {stage0_16[0], stage0_16[1], stage0_16[2], stage0_16[3], stage0_16[4], stage0_16[5]},
      {stage1_18[0],stage1_17[55],stage1_16[108],stage1_15[131],stage1_14[166]}
   );
   gpc606_5 gpc621 (
      {stage0_14[324], stage0_14[325], stage0_14[326], stage0_14[327], stage0_14[328], stage0_14[329]},
      {stage0_16[6], stage0_16[7], stage0_16[8], stage0_16[9], stage0_16[10], stage0_16[11]},
      {stage1_18[1],stage1_17[56],stage1_16[109],stage1_15[132],stage1_14[167]}
   );
   gpc606_5 gpc622 (
      {stage0_14[330], stage0_14[331], stage0_14[332], stage0_14[333], stage0_14[334], stage0_14[335]},
      {stage0_16[12], stage0_16[13], stage0_16[14], stage0_16[15], stage0_16[16], stage0_16[17]},
      {stage1_18[2],stage1_17[57],stage1_16[110],stage1_15[133],stage1_14[168]}
   );
   gpc606_5 gpc623 (
      {stage0_14[336], stage0_14[337], stage0_14[338], stage0_14[339], stage0_14[340], stage0_14[341]},
      {stage0_16[18], stage0_16[19], stage0_16[20], stage0_16[21], stage0_16[22], stage0_16[23]},
      {stage1_18[3],stage1_17[58],stage1_16[111],stage1_15[134],stage1_14[169]}
   );
   gpc606_5 gpc624 (
      {stage0_14[342], stage0_14[343], stage0_14[344], stage0_14[345], stage0_14[346], stage0_14[347]},
      {stage0_16[24], stage0_16[25], stage0_16[26], stage0_16[27], stage0_16[28], stage0_16[29]},
      {stage1_18[4],stage1_17[59],stage1_16[112],stage1_15[135],stage1_14[170]}
   );
   gpc606_5 gpc625 (
      {stage0_14[348], stage0_14[349], stage0_14[350], stage0_14[351], stage0_14[352], stage0_14[353]},
      {stage0_16[30], stage0_16[31], stage0_16[32], stage0_16[33], stage0_16[34], stage0_16[35]},
      {stage1_18[5],stage1_17[60],stage1_16[113],stage1_15[136],stage1_14[171]}
   );
   gpc606_5 gpc626 (
      {stage0_14[354], stage0_14[355], stage0_14[356], stage0_14[357], stage0_14[358], stage0_14[359]},
      {stage0_16[36], stage0_16[37], stage0_16[38], stage0_16[39], stage0_16[40], stage0_16[41]},
      {stage1_18[6],stage1_17[61],stage1_16[114],stage1_15[137],stage1_14[172]}
   );
   gpc606_5 gpc627 (
      {stage0_14[360], stage0_14[361], stage0_14[362], stage0_14[363], stage0_14[364], stage0_14[365]},
      {stage0_16[42], stage0_16[43], stage0_16[44], stage0_16[45], stage0_16[46], stage0_16[47]},
      {stage1_18[7],stage1_17[62],stage1_16[115],stage1_15[138],stage1_14[173]}
   );
   gpc606_5 gpc628 (
      {stage0_14[366], stage0_14[367], stage0_14[368], stage0_14[369], stage0_14[370], stage0_14[371]},
      {stage0_16[48], stage0_16[49], stage0_16[50], stage0_16[51], stage0_16[52], stage0_16[53]},
      {stage1_18[8],stage1_17[63],stage1_16[116],stage1_15[139],stage1_14[174]}
   );
   gpc606_5 gpc629 (
      {stage0_14[372], stage0_14[373], stage0_14[374], stage0_14[375], stage0_14[376], stage0_14[377]},
      {stage0_16[54], stage0_16[55], stage0_16[56], stage0_16[57], stage0_16[58], stage0_16[59]},
      {stage1_18[9],stage1_17[64],stage1_16[117],stage1_15[140],stage1_14[175]}
   );
   gpc606_5 gpc630 (
      {stage0_14[378], stage0_14[379], stage0_14[380], stage0_14[381], stage0_14[382], stage0_14[383]},
      {stage0_16[60], stage0_16[61], stage0_16[62], stage0_16[63], stage0_16[64], stage0_16[65]},
      {stage1_18[10],stage1_17[65],stage1_16[118],stage1_15[141],stage1_14[176]}
   );
   gpc606_5 gpc631 (
      {stage0_14[384], stage0_14[385], stage0_14[386], stage0_14[387], stage0_14[388], stage0_14[389]},
      {stage0_16[66], stage0_16[67], stage0_16[68], stage0_16[69], stage0_16[70], stage0_16[71]},
      {stage1_18[11],stage1_17[66],stage1_16[119],stage1_15[142],stage1_14[177]}
   );
   gpc606_5 gpc632 (
      {stage0_14[390], stage0_14[391], stage0_14[392], stage0_14[393], stage0_14[394], stage0_14[395]},
      {stage0_16[72], stage0_16[73], stage0_16[74], stage0_16[75], stage0_16[76], stage0_16[77]},
      {stage1_18[12],stage1_17[67],stage1_16[120],stage1_15[143],stage1_14[178]}
   );
   gpc606_5 gpc633 (
      {stage0_14[396], stage0_14[397], stage0_14[398], stage0_14[399], stage0_14[400], stage0_14[401]},
      {stage0_16[78], stage0_16[79], stage0_16[80], stage0_16[81], stage0_16[82], stage0_16[83]},
      {stage1_18[13],stage1_17[68],stage1_16[121],stage1_15[144],stage1_14[179]}
   );
   gpc606_5 gpc634 (
      {stage0_14[402], stage0_14[403], stage0_14[404], stage0_14[405], stage0_14[406], stage0_14[407]},
      {stage0_16[84], stage0_16[85], stage0_16[86], stage0_16[87], stage0_16[88], stage0_16[89]},
      {stage1_18[14],stage1_17[69],stage1_16[122],stage1_15[145],stage1_14[180]}
   );
   gpc606_5 gpc635 (
      {stage0_14[408], stage0_14[409], stage0_14[410], stage0_14[411], stage0_14[412], stage0_14[413]},
      {stage0_16[90], stage0_16[91], stage0_16[92], stage0_16[93], stage0_16[94], stage0_16[95]},
      {stage1_18[15],stage1_17[70],stage1_16[123],stage1_15[146],stage1_14[181]}
   );
   gpc606_5 gpc636 (
      {stage0_14[414], stage0_14[415], stage0_14[416], stage0_14[417], stage0_14[418], stage0_14[419]},
      {stage0_16[96], stage0_16[97], stage0_16[98], stage0_16[99], stage0_16[100], stage0_16[101]},
      {stage1_18[16],stage1_17[71],stage1_16[124],stage1_15[147],stage1_14[182]}
   );
   gpc606_5 gpc637 (
      {stage0_14[420], stage0_14[421], stage0_14[422], stage0_14[423], stage0_14[424], stage0_14[425]},
      {stage0_16[102], stage0_16[103], stage0_16[104], stage0_16[105], stage0_16[106], stage0_16[107]},
      {stage1_18[17],stage1_17[72],stage1_16[125],stage1_15[148],stage1_14[183]}
   );
   gpc606_5 gpc638 (
      {stage0_14[426], stage0_14[427], stage0_14[428], stage0_14[429], stage0_14[430], stage0_14[431]},
      {stage0_16[108], stage0_16[109], stage0_16[110], stage0_16[111], stage0_16[112], stage0_16[113]},
      {stage1_18[18],stage1_17[73],stage1_16[126],stage1_15[149],stage1_14[184]}
   );
   gpc606_5 gpc639 (
      {stage0_14[432], stage0_14[433], stage0_14[434], stage0_14[435], stage0_14[436], stage0_14[437]},
      {stage0_16[114], stage0_16[115], stage0_16[116], stage0_16[117], stage0_16[118], stage0_16[119]},
      {stage1_18[19],stage1_17[74],stage1_16[127],stage1_15[150],stage1_14[185]}
   );
   gpc606_5 gpc640 (
      {stage0_14[438], stage0_14[439], stage0_14[440], stage0_14[441], stage0_14[442], stage0_14[443]},
      {stage0_16[120], stage0_16[121], stage0_16[122], stage0_16[123], stage0_16[124], stage0_16[125]},
      {stage1_18[20],stage1_17[75],stage1_16[128],stage1_15[151],stage1_14[186]}
   );
   gpc606_5 gpc641 (
      {stage0_14[444], stage0_14[445], stage0_14[446], stage0_14[447], stage0_14[448], stage0_14[449]},
      {stage0_16[126], stage0_16[127], stage0_16[128], stage0_16[129], stage0_16[130], stage0_16[131]},
      {stage1_18[21],stage1_17[76],stage1_16[129],stage1_15[152],stage1_14[187]}
   );
   gpc606_5 gpc642 (
      {stage0_14[450], stage0_14[451], stage0_14[452], stage0_14[453], stage0_14[454], stage0_14[455]},
      {stage0_16[132], stage0_16[133], stage0_16[134], stage0_16[135], stage0_16[136], stage0_16[137]},
      {stage1_18[22],stage1_17[77],stage1_16[130],stage1_15[153],stage1_14[188]}
   );
   gpc606_5 gpc643 (
      {stage0_14[456], stage0_14[457], stage0_14[458], stage0_14[459], stage0_14[460], stage0_14[461]},
      {stage0_16[138], stage0_16[139], stage0_16[140], stage0_16[141], stage0_16[142], stage0_16[143]},
      {stage1_18[23],stage1_17[78],stage1_16[131],stage1_15[154],stage1_14[189]}
   );
   gpc615_5 gpc644 (
      {stage0_14[462], stage0_14[463], stage0_14[464], stage0_14[465], stage0_14[466]},
      {stage0_15[330]},
      {stage0_16[144], stage0_16[145], stage0_16[146], stage0_16[147], stage0_16[148], stage0_16[149]},
      {stage1_18[24],stage1_17[79],stage1_16[132],stage1_15[155],stage1_14[190]}
   );
   gpc615_5 gpc645 (
      {stage0_14[467], stage0_14[468], stage0_14[469], stage0_14[470], stage0_14[471]},
      {stage0_15[331]},
      {stage0_16[150], stage0_16[151], stage0_16[152], stage0_16[153], stage0_16[154], stage0_16[155]},
      {stage1_18[25],stage1_17[80],stage1_16[133],stage1_15[156],stage1_14[191]}
   );
   gpc606_5 gpc646 (
      {stage0_15[332], stage0_15[333], stage0_15[334], stage0_15[335], stage0_15[336], stage0_15[337]},
      {stage0_17[0], stage0_17[1], stage0_17[2], stage0_17[3], stage0_17[4], stage0_17[5]},
      {stage1_19[0],stage1_18[26],stage1_17[81],stage1_16[134],stage1_15[157]}
   );
   gpc606_5 gpc647 (
      {stage0_15[338], stage0_15[339], stage0_15[340], stage0_15[341], stage0_15[342], stage0_15[343]},
      {stage0_17[6], stage0_17[7], stage0_17[8], stage0_17[9], stage0_17[10], stage0_17[11]},
      {stage1_19[1],stage1_18[27],stage1_17[82],stage1_16[135],stage1_15[158]}
   );
   gpc606_5 gpc648 (
      {stage0_15[344], stage0_15[345], stage0_15[346], stage0_15[347], stage0_15[348], stage0_15[349]},
      {stage0_17[12], stage0_17[13], stage0_17[14], stage0_17[15], stage0_17[16], stage0_17[17]},
      {stage1_19[2],stage1_18[28],stage1_17[83],stage1_16[136],stage1_15[159]}
   );
   gpc606_5 gpc649 (
      {stage0_15[350], stage0_15[351], stage0_15[352], stage0_15[353], stage0_15[354], stage0_15[355]},
      {stage0_17[18], stage0_17[19], stage0_17[20], stage0_17[21], stage0_17[22], stage0_17[23]},
      {stage1_19[3],stage1_18[29],stage1_17[84],stage1_16[137],stage1_15[160]}
   );
   gpc615_5 gpc650 (
      {stage0_15[356], stage0_15[357], stage0_15[358], stage0_15[359], stage0_15[360]},
      {stage0_16[156]},
      {stage0_17[24], stage0_17[25], stage0_17[26], stage0_17[27], stage0_17[28], stage0_17[29]},
      {stage1_19[4],stage1_18[30],stage1_17[85],stage1_16[138],stage1_15[161]}
   );
   gpc615_5 gpc651 (
      {stage0_15[361], stage0_15[362], stage0_15[363], stage0_15[364], stage0_15[365]},
      {stage0_16[157]},
      {stage0_17[30], stage0_17[31], stage0_17[32], stage0_17[33], stage0_17[34], stage0_17[35]},
      {stage1_19[5],stage1_18[31],stage1_17[86],stage1_16[139],stage1_15[162]}
   );
   gpc615_5 gpc652 (
      {stage0_15[366], stage0_15[367], stage0_15[368], stage0_15[369], stage0_15[370]},
      {stage0_16[158]},
      {stage0_17[36], stage0_17[37], stage0_17[38], stage0_17[39], stage0_17[40], stage0_17[41]},
      {stage1_19[6],stage1_18[32],stage1_17[87],stage1_16[140],stage1_15[163]}
   );
   gpc615_5 gpc653 (
      {stage0_15[371], stage0_15[372], stage0_15[373], stage0_15[374], stage0_15[375]},
      {stage0_16[159]},
      {stage0_17[42], stage0_17[43], stage0_17[44], stage0_17[45], stage0_17[46], stage0_17[47]},
      {stage1_19[7],stage1_18[33],stage1_17[88],stage1_16[141],stage1_15[164]}
   );
   gpc615_5 gpc654 (
      {stage0_15[376], stage0_15[377], stage0_15[378], stage0_15[379], stage0_15[380]},
      {stage0_16[160]},
      {stage0_17[48], stage0_17[49], stage0_17[50], stage0_17[51], stage0_17[52], stage0_17[53]},
      {stage1_19[8],stage1_18[34],stage1_17[89],stage1_16[142],stage1_15[165]}
   );
   gpc615_5 gpc655 (
      {stage0_15[381], stage0_15[382], stage0_15[383], stage0_15[384], stage0_15[385]},
      {stage0_16[161]},
      {stage0_17[54], stage0_17[55], stage0_17[56], stage0_17[57], stage0_17[58], stage0_17[59]},
      {stage1_19[9],stage1_18[35],stage1_17[90],stage1_16[143],stage1_15[166]}
   );
   gpc615_5 gpc656 (
      {stage0_15[386], stage0_15[387], stage0_15[388], stage0_15[389], stage0_15[390]},
      {stage0_16[162]},
      {stage0_17[60], stage0_17[61], stage0_17[62], stage0_17[63], stage0_17[64], stage0_17[65]},
      {stage1_19[10],stage1_18[36],stage1_17[91],stage1_16[144],stage1_15[167]}
   );
   gpc615_5 gpc657 (
      {stage0_15[391], stage0_15[392], stage0_15[393], stage0_15[394], stage0_15[395]},
      {stage0_16[163]},
      {stage0_17[66], stage0_17[67], stage0_17[68], stage0_17[69], stage0_17[70], stage0_17[71]},
      {stage1_19[11],stage1_18[37],stage1_17[92],stage1_16[145],stage1_15[168]}
   );
   gpc615_5 gpc658 (
      {stage0_15[396], stage0_15[397], stage0_15[398], stage0_15[399], stage0_15[400]},
      {stage0_16[164]},
      {stage0_17[72], stage0_17[73], stage0_17[74], stage0_17[75], stage0_17[76], stage0_17[77]},
      {stage1_19[12],stage1_18[38],stage1_17[93],stage1_16[146],stage1_15[169]}
   );
   gpc615_5 gpc659 (
      {stage0_15[401], stage0_15[402], stage0_15[403], stage0_15[404], stage0_15[405]},
      {stage0_16[165]},
      {stage0_17[78], stage0_17[79], stage0_17[80], stage0_17[81], stage0_17[82], stage0_17[83]},
      {stage1_19[13],stage1_18[39],stage1_17[94],stage1_16[147],stage1_15[170]}
   );
   gpc615_5 gpc660 (
      {stage0_15[406], stage0_15[407], stage0_15[408], stage0_15[409], stage0_15[410]},
      {stage0_16[166]},
      {stage0_17[84], stage0_17[85], stage0_17[86], stage0_17[87], stage0_17[88], stage0_17[89]},
      {stage1_19[14],stage1_18[40],stage1_17[95],stage1_16[148],stage1_15[171]}
   );
   gpc615_5 gpc661 (
      {stage0_15[411], stage0_15[412], stage0_15[413], stage0_15[414], stage0_15[415]},
      {stage0_16[167]},
      {stage0_17[90], stage0_17[91], stage0_17[92], stage0_17[93], stage0_17[94], stage0_17[95]},
      {stage1_19[15],stage1_18[41],stage1_17[96],stage1_16[149],stage1_15[172]}
   );
   gpc615_5 gpc662 (
      {stage0_15[416], stage0_15[417], stage0_15[418], stage0_15[419], stage0_15[420]},
      {stage0_16[168]},
      {stage0_17[96], stage0_17[97], stage0_17[98], stage0_17[99], stage0_17[100], stage0_17[101]},
      {stage1_19[16],stage1_18[42],stage1_17[97],stage1_16[150],stage1_15[173]}
   );
   gpc615_5 gpc663 (
      {stage0_15[421], stage0_15[422], stage0_15[423], stage0_15[424], stage0_15[425]},
      {stage0_16[169]},
      {stage0_17[102], stage0_17[103], stage0_17[104], stage0_17[105], stage0_17[106], stage0_17[107]},
      {stage1_19[17],stage1_18[43],stage1_17[98],stage1_16[151],stage1_15[174]}
   );
   gpc615_5 gpc664 (
      {stage0_15[426], stage0_15[427], stage0_15[428], stage0_15[429], stage0_15[430]},
      {stage0_16[170]},
      {stage0_17[108], stage0_17[109], stage0_17[110], stage0_17[111], stage0_17[112], stage0_17[113]},
      {stage1_19[18],stage1_18[44],stage1_17[99],stage1_16[152],stage1_15[175]}
   );
   gpc615_5 gpc665 (
      {stage0_15[431], stage0_15[432], stage0_15[433], stage0_15[434], stage0_15[435]},
      {stage0_16[171]},
      {stage0_17[114], stage0_17[115], stage0_17[116], stage0_17[117], stage0_17[118], stage0_17[119]},
      {stage1_19[19],stage1_18[45],stage1_17[100],stage1_16[153],stage1_15[176]}
   );
   gpc615_5 gpc666 (
      {stage0_15[436], stage0_15[437], stage0_15[438], stage0_15[439], stage0_15[440]},
      {stage0_16[172]},
      {stage0_17[120], stage0_17[121], stage0_17[122], stage0_17[123], stage0_17[124], stage0_17[125]},
      {stage1_19[20],stage1_18[46],stage1_17[101],stage1_16[154],stage1_15[177]}
   );
   gpc615_5 gpc667 (
      {stage0_15[441], stage0_15[442], stage0_15[443], stage0_15[444], stage0_15[445]},
      {stage0_16[173]},
      {stage0_17[126], stage0_17[127], stage0_17[128], stage0_17[129], stage0_17[130], stage0_17[131]},
      {stage1_19[21],stage1_18[47],stage1_17[102],stage1_16[155],stage1_15[178]}
   );
   gpc615_5 gpc668 (
      {stage0_15[446], stage0_15[447], stage0_15[448], stage0_15[449], stage0_15[450]},
      {stage0_16[174]},
      {stage0_17[132], stage0_17[133], stage0_17[134], stage0_17[135], stage0_17[136], stage0_17[137]},
      {stage1_19[22],stage1_18[48],stage1_17[103],stage1_16[156],stage1_15[179]}
   );
   gpc615_5 gpc669 (
      {stage0_15[451], stage0_15[452], stage0_15[453], stage0_15[454], stage0_15[455]},
      {stage0_16[175]},
      {stage0_17[138], stage0_17[139], stage0_17[140], stage0_17[141], stage0_17[142], stage0_17[143]},
      {stage1_19[23],stage1_18[49],stage1_17[104],stage1_16[157],stage1_15[180]}
   );
   gpc606_5 gpc670 (
      {stage0_16[176], stage0_16[177], stage0_16[178], stage0_16[179], stage0_16[180], stage0_16[181]},
      {stage0_18[0], stage0_18[1], stage0_18[2], stage0_18[3], stage0_18[4], stage0_18[5]},
      {stage1_20[0],stage1_19[24],stage1_18[50],stage1_17[105],stage1_16[158]}
   );
   gpc606_5 gpc671 (
      {stage0_16[182], stage0_16[183], stage0_16[184], stage0_16[185], stage0_16[186], stage0_16[187]},
      {stage0_18[6], stage0_18[7], stage0_18[8], stage0_18[9], stage0_18[10], stage0_18[11]},
      {stage1_20[1],stage1_19[25],stage1_18[51],stage1_17[106],stage1_16[159]}
   );
   gpc606_5 gpc672 (
      {stage0_16[188], stage0_16[189], stage0_16[190], stage0_16[191], stage0_16[192], stage0_16[193]},
      {stage0_18[12], stage0_18[13], stage0_18[14], stage0_18[15], stage0_18[16], stage0_18[17]},
      {stage1_20[2],stage1_19[26],stage1_18[52],stage1_17[107],stage1_16[160]}
   );
   gpc606_5 gpc673 (
      {stage0_16[194], stage0_16[195], stage0_16[196], stage0_16[197], stage0_16[198], stage0_16[199]},
      {stage0_18[18], stage0_18[19], stage0_18[20], stage0_18[21], stage0_18[22], stage0_18[23]},
      {stage1_20[3],stage1_19[27],stage1_18[53],stage1_17[108],stage1_16[161]}
   );
   gpc606_5 gpc674 (
      {stage0_16[200], stage0_16[201], stage0_16[202], stage0_16[203], stage0_16[204], stage0_16[205]},
      {stage0_18[24], stage0_18[25], stage0_18[26], stage0_18[27], stage0_18[28], stage0_18[29]},
      {stage1_20[4],stage1_19[28],stage1_18[54],stage1_17[109],stage1_16[162]}
   );
   gpc606_5 gpc675 (
      {stage0_16[206], stage0_16[207], stage0_16[208], stage0_16[209], stage0_16[210], stage0_16[211]},
      {stage0_18[30], stage0_18[31], stage0_18[32], stage0_18[33], stage0_18[34], stage0_18[35]},
      {stage1_20[5],stage1_19[29],stage1_18[55],stage1_17[110],stage1_16[163]}
   );
   gpc606_5 gpc676 (
      {stage0_16[212], stage0_16[213], stage0_16[214], stage0_16[215], stage0_16[216], stage0_16[217]},
      {stage0_18[36], stage0_18[37], stage0_18[38], stage0_18[39], stage0_18[40], stage0_18[41]},
      {stage1_20[6],stage1_19[30],stage1_18[56],stage1_17[111],stage1_16[164]}
   );
   gpc606_5 gpc677 (
      {stage0_16[218], stage0_16[219], stage0_16[220], stage0_16[221], stage0_16[222], stage0_16[223]},
      {stage0_18[42], stage0_18[43], stage0_18[44], stage0_18[45], stage0_18[46], stage0_18[47]},
      {stage1_20[7],stage1_19[31],stage1_18[57],stage1_17[112],stage1_16[165]}
   );
   gpc606_5 gpc678 (
      {stage0_16[224], stage0_16[225], stage0_16[226], stage0_16[227], stage0_16[228], stage0_16[229]},
      {stage0_18[48], stage0_18[49], stage0_18[50], stage0_18[51], stage0_18[52], stage0_18[53]},
      {stage1_20[8],stage1_19[32],stage1_18[58],stage1_17[113],stage1_16[166]}
   );
   gpc606_5 gpc679 (
      {stage0_16[230], stage0_16[231], stage0_16[232], stage0_16[233], stage0_16[234], stage0_16[235]},
      {stage0_18[54], stage0_18[55], stage0_18[56], stage0_18[57], stage0_18[58], stage0_18[59]},
      {stage1_20[9],stage1_19[33],stage1_18[59],stage1_17[114],stage1_16[167]}
   );
   gpc606_5 gpc680 (
      {stage0_16[236], stage0_16[237], stage0_16[238], stage0_16[239], stage0_16[240], stage0_16[241]},
      {stage0_18[60], stage0_18[61], stage0_18[62], stage0_18[63], stage0_18[64], stage0_18[65]},
      {stage1_20[10],stage1_19[34],stage1_18[60],stage1_17[115],stage1_16[168]}
   );
   gpc606_5 gpc681 (
      {stage0_16[242], stage0_16[243], stage0_16[244], stage0_16[245], stage0_16[246], stage0_16[247]},
      {stage0_18[66], stage0_18[67], stage0_18[68], stage0_18[69], stage0_18[70], stage0_18[71]},
      {stage1_20[11],stage1_19[35],stage1_18[61],stage1_17[116],stage1_16[169]}
   );
   gpc606_5 gpc682 (
      {stage0_16[248], stage0_16[249], stage0_16[250], stage0_16[251], stage0_16[252], stage0_16[253]},
      {stage0_18[72], stage0_18[73], stage0_18[74], stage0_18[75], stage0_18[76], stage0_18[77]},
      {stage1_20[12],stage1_19[36],stage1_18[62],stage1_17[117],stage1_16[170]}
   );
   gpc606_5 gpc683 (
      {stage0_16[254], stage0_16[255], stage0_16[256], stage0_16[257], stage0_16[258], stage0_16[259]},
      {stage0_18[78], stage0_18[79], stage0_18[80], stage0_18[81], stage0_18[82], stage0_18[83]},
      {stage1_20[13],stage1_19[37],stage1_18[63],stage1_17[118],stage1_16[171]}
   );
   gpc606_5 gpc684 (
      {stage0_16[260], stage0_16[261], stage0_16[262], stage0_16[263], stage0_16[264], stage0_16[265]},
      {stage0_18[84], stage0_18[85], stage0_18[86], stage0_18[87], stage0_18[88], stage0_18[89]},
      {stage1_20[14],stage1_19[38],stage1_18[64],stage1_17[119],stage1_16[172]}
   );
   gpc606_5 gpc685 (
      {stage0_16[266], stage0_16[267], stage0_16[268], stage0_16[269], stage0_16[270], stage0_16[271]},
      {stage0_18[90], stage0_18[91], stage0_18[92], stage0_18[93], stage0_18[94], stage0_18[95]},
      {stage1_20[15],stage1_19[39],stage1_18[65],stage1_17[120],stage1_16[173]}
   );
   gpc606_5 gpc686 (
      {stage0_16[272], stage0_16[273], stage0_16[274], stage0_16[275], stage0_16[276], stage0_16[277]},
      {stage0_18[96], stage0_18[97], stage0_18[98], stage0_18[99], stage0_18[100], stage0_18[101]},
      {stage1_20[16],stage1_19[40],stage1_18[66],stage1_17[121],stage1_16[174]}
   );
   gpc606_5 gpc687 (
      {stage0_16[278], stage0_16[279], stage0_16[280], stage0_16[281], stage0_16[282], stage0_16[283]},
      {stage0_18[102], stage0_18[103], stage0_18[104], stage0_18[105], stage0_18[106], stage0_18[107]},
      {stage1_20[17],stage1_19[41],stage1_18[67],stage1_17[122],stage1_16[175]}
   );
   gpc606_5 gpc688 (
      {stage0_16[284], stage0_16[285], stage0_16[286], stage0_16[287], stage0_16[288], stage0_16[289]},
      {stage0_18[108], stage0_18[109], stage0_18[110], stage0_18[111], stage0_18[112], stage0_18[113]},
      {stage1_20[18],stage1_19[42],stage1_18[68],stage1_17[123],stage1_16[176]}
   );
   gpc606_5 gpc689 (
      {stage0_16[290], stage0_16[291], stage0_16[292], stage0_16[293], stage0_16[294], stage0_16[295]},
      {stage0_18[114], stage0_18[115], stage0_18[116], stage0_18[117], stage0_18[118], stage0_18[119]},
      {stage1_20[19],stage1_19[43],stage1_18[69],stage1_17[124],stage1_16[177]}
   );
   gpc606_5 gpc690 (
      {stage0_16[296], stage0_16[297], stage0_16[298], stage0_16[299], stage0_16[300], stage0_16[301]},
      {stage0_18[120], stage0_18[121], stage0_18[122], stage0_18[123], stage0_18[124], stage0_18[125]},
      {stage1_20[20],stage1_19[44],stage1_18[70],stage1_17[125],stage1_16[178]}
   );
   gpc606_5 gpc691 (
      {stage0_16[302], stage0_16[303], stage0_16[304], stage0_16[305], stage0_16[306], stage0_16[307]},
      {stage0_18[126], stage0_18[127], stage0_18[128], stage0_18[129], stage0_18[130], stage0_18[131]},
      {stage1_20[21],stage1_19[45],stage1_18[71],stage1_17[126],stage1_16[179]}
   );
   gpc606_5 gpc692 (
      {stage0_16[308], stage0_16[309], stage0_16[310], stage0_16[311], stage0_16[312], stage0_16[313]},
      {stage0_18[132], stage0_18[133], stage0_18[134], stage0_18[135], stage0_18[136], stage0_18[137]},
      {stage1_20[22],stage1_19[46],stage1_18[72],stage1_17[127],stage1_16[180]}
   );
   gpc606_5 gpc693 (
      {stage0_16[314], stage0_16[315], stage0_16[316], stage0_16[317], stage0_16[318], stage0_16[319]},
      {stage0_18[138], stage0_18[139], stage0_18[140], stage0_18[141], stage0_18[142], stage0_18[143]},
      {stage1_20[23],stage1_19[47],stage1_18[73],stage1_17[128],stage1_16[181]}
   );
   gpc606_5 gpc694 (
      {stage0_16[320], stage0_16[321], stage0_16[322], stage0_16[323], stage0_16[324], stage0_16[325]},
      {stage0_18[144], stage0_18[145], stage0_18[146], stage0_18[147], stage0_18[148], stage0_18[149]},
      {stage1_20[24],stage1_19[48],stage1_18[74],stage1_17[129],stage1_16[182]}
   );
   gpc606_5 gpc695 (
      {stage0_16[326], stage0_16[327], stage0_16[328], stage0_16[329], stage0_16[330], stage0_16[331]},
      {stage0_18[150], stage0_18[151], stage0_18[152], stage0_18[153], stage0_18[154], stage0_18[155]},
      {stage1_20[25],stage1_19[49],stage1_18[75],stage1_17[130],stage1_16[183]}
   );
   gpc606_5 gpc696 (
      {stage0_16[332], stage0_16[333], stage0_16[334], stage0_16[335], stage0_16[336], stage0_16[337]},
      {stage0_18[156], stage0_18[157], stage0_18[158], stage0_18[159], stage0_18[160], stage0_18[161]},
      {stage1_20[26],stage1_19[50],stage1_18[76],stage1_17[131],stage1_16[184]}
   );
   gpc606_5 gpc697 (
      {stage0_16[338], stage0_16[339], stage0_16[340], stage0_16[341], stage0_16[342], stage0_16[343]},
      {stage0_18[162], stage0_18[163], stage0_18[164], stage0_18[165], stage0_18[166], stage0_18[167]},
      {stage1_20[27],stage1_19[51],stage1_18[77],stage1_17[132],stage1_16[185]}
   );
   gpc606_5 gpc698 (
      {stage0_16[344], stage0_16[345], stage0_16[346], stage0_16[347], stage0_16[348], stage0_16[349]},
      {stage0_18[168], stage0_18[169], stage0_18[170], stage0_18[171], stage0_18[172], stage0_18[173]},
      {stage1_20[28],stage1_19[52],stage1_18[78],stage1_17[133],stage1_16[186]}
   );
   gpc606_5 gpc699 (
      {stage0_16[350], stage0_16[351], stage0_16[352], stage0_16[353], stage0_16[354], stage0_16[355]},
      {stage0_18[174], stage0_18[175], stage0_18[176], stage0_18[177], stage0_18[178], stage0_18[179]},
      {stage1_20[29],stage1_19[53],stage1_18[79],stage1_17[134],stage1_16[187]}
   );
   gpc606_5 gpc700 (
      {stage0_16[356], stage0_16[357], stage0_16[358], stage0_16[359], stage0_16[360], stage0_16[361]},
      {stage0_18[180], stage0_18[181], stage0_18[182], stage0_18[183], stage0_18[184], stage0_18[185]},
      {stage1_20[30],stage1_19[54],stage1_18[80],stage1_17[135],stage1_16[188]}
   );
   gpc606_5 gpc701 (
      {stage0_16[362], stage0_16[363], stage0_16[364], stage0_16[365], stage0_16[366], stage0_16[367]},
      {stage0_18[186], stage0_18[187], stage0_18[188], stage0_18[189], stage0_18[190], stage0_18[191]},
      {stage1_20[31],stage1_19[55],stage1_18[81],stage1_17[136],stage1_16[189]}
   );
   gpc606_5 gpc702 (
      {stage0_16[368], stage0_16[369], stage0_16[370], stage0_16[371], stage0_16[372], stage0_16[373]},
      {stage0_18[192], stage0_18[193], stage0_18[194], stage0_18[195], stage0_18[196], stage0_18[197]},
      {stage1_20[32],stage1_19[56],stage1_18[82],stage1_17[137],stage1_16[190]}
   );
   gpc606_5 gpc703 (
      {stage0_16[374], stage0_16[375], stage0_16[376], stage0_16[377], stage0_16[378], stage0_16[379]},
      {stage0_18[198], stage0_18[199], stage0_18[200], stage0_18[201], stage0_18[202], stage0_18[203]},
      {stage1_20[33],stage1_19[57],stage1_18[83],stage1_17[138],stage1_16[191]}
   );
   gpc606_5 gpc704 (
      {stage0_16[380], stage0_16[381], stage0_16[382], stage0_16[383], stage0_16[384], stage0_16[385]},
      {stage0_18[204], stage0_18[205], stage0_18[206], stage0_18[207], stage0_18[208], stage0_18[209]},
      {stage1_20[34],stage1_19[58],stage1_18[84],stage1_17[139],stage1_16[192]}
   );
   gpc606_5 gpc705 (
      {stage0_16[386], stage0_16[387], stage0_16[388], stage0_16[389], stage0_16[390], stage0_16[391]},
      {stage0_18[210], stage0_18[211], stage0_18[212], stage0_18[213], stage0_18[214], stage0_18[215]},
      {stage1_20[35],stage1_19[59],stage1_18[85],stage1_17[140],stage1_16[193]}
   );
   gpc606_5 gpc706 (
      {stage0_16[392], stage0_16[393], stage0_16[394], stage0_16[395], stage0_16[396], stage0_16[397]},
      {stage0_18[216], stage0_18[217], stage0_18[218], stage0_18[219], stage0_18[220], stage0_18[221]},
      {stage1_20[36],stage1_19[60],stage1_18[86],stage1_17[141],stage1_16[194]}
   );
   gpc606_5 gpc707 (
      {stage0_16[398], stage0_16[399], stage0_16[400], stage0_16[401], stage0_16[402], stage0_16[403]},
      {stage0_18[222], stage0_18[223], stage0_18[224], stage0_18[225], stage0_18[226], stage0_18[227]},
      {stage1_20[37],stage1_19[61],stage1_18[87],stage1_17[142],stage1_16[195]}
   );
   gpc606_5 gpc708 (
      {stage0_16[404], stage0_16[405], stage0_16[406], stage0_16[407], stage0_16[408], stage0_16[409]},
      {stage0_18[228], stage0_18[229], stage0_18[230], stage0_18[231], stage0_18[232], stage0_18[233]},
      {stage1_20[38],stage1_19[62],stage1_18[88],stage1_17[143],stage1_16[196]}
   );
   gpc606_5 gpc709 (
      {stage0_16[410], stage0_16[411], stage0_16[412], stage0_16[413], stage0_16[414], stage0_16[415]},
      {stage0_18[234], stage0_18[235], stage0_18[236], stage0_18[237], stage0_18[238], stage0_18[239]},
      {stage1_20[39],stage1_19[63],stage1_18[89],stage1_17[144],stage1_16[197]}
   );
   gpc606_5 gpc710 (
      {stage0_16[416], stage0_16[417], stage0_16[418], stage0_16[419], stage0_16[420], stage0_16[421]},
      {stage0_18[240], stage0_18[241], stage0_18[242], stage0_18[243], stage0_18[244], stage0_18[245]},
      {stage1_20[40],stage1_19[64],stage1_18[90],stage1_17[145],stage1_16[198]}
   );
   gpc606_5 gpc711 (
      {stage0_16[422], stage0_16[423], stage0_16[424], stage0_16[425], stage0_16[426], stage0_16[427]},
      {stage0_18[246], stage0_18[247], stage0_18[248], stage0_18[249], stage0_18[250], stage0_18[251]},
      {stage1_20[41],stage1_19[65],stage1_18[91],stage1_17[146],stage1_16[199]}
   );
   gpc606_5 gpc712 (
      {stage0_16[428], stage0_16[429], stage0_16[430], stage0_16[431], stage0_16[432], stage0_16[433]},
      {stage0_18[252], stage0_18[253], stage0_18[254], stage0_18[255], stage0_18[256], stage0_18[257]},
      {stage1_20[42],stage1_19[66],stage1_18[92],stage1_17[147],stage1_16[200]}
   );
   gpc606_5 gpc713 (
      {stage0_16[434], stage0_16[435], stage0_16[436], stage0_16[437], stage0_16[438], stage0_16[439]},
      {stage0_18[258], stage0_18[259], stage0_18[260], stage0_18[261], stage0_18[262], stage0_18[263]},
      {stage1_20[43],stage1_19[67],stage1_18[93],stage1_17[148],stage1_16[201]}
   );
   gpc606_5 gpc714 (
      {stage0_16[440], stage0_16[441], stage0_16[442], stage0_16[443], stage0_16[444], stage0_16[445]},
      {stage0_18[264], stage0_18[265], stage0_18[266], stage0_18[267], stage0_18[268], stage0_18[269]},
      {stage1_20[44],stage1_19[68],stage1_18[94],stage1_17[149],stage1_16[202]}
   );
   gpc606_5 gpc715 (
      {stage0_16[446], stage0_16[447], stage0_16[448], stage0_16[449], stage0_16[450], stage0_16[451]},
      {stage0_18[270], stage0_18[271], stage0_18[272], stage0_18[273], stage0_18[274], stage0_18[275]},
      {stage1_20[45],stage1_19[69],stage1_18[95],stage1_17[150],stage1_16[203]}
   );
   gpc606_5 gpc716 (
      {stage0_16[452], stage0_16[453], stage0_16[454], stage0_16[455], stage0_16[456], stage0_16[457]},
      {stage0_18[276], stage0_18[277], stage0_18[278], stage0_18[279], stage0_18[280], stage0_18[281]},
      {stage1_20[46],stage1_19[70],stage1_18[96],stage1_17[151],stage1_16[204]}
   );
   gpc606_5 gpc717 (
      {stage0_16[458], stage0_16[459], stage0_16[460], stage0_16[461], stage0_16[462], stage0_16[463]},
      {stage0_18[282], stage0_18[283], stage0_18[284], stage0_18[285], stage0_18[286], stage0_18[287]},
      {stage1_20[47],stage1_19[71],stage1_18[97],stage1_17[152],stage1_16[205]}
   );
   gpc606_5 gpc718 (
      {stage0_16[464], stage0_16[465], stage0_16[466], stage0_16[467], stage0_16[468], stage0_16[469]},
      {stage0_18[288], stage0_18[289], stage0_18[290], stage0_18[291], stage0_18[292], stage0_18[293]},
      {stage1_20[48],stage1_19[72],stage1_18[98],stage1_17[153],stage1_16[206]}
   );
   gpc606_5 gpc719 (
      {stage0_16[470], stage0_16[471], stage0_16[472], stage0_16[473], stage0_16[474], stage0_16[475]},
      {stage0_18[294], stage0_18[295], stage0_18[296], stage0_18[297], stage0_18[298], stage0_18[299]},
      {stage1_20[49],stage1_19[73],stage1_18[99],stage1_17[154],stage1_16[207]}
   );
   gpc606_5 gpc720 (
      {stage0_16[476], stage0_16[477], stage0_16[478], stage0_16[479], stage0_16[480], stage0_16[481]},
      {stage0_18[300], stage0_18[301], stage0_18[302], stage0_18[303], stage0_18[304], stage0_18[305]},
      {stage1_20[50],stage1_19[74],stage1_18[100],stage1_17[155],stage1_16[208]}
   );
   gpc606_5 gpc721 (
      {stage0_16[482], stage0_16[483], stage0_16[484], stage0_16[485], stage0_16[486], stage0_16[487]},
      {stage0_18[306], stage0_18[307], stage0_18[308], stage0_18[309], stage0_18[310], stage0_18[311]},
      {stage1_20[51],stage1_19[75],stage1_18[101],stage1_17[156],stage1_16[209]}
   );
   gpc606_5 gpc722 (
      {stage0_16[488], stage0_16[489], stage0_16[490], stage0_16[491], stage0_16[492], stage0_16[493]},
      {stage0_18[312], stage0_18[313], stage0_18[314], stage0_18[315], stage0_18[316], stage0_18[317]},
      {stage1_20[52],stage1_19[76],stage1_18[102],stage1_17[157],stage1_16[210]}
   );
   gpc606_5 gpc723 (
      {stage0_16[494], stage0_16[495], stage0_16[496], stage0_16[497], stage0_16[498], stage0_16[499]},
      {stage0_18[318], stage0_18[319], stage0_18[320], stage0_18[321], stage0_18[322], stage0_18[323]},
      {stage1_20[53],stage1_19[77],stage1_18[103],stage1_17[158],stage1_16[211]}
   );
   gpc606_5 gpc724 (
      {stage0_16[500], stage0_16[501], stage0_16[502], stage0_16[503], stage0_16[504], stage0_16[505]},
      {stage0_18[324], stage0_18[325], stage0_18[326], stage0_18[327], stage0_18[328], stage0_18[329]},
      {stage1_20[54],stage1_19[78],stage1_18[104],stage1_17[159],stage1_16[212]}
   );
   gpc606_5 gpc725 (
      {stage0_16[506], stage0_16[507], stage0_16[508], stage0_16[509], stage0_16[510], stage0_16[511]},
      {stage0_18[330], stage0_18[331], stage0_18[332], stage0_18[333], stage0_18[334], stage0_18[335]},
      {stage1_20[55],stage1_19[79],stage1_18[105],stage1_17[160],stage1_16[213]}
   );
   gpc606_5 gpc726 (
      {stage0_17[144], stage0_17[145], stage0_17[146], stage0_17[147], stage0_17[148], stage0_17[149]},
      {stage0_19[0], stage0_19[1], stage0_19[2], stage0_19[3], stage0_19[4], stage0_19[5]},
      {stage1_21[0],stage1_20[56],stage1_19[80],stage1_18[106],stage1_17[161]}
   );
   gpc606_5 gpc727 (
      {stage0_17[150], stage0_17[151], stage0_17[152], stage0_17[153], stage0_17[154], stage0_17[155]},
      {stage0_19[6], stage0_19[7], stage0_19[8], stage0_19[9], stage0_19[10], stage0_19[11]},
      {stage1_21[1],stage1_20[57],stage1_19[81],stage1_18[107],stage1_17[162]}
   );
   gpc606_5 gpc728 (
      {stage0_17[156], stage0_17[157], stage0_17[158], stage0_17[159], stage0_17[160], stage0_17[161]},
      {stage0_19[12], stage0_19[13], stage0_19[14], stage0_19[15], stage0_19[16], stage0_19[17]},
      {stage1_21[2],stage1_20[58],stage1_19[82],stage1_18[108],stage1_17[163]}
   );
   gpc606_5 gpc729 (
      {stage0_17[162], stage0_17[163], stage0_17[164], stage0_17[165], stage0_17[166], stage0_17[167]},
      {stage0_19[18], stage0_19[19], stage0_19[20], stage0_19[21], stage0_19[22], stage0_19[23]},
      {stage1_21[3],stage1_20[59],stage1_19[83],stage1_18[109],stage1_17[164]}
   );
   gpc606_5 gpc730 (
      {stage0_17[168], stage0_17[169], stage0_17[170], stage0_17[171], stage0_17[172], stage0_17[173]},
      {stage0_19[24], stage0_19[25], stage0_19[26], stage0_19[27], stage0_19[28], stage0_19[29]},
      {stage1_21[4],stage1_20[60],stage1_19[84],stage1_18[110],stage1_17[165]}
   );
   gpc606_5 gpc731 (
      {stage0_17[174], stage0_17[175], stage0_17[176], stage0_17[177], stage0_17[178], stage0_17[179]},
      {stage0_19[30], stage0_19[31], stage0_19[32], stage0_19[33], stage0_19[34], stage0_19[35]},
      {stage1_21[5],stage1_20[61],stage1_19[85],stage1_18[111],stage1_17[166]}
   );
   gpc606_5 gpc732 (
      {stage0_17[180], stage0_17[181], stage0_17[182], stage0_17[183], stage0_17[184], stage0_17[185]},
      {stage0_19[36], stage0_19[37], stage0_19[38], stage0_19[39], stage0_19[40], stage0_19[41]},
      {stage1_21[6],stage1_20[62],stage1_19[86],stage1_18[112],stage1_17[167]}
   );
   gpc606_5 gpc733 (
      {stage0_17[186], stage0_17[187], stage0_17[188], stage0_17[189], stage0_17[190], stage0_17[191]},
      {stage0_19[42], stage0_19[43], stage0_19[44], stage0_19[45], stage0_19[46], stage0_19[47]},
      {stage1_21[7],stage1_20[63],stage1_19[87],stage1_18[113],stage1_17[168]}
   );
   gpc606_5 gpc734 (
      {stage0_17[192], stage0_17[193], stage0_17[194], stage0_17[195], stage0_17[196], stage0_17[197]},
      {stage0_19[48], stage0_19[49], stage0_19[50], stage0_19[51], stage0_19[52], stage0_19[53]},
      {stage1_21[8],stage1_20[64],stage1_19[88],stage1_18[114],stage1_17[169]}
   );
   gpc606_5 gpc735 (
      {stage0_17[198], stage0_17[199], stage0_17[200], stage0_17[201], stage0_17[202], stage0_17[203]},
      {stage0_19[54], stage0_19[55], stage0_19[56], stage0_19[57], stage0_19[58], stage0_19[59]},
      {stage1_21[9],stage1_20[65],stage1_19[89],stage1_18[115],stage1_17[170]}
   );
   gpc606_5 gpc736 (
      {stage0_17[204], stage0_17[205], stage0_17[206], stage0_17[207], stage0_17[208], stage0_17[209]},
      {stage0_19[60], stage0_19[61], stage0_19[62], stage0_19[63], stage0_19[64], stage0_19[65]},
      {stage1_21[10],stage1_20[66],stage1_19[90],stage1_18[116],stage1_17[171]}
   );
   gpc606_5 gpc737 (
      {stage0_17[210], stage0_17[211], stage0_17[212], stage0_17[213], stage0_17[214], stage0_17[215]},
      {stage0_19[66], stage0_19[67], stage0_19[68], stage0_19[69], stage0_19[70], stage0_19[71]},
      {stage1_21[11],stage1_20[67],stage1_19[91],stage1_18[117],stage1_17[172]}
   );
   gpc606_5 gpc738 (
      {stage0_17[216], stage0_17[217], stage0_17[218], stage0_17[219], stage0_17[220], stage0_17[221]},
      {stage0_19[72], stage0_19[73], stage0_19[74], stage0_19[75], stage0_19[76], stage0_19[77]},
      {stage1_21[12],stage1_20[68],stage1_19[92],stage1_18[118],stage1_17[173]}
   );
   gpc606_5 gpc739 (
      {stage0_17[222], stage0_17[223], stage0_17[224], stage0_17[225], stage0_17[226], stage0_17[227]},
      {stage0_19[78], stage0_19[79], stage0_19[80], stage0_19[81], stage0_19[82], stage0_19[83]},
      {stage1_21[13],stage1_20[69],stage1_19[93],stage1_18[119],stage1_17[174]}
   );
   gpc606_5 gpc740 (
      {stage0_17[228], stage0_17[229], stage0_17[230], stage0_17[231], stage0_17[232], stage0_17[233]},
      {stage0_19[84], stage0_19[85], stage0_19[86], stage0_19[87], stage0_19[88], stage0_19[89]},
      {stage1_21[14],stage1_20[70],stage1_19[94],stage1_18[120],stage1_17[175]}
   );
   gpc606_5 gpc741 (
      {stage0_17[234], stage0_17[235], stage0_17[236], stage0_17[237], stage0_17[238], stage0_17[239]},
      {stage0_19[90], stage0_19[91], stage0_19[92], stage0_19[93], stage0_19[94], stage0_19[95]},
      {stage1_21[15],stage1_20[71],stage1_19[95],stage1_18[121],stage1_17[176]}
   );
   gpc606_5 gpc742 (
      {stage0_17[240], stage0_17[241], stage0_17[242], stage0_17[243], stage0_17[244], stage0_17[245]},
      {stage0_19[96], stage0_19[97], stage0_19[98], stage0_19[99], stage0_19[100], stage0_19[101]},
      {stage1_21[16],stage1_20[72],stage1_19[96],stage1_18[122],stage1_17[177]}
   );
   gpc606_5 gpc743 (
      {stage0_17[246], stage0_17[247], stage0_17[248], stage0_17[249], stage0_17[250], stage0_17[251]},
      {stage0_19[102], stage0_19[103], stage0_19[104], stage0_19[105], stage0_19[106], stage0_19[107]},
      {stage1_21[17],stage1_20[73],stage1_19[97],stage1_18[123],stage1_17[178]}
   );
   gpc606_5 gpc744 (
      {stage0_17[252], stage0_17[253], stage0_17[254], stage0_17[255], stage0_17[256], stage0_17[257]},
      {stage0_19[108], stage0_19[109], stage0_19[110], stage0_19[111], stage0_19[112], stage0_19[113]},
      {stage1_21[18],stage1_20[74],stage1_19[98],stage1_18[124],stage1_17[179]}
   );
   gpc606_5 gpc745 (
      {stage0_17[258], stage0_17[259], stage0_17[260], stage0_17[261], stage0_17[262], stage0_17[263]},
      {stage0_19[114], stage0_19[115], stage0_19[116], stage0_19[117], stage0_19[118], stage0_19[119]},
      {stage1_21[19],stage1_20[75],stage1_19[99],stage1_18[125],stage1_17[180]}
   );
   gpc606_5 gpc746 (
      {stage0_17[264], stage0_17[265], stage0_17[266], stage0_17[267], stage0_17[268], stage0_17[269]},
      {stage0_19[120], stage0_19[121], stage0_19[122], stage0_19[123], stage0_19[124], stage0_19[125]},
      {stage1_21[20],stage1_20[76],stage1_19[100],stage1_18[126],stage1_17[181]}
   );
   gpc606_5 gpc747 (
      {stage0_17[270], stage0_17[271], stage0_17[272], stage0_17[273], stage0_17[274], stage0_17[275]},
      {stage0_19[126], stage0_19[127], stage0_19[128], stage0_19[129], stage0_19[130], stage0_19[131]},
      {stage1_21[21],stage1_20[77],stage1_19[101],stage1_18[127],stage1_17[182]}
   );
   gpc606_5 gpc748 (
      {stage0_17[276], stage0_17[277], stage0_17[278], stage0_17[279], stage0_17[280], stage0_17[281]},
      {stage0_19[132], stage0_19[133], stage0_19[134], stage0_19[135], stage0_19[136], stage0_19[137]},
      {stage1_21[22],stage1_20[78],stage1_19[102],stage1_18[128],stage1_17[183]}
   );
   gpc606_5 gpc749 (
      {stage0_17[282], stage0_17[283], stage0_17[284], stage0_17[285], stage0_17[286], stage0_17[287]},
      {stage0_19[138], stage0_19[139], stage0_19[140], stage0_19[141], stage0_19[142], stage0_19[143]},
      {stage1_21[23],stage1_20[79],stage1_19[103],stage1_18[129],stage1_17[184]}
   );
   gpc606_5 gpc750 (
      {stage0_17[288], stage0_17[289], stage0_17[290], stage0_17[291], stage0_17[292], stage0_17[293]},
      {stage0_19[144], stage0_19[145], stage0_19[146], stage0_19[147], stage0_19[148], stage0_19[149]},
      {stage1_21[24],stage1_20[80],stage1_19[104],stage1_18[130],stage1_17[185]}
   );
   gpc606_5 gpc751 (
      {stage0_17[294], stage0_17[295], stage0_17[296], stage0_17[297], stage0_17[298], stage0_17[299]},
      {stage0_19[150], stage0_19[151], stage0_19[152], stage0_19[153], stage0_19[154], stage0_19[155]},
      {stage1_21[25],stage1_20[81],stage1_19[105],stage1_18[131],stage1_17[186]}
   );
   gpc606_5 gpc752 (
      {stage0_17[300], stage0_17[301], stage0_17[302], stage0_17[303], stage0_17[304], stage0_17[305]},
      {stage0_19[156], stage0_19[157], stage0_19[158], stage0_19[159], stage0_19[160], stage0_19[161]},
      {stage1_21[26],stage1_20[82],stage1_19[106],stage1_18[132],stage1_17[187]}
   );
   gpc606_5 gpc753 (
      {stage0_17[306], stage0_17[307], stage0_17[308], stage0_17[309], stage0_17[310], stage0_17[311]},
      {stage0_19[162], stage0_19[163], stage0_19[164], stage0_19[165], stage0_19[166], stage0_19[167]},
      {stage1_21[27],stage1_20[83],stage1_19[107],stage1_18[133],stage1_17[188]}
   );
   gpc606_5 gpc754 (
      {stage0_17[312], stage0_17[313], stage0_17[314], stage0_17[315], stage0_17[316], stage0_17[317]},
      {stage0_19[168], stage0_19[169], stage0_19[170], stage0_19[171], stage0_19[172], stage0_19[173]},
      {stage1_21[28],stage1_20[84],stage1_19[108],stage1_18[134],stage1_17[189]}
   );
   gpc606_5 gpc755 (
      {stage0_17[318], stage0_17[319], stage0_17[320], stage0_17[321], stage0_17[322], stage0_17[323]},
      {stage0_19[174], stage0_19[175], stage0_19[176], stage0_19[177], stage0_19[178], stage0_19[179]},
      {stage1_21[29],stage1_20[85],stage1_19[109],stage1_18[135],stage1_17[190]}
   );
   gpc606_5 gpc756 (
      {stage0_17[324], stage0_17[325], stage0_17[326], stage0_17[327], stage0_17[328], stage0_17[329]},
      {stage0_19[180], stage0_19[181], stage0_19[182], stage0_19[183], stage0_19[184], stage0_19[185]},
      {stage1_21[30],stage1_20[86],stage1_19[110],stage1_18[136],stage1_17[191]}
   );
   gpc606_5 gpc757 (
      {stage0_17[330], stage0_17[331], stage0_17[332], stage0_17[333], stage0_17[334], stage0_17[335]},
      {stage0_19[186], stage0_19[187], stage0_19[188], stage0_19[189], stage0_19[190], stage0_19[191]},
      {stage1_21[31],stage1_20[87],stage1_19[111],stage1_18[137],stage1_17[192]}
   );
   gpc606_5 gpc758 (
      {stage0_17[336], stage0_17[337], stage0_17[338], stage0_17[339], stage0_17[340], stage0_17[341]},
      {stage0_19[192], stage0_19[193], stage0_19[194], stage0_19[195], stage0_19[196], stage0_19[197]},
      {stage1_21[32],stage1_20[88],stage1_19[112],stage1_18[138],stage1_17[193]}
   );
   gpc606_5 gpc759 (
      {stage0_17[342], stage0_17[343], stage0_17[344], stage0_17[345], stage0_17[346], stage0_17[347]},
      {stage0_19[198], stage0_19[199], stage0_19[200], stage0_19[201], stage0_19[202], stage0_19[203]},
      {stage1_21[33],stage1_20[89],stage1_19[113],stage1_18[139],stage1_17[194]}
   );
   gpc606_5 gpc760 (
      {stage0_17[348], stage0_17[349], stage0_17[350], stage0_17[351], stage0_17[352], stage0_17[353]},
      {stage0_19[204], stage0_19[205], stage0_19[206], stage0_19[207], stage0_19[208], stage0_19[209]},
      {stage1_21[34],stage1_20[90],stage1_19[114],stage1_18[140],stage1_17[195]}
   );
   gpc606_5 gpc761 (
      {stage0_17[354], stage0_17[355], stage0_17[356], stage0_17[357], stage0_17[358], stage0_17[359]},
      {stage0_19[210], stage0_19[211], stage0_19[212], stage0_19[213], stage0_19[214], stage0_19[215]},
      {stage1_21[35],stage1_20[91],stage1_19[115],stage1_18[141],stage1_17[196]}
   );
   gpc606_5 gpc762 (
      {stage0_17[360], stage0_17[361], stage0_17[362], stage0_17[363], stage0_17[364], stage0_17[365]},
      {stage0_19[216], stage0_19[217], stage0_19[218], stage0_19[219], stage0_19[220], stage0_19[221]},
      {stage1_21[36],stage1_20[92],stage1_19[116],stage1_18[142],stage1_17[197]}
   );
   gpc606_5 gpc763 (
      {stage0_17[366], stage0_17[367], stage0_17[368], stage0_17[369], stage0_17[370], stage0_17[371]},
      {stage0_19[222], stage0_19[223], stage0_19[224], stage0_19[225], stage0_19[226], stage0_19[227]},
      {stage1_21[37],stage1_20[93],stage1_19[117],stage1_18[143],stage1_17[198]}
   );
   gpc606_5 gpc764 (
      {stage0_17[372], stage0_17[373], stage0_17[374], stage0_17[375], stage0_17[376], stage0_17[377]},
      {stage0_19[228], stage0_19[229], stage0_19[230], stage0_19[231], stage0_19[232], stage0_19[233]},
      {stage1_21[38],stage1_20[94],stage1_19[118],stage1_18[144],stage1_17[199]}
   );
   gpc606_5 gpc765 (
      {stage0_17[378], stage0_17[379], stage0_17[380], stage0_17[381], stage0_17[382], stage0_17[383]},
      {stage0_19[234], stage0_19[235], stage0_19[236], stage0_19[237], stage0_19[238], stage0_19[239]},
      {stage1_21[39],stage1_20[95],stage1_19[119],stage1_18[145],stage1_17[200]}
   );
   gpc606_5 gpc766 (
      {stage0_17[384], stage0_17[385], stage0_17[386], stage0_17[387], stage0_17[388], stage0_17[389]},
      {stage0_19[240], stage0_19[241], stage0_19[242], stage0_19[243], stage0_19[244], stage0_19[245]},
      {stage1_21[40],stage1_20[96],stage1_19[120],stage1_18[146],stage1_17[201]}
   );
   gpc606_5 gpc767 (
      {stage0_17[390], stage0_17[391], stage0_17[392], stage0_17[393], stage0_17[394], stage0_17[395]},
      {stage0_19[246], stage0_19[247], stage0_19[248], stage0_19[249], stage0_19[250], stage0_19[251]},
      {stage1_21[41],stage1_20[97],stage1_19[121],stage1_18[147],stage1_17[202]}
   );
   gpc606_5 gpc768 (
      {stage0_17[396], stage0_17[397], stage0_17[398], stage0_17[399], stage0_17[400], stage0_17[401]},
      {stage0_19[252], stage0_19[253], stage0_19[254], stage0_19[255], stage0_19[256], stage0_19[257]},
      {stage1_21[42],stage1_20[98],stage1_19[122],stage1_18[148],stage1_17[203]}
   );
   gpc606_5 gpc769 (
      {stage0_17[402], stage0_17[403], stage0_17[404], stage0_17[405], stage0_17[406], stage0_17[407]},
      {stage0_19[258], stage0_19[259], stage0_19[260], stage0_19[261], stage0_19[262], stage0_19[263]},
      {stage1_21[43],stage1_20[99],stage1_19[123],stage1_18[149],stage1_17[204]}
   );
   gpc606_5 gpc770 (
      {stage0_17[408], stage0_17[409], stage0_17[410], stage0_17[411], stage0_17[412], stage0_17[413]},
      {stage0_19[264], stage0_19[265], stage0_19[266], stage0_19[267], stage0_19[268], stage0_19[269]},
      {stage1_21[44],stage1_20[100],stage1_19[124],stage1_18[150],stage1_17[205]}
   );
   gpc606_5 gpc771 (
      {stage0_17[414], stage0_17[415], stage0_17[416], stage0_17[417], stage0_17[418], stage0_17[419]},
      {stage0_19[270], stage0_19[271], stage0_19[272], stage0_19[273], stage0_19[274], stage0_19[275]},
      {stage1_21[45],stage1_20[101],stage1_19[125],stage1_18[151],stage1_17[206]}
   );
   gpc606_5 gpc772 (
      {stage0_17[420], stage0_17[421], stage0_17[422], stage0_17[423], stage0_17[424], stage0_17[425]},
      {stage0_19[276], stage0_19[277], stage0_19[278], stage0_19[279], stage0_19[280], stage0_19[281]},
      {stage1_21[46],stage1_20[102],stage1_19[126],stage1_18[152],stage1_17[207]}
   );
   gpc606_5 gpc773 (
      {stage0_17[426], stage0_17[427], stage0_17[428], stage0_17[429], stage0_17[430], stage0_17[431]},
      {stage0_19[282], stage0_19[283], stage0_19[284], stage0_19[285], stage0_19[286], stage0_19[287]},
      {stage1_21[47],stage1_20[103],stage1_19[127],stage1_18[153],stage1_17[208]}
   );
   gpc606_5 gpc774 (
      {stage0_17[432], stage0_17[433], stage0_17[434], stage0_17[435], stage0_17[436], stage0_17[437]},
      {stage0_19[288], stage0_19[289], stage0_19[290], stage0_19[291], stage0_19[292], stage0_19[293]},
      {stage1_21[48],stage1_20[104],stage1_19[128],stage1_18[154],stage1_17[209]}
   );
   gpc606_5 gpc775 (
      {stage0_17[438], stage0_17[439], stage0_17[440], stage0_17[441], stage0_17[442], stage0_17[443]},
      {stage0_19[294], stage0_19[295], stage0_19[296], stage0_19[297], stage0_19[298], stage0_19[299]},
      {stage1_21[49],stage1_20[105],stage1_19[129],stage1_18[155],stage1_17[210]}
   );
   gpc606_5 gpc776 (
      {stage0_17[444], stage0_17[445], stage0_17[446], stage0_17[447], stage0_17[448], stage0_17[449]},
      {stage0_19[300], stage0_19[301], stage0_19[302], stage0_19[303], stage0_19[304], stage0_19[305]},
      {stage1_21[50],stage1_20[106],stage1_19[130],stage1_18[156],stage1_17[211]}
   );
   gpc606_5 gpc777 (
      {stage0_17[450], stage0_17[451], stage0_17[452], stage0_17[453], stage0_17[454], stage0_17[455]},
      {stage0_19[306], stage0_19[307], stage0_19[308], stage0_19[309], stage0_19[310], stage0_19[311]},
      {stage1_21[51],stage1_20[107],stage1_19[131],stage1_18[157],stage1_17[212]}
   );
   gpc606_5 gpc778 (
      {stage0_17[456], stage0_17[457], stage0_17[458], stage0_17[459], stage0_17[460], stage0_17[461]},
      {stage0_19[312], stage0_19[313], stage0_19[314], stage0_19[315], stage0_19[316], stage0_19[317]},
      {stage1_21[52],stage1_20[108],stage1_19[132],stage1_18[158],stage1_17[213]}
   );
   gpc606_5 gpc779 (
      {stage0_17[462], stage0_17[463], stage0_17[464], stage0_17[465], stage0_17[466], stage0_17[467]},
      {stage0_19[318], stage0_19[319], stage0_19[320], stage0_19[321], stage0_19[322], stage0_19[323]},
      {stage1_21[53],stage1_20[109],stage1_19[133],stage1_18[159],stage1_17[214]}
   );
   gpc606_5 gpc780 (
      {stage0_17[468], stage0_17[469], stage0_17[470], stage0_17[471], stage0_17[472], stage0_17[473]},
      {stage0_19[324], stage0_19[325], stage0_19[326], stage0_19[327], stage0_19[328], stage0_19[329]},
      {stage1_21[54],stage1_20[110],stage1_19[134],stage1_18[160],stage1_17[215]}
   );
   gpc606_5 gpc781 (
      {stage0_17[474], stage0_17[475], stage0_17[476], stage0_17[477], stage0_17[478], stage0_17[479]},
      {stage0_19[330], stage0_19[331], stage0_19[332], stage0_19[333], stage0_19[334], stage0_19[335]},
      {stage1_21[55],stage1_20[111],stage1_19[135],stage1_18[161],stage1_17[216]}
   );
   gpc606_5 gpc782 (
      {stage0_17[480], stage0_17[481], stage0_17[482], stage0_17[483], stage0_17[484], stage0_17[485]},
      {stage0_19[336], stage0_19[337], stage0_19[338], stage0_19[339], stage0_19[340], stage0_19[341]},
      {stage1_21[56],stage1_20[112],stage1_19[136],stage1_18[162],stage1_17[217]}
   );
   gpc606_5 gpc783 (
      {stage0_17[486], stage0_17[487], stage0_17[488], stage0_17[489], stage0_17[490], stage0_17[491]},
      {stage0_19[342], stage0_19[343], stage0_19[344], stage0_19[345], stage0_19[346], stage0_19[347]},
      {stage1_21[57],stage1_20[113],stage1_19[137],stage1_18[163],stage1_17[218]}
   );
   gpc606_5 gpc784 (
      {stage0_17[492], stage0_17[493], stage0_17[494], stage0_17[495], stage0_17[496], stage0_17[497]},
      {stage0_19[348], stage0_19[349], stage0_19[350], stage0_19[351], stage0_19[352], stage0_19[353]},
      {stage1_21[58],stage1_20[114],stage1_19[138],stage1_18[164],stage1_17[219]}
   );
   gpc606_5 gpc785 (
      {stage0_17[498], stage0_17[499], stage0_17[500], stage0_17[501], stage0_17[502], stage0_17[503]},
      {stage0_19[354], stage0_19[355], stage0_19[356], stage0_19[357], stage0_19[358], stage0_19[359]},
      {stage1_21[59],stage1_20[115],stage1_19[139],stage1_18[165],stage1_17[220]}
   );
   gpc606_5 gpc786 (
      {stage0_17[504], stage0_17[505], stage0_17[506], stage0_17[507], stage0_17[508], stage0_17[509]},
      {stage0_19[360], stage0_19[361], stage0_19[362], stage0_19[363], stage0_19[364], stage0_19[365]},
      {stage1_21[60],stage1_20[116],stage1_19[140],stage1_18[166],stage1_17[221]}
   );
   gpc615_5 gpc787 (
      {stage0_18[336], stage0_18[337], stage0_18[338], stage0_18[339], stage0_18[340]},
      {stage0_19[366]},
      {stage0_20[0], stage0_20[1], stage0_20[2], stage0_20[3], stage0_20[4], stage0_20[5]},
      {stage1_22[0],stage1_21[61],stage1_20[117],stage1_19[141],stage1_18[167]}
   );
   gpc615_5 gpc788 (
      {stage0_18[341], stage0_18[342], stage0_18[343], stage0_18[344], stage0_18[345]},
      {stage0_19[367]},
      {stage0_20[6], stage0_20[7], stage0_20[8], stage0_20[9], stage0_20[10], stage0_20[11]},
      {stage1_22[1],stage1_21[62],stage1_20[118],stage1_19[142],stage1_18[168]}
   );
   gpc615_5 gpc789 (
      {stage0_18[346], stage0_18[347], stage0_18[348], stage0_18[349], stage0_18[350]},
      {stage0_19[368]},
      {stage0_20[12], stage0_20[13], stage0_20[14], stage0_20[15], stage0_20[16], stage0_20[17]},
      {stage1_22[2],stage1_21[63],stage1_20[119],stage1_19[143],stage1_18[169]}
   );
   gpc615_5 gpc790 (
      {stage0_18[351], stage0_18[352], stage0_18[353], stage0_18[354], stage0_18[355]},
      {stage0_19[369]},
      {stage0_20[18], stage0_20[19], stage0_20[20], stage0_20[21], stage0_20[22], stage0_20[23]},
      {stage1_22[3],stage1_21[64],stage1_20[120],stage1_19[144],stage1_18[170]}
   );
   gpc615_5 gpc791 (
      {stage0_18[356], stage0_18[357], stage0_18[358], stage0_18[359], stage0_18[360]},
      {stage0_19[370]},
      {stage0_20[24], stage0_20[25], stage0_20[26], stage0_20[27], stage0_20[28], stage0_20[29]},
      {stage1_22[4],stage1_21[65],stage1_20[121],stage1_19[145],stage1_18[171]}
   );
   gpc615_5 gpc792 (
      {stage0_18[361], stage0_18[362], stage0_18[363], stage0_18[364], stage0_18[365]},
      {stage0_19[371]},
      {stage0_20[30], stage0_20[31], stage0_20[32], stage0_20[33], stage0_20[34], stage0_20[35]},
      {stage1_22[5],stage1_21[66],stage1_20[122],stage1_19[146],stage1_18[172]}
   );
   gpc615_5 gpc793 (
      {stage0_18[366], stage0_18[367], stage0_18[368], stage0_18[369], stage0_18[370]},
      {stage0_19[372]},
      {stage0_20[36], stage0_20[37], stage0_20[38], stage0_20[39], stage0_20[40], stage0_20[41]},
      {stage1_22[6],stage1_21[67],stage1_20[123],stage1_19[147],stage1_18[173]}
   );
   gpc615_5 gpc794 (
      {stage0_18[371], stage0_18[372], stage0_18[373], stage0_18[374], stage0_18[375]},
      {stage0_19[373]},
      {stage0_20[42], stage0_20[43], stage0_20[44], stage0_20[45], stage0_20[46], stage0_20[47]},
      {stage1_22[7],stage1_21[68],stage1_20[124],stage1_19[148],stage1_18[174]}
   );
   gpc615_5 gpc795 (
      {stage0_18[376], stage0_18[377], stage0_18[378], stage0_18[379], stage0_18[380]},
      {stage0_19[374]},
      {stage0_20[48], stage0_20[49], stage0_20[50], stage0_20[51], stage0_20[52], stage0_20[53]},
      {stage1_22[8],stage1_21[69],stage1_20[125],stage1_19[149],stage1_18[175]}
   );
   gpc615_5 gpc796 (
      {stage0_18[381], stage0_18[382], stage0_18[383], stage0_18[384], stage0_18[385]},
      {stage0_19[375]},
      {stage0_20[54], stage0_20[55], stage0_20[56], stage0_20[57], stage0_20[58], stage0_20[59]},
      {stage1_22[9],stage1_21[70],stage1_20[126],stage1_19[150],stage1_18[176]}
   );
   gpc615_5 gpc797 (
      {stage0_18[386], stage0_18[387], stage0_18[388], stage0_18[389], stage0_18[390]},
      {stage0_19[376]},
      {stage0_20[60], stage0_20[61], stage0_20[62], stage0_20[63], stage0_20[64], stage0_20[65]},
      {stage1_22[10],stage1_21[71],stage1_20[127],stage1_19[151],stage1_18[177]}
   );
   gpc615_5 gpc798 (
      {stage0_18[391], stage0_18[392], stage0_18[393], stage0_18[394], stage0_18[395]},
      {stage0_19[377]},
      {stage0_20[66], stage0_20[67], stage0_20[68], stage0_20[69], stage0_20[70], stage0_20[71]},
      {stage1_22[11],stage1_21[72],stage1_20[128],stage1_19[152],stage1_18[178]}
   );
   gpc615_5 gpc799 (
      {stage0_18[396], stage0_18[397], stage0_18[398], stage0_18[399], stage0_18[400]},
      {stage0_19[378]},
      {stage0_20[72], stage0_20[73], stage0_20[74], stage0_20[75], stage0_20[76], stage0_20[77]},
      {stage1_22[12],stage1_21[73],stage1_20[129],stage1_19[153],stage1_18[179]}
   );
   gpc615_5 gpc800 (
      {stage0_18[401], stage0_18[402], stage0_18[403], stage0_18[404], stage0_18[405]},
      {stage0_19[379]},
      {stage0_20[78], stage0_20[79], stage0_20[80], stage0_20[81], stage0_20[82], stage0_20[83]},
      {stage1_22[13],stage1_21[74],stage1_20[130],stage1_19[154],stage1_18[180]}
   );
   gpc615_5 gpc801 (
      {stage0_18[406], stage0_18[407], stage0_18[408], stage0_18[409], stage0_18[410]},
      {stage0_19[380]},
      {stage0_20[84], stage0_20[85], stage0_20[86], stage0_20[87], stage0_20[88], stage0_20[89]},
      {stage1_22[14],stage1_21[75],stage1_20[131],stage1_19[155],stage1_18[181]}
   );
   gpc615_5 gpc802 (
      {stage0_18[411], stage0_18[412], stage0_18[413], stage0_18[414], stage0_18[415]},
      {stage0_19[381]},
      {stage0_20[90], stage0_20[91], stage0_20[92], stage0_20[93], stage0_20[94], stage0_20[95]},
      {stage1_22[15],stage1_21[76],stage1_20[132],stage1_19[156],stage1_18[182]}
   );
   gpc615_5 gpc803 (
      {stage0_18[416], stage0_18[417], stage0_18[418], stage0_18[419], stage0_18[420]},
      {stage0_19[382]},
      {stage0_20[96], stage0_20[97], stage0_20[98], stage0_20[99], stage0_20[100], stage0_20[101]},
      {stage1_22[16],stage1_21[77],stage1_20[133],stage1_19[157],stage1_18[183]}
   );
   gpc615_5 gpc804 (
      {stage0_18[421], stage0_18[422], stage0_18[423], stage0_18[424], stage0_18[425]},
      {stage0_19[383]},
      {stage0_20[102], stage0_20[103], stage0_20[104], stage0_20[105], stage0_20[106], stage0_20[107]},
      {stage1_22[17],stage1_21[78],stage1_20[134],stage1_19[158],stage1_18[184]}
   );
   gpc615_5 gpc805 (
      {stage0_18[426], stage0_18[427], stage0_18[428], stage0_18[429], stage0_18[430]},
      {stage0_19[384]},
      {stage0_20[108], stage0_20[109], stage0_20[110], stage0_20[111], stage0_20[112], stage0_20[113]},
      {stage1_22[18],stage1_21[79],stage1_20[135],stage1_19[159],stage1_18[185]}
   );
   gpc615_5 gpc806 (
      {stage0_18[431], stage0_18[432], stage0_18[433], stage0_18[434], stage0_18[435]},
      {stage0_19[385]},
      {stage0_20[114], stage0_20[115], stage0_20[116], stage0_20[117], stage0_20[118], stage0_20[119]},
      {stage1_22[19],stage1_21[80],stage1_20[136],stage1_19[160],stage1_18[186]}
   );
   gpc615_5 gpc807 (
      {stage0_18[436], stage0_18[437], stage0_18[438], stage0_18[439], stage0_18[440]},
      {stage0_19[386]},
      {stage0_20[120], stage0_20[121], stage0_20[122], stage0_20[123], stage0_20[124], stage0_20[125]},
      {stage1_22[20],stage1_21[81],stage1_20[137],stage1_19[161],stage1_18[187]}
   );
   gpc615_5 gpc808 (
      {stage0_18[441], stage0_18[442], stage0_18[443], stage0_18[444], stage0_18[445]},
      {stage0_19[387]},
      {stage0_20[126], stage0_20[127], stage0_20[128], stage0_20[129], stage0_20[130], stage0_20[131]},
      {stage1_22[21],stage1_21[82],stage1_20[138],stage1_19[162],stage1_18[188]}
   );
   gpc615_5 gpc809 (
      {stage0_18[446], stage0_18[447], stage0_18[448], stage0_18[449], stage0_18[450]},
      {stage0_19[388]},
      {stage0_20[132], stage0_20[133], stage0_20[134], stage0_20[135], stage0_20[136], stage0_20[137]},
      {stage1_22[22],stage1_21[83],stage1_20[139],stage1_19[163],stage1_18[189]}
   );
   gpc615_5 gpc810 (
      {stage0_18[451], stage0_18[452], stage0_18[453], stage0_18[454], stage0_18[455]},
      {stage0_19[389]},
      {stage0_20[138], stage0_20[139], stage0_20[140], stage0_20[141], stage0_20[142], stage0_20[143]},
      {stage1_22[23],stage1_21[84],stage1_20[140],stage1_19[164],stage1_18[190]}
   );
   gpc615_5 gpc811 (
      {stage0_18[456], stage0_18[457], stage0_18[458], stage0_18[459], stage0_18[460]},
      {stage0_19[390]},
      {stage0_20[144], stage0_20[145], stage0_20[146], stage0_20[147], stage0_20[148], stage0_20[149]},
      {stage1_22[24],stage1_21[85],stage1_20[141],stage1_19[165],stage1_18[191]}
   );
   gpc615_5 gpc812 (
      {stage0_18[461], stage0_18[462], stage0_18[463], stage0_18[464], stage0_18[465]},
      {stage0_19[391]},
      {stage0_20[150], stage0_20[151], stage0_20[152], stage0_20[153], stage0_20[154], stage0_20[155]},
      {stage1_22[25],stage1_21[86],stage1_20[142],stage1_19[166],stage1_18[192]}
   );
   gpc615_5 gpc813 (
      {stage0_18[466], stage0_18[467], stage0_18[468], stage0_18[469], stage0_18[470]},
      {stage0_19[392]},
      {stage0_20[156], stage0_20[157], stage0_20[158], stage0_20[159], stage0_20[160], stage0_20[161]},
      {stage1_22[26],stage1_21[87],stage1_20[143],stage1_19[167],stage1_18[193]}
   );
   gpc615_5 gpc814 (
      {stage0_18[471], stage0_18[472], stage0_18[473], stage0_18[474], stage0_18[475]},
      {stage0_19[393]},
      {stage0_20[162], stage0_20[163], stage0_20[164], stage0_20[165], stage0_20[166], stage0_20[167]},
      {stage1_22[27],stage1_21[88],stage1_20[144],stage1_19[168],stage1_18[194]}
   );
   gpc615_5 gpc815 (
      {stage0_18[476], stage0_18[477], stage0_18[478], stage0_18[479], stage0_18[480]},
      {stage0_19[394]},
      {stage0_20[168], stage0_20[169], stage0_20[170], stage0_20[171], stage0_20[172], stage0_20[173]},
      {stage1_22[28],stage1_21[89],stage1_20[145],stage1_19[169],stage1_18[195]}
   );
   gpc615_5 gpc816 (
      {stage0_18[481], stage0_18[482], stage0_18[483], stage0_18[484], stage0_18[485]},
      {stage0_19[395]},
      {stage0_20[174], stage0_20[175], stage0_20[176], stage0_20[177], stage0_20[178], stage0_20[179]},
      {stage1_22[29],stage1_21[90],stage1_20[146],stage1_19[170],stage1_18[196]}
   );
   gpc615_5 gpc817 (
      {stage0_18[486], stage0_18[487], stage0_18[488], stage0_18[489], stage0_18[490]},
      {stage0_19[396]},
      {stage0_20[180], stage0_20[181], stage0_20[182], stage0_20[183], stage0_20[184], stage0_20[185]},
      {stage1_22[30],stage1_21[91],stage1_20[147],stage1_19[171],stage1_18[197]}
   );
   gpc615_5 gpc818 (
      {stage0_18[491], stage0_18[492], stage0_18[493], stage0_18[494], stage0_18[495]},
      {stage0_19[397]},
      {stage0_20[186], stage0_20[187], stage0_20[188], stage0_20[189], stage0_20[190], stage0_20[191]},
      {stage1_22[31],stage1_21[92],stage1_20[148],stage1_19[172],stage1_18[198]}
   );
   gpc615_5 gpc819 (
      {stage0_18[496], stage0_18[497], stage0_18[498], stage0_18[499], stage0_18[500]},
      {stage0_19[398]},
      {stage0_20[192], stage0_20[193], stage0_20[194], stage0_20[195], stage0_20[196], stage0_20[197]},
      {stage1_22[32],stage1_21[93],stage1_20[149],stage1_19[173],stage1_18[199]}
   );
   gpc615_5 gpc820 (
      {stage0_18[501], stage0_18[502], stage0_18[503], stage0_18[504], stage0_18[505]},
      {stage0_19[399]},
      {stage0_20[198], stage0_20[199], stage0_20[200], stage0_20[201], stage0_20[202], stage0_20[203]},
      {stage1_22[33],stage1_21[94],stage1_20[150],stage1_19[174],stage1_18[200]}
   );
   gpc615_5 gpc821 (
      {stage0_18[506], stage0_18[507], stage0_18[508], stage0_18[509], stage0_18[510]},
      {stage0_19[400]},
      {stage0_20[204], stage0_20[205], stage0_20[206], stage0_20[207], stage0_20[208], stage0_20[209]},
      {stage1_22[34],stage1_21[95],stage1_20[151],stage1_19[175],stage1_18[201]}
   );
   gpc615_5 gpc822 (
      {stage0_19[401], stage0_19[402], stage0_19[403], stage0_19[404], stage0_19[405]},
      {stage0_20[210]},
      {stage0_21[0], stage0_21[1], stage0_21[2], stage0_21[3], stage0_21[4], stage0_21[5]},
      {stage1_23[0],stage1_22[35],stage1_21[96],stage1_20[152],stage1_19[176]}
   );
   gpc615_5 gpc823 (
      {stage0_19[406], stage0_19[407], stage0_19[408], stage0_19[409], stage0_19[410]},
      {stage0_20[211]},
      {stage0_21[6], stage0_21[7], stage0_21[8], stage0_21[9], stage0_21[10], stage0_21[11]},
      {stage1_23[1],stage1_22[36],stage1_21[97],stage1_20[153],stage1_19[177]}
   );
   gpc615_5 gpc824 (
      {stage0_19[411], stage0_19[412], stage0_19[413], stage0_19[414], stage0_19[415]},
      {stage0_20[212]},
      {stage0_21[12], stage0_21[13], stage0_21[14], stage0_21[15], stage0_21[16], stage0_21[17]},
      {stage1_23[2],stage1_22[37],stage1_21[98],stage1_20[154],stage1_19[178]}
   );
   gpc615_5 gpc825 (
      {stage0_19[416], stage0_19[417], stage0_19[418], stage0_19[419], stage0_19[420]},
      {stage0_20[213]},
      {stage0_21[18], stage0_21[19], stage0_21[20], stage0_21[21], stage0_21[22], stage0_21[23]},
      {stage1_23[3],stage1_22[38],stage1_21[99],stage1_20[155],stage1_19[179]}
   );
   gpc615_5 gpc826 (
      {stage0_19[421], stage0_19[422], stage0_19[423], stage0_19[424], stage0_19[425]},
      {stage0_20[214]},
      {stage0_21[24], stage0_21[25], stage0_21[26], stage0_21[27], stage0_21[28], stage0_21[29]},
      {stage1_23[4],stage1_22[39],stage1_21[100],stage1_20[156],stage1_19[180]}
   );
   gpc615_5 gpc827 (
      {stage0_19[426], stage0_19[427], stage0_19[428], stage0_19[429], stage0_19[430]},
      {stage0_20[215]},
      {stage0_21[30], stage0_21[31], stage0_21[32], stage0_21[33], stage0_21[34], stage0_21[35]},
      {stage1_23[5],stage1_22[40],stage1_21[101],stage1_20[157],stage1_19[181]}
   );
   gpc606_5 gpc828 (
      {stage0_20[216], stage0_20[217], stage0_20[218], stage0_20[219], stage0_20[220], stage0_20[221]},
      {stage0_22[0], stage0_22[1], stage0_22[2], stage0_22[3], stage0_22[4], stage0_22[5]},
      {stage1_24[0],stage1_23[6],stage1_22[41],stage1_21[102],stage1_20[158]}
   );
   gpc606_5 gpc829 (
      {stage0_20[222], stage0_20[223], stage0_20[224], stage0_20[225], stage0_20[226], stage0_20[227]},
      {stage0_22[6], stage0_22[7], stage0_22[8], stage0_22[9], stage0_22[10], stage0_22[11]},
      {stage1_24[1],stage1_23[7],stage1_22[42],stage1_21[103],stage1_20[159]}
   );
   gpc606_5 gpc830 (
      {stage0_20[228], stage0_20[229], stage0_20[230], stage0_20[231], stage0_20[232], stage0_20[233]},
      {stage0_22[12], stage0_22[13], stage0_22[14], stage0_22[15], stage0_22[16], stage0_22[17]},
      {stage1_24[2],stage1_23[8],stage1_22[43],stage1_21[104],stage1_20[160]}
   );
   gpc606_5 gpc831 (
      {stage0_20[234], stage0_20[235], stage0_20[236], stage0_20[237], stage0_20[238], stage0_20[239]},
      {stage0_22[18], stage0_22[19], stage0_22[20], stage0_22[21], stage0_22[22], stage0_22[23]},
      {stage1_24[3],stage1_23[9],stage1_22[44],stage1_21[105],stage1_20[161]}
   );
   gpc606_5 gpc832 (
      {stage0_20[240], stage0_20[241], stage0_20[242], stage0_20[243], stage0_20[244], stage0_20[245]},
      {stage0_22[24], stage0_22[25], stage0_22[26], stage0_22[27], stage0_22[28], stage0_22[29]},
      {stage1_24[4],stage1_23[10],stage1_22[45],stage1_21[106],stage1_20[162]}
   );
   gpc606_5 gpc833 (
      {stage0_20[246], stage0_20[247], stage0_20[248], stage0_20[249], stage0_20[250], stage0_20[251]},
      {stage0_22[30], stage0_22[31], stage0_22[32], stage0_22[33], stage0_22[34], stage0_22[35]},
      {stage1_24[5],stage1_23[11],stage1_22[46],stage1_21[107],stage1_20[163]}
   );
   gpc606_5 gpc834 (
      {stage0_20[252], stage0_20[253], stage0_20[254], stage0_20[255], stage0_20[256], stage0_20[257]},
      {stage0_22[36], stage0_22[37], stage0_22[38], stage0_22[39], stage0_22[40], stage0_22[41]},
      {stage1_24[6],stage1_23[12],stage1_22[47],stage1_21[108],stage1_20[164]}
   );
   gpc606_5 gpc835 (
      {stage0_20[258], stage0_20[259], stage0_20[260], stage0_20[261], stage0_20[262], stage0_20[263]},
      {stage0_22[42], stage0_22[43], stage0_22[44], stage0_22[45], stage0_22[46], stage0_22[47]},
      {stage1_24[7],stage1_23[13],stage1_22[48],stage1_21[109],stage1_20[165]}
   );
   gpc606_5 gpc836 (
      {stage0_20[264], stage0_20[265], stage0_20[266], stage0_20[267], stage0_20[268], stage0_20[269]},
      {stage0_22[48], stage0_22[49], stage0_22[50], stage0_22[51], stage0_22[52], stage0_22[53]},
      {stage1_24[8],stage1_23[14],stage1_22[49],stage1_21[110],stage1_20[166]}
   );
   gpc606_5 gpc837 (
      {stage0_20[270], stage0_20[271], stage0_20[272], stage0_20[273], stage0_20[274], stage0_20[275]},
      {stage0_22[54], stage0_22[55], stage0_22[56], stage0_22[57], stage0_22[58], stage0_22[59]},
      {stage1_24[9],stage1_23[15],stage1_22[50],stage1_21[111],stage1_20[167]}
   );
   gpc606_5 gpc838 (
      {stage0_20[276], stage0_20[277], stage0_20[278], stage0_20[279], stage0_20[280], stage0_20[281]},
      {stage0_22[60], stage0_22[61], stage0_22[62], stage0_22[63], stage0_22[64], stage0_22[65]},
      {stage1_24[10],stage1_23[16],stage1_22[51],stage1_21[112],stage1_20[168]}
   );
   gpc606_5 gpc839 (
      {stage0_20[282], stage0_20[283], stage0_20[284], stage0_20[285], stage0_20[286], stage0_20[287]},
      {stage0_22[66], stage0_22[67], stage0_22[68], stage0_22[69], stage0_22[70], stage0_22[71]},
      {stage1_24[11],stage1_23[17],stage1_22[52],stage1_21[113],stage1_20[169]}
   );
   gpc606_5 gpc840 (
      {stage0_20[288], stage0_20[289], stage0_20[290], stage0_20[291], stage0_20[292], stage0_20[293]},
      {stage0_22[72], stage0_22[73], stage0_22[74], stage0_22[75], stage0_22[76], stage0_22[77]},
      {stage1_24[12],stage1_23[18],stage1_22[53],stage1_21[114],stage1_20[170]}
   );
   gpc606_5 gpc841 (
      {stage0_20[294], stage0_20[295], stage0_20[296], stage0_20[297], stage0_20[298], stage0_20[299]},
      {stage0_22[78], stage0_22[79], stage0_22[80], stage0_22[81], stage0_22[82], stage0_22[83]},
      {stage1_24[13],stage1_23[19],stage1_22[54],stage1_21[115],stage1_20[171]}
   );
   gpc606_5 gpc842 (
      {stage0_20[300], stage0_20[301], stage0_20[302], stage0_20[303], stage0_20[304], stage0_20[305]},
      {stage0_22[84], stage0_22[85], stage0_22[86], stage0_22[87], stage0_22[88], stage0_22[89]},
      {stage1_24[14],stage1_23[20],stage1_22[55],stage1_21[116],stage1_20[172]}
   );
   gpc606_5 gpc843 (
      {stage0_20[306], stage0_20[307], stage0_20[308], stage0_20[309], stage0_20[310], stage0_20[311]},
      {stage0_22[90], stage0_22[91], stage0_22[92], stage0_22[93], stage0_22[94], stage0_22[95]},
      {stage1_24[15],stage1_23[21],stage1_22[56],stage1_21[117],stage1_20[173]}
   );
   gpc606_5 gpc844 (
      {stage0_20[312], stage0_20[313], stage0_20[314], stage0_20[315], stage0_20[316], stage0_20[317]},
      {stage0_22[96], stage0_22[97], stage0_22[98], stage0_22[99], stage0_22[100], stage0_22[101]},
      {stage1_24[16],stage1_23[22],stage1_22[57],stage1_21[118],stage1_20[174]}
   );
   gpc606_5 gpc845 (
      {stage0_20[318], stage0_20[319], stage0_20[320], stage0_20[321], stage0_20[322], stage0_20[323]},
      {stage0_22[102], stage0_22[103], stage0_22[104], stage0_22[105], stage0_22[106], stage0_22[107]},
      {stage1_24[17],stage1_23[23],stage1_22[58],stage1_21[119],stage1_20[175]}
   );
   gpc606_5 gpc846 (
      {stage0_20[324], stage0_20[325], stage0_20[326], stage0_20[327], stage0_20[328], stage0_20[329]},
      {stage0_22[108], stage0_22[109], stage0_22[110], stage0_22[111], stage0_22[112], stage0_22[113]},
      {stage1_24[18],stage1_23[24],stage1_22[59],stage1_21[120],stage1_20[176]}
   );
   gpc606_5 gpc847 (
      {stage0_20[330], stage0_20[331], stage0_20[332], stage0_20[333], stage0_20[334], stage0_20[335]},
      {stage0_22[114], stage0_22[115], stage0_22[116], stage0_22[117], stage0_22[118], stage0_22[119]},
      {stage1_24[19],stage1_23[25],stage1_22[60],stage1_21[121],stage1_20[177]}
   );
   gpc606_5 gpc848 (
      {stage0_20[336], stage0_20[337], stage0_20[338], stage0_20[339], stage0_20[340], stage0_20[341]},
      {stage0_22[120], stage0_22[121], stage0_22[122], stage0_22[123], stage0_22[124], stage0_22[125]},
      {stage1_24[20],stage1_23[26],stage1_22[61],stage1_21[122],stage1_20[178]}
   );
   gpc606_5 gpc849 (
      {stage0_20[342], stage0_20[343], stage0_20[344], stage0_20[345], stage0_20[346], stage0_20[347]},
      {stage0_22[126], stage0_22[127], stage0_22[128], stage0_22[129], stage0_22[130], stage0_22[131]},
      {stage1_24[21],stage1_23[27],stage1_22[62],stage1_21[123],stage1_20[179]}
   );
   gpc606_5 gpc850 (
      {stage0_20[348], stage0_20[349], stage0_20[350], stage0_20[351], stage0_20[352], stage0_20[353]},
      {stage0_22[132], stage0_22[133], stage0_22[134], stage0_22[135], stage0_22[136], stage0_22[137]},
      {stage1_24[22],stage1_23[28],stage1_22[63],stage1_21[124],stage1_20[180]}
   );
   gpc606_5 gpc851 (
      {stage0_20[354], stage0_20[355], stage0_20[356], stage0_20[357], stage0_20[358], stage0_20[359]},
      {stage0_22[138], stage0_22[139], stage0_22[140], stage0_22[141], stage0_22[142], stage0_22[143]},
      {stage1_24[23],stage1_23[29],stage1_22[64],stage1_21[125],stage1_20[181]}
   );
   gpc606_5 gpc852 (
      {stage0_20[360], stage0_20[361], stage0_20[362], stage0_20[363], stage0_20[364], stage0_20[365]},
      {stage0_22[144], stage0_22[145], stage0_22[146], stage0_22[147], stage0_22[148], stage0_22[149]},
      {stage1_24[24],stage1_23[30],stage1_22[65],stage1_21[126],stage1_20[182]}
   );
   gpc606_5 gpc853 (
      {stage0_20[366], stage0_20[367], stage0_20[368], stage0_20[369], stage0_20[370], stage0_20[371]},
      {stage0_22[150], stage0_22[151], stage0_22[152], stage0_22[153], stage0_22[154], stage0_22[155]},
      {stage1_24[25],stage1_23[31],stage1_22[66],stage1_21[127],stage1_20[183]}
   );
   gpc606_5 gpc854 (
      {stage0_20[372], stage0_20[373], stage0_20[374], stage0_20[375], stage0_20[376], stage0_20[377]},
      {stage0_22[156], stage0_22[157], stage0_22[158], stage0_22[159], stage0_22[160], stage0_22[161]},
      {stage1_24[26],stage1_23[32],stage1_22[67],stage1_21[128],stage1_20[184]}
   );
   gpc606_5 gpc855 (
      {stage0_20[378], stage0_20[379], stage0_20[380], stage0_20[381], stage0_20[382], stage0_20[383]},
      {stage0_22[162], stage0_22[163], stage0_22[164], stage0_22[165], stage0_22[166], stage0_22[167]},
      {stage1_24[27],stage1_23[33],stage1_22[68],stage1_21[129],stage1_20[185]}
   );
   gpc606_5 gpc856 (
      {stage0_20[384], stage0_20[385], stage0_20[386], stage0_20[387], stage0_20[388], stage0_20[389]},
      {stage0_22[168], stage0_22[169], stage0_22[170], stage0_22[171], stage0_22[172], stage0_22[173]},
      {stage1_24[28],stage1_23[34],stage1_22[69],stage1_21[130],stage1_20[186]}
   );
   gpc606_5 gpc857 (
      {stage0_20[390], stage0_20[391], stage0_20[392], stage0_20[393], stage0_20[394], stage0_20[395]},
      {stage0_22[174], stage0_22[175], stage0_22[176], stage0_22[177], stage0_22[178], stage0_22[179]},
      {stage1_24[29],stage1_23[35],stage1_22[70],stage1_21[131],stage1_20[187]}
   );
   gpc606_5 gpc858 (
      {stage0_20[396], stage0_20[397], stage0_20[398], stage0_20[399], stage0_20[400], stage0_20[401]},
      {stage0_22[180], stage0_22[181], stage0_22[182], stage0_22[183], stage0_22[184], stage0_22[185]},
      {stage1_24[30],stage1_23[36],stage1_22[71],stage1_21[132],stage1_20[188]}
   );
   gpc606_5 gpc859 (
      {stage0_20[402], stage0_20[403], stage0_20[404], stage0_20[405], stage0_20[406], stage0_20[407]},
      {stage0_22[186], stage0_22[187], stage0_22[188], stage0_22[189], stage0_22[190], stage0_22[191]},
      {stage1_24[31],stage1_23[37],stage1_22[72],stage1_21[133],stage1_20[189]}
   );
   gpc606_5 gpc860 (
      {stage0_20[408], stage0_20[409], stage0_20[410], stage0_20[411], stage0_20[412], stage0_20[413]},
      {stage0_22[192], stage0_22[193], stage0_22[194], stage0_22[195], stage0_22[196], stage0_22[197]},
      {stage1_24[32],stage1_23[38],stage1_22[73],stage1_21[134],stage1_20[190]}
   );
   gpc606_5 gpc861 (
      {stage0_20[414], stage0_20[415], stage0_20[416], stage0_20[417], stage0_20[418], stage0_20[419]},
      {stage0_22[198], stage0_22[199], stage0_22[200], stage0_22[201], stage0_22[202], stage0_22[203]},
      {stage1_24[33],stage1_23[39],stage1_22[74],stage1_21[135],stage1_20[191]}
   );
   gpc606_5 gpc862 (
      {stage0_20[420], stage0_20[421], stage0_20[422], stage0_20[423], stage0_20[424], stage0_20[425]},
      {stage0_22[204], stage0_22[205], stage0_22[206], stage0_22[207], stage0_22[208], stage0_22[209]},
      {stage1_24[34],stage1_23[40],stage1_22[75],stage1_21[136],stage1_20[192]}
   );
   gpc606_5 gpc863 (
      {stage0_20[426], stage0_20[427], stage0_20[428], stage0_20[429], stage0_20[430], stage0_20[431]},
      {stage0_22[210], stage0_22[211], stage0_22[212], stage0_22[213], stage0_22[214], stage0_22[215]},
      {stage1_24[35],stage1_23[41],stage1_22[76],stage1_21[137],stage1_20[193]}
   );
   gpc606_5 gpc864 (
      {stage0_20[432], stage0_20[433], stage0_20[434], stage0_20[435], stage0_20[436], stage0_20[437]},
      {stage0_22[216], stage0_22[217], stage0_22[218], stage0_22[219], stage0_22[220], stage0_22[221]},
      {stage1_24[36],stage1_23[42],stage1_22[77],stage1_21[138],stage1_20[194]}
   );
   gpc606_5 gpc865 (
      {stage0_20[438], stage0_20[439], stage0_20[440], stage0_20[441], stage0_20[442], stage0_20[443]},
      {stage0_22[222], stage0_22[223], stage0_22[224], stage0_22[225], stage0_22[226], stage0_22[227]},
      {stage1_24[37],stage1_23[43],stage1_22[78],stage1_21[139],stage1_20[195]}
   );
   gpc606_5 gpc866 (
      {stage0_20[444], stage0_20[445], stage0_20[446], stage0_20[447], stage0_20[448], stage0_20[449]},
      {stage0_22[228], stage0_22[229], stage0_22[230], stage0_22[231], stage0_22[232], stage0_22[233]},
      {stage1_24[38],stage1_23[44],stage1_22[79],stage1_21[140],stage1_20[196]}
   );
   gpc606_5 gpc867 (
      {stage0_20[450], stage0_20[451], stage0_20[452], stage0_20[453], stage0_20[454], stage0_20[455]},
      {stage0_22[234], stage0_22[235], stage0_22[236], stage0_22[237], stage0_22[238], stage0_22[239]},
      {stage1_24[39],stage1_23[45],stage1_22[80],stage1_21[141],stage1_20[197]}
   );
   gpc606_5 gpc868 (
      {stage0_20[456], stage0_20[457], stage0_20[458], stage0_20[459], stage0_20[460], stage0_20[461]},
      {stage0_22[240], stage0_22[241], stage0_22[242], stage0_22[243], stage0_22[244], stage0_22[245]},
      {stage1_24[40],stage1_23[46],stage1_22[81],stage1_21[142],stage1_20[198]}
   );
   gpc606_5 gpc869 (
      {stage0_20[462], stage0_20[463], stage0_20[464], stage0_20[465], stage0_20[466], stage0_20[467]},
      {stage0_22[246], stage0_22[247], stage0_22[248], stage0_22[249], stage0_22[250], stage0_22[251]},
      {stage1_24[41],stage1_23[47],stage1_22[82],stage1_21[143],stage1_20[199]}
   );
   gpc606_5 gpc870 (
      {stage0_20[468], stage0_20[469], stage0_20[470], stage0_20[471], stage0_20[472], stage0_20[473]},
      {stage0_22[252], stage0_22[253], stage0_22[254], stage0_22[255], stage0_22[256], stage0_22[257]},
      {stage1_24[42],stage1_23[48],stage1_22[83],stage1_21[144],stage1_20[200]}
   );
   gpc606_5 gpc871 (
      {stage0_20[474], stage0_20[475], stage0_20[476], stage0_20[477], stage0_20[478], stage0_20[479]},
      {stage0_22[258], stage0_22[259], stage0_22[260], stage0_22[261], stage0_22[262], stage0_22[263]},
      {stage1_24[43],stage1_23[49],stage1_22[84],stage1_21[145],stage1_20[201]}
   );
   gpc606_5 gpc872 (
      {stage0_20[480], stage0_20[481], stage0_20[482], stage0_20[483], stage0_20[484], stage0_20[485]},
      {stage0_22[264], stage0_22[265], stage0_22[266], stage0_22[267], stage0_22[268], stage0_22[269]},
      {stage1_24[44],stage1_23[50],stage1_22[85],stage1_21[146],stage1_20[202]}
   );
   gpc606_5 gpc873 (
      {stage0_20[486], stage0_20[487], stage0_20[488], stage0_20[489], stage0_20[490], stage0_20[491]},
      {stage0_22[270], stage0_22[271], stage0_22[272], stage0_22[273], stage0_22[274], stage0_22[275]},
      {stage1_24[45],stage1_23[51],stage1_22[86],stage1_21[147],stage1_20[203]}
   );
   gpc606_5 gpc874 (
      {stage0_20[492], stage0_20[493], stage0_20[494], stage0_20[495], stage0_20[496], stage0_20[497]},
      {stage0_22[276], stage0_22[277], stage0_22[278], stage0_22[279], stage0_22[280], stage0_22[281]},
      {stage1_24[46],stage1_23[52],stage1_22[87],stage1_21[148],stage1_20[204]}
   );
   gpc606_5 gpc875 (
      {stage0_20[498], stage0_20[499], stage0_20[500], stage0_20[501], stage0_20[502], stage0_20[503]},
      {stage0_22[282], stage0_22[283], stage0_22[284], stage0_22[285], stage0_22[286], stage0_22[287]},
      {stage1_24[47],stage1_23[53],stage1_22[88],stage1_21[149],stage1_20[205]}
   );
   gpc606_5 gpc876 (
      {stage0_21[36], stage0_21[37], stage0_21[38], stage0_21[39], stage0_21[40], stage0_21[41]},
      {stage0_23[0], stage0_23[1], stage0_23[2], stage0_23[3], stage0_23[4], stage0_23[5]},
      {stage1_25[0],stage1_24[48],stage1_23[54],stage1_22[89],stage1_21[150]}
   );
   gpc606_5 gpc877 (
      {stage0_21[42], stage0_21[43], stage0_21[44], stage0_21[45], stage0_21[46], stage0_21[47]},
      {stage0_23[6], stage0_23[7], stage0_23[8], stage0_23[9], stage0_23[10], stage0_23[11]},
      {stage1_25[1],stage1_24[49],stage1_23[55],stage1_22[90],stage1_21[151]}
   );
   gpc606_5 gpc878 (
      {stage0_21[48], stage0_21[49], stage0_21[50], stage0_21[51], stage0_21[52], stage0_21[53]},
      {stage0_23[12], stage0_23[13], stage0_23[14], stage0_23[15], stage0_23[16], stage0_23[17]},
      {stage1_25[2],stage1_24[50],stage1_23[56],stage1_22[91],stage1_21[152]}
   );
   gpc606_5 gpc879 (
      {stage0_21[54], stage0_21[55], stage0_21[56], stage0_21[57], stage0_21[58], stage0_21[59]},
      {stage0_23[18], stage0_23[19], stage0_23[20], stage0_23[21], stage0_23[22], stage0_23[23]},
      {stage1_25[3],stage1_24[51],stage1_23[57],stage1_22[92],stage1_21[153]}
   );
   gpc606_5 gpc880 (
      {stage0_21[60], stage0_21[61], stage0_21[62], stage0_21[63], stage0_21[64], stage0_21[65]},
      {stage0_23[24], stage0_23[25], stage0_23[26], stage0_23[27], stage0_23[28], stage0_23[29]},
      {stage1_25[4],stage1_24[52],stage1_23[58],stage1_22[93],stage1_21[154]}
   );
   gpc606_5 gpc881 (
      {stage0_21[66], stage0_21[67], stage0_21[68], stage0_21[69], stage0_21[70], stage0_21[71]},
      {stage0_23[30], stage0_23[31], stage0_23[32], stage0_23[33], stage0_23[34], stage0_23[35]},
      {stage1_25[5],stage1_24[53],stage1_23[59],stage1_22[94],stage1_21[155]}
   );
   gpc606_5 gpc882 (
      {stage0_21[72], stage0_21[73], stage0_21[74], stage0_21[75], stage0_21[76], stage0_21[77]},
      {stage0_23[36], stage0_23[37], stage0_23[38], stage0_23[39], stage0_23[40], stage0_23[41]},
      {stage1_25[6],stage1_24[54],stage1_23[60],stage1_22[95],stage1_21[156]}
   );
   gpc606_5 gpc883 (
      {stage0_21[78], stage0_21[79], stage0_21[80], stage0_21[81], stage0_21[82], stage0_21[83]},
      {stage0_23[42], stage0_23[43], stage0_23[44], stage0_23[45], stage0_23[46], stage0_23[47]},
      {stage1_25[7],stage1_24[55],stage1_23[61],stage1_22[96],stage1_21[157]}
   );
   gpc606_5 gpc884 (
      {stage0_21[84], stage0_21[85], stage0_21[86], stage0_21[87], stage0_21[88], stage0_21[89]},
      {stage0_23[48], stage0_23[49], stage0_23[50], stage0_23[51], stage0_23[52], stage0_23[53]},
      {stage1_25[8],stage1_24[56],stage1_23[62],stage1_22[97],stage1_21[158]}
   );
   gpc606_5 gpc885 (
      {stage0_21[90], stage0_21[91], stage0_21[92], stage0_21[93], stage0_21[94], stage0_21[95]},
      {stage0_23[54], stage0_23[55], stage0_23[56], stage0_23[57], stage0_23[58], stage0_23[59]},
      {stage1_25[9],stage1_24[57],stage1_23[63],stage1_22[98],stage1_21[159]}
   );
   gpc606_5 gpc886 (
      {stage0_21[96], stage0_21[97], stage0_21[98], stage0_21[99], stage0_21[100], stage0_21[101]},
      {stage0_23[60], stage0_23[61], stage0_23[62], stage0_23[63], stage0_23[64], stage0_23[65]},
      {stage1_25[10],stage1_24[58],stage1_23[64],stage1_22[99],stage1_21[160]}
   );
   gpc606_5 gpc887 (
      {stage0_21[102], stage0_21[103], stage0_21[104], stage0_21[105], stage0_21[106], stage0_21[107]},
      {stage0_23[66], stage0_23[67], stage0_23[68], stage0_23[69], stage0_23[70], stage0_23[71]},
      {stage1_25[11],stage1_24[59],stage1_23[65],stage1_22[100],stage1_21[161]}
   );
   gpc606_5 gpc888 (
      {stage0_21[108], stage0_21[109], stage0_21[110], stage0_21[111], stage0_21[112], stage0_21[113]},
      {stage0_23[72], stage0_23[73], stage0_23[74], stage0_23[75], stage0_23[76], stage0_23[77]},
      {stage1_25[12],stage1_24[60],stage1_23[66],stage1_22[101],stage1_21[162]}
   );
   gpc606_5 gpc889 (
      {stage0_21[114], stage0_21[115], stage0_21[116], stage0_21[117], stage0_21[118], stage0_21[119]},
      {stage0_23[78], stage0_23[79], stage0_23[80], stage0_23[81], stage0_23[82], stage0_23[83]},
      {stage1_25[13],stage1_24[61],stage1_23[67],stage1_22[102],stage1_21[163]}
   );
   gpc606_5 gpc890 (
      {stage0_21[120], stage0_21[121], stage0_21[122], stage0_21[123], stage0_21[124], stage0_21[125]},
      {stage0_23[84], stage0_23[85], stage0_23[86], stage0_23[87], stage0_23[88], stage0_23[89]},
      {stage1_25[14],stage1_24[62],stage1_23[68],stage1_22[103],stage1_21[164]}
   );
   gpc606_5 gpc891 (
      {stage0_21[126], stage0_21[127], stage0_21[128], stage0_21[129], stage0_21[130], stage0_21[131]},
      {stage0_23[90], stage0_23[91], stage0_23[92], stage0_23[93], stage0_23[94], stage0_23[95]},
      {stage1_25[15],stage1_24[63],stage1_23[69],stage1_22[104],stage1_21[165]}
   );
   gpc606_5 gpc892 (
      {stage0_21[132], stage0_21[133], stage0_21[134], stage0_21[135], stage0_21[136], stage0_21[137]},
      {stage0_23[96], stage0_23[97], stage0_23[98], stage0_23[99], stage0_23[100], stage0_23[101]},
      {stage1_25[16],stage1_24[64],stage1_23[70],stage1_22[105],stage1_21[166]}
   );
   gpc606_5 gpc893 (
      {stage0_21[138], stage0_21[139], stage0_21[140], stage0_21[141], stage0_21[142], stage0_21[143]},
      {stage0_23[102], stage0_23[103], stage0_23[104], stage0_23[105], stage0_23[106], stage0_23[107]},
      {stage1_25[17],stage1_24[65],stage1_23[71],stage1_22[106],stage1_21[167]}
   );
   gpc606_5 gpc894 (
      {stage0_21[144], stage0_21[145], stage0_21[146], stage0_21[147], stage0_21[148], stage0_21[149]},
      {stage0_23[108], stage0_23[109], stage0_23[110], stage0_23[111], stage0_23[112], stage0_23[113]},
      {stage1_25[18],stage1_24[66],stage1_23[72],stage1_22[107],stage1_21[168]}
   );
   gpc606_5 gpc895 (
      {stage0_21[150], stage0_21[151], stage0_21[152], stage0_21[153], stage0_21[154], stage0_21[155]},
      {stage0_23[114], stage0_23[115], stage0_23[116], stage0_23[117], stage0_23[118], stage0_23[119]},
      {stage1_25[19],stage1_24[67],stage1_23[73],stage1_22[108],stage1_21[169]}
   );
   gpc606_5 gpc896 (
      {stage0_21[156], stage0_21[157], stage0_21[158], stage0_21[159], stage0_21[160], stage0_21[161]},
      {stage0_23[120], stage0_23[121], stage0_23[122], stage0_23[123], stage0_23[124], stage0_23[125]},
      {stage1_25[20],stage1_24[68],stage1_23[74],stage1_22[109],stage1_21[170]}
   );
   gpc606_5 gpc897 (
      {stage0_21[162], stage0_21[163], stage0_21[164], stage0_21[165], stage0_21[166], stage0_21[167]},
      {stage0_23[126], stage0_23[127], stage0_23[128], stage0_23[129], stage0_23[130], stage0_23[131]},
      {stage1_25[21],stage1_24[69],stage1_23[75],stage1_22[110],stage1_21[171]}
   );
   gpc606_5 gpc898 (
      {stage0_21[168], stage0_21[169], stage0_21[170], stage0_21[171], stage0_21[172], stage0_21[173]},
      {stage0_23[132], stage0_23[133], stage0_23[134], stage0_23[135], stage0_23[136], stage0_23[137]},
      {stage1_25[22],stage1_24[70],stage1_23[76],stage1_22[111],stage1_21[172]}
   );
   gpc606_5 gpc899 (
      {stage0_21[174], stage0_21[175], stage0_21[176], stage0_21[177], stage0_21[178], stage0_21[179]},
      {stage0_23[138], stage0_23[139], stage0_23[140], stage0_23[141], stage0_23[142], stage0_23[143]},
      {stage1_25[23],stage1_24[71],stage1_23[77],stage1_22[112],stage1_21[173]}
   );
   gpc606_5 gpc900 (
      {stage0_21[180], stage0_21[181], stage0_21[182], stage0_21[183], stage0_21[184], stage0_21[185]},
      {stage0_23[144], stage0_23[145], stage0_23[146], stage0_23[147], stage0_23[148], stage0_23[149]},
      {stage1_25[24],stage1_24[72],stage1_23[78],stage1_22[113],stage1_21[174]}
   );
   gpc606_5 gpc901 (
      {stage0_21[186], stage0_21[187], stage0_21[188], stage0_21[189], stage0_21[190], stage0_21[191]},
      {stage0_23[150], stage0_23[151], stage0_23[152], stage0_23[153], stage0_23[154], stage0_23[155]},
      {stage1_25[25],stage1_24[73],stage1_23[79],stage1_22[114],stage1_21[175]}
   );
   gpc606_5 gpc902 (
      {stage0_21[192], stage0_21[193], stage0_21[194], stage0_21[195], stage0_21[196], stage0_21[197]},
      {stage0_23[156], stage0_23[157], stage0_23[158], stage0_23[159], stage0_23[160], stage0_23[161]},
      {stage1_25[26],stage1_24[74],stage1_23[80],stage1_22[115],stage1_21[176]}
   );
   gpc606_5 gpc903 (
      {stage0_21[198], stage0_21[199], stage0_21[200], stage0_21[201], stage0_21[202], stage0_21[203]},
      {stage0_23[162], stage0_23[163], stage0_23[164], stage0_23[165], stage0_23[166], stage0_23[167]},
      {stage1_25[27],stage1_24[75],stage1_23[81],stage1_22[116],stage1_21[177]}
   );
   gpc606_5 gpc904 (
      {stage0_21[204], stage0_21[205], stage0_21[206], stage0_21[207], stage0_21[208], stage0_21[209]},
      {stage0_23[168], stage0_23[169], stage0_23[170], stage0_23[171], stage0_23[172], stage0_23[173]},
      {stage1_25[28],stage1_24[76],stage1_23[82],stage1_22[117],stage1_21[178]}
   );
   gpc606_5 gpc905 (
      {stage0_21[210], stage0_21[211], stage0_21[212], stage0_21[213], stage0_21[214], stage0_21[215]},
      {stage0_23[174], stage0_23[175], stage0_23[176], stage0_23[177], stage0_23[178], stage0_23[179]},
      {stage1_25[29],stage1_24[77],stage1_23[83],stage1_22[118],stage1_21[179]}
   );
   gpc606_5 gpc906 (
      {stage0_21[216], stage0_21[217], stage0_21[218], stage0_21[219], stage0_21[220], stage0_21[221]},
      {stage0_23[180], stage0_23[181], stage0_23[182], stage0_23[183], stage0_23[184], stage0_23[185]},
      {stage1_25[30],stage1_24[78],stage1_23[84],stage1_22[119],stage1_21[180]}
   );
   gpc606_5 gpc907 (
      {stage0_21[222], stage0_21[223], stage0_21[224], stage0_21[225], stage0_21[226], stage0_21[227]},
      {stage0_23[186], stage0_23[187], stage0_23[188], stage0_23[189], stage0_23[190], stage0_23[191]},
      {stage1_25[31],stage1_24[79],stage1_23[85],stage1_22[120],stage1_21[181]}
   );
   gpc606_5 gpc908 (
      {stage0_21[228], stage0_21[229], stage0_21[230], stage0_21[231], stage0_21[232], stage0_21[233]},
      {stage0_23[192], stage0_23[193], stage0_23[194], stage0_23[195], stage0_23[196], stage0_23[197]},
      {stage1_25[32],stage1_24[80],stage1_23[86],stage1_22[121],stage1_21[182]}
   );
   gpc606_5 gpc909 (
      {stage0_21[234], stage0_21[235], stage0_21[236], stage0_21[237], stage0_21[238], stage0_21[239]},
      {stage0_23[198], stage0_23[199], stage0_23[200], stage0_23[201], stage0_23[202], stage0_23[203]},
      {stage1_25[33],stage1_24[81],stage1_23[87],stage1_22[122],stage1_21[183]}
   );
   gpc606_5 gpc910 (
      {stage0_21[240], stage0_21[241], stage0_21[242], stage0_21[243], stage0_21[244], stage0_21[245]},
      {stage0_23[204], stage0_23[205], stage0_23[206], stage0_23[207], stage0_23[208], stage0_23[209]},
      {stage1_25[34],stage1_24[82],stage1_23[88],stage1_22[123],stage1_21[184]}
   );
   gpc606_5 gpc911 (
      {stage0_21[246], stage0_21[247], stage0_21[248], stage0_21[249], stage0_21[250], stage0_21[251]},
      {stage0_23[210], stage0_23[211], stage0_23[212], stage0_23[213], stage0_23[214], stage0_23[215]},
      {stage1_25[35],stage1_24[83],stage1_23[89],stage1_22[124],stage1_21[185]}
   );
   gpc606_5 gpc912 (
      {stage0_21[252], stage0_21[253], stage0_21[254], stage0_21[255], stage0_21[256], stage0_21[257]},
      {stage0_23[216], stage0_23[217], stage0_23[218], stage0_23[219], stage0_23[220], stage0_23[221]},
      {stage1_25[36],stage1_24[84],stage1_23[90],stage1_22[125],stage1_21[186]}
   );
   gpc606_5 gpc913 (
      {stage0_21[258], stage0_21[259], stage0_21[260], stage0_21[261], stage0_21[262], stage0_21[263]},
      {stage0_23[222], stage0_23[223], stage0_23[224], stage0_23[225], stage0_23[226], stage0_23[227]},
      {stage1_25[37],stage1_24[85],stage1_23[91],stage1_22[126],stage1_21[187]}
   );
   gpc606_5 gpc914 (
      {stage0_21[264], stage0_21[265], stage0_21[266], stage0_21[267], stage0_21[268], stage0_21[269]},
      {stage0_23[228], stage0_23[229], stage0_23[230], stage0_23[231], stage0_23[232], stage0_23[233]},
      {stage1_25[38],stage1_24[86],stage1_23[92],stage1_22[127],stage1_21[188]}
   );
   gpc606_5 gpc915 (
      {stage0_21[270], stage0_21[271], stage0_21[272], stage0_21[273], stage0_21[274], stage0_21[275]},
      {stage0_23[234], stage0_23[235], stage0_23[236], stage0_23[237], stage0_23[238], stage0_23[239]},
      {stage1_25[39],stage1_24[87],stage1_23[93],stage1_22[128],stage1_21[189]}
   );
   gpc615_5 gpc916 (
      {stage0_21[276], stage0_21[277], stage0_21[278], stage0_21[279], stage0_21[280]},
      {stage0_22[288]},
      {stage0_23[240], stage0_23[241], stage0_23[242], stage0_23[243], stage0_23[244], stage0_23[245]},
      {stage1_25[40],stage1_24[88],stage1_23[94],stage1_22[129],stage1_21[190]}
   );
   gpc615_5 gpc917 (
      {stage0_21[281], stage0_21[282], stage0_21[283], stage0_21[284], stage0_21[285]},
      {stage0_22[289]},
      {stage0_23[246], stage0_23[247], stage0_23[248], stage0_23[249], stage0_23[250], stage0_23[251]},
      {stage1_25[41],stage1_24[89],stage1_23[95],stage1_22[130],stage1_21[191]}
   );
   gpc615_5 gpc918 (
      {stage0_21[286], stage0_21[287], stage0_21[288], stage0_21[289], stage0_21[290]},
      {stage0_22[290]},
      {stage0_23[252], stage0_23[253], stage0_23[254], stage0_23[255], stage0_23[256], stage0_23[257]},
      {stage1_25[42],stage1_24[90],stage1_23[96],stage1_22[131],stage1_21[192]}
   );
   gpc615_5 gpc919 (
      {stage0_21[291], stage0_21[292], stage0_21[293], stage0_21[294], stage0_21[295]},
      {stage0_22[291]},
      {stage0_23[258], stage0_23[259], stage0_23[260], stage0_23[261], stage0_23[262], stage0_23[263]},
      {stage1_25[43],stage1_24[91],stage1_23[97],stage1_22[132],stage1_21[193]}
   );
   gpc615_5 gpc920 (
      {stage0_21[296], stage0_21[297], stage0_21[298], stage0_21[299], stage0_21[300]},
      {stage0_22[292]},
      {stage0_23[264], stage0_23[265], stage0_23[266], stage0_23[267], stage0_23[268], stage0_23[269]},
      {stage1_25[44],stage1_24[92],stage1_23[98],stage1_22[133],stage1_21[194]}
   );
   gpc615_5 gpc921 (
      {stage0_21[301], stage0_21[302], stage0_21[303], stage0_21[304], stage0_21[305]},
      {stage0_22[293]},
      {stage0_23[270], stage0_23[271], stage0_23[272], stage0_23[273], stage0_23[274], stage0_23[275]},
      {stage1_25[45],stage1_24[93],stage1_23[99],stage1_22[134],stage1_21[195]}
   );
   gpc615_5 gpc922 (
      {stage0_21[306], stage0_21[307], stage0_21[308], stage0_21[309], stage0_21[310]},
      {stage0_22[294]},
      {stage0_23[276], stage0_23[277], stage0_23[278], stage0_23[279], stage0_23[280], stage0_23[281]},
      {stage1_25[46],stage1_24[94],stage1_23[100],stage1_22[135],stage1_21[196]}
   );
   gpc615_5 gpc923 (
      {stage0_21[311], stage0_21[312], stage0_21[313], stage0_21[314], stage0_21[315]},
      {stage0_22[295]},
      {stage0_23[282], stage0_23[283], stage0_23[284], stage0_23[285], stage0_23[286], stage0_23[287]},
      {stage1_25[47],stage1_24[95],stage1_23[101],stage1_22[136],stage1_21[197]}
   );
   gpc615_5 gpc924 (
      {stage0_21[316], stage0_21[317], stage0_21[318], stage0_21[319], stage0_21[320]},
      {stage0_22[296]},
      {stage0_23[288], stage0_23[289], stage0_23[290], stage0_23[291], stage0_23[292], stage0_23[293]},
      {stage1_25[48],stage1_24[96],stage1_23[102],stage1_22[137],stage1_21[198]}
   );
   gpc615_5 gpc925 (
      {stage0_21[321], stage0_21[322], stage0_21[323], stage0_21[324], stage0_21[325]},
      {stage0_22[297]},
      {stage0_23[294], stage0_23[295], stage0_23[296], stage0_23[297], stage0_23[298], stage0_23[299]},
      {stage1_25[49],stage1_24[97],stage1_23[103],stage1_22[138],stage1_21[199]}
   );
   gpc615_5 gpc926 (
      {stage0_21[326], stage0_21[327], stage0_21[328], stage0_21[329], stage0_21[330]},
      {stage0_22[298]},
      {stage0_23[300], stage0_23[301], stage0_23[302], stage0_23[303], stage0_23[304], stage0_23[305]},
      {stage1_25[50],stage1_24[98],stage1_23[104],stage1_22[139],stage1_21[200]}
   );
   gpc615_5 gpc927 (
      {stage0_21[331], stage0_21[332], stage0_21[333], stage0_21[334], stage0_21[335]},
      {stage0_22[299]},
      {stage0_23[306], stage0_23[307], stage0_23[308], stage0_23[309], stage0_23[310], stage0_23[311]},
      {stage1_25[51],stage1_24[99],stage1_23[105],stage1_22[140],stage1_21[201]}
   );
   gpc615_5 gpc928 (
      {stage0_21[336], stage0_21[337], stage0_21[338], stage0_21[339], stage0_21[340]},
      {stage0_22[300]},
      {stage0_23[312], stage0_23[313], stage0_23[314], stage0_23[315], stage0_23[316], stage0_23[317]},
      {stage1_25[52],stage1_24[100],stage1_23[106],stage1_22[141],stage1_21[202]}
   );
   gpc615_5 gpc929 (
      {stage0_21[341], stage0_21[342], stage0_21[343], stage0_21[344], stage0_21[345]},
      {stage0_22[301]},
      {stage0_23[318], stage0_23[319], stage0_23[320], stage0_23[321], stage0_23[322], stage0_23[323]},
      {stage1_25[53],stage1_24[101],stage1_23[107],stage1_22[142],stage1_21[203]}
   );
   gpc615_5 gpc930 (
      {stage0_21[346], stage0_21[347], stage0_21[348], stage0_21[349], stage0_21[350]},
      {stage0_22[302]},
      {stage0_23[324], stage0_23[325], stage0_23[326], stage0_23[327], stage0_23[328], stage0_23[329]},
      {stage1_25[54],stage1_24[102],stage1_23[108],stage1_22[143],stage1_21[204]}
   );
   gpc615_5 gpc931 (
      {stage0_21[351], stage0_21[352], stage0_21[353], stage0_21[354], stage0_21[355]},
      {stage0_22[303]},
      {stage0_23[330], stage0_23[331], stage0_23[332], stage0_23[333], stage0_23[334], stage0_23[335]},
      {stage1_25[55],stage1_24[103],stage1_23[109],stage1_22[144],stage1_21[205]}
   );
   gpc615_5 gpc932 (
      {stage0_21[356], stage0_21[357], stage0_21[358], stage0_21[359], stage0_21[360]},
      {stage0_22[304]},
      {stage0_23[336], stage0_23[337], stage0_23[338], stage0_23[339], stage0_23[340], stage0_23[341]},
      {stage1_25[56],stage1_24[104],stage1_23[110],stage1_22[145],stage1_21[206]}
   );
   gpc615_5 gpc933 (
      {stage0_21[361], stage0_21[362], stage0_21[363], stage0_21[364], stage0_21[365]},
      {stage0_22[305]},
      {stage0_23[342], stage0_23[343], stage0_23[344], stage0_23[345], stage0_23[346], stage0_23[347]},
      {stage1_25[57],stage1_24[105],stage1_23[111],stage1_22[146],stage1_21[207]}
   );
   gpc615_5 gpc934 (
      {stage0_21[366], stage0_21[367], stage0_21[368], stage0_21[369], stage0_21[370]},
      {stage0_22[306]},
      {stage0_23[348], stage0_23[349], stage0_23[350], stage0_23[351], stage0_23[352], stage0_23[353]},
      {stage1_25[58],stage1_24[106],stage1_23[112],stage1_22[147],stage1_21[208]}
   );
   gpc615_5 gpc935 (
      {stage0_21[371], stage0_21[372], stage0_21[373], stage0_21[374], stage0_21[375]},
      {stage0_22[307]},
      {stage0_23[354], stage0_23[355], stage0_23[356], stage0_23[357], stage0_23[358], stage0_23[359]},
      {stage1_25[59],stage1_24[107],stage1_23[113],stage1_22[148],stage1_21[209]}
   );
   gpc615_5 gpc936 (
      {stage0_21[376], stage0_21[377], stage0_21[378], stage0_21[379], stage0_21[380]},
      {stage0_22[308]},
      {stage0_23[360], stage0_23[361], stage0_23[362], stage0_23[363], stage0_23[364], stage0_23[365]},
      {stage1_25[60],stage1_24[108],stage1_23[114],stage1_22[149],stage1_21[210]}
   );
   gpc615_5 gpc937 (
      {stage0_21[381], stage0_21[382], stage0_21[383], stage0_21[384], stage0_21[385]},
      {stage0_22[309]},
      {stage0_23[366], stage0_23[367], stage0_23[368], stage0_23[369], stage0_23[370], stage0_23[371]},
      {stage1_25[61],stage1_24[109],stage1_23[115],stage1_22[150],stage1_21[211]}
   );
   gpc615_5 gpc938 (
      {stage0_21[386], stage0_21[387], stage0_21[388], stage0_21[389], stage0_21[390]},
      {stage0_22[310]},
      {stage0_23[372], stage0_23[373], stage0_23[374], stage0_23[375], stage0_23[376], stage0_23[377]},
      {stage1_25[62],stage1_24[110],stage1_23[116],stage1_22[151],stage1_21[212]}
   );
   gpc615_5 gpc939 (
      {stage0_21[391], stage0_21[392], stage0_21[393], stage0_21[394], stage0_21[395]},
      {stage0_22[311]},
      {stage0_23[378], stage0_23[379], stage0_23[380], stage0_23[381], stage0_23[382], stage0_23[383]},
      {stage1_25[63],stage1_24[111],stage1_23[117],stage1_22[152],stage1_21[213]}
   );
   gpc615_5 gpc940 (
      {stage0_21[396], stage0_21[397], stage0_21[398], stage0_21[399], stage0_21[400]},
      {stage0_22[312]},
      {stage0_23[384], stage0_23[385], stage0_23[386], stage0_23[387], stage0_23[388], stage0_23[389]},
      {stage1_25[64],stage1_24[112],stage1_23[118],stage1_22[153],stage1_21[214]}
   );
   gpc615_5 gpc941 (
      {stage0_21[401], stage0_21[402], stage0_21[403], stage0_21[404], stage0_21[405]},
      {stage0_22[313]},
      {stage0_23[390], stage0_23[391], stage0_23[392], stage0_23[393], stage0_23[394], stage0_23[395]},
      {stage1_25[65],stage1_24[113],stage1_23[119],stage1_22[154],stage1_21[215]}
   );
   gpc615_5 gpc942 (
      {stage0_21[406], stage0_21[407], stage0_21[408], stage0_21[409], stage0_21[410]},
      {stage0_22[314]},
      {stage0_23[396], stage0_23[397], stage0_23[398], stage0_23[399], stage0_23[400], stage0_23[401]},
      {stage1_25[66],stage1_24[114],stage1_23[120],stage1_22[155],stage1_21[216]}
   );
   gpc615_5 gpc943 (
      {stage0_21[411], stage0_21[412], stage0_21[413], stage0_21[414], stage0_21[415]},
      {stage0_22[315]},
      {stage0_23[402], stage0_23[403], stage0_23[404], stage0_23[405], stage0_23[406], stage0_23[407]},
      {stage1_25[67],stage1_24[115],stage1_23[121],stage1_22[156],stage1_21[217]}
   );
   gpc615_5 gpc944 (
      {stage0_21[416], stage0_21[417], stage0_21[418], stage0_21[419], stage0_21[420]},
      {stage0_22[316]},
      {stage0_23[408], stage0_23[409], stage0_23[410], stage0_23[411], stage0_23[412], stage0_23[413]},
      {stage1_25[68],stage1_24[116],stage1_23[122],stage1_22[157],stage1_21[218]}
   );
   gpc615_5 gpc945 (
      {stage0_21[421], stage0_21[422], stage0_21[423], stage0_21[424], stage0_21[425]},
      {stage0_22[317]},
      {stage0_23[414], stage0_23[415], stage0_23[416], stage0_23[417], stage0_23[418], stage0_23[419]},
      {stage1_25[69],stage1_24[117],stage1_23[123],stage1_22[158],stage1_21[219]}
   );
   gpc615_5 gpc946 (
      {stage0_21[426], stage0_21[427], stage0_21[428], stage0_21[429], stage0_21[430]},
      {stage0_22[318]},
      {stage0_23[420], stage0_23[421], stage0_23[422], stage0_23[423], stage0_23[424], stage0_23[425]},
      {stage1_25[70],stage1_24[118],stage1_23[124],stage1_22[159],stage1_21[220]}
   );
   gpc615_5 gpc947 (
      {stage0_21[431], stage0_21[432], stage0_21[433], stage0_21[434], stage0_21[435]},
      {stage0_22[319]},
      {stage0_23[426], stage0_23[427], stage0_23[428], stage0_23[429], stage0_23[430], stage0_23[431]},
      {stage1_25[71],stage1_24[119],stage1_23[125],stage1_22[160],stage1_21[221]}
   );
   gpc615_5 gpc948 (
      {stage0_21[436], stage0_21[437], stage0_21[438], stage0_21[439], stage0_21[440]},
      {stage0_22[320]},
      {stage0_23[432], stage0_23[433], stage0_23[434], stage0_23[435], stage0_23[436], stage0_23[437]},
      {stage1_25[72],stage1_24[120],stage1_23[126],stage1_22[161],stage1_21[222]}
   );
   gpc615_5 gpc949 (
      {stage0_21[441], stage0_21[442], stage0_21[443], stage0_21[444], stage0_21[445]},
      {stage0_22[321]},
      {stage0_23[438], stage0_23[439], stage0_23[440], stage0_23[441], stage0_23[442], stage0_23[443]},
      {stage1_25[73],stage1_24[121],stage1_23[127],stage1_22[162],stage1_21[223]}
   );
   gpc615_5 gpc950 (
      {stage0_21[446], stage0_21[447], stage0_21[448], stage0_21[449], stage0_21[450]},
      {stage0_22[322]},
      {stage0_23[444], stage0_23[445], stage0_23[446], stage0_23[447], stage0_23[448], stage0_23[449]},
      {stage1_25[74],stage1_24[122],stage1_23[128],stage1_22[163],stage1_21[224]}
   );
   gpc615_5 gpc951 (
      {stage0_21[451], stage0_21[452], stage0_21[453], stage0_21[454], stage0_21[455]},
      {stage0_22[323]},
      {stage0_23[450], stage0_23[451], stage0_23[452], stage0_23[453], stage0_23[454], stage0_23[455]},
      {stage1_25[75],stage1_24[123],stage1_23[129],stage1_22[164],stage1_21[225]}
   );
   gpc615_5 gpc952 (
      {stage0_21[456], stage0_21[457], stage0_21[458], stage0_21[459], stage0_21[460]},
      {stage0_22[324]},
      {stage0_23[456], stage0_23[457], stage0_23[458], stage0_23[459], stage0_23[460], stage0_23[461]},
      {stage1_25[76],stage1_24[124],stage1_23[130],stage1_22[165],stage1_21[226]}
   );
   gpc615_5 gpc953 (
      {stage0_21[461], stage0_21[462], stage0_21[463], stage0_21[464], stage0_21[465]},
      {stage0_22[325]},
      {stage0_23[462], stage0_23[463], stage0_23[464], stage0_23[465], stage0_23[466], stage0_23[467]},
      {stage1_25[77],stage1_24[125],stage1_23[131],stage1_22[166],stage1_21[227]}
   );
   gpc615_5 gpc954 (
      {stage0_21[466], stage0_21[467], stage0_21[468], stage0_21[469], stage0_21[470]},
      {stage0_22[326]},
      {stage0_23[468], stage0_23[469], stage0_23[470], stage0_23[471], stage0_23[472], stage0_23[473]},
      {stage1_25[78],stage1_24[126],stage1_23[132],stage1_22[167],stage1_21[228]}
   );
   gpc606_5 gpc955 (
      {stage0_22[327], stage0_22[328], stage0_22[329], stage0_22[330], stage0_22[331], stage0_22[332]},
      {stage0_24[0], stage0_24[1], stage0_24[2], stage0_24[3], stage0_24[4], stage0_24[5]},
      {stage1_26[0],stage1_25[79],stage1_24[127],stage1_23[133],stage1_22[168]}
   );
   gpc606_5 gpc956 (
      {stage0_22[333], stage0_22[334], stage0_22[335], stage0_22[336], stage0_22[337], stage0_22[338]},
      {stage0_24[6], stage0_24[7], stage0_24[8], stage0_24[9], stage0_24[10], stage0_24[11]},
      {stage1_26[1],stage1_25[80],stage1_24[128],stage1_23[134],stage1_22[169]}
   );
   gpc606_5 gpc957 (
      {stage0_22[339], stage0_22[340], stage0_22[341], stage0_22[342], stage0_22[343], stage0_22[344]},
      {stage0_24[12], stage0_24[13], stage0_24[14], stage0_24[15], stage0_24[16], stage0_24[17]},
      {stage1_26[2],stage1_25[81],stage1_24[129],stage1_23[135],stage1_22[170]}
   );
   gpc606_5 gpc958 (
      {stage0_22[345], stage0_22[346], stage0_22[347], stage0_22[348], stage0_22[349], stage0_22[350]},
      {stage0_24[18], stage0_24[19], stage0_24[20], stage0_24[21], stage0_24[22], stage0_24[23]},
      {stage1_26[3],stage1_25[82],stage1_24[130],stage1_23[136],stage1_22[171]}
   );
   gpc606_5 gpc959 (
      {stage0_22[351], stage0_22[352], stage0_22[353], stage0_22[354], stage0_22[355], stage0_22[356]},
      {stage0_24[24], stage0_24[25], stage0_24[26], stage0_24[27], stage0_24[28], stage0_24[29]},
      {stage1_26[4],stage1_25[83],stage1_24[131],stage1_23[137],stage1_22[172]}
   );
   gpc606_5 gpc960 (
      {stage0_22[357], stage0_22[358], stage0_22[359], stage0_22[360], stage0_22[361], stage0_22[362]},
      {stage0_24[30], stage0_24[31], stage0_24[32], stage0_24[33], stage0_24[34], stage0_24[35]},
      {stage1_26[5],stage1_25[84],stage1_24[132],stage1_23[138],stage1_22[173]}
   );
   gpc606_5 gpc961 (
      {stage0_22[363], stage0_22[364], stage0_22[365], stage0_22[366], stage0_22[367], stage0_22[368]},
      {stage0_24[36], stage0_24[37], stage0_24[38], stage0_24[39], stage0_24[40], stage0_24[41]},
      {stage1_26[6],stage1_25[85],stage1_24[133],stage1_23[139],stage1_22[174]}
   );
   gpc606_5 gpc962 (
      {stage0_22[369], stage0_22[370], stage0_22[371], stage0_22[372], stage0_22[373], stage0_22[374]},
      {stage0_24[42], stage0_24[43], stage0_24[44], stage0_24[45], stage0_24[46], stage0_24[47]},
      {stage1_26[7],stage1_25[86],stage1_24[134],stage1_23[140],stage1_22[175]}
   );
   gpc606_5 gpc963 (
      {stage0_22[375], stage0_22[376], stage0_22[377], stage0_22[378], stage0_22[379], stage0_22[380]},
      {stage0_24[48], stage0_24[49], stage0_24[50], stage0_24[51], stage0_24[52], stage0_24[53]},
      {stage1_26[8],stage1_25[87],stage1_24[135],stage1_23[141],stage1_22[176]}
   );
   gpc606_5 gpc964 (
      {stage0_22[381], stage0_22[382], stage0_22[383], stage0_22[384], stage0_22[385], stage0_22[386]},
      {stage0_24[54], stage0_24[55], stage0_24[56], stage0_24[57], stage0_24[58], stage0_24[59]},
      {stage1_26[9],stage1_25[88],stage1_24[136],stage1_23[142],stage1_22[177]}
   );
   gpc606_5 gpc965 (
      {stage0_22[387], stage0_22[388], stage0_22[389], stage0_22[390], stage0_22[391], stage0_22[392]},
      {stage0_24[60], stage0_24[61], stage0_24[62], stage0_24[63], stage0_24[64], stage0_24[65]},
      {stage1_26[10],stage1_25[89],stage1_24[137],stage1_23[143],stage1_22[178]}
   );
   gpc615_5 gpc966 (
      {stage0_22[393], stage0_22[394], stage0_22[395], stage0_22[396], stage0_22[397]},
      {stage0_23[474]},
      {stage0_24[66], stage0_24[67], stage0_24[68], stage0_24[69], stage0_24[70], stage0_24[71]},
      {stage1_26[11],stage1_25[90],stage1_24[138],stage1_23[144],stage1_22[179]}
   );
   gpc615_5 gpc967 (
      {stage0_22[398], stage0_22[399], stage0_22[400], stage0_22[401], stage0_22[402]},
      {stage0_23[475]},
      {stage0_24[72], stage0_24[73], stage0_24[74], stage0_24[75], stage0_24[76], stage0_24[77]},
      {stage1_26[12],stage1_25[91],stage1_24[139],stage1_23[145],stage1_22[180]}
   );
   gpc615_5 gpc968 (
      {stage0_22[403], stage0_22[404], stage0_22[405], stage0_22[406], stage0_22[407]},
      {stage0_23[476]},
      {stage0_24[78], stage0_24[79], stage0_24[80], stage0_24[81], stage0_24[82], stage0_24[83]},
      {stage1_26[13],stage1_25[92],stage1_24[140],stage1_23[146],stage1_22[181]}
   );
   gpc615_5 gpc969 (
      {stage0_22[408], stage0_22[409], stage0_22[410], stage0_22[411], stage0_22[412]},
      {stage0_23[477]},
      {stage0_24[84], stage0_24[85], stage0_24[86], stage0_24[87], stage0_24[88], stage0_24[89]},
      {stage1_26[14],stage1_25[93],stage1_24[141],stage1_23[147],stage1_22[182]}
   );
   gpc615_5 gpc970 (
      {stage0_22[413], stage0_22[414], stage0_22[415], stage0_22[416], stage0_22[417]},
      {stage0_23[478]},
      {stage0_24[90], stage0_24[91], stage0_24[92], stage0_24[93], stage0_24[94], stage0_24[95]},
      {stage1_26[15],stage1_25[94],stage1_24[142],stage1_23[148],stage1_22[183]}
   );
   gpc615_5 gpc971 (
      {stage0_22[418], stage0_22[419], stage0_22[420], stage0_22[421], stage0_22[422]},
      {stage0_23[479]},
      {stage0_24[96], stage0_24[97], stage0_24[98], stage0_24[99], stage0_24[100], stage0_24[101]},
      {stage1_26[16],stage1_25[95],stage1_24[143],stage1_23[149],stage1_22[184]}
   );
   gpc615_5 gpc972 (
      {stage0_23[480], stage0_23[481], stage0_23[482], stage0_23[483], stage0_23[484]},
      {stage0_24[102]},
      {stage0_25[0], stage0_25[1], stage0_25[2], stage0_25[3], stage0_25[4], stage0_25[5]},
      {stage1_27[0],stage1_26[17],stage1_25[96],stage1_24[144],stage1_23[150]}
   );
   gpc615_5 gpc973 (
      {stage0_23[485], stage0_23[486], stage0_23[487], stage0_23[488], stage0_23[489]},
      {stage0_24[103]},
      {stage0_25[6], stage0_25[7], stage0_25[8], stage0_25[9], stage0_25[10], stage0_25[11]},
      {stage1_27[1],stage1_26[18],stage1_25[97],stage1_24[145],stage1_23[151]}
   );
   gpc615_5 gpc974 (
      {stage0_23[490], stage0_23[491], stage0_23[492], stage0_23[493], stage0_23[494]},
      {stage0_24[104]},
      {stage0_25[12], stage0_25[13], stage0_25[14], stage0_25[15], stage0_25[16], stage0_25[17]},
      {stage1_27[2],stage1_26[19],stage1_25[98],stage1_24[146],stage1_23[152]}
   );
   gpc615_5 gpc975 (
      {stage0_23[495], stage0_23[496], stage0_23[497], stage0_23[498], stage0_23[499]},
      {stage0_24[105]},
      {stage0_25[18], stage0_25[19], stage0_25[20], stage0_25[21], stage0_25[22], stage0_25[23]},
      {stage1_27[3],stage1_26[20],stage1_25[99],stage1_24[147],stage1_23[153]}
   );
   gpc606_5 gpc976 (
      {stage0_24[106], stage0_24[107], stage0_24[108], stage0_24[109], stage0_24[110], stage0_24[111]},
      {stage0_26[0], stage0_26[1], stage0_26[2], stage0_26[3], stage0_26[4], stage0_26[5]},
      {stage1_28[0],stage1_27[4],stage1_26[21],stage1_25[100],stage1_24[148]}
   );
   gpc606_5 gpc977 (
      {stage0_24[112], stage0_24[113], stage0_24[114], stage0_24[115], stage0_24[116], stage0_24[117]},
      {stage0_26[6], stage0_26[7], stage0_26[8], stage0_26[9], stage0_26[10], stage0_26[11]},
      {stage1_28[1],stage1_27[5],stage1_26[22],stage1_25[101],stage1_24[149]}
   );
   gpc606_5 gpc978 (
      {stage0_24[118], stage0_24[119], stage0_24[120], stage0_24[121], stage0_24[122], stage0_24[123]},
      {stage0_26[12], stage0_26[13], stage0_26[14], stage0_26[15], stage0_26[16], stage0_26[17]},
      {stage1_28[2],stage1_27[6],stage1_26[23],stage1_25[102],stage1_24[150]}
   );
   gpc606_5 gpc979 (
      {stage0_24[124], stage0_24[125], stage0_24[126], stage0_24[127], stage0_24[128], stage0_24[129]},
      {stage0_26[18], stage0_26[19], stage0_26[20], stage0_26[21], stage0_26[22], stage0_26[23]},
      {stage1_28[3],stage1_27[7],stage1_26[24],stage1_25[103],stage1_24[151]}
   );
   gpc606_5 gpc980 (
      {stage0_24[130], stage0_24[131], stage0_24[132], stage0_24[133], stage0_24[134], stage0_24[135]},
      {stage0_26[24], stage0_26[25], stage0_26[26], stage0_26[27], stage0_26[28], stage0_26[29]},
      {stage1_28[4],stage1_27[8],stage1_26[25],stage1_25[104],stage1_24[152]}
   );
   gpc606_5 gpc981 (
      {stage0_24[136], stage0_24[137], stage0_24[138], stage0_24[139], stage0_24[140], stage0_24[141]},
      {stage0_26[30], stage0_26[31], stage0_26[32], stage0_26[33], stage0_26[34], stage0_26[35]},
      {stage1_28[5],stage1_27[9],stage1_26[26],stage1_25[105],stage1_24[153]}
   );
   gpc606_5 gpc982 (
      {stage0_24[142], stage0_24[143], stage0_24[144], stage0_24[145], stage0_24[146], stage0_24[147]},
      {stage0_26[36], stage0_26[37], stage0_26[38], stage0_26[39], stage0_26[40], stage0_26[41]},
      {stage1_28[6],stage1_27[10],stage1_26[27],stage1_25[106],stage1_24[154]}
   );
   gpc606_5 gpc983 (
      {stage0_24[148], stage0_24[149], stage0_24[150], stage0_24[151], stage0_24[152], stage0_24[153]},
      {stage0_26[42], stage0_26[43], stage0_26[44], stage0_26[45], stage0_26[46], stage0_26[47]},
      {stage1_28[7],stage1_27[11],stage1_26[28],stage1_25[107],stage1_24[155]}
   );
   gpc606_5 gpc984 (
      {stage0_24[154], stage0_24[155], stage0_24[156], stage0_24[157], stage0_24[158], stage0_24[159]},
      {stage0_26[48], stage0_26[49], stage0_26[50], stage0_26[51], stage0_26[52], stage0_26[53]},
      {stage1_28[8],stage1_27[12],stage1_26[29],stage1_25[108],stage1_24[156]}
   );
   gpc606_5 gpc985 (
      {stage0_24[160], stage0_24[161], stage0_24[162], stage0_24[163], stage0_24[164], stage0_24[165]},
      {stage0_26[54], stage0_26[55], stage0_26[56], stage0_26[57], stage0_26[58], stage0_26[59]},
      {stage1_28[9],stage1_27[13],stage1_26[30],stage1_25[109],stage1_24[157]}
   );
   gpc606_5 gpc986 (
      {stage0_24[166], stage0_24[167], stage0_24[168], stage0_24[169], stage0_24[170], stage0_24[171]},
      {stage0_26[60], stage0_26[61], stage0_26[62], stage0_26[63], stage0_26[64], stage0_26[65]},
      {stage1_28[10],stage1_27[14],stage1_26[31],stage1_25[110],stage1_24[158]}
   );
   gpc606_5 gpc987 (
      {stage0_24[172], stage0_24[173], stage0_24[174], stage0_24[175], stage0_24[176], stage0_24[177]},
      {stage0_26[66], stage0_26[67], stage0_26[68], stage0_26[69], stage0_26[70], stage0_26[71]},
      {stage1_28[11],stage1_27[15],stage1_26[32],stage1_25[111],stage1_24[159]}
   );
   gpc606_5 gpc988 (
      {stage0_24[178], stage0_24[179], stage0_24[180], stage0_24[181], stage0_24[182], stage0_24[183]},
      {stage0_26[72], stage0_26[73], stage0_26[74], stage0_26[75], stage0_26[76], stage0_26[77]},
      {stage1_28[12],stage1_27[16],stage1_26[33],stage1_25[112],stage1_24[160]}
   );
   gpc606_5 gpc989 (
      {stage0_24[184], stage0_24[185], stage0_24[186], stage0_24[187], stage0_24[188], stage0_24[189]},
      {stage0_26[78], stage0_26[79], stage0_26[80], stage0_26[81], stage0_26[82], stage0_26[83]},
      {stage1_28[13],stage1_27[17],stage1_26[34],stage1_25[113],stage1_24[161]}
   );
   gpc606_5 gpc990 (
      {stage0_24[190], stage0_24[191], stage0_24[192], stage0_24[193], stage0_24[194], stage0_24[195]},
      {stage0_26[84], stage0_26[85], stage0_26[86], stage0_26[87], stage0_26[88], stage0_26[89]},
      {stage1_28[14],stage1_27[18],stage1_26[35],stage1_25[114],stage1_24[162]}
   );
   gpc606_5 gpc991 (
      {stage0_24[196], stage0_24[197], stage0_24[198], stage0_24[199], stage0_24[200], stage0_24[201]},
      {stage0_26[90], stage0_26[91], stage0_26[92], stage0_26[93], stage0_26[94], stage0_26[95]},
      {stage1_28[15],stage1_27[19],stage1_26[36],stage1_25[115],stage1_24[163]}
   );
   gpc606_5 gpc992 (
      {stage0_24[202], stage0_24[203], stage0_24[204], stage0_24[205], stage0_24[206], stage0_24[207]},
      {stage0_26[96], stage0_26[97], stage0_26[98], stage0_26[99], stage0_26[100], stage0_26[101]},
      {stage1_28[16],stage1_27[20],stage1_26[37],stage1_25[116],stage1_24[164]}
   );
   gpc606_5 gpc993 (
      {stage0_24[208], stage0_24[209], stage0_24[210], stage0_24[211], stage0_24[212], stage0_24[213]},
      {stage0_26[102], stage0_26[103], stage0_26[104], stage0_26[105], stage0_26[106], stage0_26[107]},
      {stage1_28[17],stage1_27[21],stage1_26[38],stage1_25[117],stage1_24[165]}
   );
   gpc606_5 gpc994 (
      {stage0_24[214], stage0_24[215], stage0_24[216], stage0_24[217], stage0_24[218], stage0_24[219]},
      {stage0_26[108], stage0_26[109], stage0_26[110], stage0_26[111], stage0_26[112], stage0_26[113]},
      {stage1_28[18],stage1_27[22],stage1_26[39],stage1_25[118],stage1_24[166]}
   );
   gpc606_5 gpc995 (
      {stage0_24[220], stage0_24[221], stage0_24[222], stage0_24[223], stage0_24[224], stage0_24[225]},
      {stage0_26[114], stage0_26[115], stage0_26[116], stage0_26[117], stage0_26[118], stage0_26[119]},
      {stage1_28[19],stage1_27[23],stage1_26[40],stage1_25[119],stage1_24[167]}
   );
   gpc606_5 gpc996 (
      {stage0_24[226], stage0_24[227], stage0_24[228], stage0_24[229], stage0_24[230], stage0_24[231]},
      {stage0_26[120], stage0_26[121], stage0_26[122], stage0_26[123], stage0_26[124], stage0_26[125]},
      {stage1_28[20],stage1_27[24],stage1_26[41],stage1_25[120],stage1_24[168]}
   );
   gpc606_5 gpc997 (
      {stage0_24[232], stage0_24[233], stage0_24[234], stage0_24[235], stage0_24[236], stage0_24[237]},
      {stage0_26[126], stage0_26[127], stage0_26[128], stage0_26[129], stage0_26[130], stage0_26[131]},
      {stage1_28[21],stage1_27[25],stage1_26[42],stage1_25[121],stage1_24[169]}
   );
   gpc606_5 gpc998 (
      {stage0_24[238], stage0_24[239], stage0_24[240], stage0_24[241], stage0_24[242], stage0_24[243]},
      {stage0_26[132], stage0_26[133], stage0_26[134], stage0_26[135], stage0_26[136], stage0_26[137]},
      {stage1_28[22],stage1_27[26],stage1_26[43],stage1_25[122],stage1_24[170]}
   );
   gpc606_5 gpc999 (
      {stage0_24[244], stage0_24[245], stage0_24[246], stage0_24[247], stage0_24[248], stage0_24[249]},
      {stage0_26[138], stage0_26[139], stage0_26[140], stage0_26[141], stage0_26[142], stage0_26[143]},
      {stage1_28[23],stage1_27[27],stage1_26[44],stage1_25[123],stage1_24[171]}
   );
   gpc606_5 gpc1000 (
      {stage0_24[250], stage0_24[251], stage0_24[252], stage0_24[253], stage0_24[254], stage0_24[255]},
      {stage0_26[144], stage0_26[145], stage0_26[146], stage0_26[147], stage0_26[148], stage0_26[149]},
      {stage1_28[24],stage1_27[28],stage1_26[45],stage1_25[124],stage1_24[172]}
   );
   gpc606_5 gpc1001 (
      {stage0_24[256], stage0_24[257], stage0_24[258], stage0_24[259], stage0_24[260], stage0_24[261]},
      {stage0_26[150], stage0_26[151], stage0_26[152], stage0_26[153], stage0_26[154], stage0_26[155]},
      {stage1_28[25],stage1_27[29],stage1_26[46],stage1_25[125],stage1_24[173]}
   );
   gpc606_5 gpc1002 (
      {stage0_24[262], stage0_24[263], stage0_24[264], stage0_24[265], stage0_24[266], stage0_24[267]},
      {stage0_26[156], stage0_26[157], stage0_26[158], stage0_26[159], stage0_26[160], stage0_26[161]},
      {stage1_28[26],stage1_27[30],stage1_26[47],stage1_25[126],stage1_24[174]}
   );
   gpc606_5 gpc1003 (
      {stage0_24[268], stage0_24[269], stage0_24[270], stage0_24[271], stage0_24[272], stage0_24[273]},
      {stage0_26[162], stage0_26[163], stage0_26[164], stage0_26[165], stage0_26[166], stage0_26[167]},
      {stage1_28[27],stage1_27[31],stage1_26[48],stage1_25[127],stage1_24[175]}
   );
   gpc606_5 gpc1004 (
      {stage0_24[274], stage0_24[275], stage0_24[276], stage0_24[277], stage0_24[278], stage0_24[279]},
      {stage0_26[168], stage0_26[169], stage0_26[170], stage0_26[171], stage0_26[172], stage0_26[173]},
      {stage1_28[28],stage1_27[32],stage1_26[49],stage1_25[128],stage1_24[176]}
   );
   gpc606_5 gpc1005 (
      {stage0_24[280], stage0_24[281], stage0_24[282], stage0_24[283], stage0_24[284], stage0_24[285]},
      {stage0_26[174], stage0_26[175], stage0_26[176], stage0_26[177], stage0_26[178], stage0_26[179]},
      {stage1_28[29],stage1_27[33],stage1_26[50],stage1_25[129],stage1_24[177]}
   );
   gpc606_5 gpc1006 (
      {stage0_24[286], stage0_24[287], stage0_24[288], stage0_24[289], stage0_24[290], stage0_24[291]},
      {stage0_26[180], stage0_26[181], stage0_26[182], stage0_26[183], stage0_26[184], stage0_26[185]},
      {stage1_28[30],stage1_27[34],stage1_26[51],stage1_25[130],stage1_24[178]}
   );
   gpc606_5 gpc1007 (
      {stage0_24[292], stage0_24[293], stage0_24[294], stage0_24[295], stage0_24[296], stage0_24[297]},
      {stage0_26[186], stage0_26[187], stage0_26[188], stage0_26[189], stage0_26[190], stage0_26[191]},
      {stage1_28[31],stage1_27[35],stage1_26[52],stage1_25[131],stage1_24[179]}
   );
   gpc606_5 gpc1008 (
      {stage0_24[298], stage0_24[299], stage0_24[300], stage0_24[301], stage0_24[302], stage0_24[303]},
      {stage0_26[192], stage0_26[193], stage0_26[194], stage0_26[195], stage0_26[196], stage0_26[197]},
      {stage1_28[32],stage1_27[36],stage1_26[53],stage1_25[132],stage1_24[180]}
   );
   gpc606_5 gpc1009 (
      {stage0_24[304], stage0_24[305], stage0_24[306], stage0_24[307], stage0_24[308], stage0_24[309]},
      {stage0_26[198], stage0_26[199], stage0_26[200], stage0_26[201], stage0_26[202], stage0_26[203]},
      {stage1_28[33],stage1_27[37],stage1_26[54],stage1_25[133],stage1_24[181]}
   );
   gpc606_5 gpc1010 (
      {stage0_24[310], stage0_24[311], stage0_24[312], stage0_24[313], stage0_24[314], stage0_24[315]},
      {stage0_26[204], stage0_26[205], stage0_26[206], stage0_26[207], stage0_26[208], stage0_26[209]},
      {stage1_28[34],stage1_27[38],stage1_26[55],stage1_25[134],stage1_24[182]}
   );
   gpc606_5 gpc1011 (
      {stage0_24[316], stage0_24[317], stage0_24[318], stage0_24[319], stage0_24[320], stage0_24[321]},
      {stage0_26[210], stage0_26[211], stage0_26[212], stage0_26[213], stage0_26[214], stage0_26[215]},
      {stage1_28[35],stage1_27[39],stage1_26[56],stage1_25[135],stage1_24[183]}
   );
   gpc606_5 gpc1012 (
      {stage0_24[322], stage0_24[323], stage0_24[324], stage0_24[325], stage0_24[326], stage0_24[327]},
      {stage0_26[216], stage0_26[217], stage0_26[218], stage0_26[219], stage0_26[220], stage0_26[221]},
      {stage1_28[36],stage1_27[40],stage1_26[57],stage1_25[136],stage1_24[184]}
   );
   gpc606_5 gpc1013 (
      {stage0_24[328], stage0_24[329], stage0_24[330], stage0_24[331], stage0_24[332], stage0_24[333]},
      {stage0_26[222], stage0_26[223], stage0_26[224], stage0_26[225], stage0_26[226], stage0_26[227]},
      {stage1_28[37],stage1_27[41],stage1_26[58],stage1_25[137],stage1_24[185]}
   );
   gpc606_5 gpc1014 (
      {stage0_24[334], stage0_24[335], stage0_24[336], stage0_24[337], stage0_24[338], stage0_24[339]},
      {stage0_26[228], stage0_26[229], stage0_26[230], stage0_26[231], stage0_26[232], stage0_26[233]},
      {stage1_28[38],stage1_27[42],stage1_26[59],stage1_25[138],stage1_24[186]}
   );
   gpc606_5 gpc1015 (
      {stage0_24[340], stage0_24[341], stage0_24[342], stage0_24[343], stage0_24[344], stage0_24[345]},
      {stage0_26[234], stage0_26[235], stage0_26[236], stage0_26[237], stage0_26[238], stage0_26[239]},
      {stage1_28[39],stage1_27[43],stage1_26[60],stage1_25[139],stage1_24[187]}
   );
   gpc606_5 gpc1016 (
      {stage0_24[346], stage0_24[347], stage0_24[348], stage0_24[349], stage0_24[350], stage0_24[351]},
      {stage0_26[240], stage0_26[241], stage0_26[242], stage0_26[243], stage0_26[244], stage0_26[245]},
      {stage1_28[40],stage1_27[44],stage1_26[61],stage1_25[140],stage1_24[188]}
   );
   gpc615_5 gpc1017 (
      {stage0_24[352], stage0_24[353], stage0_24[354], stage0_24[355], stage0_24[356]},
      {stage0_25[24]},
      {stage0_26[246], stage0_26[247], stage0_26[248], stage0_26[249], stage0_26[250], stage0_26[251]},
      {stage1_28[41],stage1_27[45],stage1_26[62],stage1_25[141],stage1_24[189]}
   );
   gpc615_5 gpc1018 (
      {stage0_24[357], stage0_24[358], stage0_24[359], stage0_24[360], stage0_24[361]},
      {stage0_25[25]},
      {stage0_26[252], stage0_26[253], stage0_26[254], stage0_26[255], stage0_26[256], stage0_26[257]},
      {stage1_28[42],stage1_27[46],stage1_26[63],stage1_25[142],stage1_24[190]}
   );
   gpc615_5 gpc1019 (
      {stage0_24[362], stage0_24[363], stage0_24[364], stage0_24[365], stage0_24[366]},
      {stage0_25[26]},
      {stage0_26[258], stage0_26[259], stage0_26[260], stage0_26[261], stage0_26[262], stage0_26[263]},
      {stage1_28[43],stage1_27[47],stage1_26[64],stage1_25[143],stage1_24[191]}
   );
   gpc615_5 gpc1020 (
      {stage0_24[367], stage0_24[368], stage0_24[369], stage0_24[370], stage0_24[371]},
      {stage0_25[27]},
      {stage0_26[264], stage0_26[265], stage0_26[266], stage0_26[267], stage0_26[268], stage0_26[269]},
      {stage1_28[44],stage1_27[48],stage1_26[65],stage1_25[144],stage1_24[192]}
   );
   gpc615_5 gpc1021 (
      {stage0_24[372], stage0_24[373], stage0_24[374], stage0_24[375], stage0_24[376]},
      {stage0_25[28]},
      {stage0_26[270], stage0_26[271], stage0_26[272], stage0_26[273], stage0_26[274], stage0_26[275]},
      {stage1_28[45],stage1_27[49],stage1_26[66],stage1_25[145],stage1_24[193]}
   );
   gpc615_5 gpc1022 (
      {stage0_24[377], stage0_24[378], stage0_24[379], stage0_24[380], stage0_24[381]},
      {stage0_25[29]},
      {stage0_26[276], stage0_26[277], stage0_26[278], stage0_26[279], stage0_26[280], stage0_26[281]},
      {stage1_28[46],stage1_27[50],stage1_26[67],stage1_25[146],stage1_24[194]}
   );
   gpc615_5 gpc1023 (
      {stage0_24[382], stage0_24[383], stage0_24[384], stage0_24[385], stage0_24[386]},
      {stage0_25[30]},
      {stage0_26[282], stage0_26[283], stage0_26[284], stage0_26[285], stage0_26[286], stage0_26[287]},
      {stage1_28[47],stage1_27[51],stage1_26[68],stage1_25[147],stage1_24[195]}
   );
   gpc615_5 gpc1024 (
      {stage0_24[387], stage0_24[388], stage0_24[389], stage0_24[390], stage0_24[391]},
      {stage0_25[31]},
      {stage0_26[288], stage0_26[289], stage0_26[290], stage0_26[291], stage0_26[292], stage0_26[293]},
      {stage1_28[48],stage1_27[52],stage1_26[69],stage1_25[148],stage1_24[196]}
   );
   gpc615_5 gpc1025 (
      {stage0_24[392], stage0_24[393], stage0_24[394], stage0_24[395], stage0_24[396]},
      {stage0_25[32]},
      {stage0_26[294], stage0_26[295], stage0_26[296], stage0_26[297], stage0_26[298], stage0_26[299]},
      {stage1_28[49],stage1_27[53],stage1_26[70],stage1_25[149],stage1_24[197]}
   );
   gpc615_5 gpc1026 (
      {stage0_24[397], stage0_24[398], stage0_24[399], stage0_24[400], stage0_24[401]},
      {stage0_25[33]},
      {stage0_26[300], stage0_26[301], stage0_26[302], stage0_26[303], stage0_26[304], stage0_26[305]},
      {stage1_28[50],stage1_27[54],stage1_26[71],stage1_25[150],stage1_24[198]}
   );
   gpc615_5 gpc1027 (
      {stage0_24[402], stage0_24[403], stage0_24[404], stage0_24[405], stage0_24[406]},
      {stage0_25[34]},
      {stage0_26[306], stage0_26[307], stage0_26[308], stage0_26[309], stage0_26[310], stage0_26[311]},
      {stage1_28[51],stage1_27[55],stage1_26[72],stage1_25[151],stage1_24[199]}
   );
   gpc615_5 gpc1028 (
      {stage0_24[407], stage0_24[408], stage0_24[409], stage0_24[410], stage0_24[411]},
      {stage0_25[35]},
      {stage0_26[312], stage0_26[313], stage0_26[314], stage0_26[315], stage0_26[316], stage0_26[317]},
      {stage1_28[52],stage1_27[56],stage1_26[73],stage1_25[152],stage1_24[200]}
   );
   gpc615_5 gpc1029 (
      {stage0_24[412], stage0_24[413], stage0_24[414], stage0_24[415], stage0_24[416]},
      {stage0_25[36]},
      {stage0_26[318], stage0_26[319], stage0_26[320], stage0_26[321], stage0_26[322], stage0_26[323]},
      {stage1_28[53],stage1_27[57],stage1_26[74],stage1_25[153],stage1_24[201]}
   );
   gpc615_5 gpc1030 (
      {stage0_24[417], stage0_24[418], stage0_24[419], stage0_24[420], stage0_24[421]},
      {stage0_25[37]},
      {stage0_26[324], stage0_26[325], stage0_26[326], stage0_26[327], stage0_26[328], stage0_26[329]},
      {stage1_28[54],stage1_27[58],stage1_26[75],stage1_25[154],stage1_24[202]}
   );
   gpc615_5 gpc1031 (
      {stage0_24[422], stage0_24[423], stage0_24[424], stage0_24[425], stage0_24[426]},
      {stage0_25[38]},
      {stage0_26[330], stage0_26[331], stage0_26[332], stage0_26[333], stage0_26[334], stage0_26[335]},
      {stage1_28[55],stage1_27[59],stage1_26[76],stage1_25[155],stage1_24[203]}
   );
   gpc615_5 gpc1032 (
      {stage0_24[427], stage0_24[428], stage0_24[429], stage0_24[430], stage0_24[431]},
      {stage0_25[39]},
      {stage0_26[336], stage0_26[337], stage0_26[338], stage0_26[339], stage0_26[340], stage0_26[341]},
      {stage1_28[56],stage1_27[60],stage1_26[77],stage1_25[156],stage1_24[204]}
   );
   gpc615_5 gpc1033 (
      {stage0_24[432], stage0_24[433], stage0_24[434], stage0_24[435], stage0_24[436]},
      {stage0_25[40]},
      {stage0_26[342], stage0_26[343], stage0_26[344], stage0_26[345], stage0_26[346], stage0_26[347]},
      {stage1_28[57],stage1_27[61],stage1_26[78],stage1_25[157],stage1_24[205]}
   );
   gpc615_5 gpc1034 (
      {stage0_24[437], stage0_24[438], stage0_24[439], stage0_24[440], stage0_24[441]},
      {stage0_25[41]},
      {stage0_26[348], stage0_26[349], stage0_26[350], stage0_26[351], stage0_26[352], stage0_26[353]},
      {stage1_28[58],stage1_27[62],stage1_26[79],stage1_25[158],stage1_24[206]}
   );
   gpc615_5 gpc1035 (
      {stage0_24[442], stage0_24[443], stage0_24[444], stage0_24[445], stage0_24[446]},
      {stage0_25[42]},
      {stage0_26[354], stage0_26[355], stage0_26[356], stage0_26[357], stage0_26[358], stage0_26[359]},
      {stage1_28[59],stage1_27[63],stage1_26[80],stage1_25[159],stage1_24[207]}
   );
   gpc615_5 gpc1036 (
      {stage0_24[447], stage0_24[448], stage0_24[449], stage0_24[450], stage0_24[451]},
      {stage0_25[43]},
      {stage0_26[360], stage0_26[361], stage0_26[362], stage0_26[363], stage0_26[364], stage0_26[365]},
      {stage1_28[60],stage1_27[64],stage1_26[81],stage1_25[160],stage1_24[208]}
   );
   gpc615_5 gpc1037 (
      {stage0_24[452], stage0_24[453], stage0_24[454], stage0_24[455], stage0_24[456]},
      {stage0_25[44]},
      {stage0_26[366], stage0_26[367], stage0_26[368], stage0_26[369], stage0_26[370], stage0_26[371]},
      {stage1_28[61],stage1_27[65],stage1_26[82],stage1_25[161],stage1_24[209]}
   );
   gpc615_5 gpc1038 (
      {stage0_24[457], stage0_24[458], stage0_24[459], stage0_24[460], stage0_24[461]},
      {stage0_25[45]},
      {stage0_26[372], stage0_26[373], stage0_26[374], stage0_26[375], stage0_26[376], stage0_26[377]},
      {stage1_28[62],stage1_27[66],stage1_26[83],stage1_25[162],stage1_24[210]}
   );
   gpc615_5 gpc1039 (
      {stage0_24[462], stage0_24[463], stage0_24[464], stage0_24[465], stage0_24[466]},
      {stage0_25[46]},
      {stage0_26[378], stage0_26[379], stage0_26[380], stage0_26[381], stage0_26[382], stage0_26[383]},
      {stage1_28[63],stage1_27[67],stage1_26[84],stage1_25[163],stage1_24[211]}
   );
   gpc615_5 gpc1040 (
      {stage0_24[467], stage0_24[468], stage0_24[469], stage0_24[470], stage0_24[471]},
      {stage0_25[47]},
      {stage0_26[384], stage0_26[385], stage0_26[386], stage0_26[387], stage0_26[388], stage0_26[389]},
      {stage1_28[64],stage1_27[68],stage1_26[85],stage1_25[164],stage1_24[212]}
   );
   gpc615_5 gpc1041 (
      {stage0_24[472], stage0_24[473], stage0_24[474], stage0_24[475], stage0_24[476]},
      {stage0_25[48]},
      {stage0_26[390], stage0_26[391], stage0_26[392], stage0_26[393], stage0_26[394], stage0_26[395]},
      {stage1_28[65],stage1_27[69],stage1_26[86],stage1_25[165],stage1_24[213]}
   );
   gpc615_5 gpc1042 (
      {stage0_24[477], stage0_24[478], stage0_24[479], stage0_24[480], stage0_24[481]},
      {stage0_25[49]},
      {stage0_26[396], stage0_26[397], stage0_26[398], stage0_26[399], stage0_26[400], stage0_26[401]},
      {stage1_28[66],stage1_27[70],stage1_26[87],stage1_25[166],stage1_24[214]}
   );
   gpc615_5 gpc1043 (
      {stage0_24[482], stage0_24[483], stage0_24[484], stage0_24[485], stage0_24[486]},
      {stage0_25[50]},
      {stage0_26[402], stage0_26[403], stage0_26[404], stage0_26[405], stage0_26[406], stage0_26[407]},
      {stage1_28[67],stage1_27[71],stage1_26[88],stage1_25[167],stage1_24[215]}
   );
   gpc615_5 gpc1044 (
      {stage0_24[487], stage0_24[488], stage0_24[489], stage0_24[490], stage0_24[491]},
      {stage0_25[51]},
      {stage0_26[408], stage0_26[409], stage0_26[410], stage0_26[411], stage0_26[412], stage0_26[413]},
      {stage1_28[68],stage1_27[72],stage1_26[89],stage1_25[168],stage1_24[216]}
   );
   gpc615_5 gpc1045 (
      {stage0_24[492], stage0_24[493], stage0_24[494], stage0_24[495], stage0_24[496]},
      {stage0_25[52]},
      {stage0_26[414], stage0_26[415], stage0_26[416], stage0_26[417], stage0_26[418], stage0_26[419]},
      {stage1_28[69],stage1_27[73],stage1_26[90],stage1_25[169],stage1_24[217]}
   );
   gpc615_5 gpc1046 (
      {stage0_24[497], stage0_24[498], stage0_24[499], stage0_24[500], stage0_24[501]},
      {stage0_25[53]},
      {stage0_26[420], stage0_26[421], stage0_26[422], stage0_26[423], stage0_26[424], stage0_26[425]},
      {stage1_28[70],stage1_27[74],stage1_26[91],stage1_25[170],stage1_24[218]}
   );
   gpc615_5 gpc1047 (
      {stage0_24[502], stage0_24[503], stage0_24[504], stage0_24[505], stage0_24[506]},
      {stage0_25[54]},
      {stage0_26[426], stage0_26[427], stage0_26[428], stage0_26[429], stage0_26[430], stage0_26[431]},
      {stage1_28[71],stage1_27[75],stage1_26[92],stage1_25[171],stage1_24[219]}
   );
   gpc615_5 gpc1048 (
      {stage0_24[507], stage0_24[508], stage0_24[509], stage0_24[510], stage0_24[511]},
      {stage0_25[55]},
      {stage0_26[432], stage0_26[433], stage0_26[434], stage0_26[435], stage0_26[436], stage0_26[437]},
      {stage1_28[72],stage1_27[76],stage1_26[93],stage1_25[172],stage1_24[220]}
   );
   gpc606_5 gpc1049 (
      {stage0_25[56], stage0_25[57], stage0_25[58], stage0_25[59], stage0_25[60], stage0_25[61]},
      {stage0_27[0], stage0_27[1], stage0_27[2], stage0_27[3], stage0_27[4], stage0_27[5]},
      {stage1_29[0],stage1_28[73],stage1_27[77],stage1_26[94],stage1_25[173]}
   );
   gpc606_5 gpc1050 (
      {stage0_25[62], stage0_25[63], stage0_25[64], stage0_25[65], stage0_25[66], stage0_25[67]},
      {stage0_27[6], stage0_27[7], stage0_27[8], stage0_27[9], stage0_27[10], stage0_27[11]},
      {stage1_29[1],stage1_28[74],stage1_27[78],stage1_26[95],stage1_25[174]}
   );
   gpc606_5 gpc1051 (
      {stage0_25[68], stage0_25[69], stage0_25[70], stage0_25[71], stage0_25[72], stage0_25[73]},
      {stage0_27[12], stage0_27[13], stage0_27[14], stage0_27[15], stage0_27[16], stage0_27[17]},
      {stage1_29[2],stage1_28[75],stage1_27[79],stage1_26[96],stage1_25[175]}
   );
   gpc606_5 gpc1052 (
      {stage0_25[74], stage0_25[75], stage0_25[76], stage0_25[77], stage0_25[78], stage0_25[79]},
      {stage0_27[18], stage0_27[19], stage0_27[20], stage0_27[21], stage0_27[22], stage0_27[23]},
      {stage1_29[3],stage1_28[76],stage1_27[80],stage1_26[97],stage1_25[176]}
   );
   gpc606_5 gpc1053 (
      {stage0_25[80], stage0_25[81], stage0_25[82], stage0_25[83], stage0_25[84], stage0_25[85]},
      {stage0_27[24], stage0_27[25], stage0_27[26], stage0_27[27], stage0_27[28], stage0_27[29]},
      {stage1_29[4],stage1_28[77],stage1_27[81],stage1_26[98],stage1_25[177]}
   );
   gpc606_5 gpc1054 (
      {stage0_25[86], stage0_25[87], stage0_25[88], stage0_25[89], stage0_25[90], stage0_25[91]},
      {stage0_27[30], stage0_27[31], stage0_27[32], stage0_27[33], stage0_27[34], stage0_27[35]},
      {stage1_29[5],stage1_28[78],stage1_27[82],stage1_26[99],stage1_25[178]}
   );
   gpc606_5 gpc1055 (
      {stage0_25[92], stage0_25[93], stage0_25[94], stage0_25[95], stage0_25[96], stage0_25[97]},
      {stage0_27[36], stage0_27[37], stage0_27[38], stage0_27[39], stage0_27[40], stage0_27[41]},
      {stage1_29[6],stage1_28[79],stage1_27[83],stage1_26[100],stage1_25[179]}
   );
   gpc606_5 gpc1056 (
      {stage0_25[98], stage0_25[99], stage0_25[100], stage0_25[101], stage0_25[102], stage0_25[103]},
      {stage0_27[42], stage0_27[43], stage0_27[44], stage0_27[45], stage0_27[46], stage0_27[47]},
      {stage1_29[7],stage1_28[80],stage1_27[84],stage1_26[101],stage1_25[180]}
   );
   gpc606_5 gpc1057 (
      {stage0_25[104], stage0_25[105], stage0_25[106], stage0_25[107], stage0_25[108], stage0_25[109]},
      {stage0_27[48], stage0_27[49], stage0_27[50], stage0_27[51], stage0_27[52], stage0_27[53]},
      {stage1_29[8],stage1_28[81],stage1_27[85],stage1_26[102],stage1_25[181]}
   );
   gpc606_5 gpc1058 (
      {stage0_25[110], stage0_25[111], stage0_25[112], stage0_25[113], stage0_25[114], stage0_25[115]},
      {stage0_27[54], stage0_27[55], stage0_27[56], stage0_27[57], stage0_27[58], stage0_27[59]},
      {stage1_29[9],stage1_28[82],stage1_27[86],stage1_26[103],stage1_25[182]}
   );
   gpc606_5 gpc1059 (
      {stage0_25[116], stage0_25[117], stage0_25[118], stage0_25[119], stage0_25[120], stage0_25[121]},
      {stage0_27[60], stage0_27[61], stage0_27[62], stage0_27[63], stage0_27[64], stage0_27[65]},
      {stage1_29[10],stage1_28[83],stage1_27[87],stage1_26[104],stage1_25[183]}
   );
   gpc606_5 gpc1060 (
      {stage0_25[122], stage0_25[123], stage0_25[124], stage0_25[125], stage0_25[126], stage0_25[127]},
      {stage0_27[66], stage0_27[67], stage0_27[68], stage0_27[69], stage0_27[70], stage0_27[71]},
      {stage1_29[11],stage1_28[84],stage1_27[88],stage1_26[105],stage1_25[184]}
   );
   gpc606_5 gpc1061 (
      {stage0_25[128], stage0_25[129], stage0_25[130], stage0_25[131], stage0_25[132], stage0_25[133]},
      {stage0_27[72], stage0_27[73], stage0_27[74], stage0_27[75], stage0_27[76], stage0_27[77]},
      {stage1_29[12],stage1_28[85],stage1_27[89],stage1_26[106],stage1_25[185]}
   );
   gpc606_5 gpc1062 (
      {stage0_25[134], stage0_25[135], stage0_25[136], stage0_25[137], stage0_25[138], stage0_25[139]},
      {stage0_27[78], stage0_27[79], stage0_27[80], stage0_27[81], stage0_27[82], stage0_27[83]},
      {stage1_29[13],stage1_28[86],stage1_27[90],stage1_26[107],stage1_25[186]}
   );
   gpc606_5 gpc1063 (
      {stage0_25[140], stage0_25[141], stage0_25[142], stage0_25[143], stage0_25[144], stage0_25[145]},
      {stage0_27[84], stage0_27[85], stage0_27[86], stage0_27[87], stage0_27[88], stage0_27[89]},
      {stage1_29[14],stage1_28[87],stage1_27[91],stage1_26[108],stage1_25[187]}
   );
   gpc606_5 gpc1064 (
      {stage0_25[146], stage0_25[147], stage0_25[148], stage0_25[149], stage0_25[150], stage0_25[151]},
      {stage0_27[90], stage0_27[91], stage0_27[92], stage0_27[93], stage0_27[94], stage0_27[95]},
      {stage1_29[15],stage1_28[88],stage1_27[92],stage1_26[109],stage1_25[188]}
   );
   gpc606_5 gpc1065 (
      {stage0_25[152], stage0_25[153], stage0_25[154], stage0_25[155], stage0_25[156], stage0_25[157]},
      {stage0_27[96], stage0_27[97], stage0_27[98], stage0_27[99], stage0_27[100], stage0_27[101]},
      {stage1_29[16],stage1_28[89],stage1_27[93],stage1_26[110],stage1_25[189]}
   );
   gpc606_5 gpc1066 (
      {stage0_25[158], stage0_25[159], stage0_25[160], stage0_25[161], stage0_25[162], stage0_25[163]},
      {stage0_27[102], stage0_27[103], stage0_27[104], stage0_27[105], stage0_27[106], stage0_27[107]},
      {stage1_29[17],stage1_28[90],stage1_27[94],stage1_26[111],stage1_25[190]}
   );
   gpc606_5 gpc1067 (
      {stage0_25[164], stage0_25[165], stage0_25[166], stage0_25[167], stage0_25[168], stage0_25[169]},
      {stage0_27[108], stage0_27[109], stage0_27[110], stage0_27[111], stage0_27[112], stage0_27[113]},
      {stage1_29[18],stage1_28[91],stage1_27[95],stage1_26[112],stage1_25[191]}
   );
   gpc606_5 gpc1068 (
      {stage0_25[170], stage0_25[171], stage0_25[172], stage0_25[173], stage0_25[174], stage0_25[175]},
      {stage0_27[114], stage0_27[115], stage0_27[116], stage0_27[117], stage0_27[118], stage0_27[119]},
      {stage1_29[19],stage1_28[92],stage1_27[96],stage1_26[113],stage1_25[192]}
   );
   gpc606_5 gpc1069 (
      {stage0_25[176], stage0_25[177], stage0_25[178], stage0_25[179], stage0_25[180], stage0_25[181]},
      {stage0_27[120], stage0_27[121], stage0_27[122], stage0_27[123], stage0_27[124], stage0_27[125]},
      {stage1_29[20],stage1_28[93],stage1_27[97],stage1_26[114],stage1_25[193]}
   );
   gpc606_5 gpc1070 (
      {stage0_25[182], stage0_25[183], stage0_25[184], stage0_25[185], stage0_25[186], stage0_25[187]},
      {stage0_27[126], stage0_27[127], stage0_27[128], stage0_27[129], stage0_27[130], stage0_27[131]},
      {stage1_29[21],stage1_28[94],stage1_27[98],stage1_26[115],stage1_25[194]}
   );
   gpc606_5 gpc1071 (
      {stage0_25[188], stage0_25[189], stage0_25[190], stage0_25[191], stage0_25[192], stage0_25[193]},
      {stage0_27[132], stage0_27[133], stage0_27[134], stage0_27[135], stage0_27[136], stage0_27[137]},
      {stage1_29[22],stage1_28[95],stage1_27[99],stage1_26[116],stage1_25[195]}
   );
   gpc606_5 gpc1072 (
      {stage0_25[194], stage0_25[195], stage0_25[196], stage0_25[197], stage0_25[198], stage0_25[199]},
      {stage0_27[138], stage0_27[139], stage0_27[140], stage0_27[141], stage0_27[142], stage0_27[143]},
      {stage1_29[23],stage1_28[96],stage1_27[100],stage1_26[117],stage1_25[196]}
   );
   gpc606_5 gpc1073 (
      {stage0_25[200], stage0_25[201], stage0_25[202], stage0_25[203], stage0_25[204], stage0_25[205]},
      {stage0_27[144], stage0_27[145], stage0_27[146], stage0_27[147], stage0_27[148], stage0_27[149]},
      {stage1_29[24],stage1_28[97],stage1_27[101],stage1_26[118],stage1_25[197]}
   );
   gpc606_5 gpc1074 (
      {stage0_25[206], stage0_25[207], stage0_25[208], stage0_25[209], stage0_25[210], stage0_25[211]},
      {stage0_27[150], stage0_27[151], stage0_27[152], stage0_27[153], stage0_27[154], stage0_27[155]},
      {stage1_29[25],stage1_28[98],stage1_27[102],stage1_26[119],stage1_25[198]}
   );
   gpc606_5 gpc1075 (
      {stage0_25[212], stage0_25[213], stage0_25[214], stage0_25[215], stage0_25[216], stage0_25[217]},
      {stage0_27[156], stage0_27[157], stage0_27[158], stage0_27[159], stage0_27[160], stage0_27[161]},
      {stage1_29[26],stage1_28[99],stage1_27[103],stage1_26[120],stage1_25[199]}
   );
   gpc606_5 gpc1076 (
      {stage0_25[218], stage0_25[219], stage0_25[220], stage0_25[221], stage0_25[222], stage0_25[223]},
      {stage0_27[162], stage0_27[163], stage0_27[164], stage0_27[165], stage0_27[166], stage0_27[167]},
      {stage1_29[27],stage1_28[100],stage1_27[104],stage1_26[121],stage1_25[200]}
   );
   gpc606_5 gpc1077 (
      {stage0_25[224], stage0_25[225], stage0_25[226], stage0_25[227], stage0_25[228], stage0_25[229]},
      {stage0_27[168], stage0_27[169], stage0_27[170], stage0_27[171], stage0_27[172], stage0_27[173]},
      {stage1_29[28],stage1_28[101],stage1_27[105],stage1_26[122],stage1_25[201]}
   );
   gpc606_5 gpc1078 (
      {stage0_25[230], stage0_25[231], stage0_25[232], stage0_25[233], stage0_25[234], stage0_25[235]},
      {stage0_27[174], stage0_27[175], stage0_27[176], stage0_27[177], stage0_27[178], stage0_27[179]},
      {stage1_29[29],stage1_28[102],stage1_27[106],stage1_26[123],stage1_25[202]}
   );
   gpc606_5 gpc1079 (
      {stage0_25[236], stage0_25[237], stage0_25[238], stage0_25[239], stage0_25[240], stage0_25[241]},
      {stage0_27[180], stage0_27[181], stage0_27[182], stage0_27[183], stage0_27[184], stage0_27[185]},
      {stage1_29[30],stage1_28[103],stage1_27[107],stage1_26[124],stage1_25[203]}
   );
   gpc606_5 gpc1080 (
      {stage0_25[242], stage0_25[243], stage0_25[244], stage0_25[245], stage0_25[246], stage0_25[247]},
      {stage0_27[186], stage0_27[187], stage0_27[188], stage0_27[189], stage0_27[190], stage0_27[191]},
      {stage1_29[31],stage1_28[104],stage1_27[108],stage1_26[125],stage1_25[204]}
   );
   gpc606_5 gpc1081 (
      {stage0_25[248], stage0_25[249], stage0_25[250], stage0_25[251], stage0_25[252], stage0_25[253]},
      {stage0_27[192], stage0_27[193], stage0_27[194], stage0_27[195], stage0_27[196], stage0_27[197]},
      {stage1_29[32],stage1_28[105],stage1_27[109],stage1_26[126],stage1_25[205]}
   );
   gpc606_5 gpc1082 (
      {stage0_25[254], stage0_25[255], stage0_25[256], stage0_25[257], stage0_25[258], stage0_25[259]},
      {stage0_27[198], stage0_27[199], stage0_27[200], stage0_27[201], stage0_27[202], stage0_27[203]},
      {stage1_29[33],stage1_28[106],stage1_27[110],stage1_26[127],stage1_25[206]}
   );
   gpc606_5 gpc1083 (
      {stage0_25[260], stage0_25[261], stage0_25[262], stage0_25[263], stage0_25[264], stage0_25[265]},
      {stage0_27[204], stage0_27[205], stage0_27[206], stage0_27[207], stage0_27[208], stage0_27[209]},
      {stage1_29[34],stage1_28[107],stage1_27[111],stage1_26[128],stage1_25[207]}
   );
   gpc606_5 gpc1084 (
      {stage0_25[266], stage0_25[267], stage0_25[268], stage0_25[269], stage0_25[270], stage0_25[271]},
      {stage0_27[210], stage0_27[211], stage0_27[212], stage0_27[213], stage0_27[214], stage0_27[215]},
      {stage1_29[35],stage1_28[108],stage1_27[112],stage1_26[129],stage1_25[208]}
   );
   gpc606_5 gpc1085 (
      {stage0_25[272], stage0_25[273], stage0_25[274], stage0_25[275], stage0_25[276], stage0_25[277]},
      {stage0_27[216], stage0_27[217], stage0_27[218], stage0_27[219], stage0_27[220], stage0_27[221]},
      {stage1_29[36],stage1_28[109],stage1_27[113],stage1_26[130],stage1_25[209]}
   );
   gpc606_5 gpc1086 (
      {stage0_25[278], stage0_25[279], stage0_25[280], stage0_25[281], stage0_25[282], stage0_25[283]},
      {stage0_27[222], stage0_27[223], stage0_27[224], stage0_27[225], stage0_27[226], stage0_27[227]},
      {stage1_29[37],stage1_28[110],stage1_27[114],stage1_26[131],stage1_25[210]}
   );
   gpc606_5 gpc1087 (
      {stage0_25[284], stage0_25[285], stage0_25[286], stage0_25[287], stage0_25[288], stage0_25[289]},
      {stage0_27[228], stage0_27[229], stage0_27[230], stage0_27[231], stage0_27[232], stage0_27[233]},
      {stage1_29[38],stage1_28[111],stage1_27[115],stage1_26[132],stage1_25[211]}
   );
   gpc606_5 gpc1088 (
      {stage0_25[290], stage0_25[291], stage0_25[292], stage0_25[293], stage0_25[294], stage0_25[295]},
      {stage0_27[234], stage0_27[235], stage0_27[236], stage0_27[237], stage0_27[238], stage0_27[239]},
      {stage1_29[39],stage1_28[112],stage1_27[116],stage1_26[133],stage1_25[212]}
   );
   gpc606_5 gpc1089 (
      {stage0_25[296], stage0_25[297], stage0_25[298], stage0_25[299], stage0_25[300], stage0_25[301]},
      {stage0_27[240], stage0_27[241], stage0_27[242], stage0_27[243], stage0_27[244], stage0_27[245]},
      {stage1_29[40],stage1_28[113],stage1_27[117],stage1_26[134],stage1_25[213]}
   );
   gpc606_5 gpc1090 (
      {stage0_25[302], stage0_25[303], stage0_25[304], stage0_25[305], stage0_25[306], stage0_25[307]},
      {stage0_27[246], stage0_27[247], stage0_27[248], stage0_27[249], stage0_27[250], stage0_27[251]},
      {stage1_29[41],stage1_28[114],stage1_27[118],stage1_26[135],stage1_25[214]}
   );
   gpc606_5 gpc1091 (
      {stage0_25[308], stage0_25[309], stage0_25[310], stage0_25[311], stage0_25[312], stage0_25[313]},
      {stage0_27[252], stage0_27[253], stage0_27[254], stage0_27[255], stage0_27[256], stage0_27[257]},
      {stage1_29[42],stage1_28[115],stage1_27[119],stage1_26[136],stage1_25[215]}
   );
   gpc606_5 gpc1092 (
      {stage0_25[314], stage0_25[315], stage0_25[316], stage0_25[317], stage0_25[318], stage0_25[319]},
      {stage0_27[258], stage0_27[259], stage0_27[260], stage0_27[261], stage0_27[262], stage0_27[263]},
      {stage1_29[43],stage1_28[116],stage1_27[120],stage1_26[137],stage1_25[216]}
   );
   gpc606_5 gpc1093 (
      {stage0_25[320], stage0_25[321], stage0_25[322], stage0_25[323], stage0_25[324], stage0_25[325]},
      {stage0_27[264], stage0_27[265], stage0_27[266], stage0_27[267], stage0_27[268], stage0_27[269]},
      {stage1_29[44],stage1_28[117],stage1_27[121],stage1_26[138],stage1_25[217]}
   );
   gpc606_5 gpc1094 (
      {stage0_25[326], stage0_25[327], stage0_25[328], stage0_25[329], stage0_25[330], stage0_25[331]},
      {stage0_27[270], stage0_27[271], stage0_27[272], stage0_27[273], stage0_27[274], stage0_27[275]},
      {stage1_29[45],stage1_28[118],stage1_27[122],stage1_26[139],stage1_25[218]}
   );
   gpc606_5 gpc1095 (
      {stage0_25[332], stage0_25[333], stage0_25[334], stage0_25[335], stage0_25[336], stage0_25[337]},
      {stage0_27[276], stage0_27[277], stage0_27[278], stage0_27[279], stage0_27[280], stage0_27[281]},
      {stage1_29[46],stage1_28[119],stage1_27[123],stage1_26[140],stage1_25[219]}
   );
   gpc606_5 gpc1096 (
      {stage0_25[338], stage0_25[339], stage0_25[340], stage0_25[341], stage0_25[342], stage0_25[343]},
      {stage0_27[282], stage0_27[283], stage0_27[284], stage0_27[285], stage0_27[286], stage0_27[287]},
      {stage1_29[47],stage1_28[120],stage1_27[124],stage1_26[141],stage1_25[220]}
   );
   gpc606_5 gpc1097 (
      {stage0_25[344], stage0_25[345], stage0_25[346], stage0_25[347], stage0_25[348], stage0_25[349]},
      {stage0_27[288], stage0_27[289], stage0_27[290], stage0_27[291], stage0_27[292], stage0_27[293]},
      {stage1_29[48],stage1_28[121],stage1_27[125],stage1_26[142],stage1_25[221]}
   );
   gpc606_5 gpc1098 (
      {stage0_25[350], stage0_25[351], stage0_25[352], stage0_25[353], stage0_25[354], stage0_25[355]},
      {stage0_27[294], stage0_27[295], stage0_27[296], stage0_27[297], stage0_27[298], stage0_27[299]},
      {stage1_29[49],stage1_28[122],stage1_27[126],stage1_26[143],stage1_25[222]}
   );
   gpc606_5 gpc1099 (
      {stage0_25[356], stage0_25[357], stage0_25[358], stage0_25[359], stage0_25[360], stage0_25[361]},
      {stage0_27[300], stage0_27[301], stage0_27[302], stage0_27[303], stage0_27[304], stage0_27[305]},
      {stage1_29[50],stage1_28[123],stage1_27[127],stage1_26[144],stage1_25[223]}
   );
   gpc606_5 gpc1100 (
      {stage0_25[362], stage0_25[363], stage0_25[364], stage0_25[365], stage0_25[366], stage0_25[367]},
      {stage0_27[306], stage0_27[307], stage0_27[308], stage0_27[309], stage0_27[310], stage0_27[311]},
      {stage1_29[51],stage1_28[124],stage1_27[128],stage1_26[145],stage1_25[224]}
   );
   gpc606_5 gpc1101 (
      {stage0_25[368], stage0_25[369], stage0_25[370], stage0_25[371], stage0_25[372], stage0_25[373]},
      {stage0_27[312], stage0_27[313], stage0_27[314], stage0_27[315], stage0_27[316], stage0_27[317]},
      {stage1_29[52],stage1_28[125],stage1_27[129],stage1_26[146],stage1_25[225]}
   );
   gpc606_5 gpc1102 (
      {stage0_25[374], stage0_25[375], stage0_25[376], stage0_25[377], stage0_25[378], stage0_25[379]},
      {stage0_27[318], stage0_27[319], stage0_27[320], stage0_27[321], stage0_27[322], stage0_27[323]},
      {stage1_29[53],stage1_28[126],stage1_27[130],stage1_26[147],stage1_25[226]}
   );
   gpc606_5 gpc1103 (
      {stage0_25[380], stage0_25[381], stage0_25[382], stage0_25[383], stage0_25[384], stage0_25[385]},
      {stage0_27[324], stage0_27[325], stage0_27[326], stage0_27[327], stage0_27[328], stage0_27[329]},
      {stage1_29[54],stage1_28[127],stage1_27[131],stage1_26[148],stage1_25[227]}
   );
   gpc606_5 gpc1104 (
      {stage0_25[386], stage0_25[387], stage0_25[388], stage0_25[389], stage0_25[390], stage0_25[391]},
      {stage0_27[330], stage0_27[331], stage0_27[332], stage0_27[333], stage0_27[334], stage0_27[335]},
      {stage1_29[55],stage1_28[128],stage1_27[132],stage1_26[149],stage1_25[228]}
   );
   gpc606_5 gpc1105 (
      {stage0_25[392], stage0_25[393], stage0_25[394], stage0_25[395], stage0_25[396], stage0_25[397]},
      {stage0_27[336], stage0_27[337], stage0_27[338], stage0_27[339], stage0_27[340], stage0_27[341]},
      {stage1_29[56],stage1_28[129],stage1_27[133],stage1_26[150],stage1_25[229]}
   );
   gpc606_5 gpc1106 (
      {stage0_25[398], stage0_25[399], stage0_25[400], stage0_25[401], stage0_25[402], stage0_25[403]},
      {stage0_27[342], stage0_27[343], stage0_27[344], stage0_27[345], stage0_27[346], stage0_27[347]},
      {stage1_29[57],stage1_28[130],stage1_27[134],stage1_26[151],stage1_25[230]}
   );
   gpc606_5 gpc1107 (
      {stage0_25[404], stage0_25[405], stage0_25[406], stage0_25[407], stage0_25[408], stage0_25[409]},
      {stage0_27[348], stage0_27[349], stage0_27[350], stage0_27[351], stage0_27[352], stage0_27[353]},
      {stage1_29[58],stage1_28[131],stage1_27[135],stage1_26[152],stage1_25[231]}
   );
   gpc606_5 gpc1108 (
      {stage0_25[410], stage0_25[411], stage0_25[412], stage0_25[413], stage0_25[414], stage0_25[415]},
      {stage0_27[354], stage0_27[355], stage0_27[356], stage0_27[357], stage0_27[358], stage0_27[359]},
      {stage1_29[59],stage1_28[132],stage1_27[136],stage1_26[153],stage1_25[232]}
   );
   gpc606_5 gpc1109 (
      {stage0_25[416], stage0_25[417], stage0_25[418], stage0_25[419], stage0_25[420], stage0_25[421]},
      {stage0_27[360], stage0_27[361], stage0_27[362], stage0_27[363], stage0_27[364], stage0_27[365]},
      {stage1_29[60],stage1_28[133],stage1_27[137],stage1_26[154],stage1_25[233]}
   );
   gpc606_5 gpc1110 (
      {stage0_25[422], stage0_25[423], stage0_25[424], stage0_25[425], stage0_25[426], stage0_25[427]},
      {stage0_27[366], stage0_27[367], stage0_27[368], stage0_27[369], stage0_27[370], stage0_27[371]},
      {stage1_29[61],stage1_28[134],stage1_27[138],stage1_26[155],stage1_25[234]}
   );
   gpc606_5 gpc1111 (
      {stage0_25[428], stage0_25[429], stage0_25[430], stage0_25[431], stage0_25[432], stage0_25[433]},
      {stage0_27[372], stage0_27[373], stage0_27[374], stage0_27[375], stage0_27[376], stage0_27[377]},
      {stage1_29[62],stage1_28[135],stage1_27[139],stage1_26[156],stage1_25[235]}
   );
   gpc606_5 gpc1112 (
      {stage0_25[434], stage0_25[435], stage0_25[436], stage0_25[437], stage0_25[438], stage0_25[439]},
      {stage0_27[378], stage0_27[379], stage0_27[380], stage0_27[381], stage0_27[382], stage0_27[383]},
      {stage1_29[63],stage1_28[136],stage1_27[140],stage1_26[157],stage1_25[236]}
   );
   gpc606_5 gpc1113 (
      {stage0_25[440], stage0_25[441], stage0_25[442], stage0_25[443], stage0_25[444], stage0_25[445]},
      {stage0_27[384], stage0_27[385], stage0_27[386], stage0_27[387], stage0_27[388], stage0_27[389]},
      {stage1_29[64],stage1_28[137],stage1_27[141],stage1_26[158],stage1_25[237]}
   );
   gpc606_5 gpc1114 (
      {stage0_25[446], stage0_25[447], stage0_25[448], stage0_25[449], stage0_25[450], stage0_25[451]},
      {stage0_27[390], stage0_27[391], stage0_27[392], stage0_27[393], stage0_27[394], stage0_27[395]},
      {stage1_29[65],stage1_28[138],stage1_27[142],stage1_26[159],stage1_25[238]}
   );
   gpc606_5 gpc1115 (
      {stage0_25[452], stage0_25[453], stage0_25[454], stage0_25[455], stage0_25[456], stage0_25[457]},
      {stage0_27[396], stage0_27[397], stage0_27[398], stage0_27[399], stage0_27[400], stage0_27[401]},
      {stage1_29[66],stage1_28[139],stage1_27[143],stage1_26[160],stage1_25[239]}
   );
   gpc606_5 gpc1116 (
      {stage0_25[458], stage0_25[459], stage0_25[460], stage0_25[461], stage0_25[462], stage0_25[463]},
      {stage0_27[402], stage0_27[403], stage0_27[404], stage0_27[405], stage0_27[406], stage0_27[407]},
      {stage1_29[67],stage1_28[140],stage1_27[144],stage1_26[161],stage1_25[240]}
   );
   gpc606_5 gpc1117 (
      {stage0_25[464], stage0_25[465], stage0_25[466], stage0_25[467], stage0_25[468], stage0_25[469]},
      {stage0_27[408], stage0_27[409], stage0_27[410], stage0_27[411], stage0_27[412], stage0_27[413]},
      {stage1_29[68],stage1_28[141],stage1_27[145],stage1_26[162],stage1_25[241]}
   );
   gpc606_5 gpc1118 (
      {stage0_25[470], stage0_25[471], stage0_25[472], stage0_25[473], stage0_25[474], stage0_25[475]},
      {stage0_27[414], stage0_27[415], stage0_27[416], stage0_27[417], stage0_27[418], stage0_27[419]},
      {stage1_29[69],stage1_28[142],stage1_27[146],stage1_26[163],stage1_25[242]}
   );
   gpc606_5 gpc1119 (
      {stage0_25[476], stage0_25[477], stage0_25[478], stage0_25[479], stage0_25[480], stage0_25[481]},
      {stage0_27[420], stage0_27[421], stage0_27[422], stage0_27[423], stage0_27[424], stage0_27[425]},
      {stage1_29[70],stage1_28[143],stage1_27[147],stage1_26[164],stage1_25[243]}
   );
   gpc615_5 gpc1120 (
      {stage0_26[438], stage0_26[439], stage0_26[440], stage0_26[441], stage0_26[442]},
      {stage0_27[426]},
      {stage0_28[0], stage0_28[1], stage0_28[2], stage0_28[3], stage0_28[4], stage0_28[5]},
      {stage1_30[0],stage1_29[71],stage1_28[144],stage1_27[148],stage1_26[165]}
   );
   gpc615_5 gpc1121 (
      {stage0_26[443], stage0_26[444], stage0_26[445], stage0_26[446], stage0_26[447]},
      {stage0_27[427]},
      {stage0_28[6], stage0_28[7], stage0_28[8], stage0_28[9], stage0_28[10], stage0_28[11]},
      {stage1_30[1],stage1_29[72],stage1_28[145],stage1_27[149],stage1_26[166]}
   );
   gpc615_5 gpc1122 (
      {stage0_26[448], stage0_26[449], stage0_26[450], stage0_26[451], stage0_26[452]},
      {stage0_27[428]},
      {stage0_28[12], stage0_28[13], stage0_28[14], stage0_28[15], stage0_28[16], stage0_28[17]},
      {stage1_30[2],stage1_29[73],stage1_28[146],stage1_27[150],stage1_26[167]}
   );
   gpc615_5 gpc1123 (
      {stage0_26[453], stage0_26[454], stage0_26[455], stage0_26[456], stage0_26[457]},
      {stage0_27[429]},
      {stage0_28[18], stage0_28[19], stage0_28[20], stage0_28[21], stage0_28[22], stage0_28[23]},
      {stage1_30[3],stage1_29[74],stage1_28[147],stage1_27[151],stage1_26[168]}
   );
   gpc615_5 gpc1124 (
      {stage0_26[458], stage0_26[459], stage0_26[460], stage0_26[461], stage0_26[462]},
      {stage0_27[430]},
      {stage0_28[24], stage0_28[25], stage0_28[26], stage0_28[27], stage0_28[28], stage0_28[29]},
      {stage1_30[4],stage1_29[75],stage1_28[148],stage1_27[152],stage1_26[169]}
   );
   gpc615_5 gpc1125 (
      {stage0_26[463], stage0_26[464], stage0_26[465], stage0_26[466], stage0_26[467]},
      {stage0_27[431]},
      {stage0_28[30], stage0_28[31], stage0_28[32], stage0_28[33], stage0_28[34], stage0_28[35]},
      {stage1_30[5],stage1_29[76],stage1_28[149],stage1_27[153],stage1_26[170]}
   );
   gpc615_5 gpc1126 (
      {stage0_26[468], stage0_26[469], stage0_26[470], stage0_26[471], stage0_26[472]},
      {stage0_27[432]},
      {stage0_28[36], stage0_28[37], stage0_28[38], stage0_28[39], stage0_28[40], stage0_28[41]},
      {stage1_30[6],stage1_29[77],stage1_28[150],stage1_27[154],stage1_26[171]}
   );
   gpc615_5 gpc1127 (
      {stage0_26[473], stage0_26[474], stage0_26[475], stage0_26[476], stage0_26[477]},
      {stage0_27[433]},
      {stage0_28[42], stage0_28[43], stage0_28[44], stage0_28[45], stage0_28[46], stage0_28[47]},
      {stage1_30[7],stage1_29[78],stage1_28[151],stage1_27[155],stage1_26[172]}
   );
   gpc615_5 gpc1128 (
      {stage0_26[478], stage0_26[479], stage0_26[480], stage0_26[481], stage0_26[482]},
      {stage0_27[434]},
      {stage0_28[48], stage0_28[49], stage0_28[50], stage0_28[51], stage0_28[52], stage0_28[53]},
      {stage1_30[8],stage1_29[79],stage1_28[152],stage1_27[156],stage1_26[173]}
   );
   gpc615_5 gpc1129 (
      {stage0_26[483], stage0_26[484], stage0_26[485], stage0_26[486], stage0_26[487]},
      {stage0_27[435]},
      {stage0_28[54], stage0_28[55], stage0_28[56], stage0_28[57], stage0_28[58], stage0_28[59]},
      {stage1_30[9],stage1_29[80],stage1_28[153],stage1_27[157],stage1_26[174]}
   );
   gpc615_5 gpc1130 (
      {stage0_26[488], stage0_26[489], stage0_26[490], stage0_26[491], stage0_26[492]},
      {stage0_27[436]},
      {stage0_28[60], stage0_28[61], stage0_28[62], stage0_28[63], stage0_28[64], stage0_28[65]},
      {stage1_30[10],stage1_29[81],stage1_28[154],stage1_27[158],stage1_26[175]}
   );
   gpc615_5 gpc1131 (
      {stage0_26[493], stage0_26[494], stage0_26[495], stage0_26[496], stage0_26[497]},
      {stage0_27[437]},
      {stage0_28[66], stage0_28[67], stage0_28[68], stage0_28[69], stage0_28[70], stage0_28[71]},
      {stage1_30[11],stage1_29[82],stage1_28[155],stage1_27[159],stage1_26[176]}
   );
   gpc606_5 gpc1132 (
      {stage0_27[438], stage0_27[439], stage0_27[440], stage0_27[441], stage0_27[442], stage0_27[443]},
      {stage0_29[0], stage0_29[1], stage0_29[2], stage0_29[3], stage0_29[4], stage0_29[5]},
      {stage1_31[0],stage1_30[12],stage1_29[83],stage1_28[156],stage1_27[160]}
   );
   gpc606_5 gpc1133 (
      {stage0_27[444], stage0_27[445], stage0_27[446], stage0_27[447], stage0_27[448], stage0_27[449]},
      {stage0_29[6], stage0_29[7], stage0_29[8], stage0_29[9], stage0_29[10], stage0_29[11]},
      {stage1_31[1],stage1_30[13],stage1_29[84],stage1_28[157],stage1_27[161]}
   );
   gpc606_5 gpc1134 (
      {stage0_27[450], stage0_27[451], stage0_27[452], stage0_27[453], stage0_27[454], stage0_27[455]},
      {stage0_29[12], stage0_29[13], stage0_29[14], stage0_29[15], stage0_29[16], stage0_29[17]},
      {stage1_31[2],stage1_30[14],stage1_29[85],stage1_28[158],stage1_27[162]}
   );
   gpc606_5 gpc1135 (
      {stage0_27[456], stage0_27[457], stage0_27[458], stage0_27[459], stage0_27[460], stage0_27[461]},
      {stage0_29[18], stage0_29[19], stage0_29[20], stage0_29[21], stage0_29[22], stage0_29[23]},
      {stage1_31[3],stage1_30[15],stage1_29[86],stage1_28[159],stage1_27[163]}
   );
   gpc606_5 gpc1136 (
      {stage0_27[462], stage0_27[463], stage0_27[464], stage0_27[465], stage0_27[466], stage0_27[467]},
      {stage0_29[24], stage0_29[25], stage0_29[26], stage0_29[27], stage0_29[28], stage0_29[29]},
      {stage1_31[4],stage1_30[16],stage1_29[87],stage1_28[160],stage1_27[164]}
   );
   gpc606_5 gpc1137 (
      {stage0_27[468], stage0_27[469], stage0_27[470], stage0_27[471], stage0_27[472], stage0_27[473]},
      {stage0_29[30], stage0_29[31], stage0_29[32], stage0_29[33], stage0_29[34], stage0_29[35]},
      {stage1_31[5],stage1_30[17],stage1_29[88],stage1_28[161],stage1_27[165]}
   );
   gpc615_5 gpc1138 (
      {stage0_27[474], stage0_27[475], stage0_27[476], stage0_27[477], stage0_27[478]},
      {stage0_28[72]},
      {stage0_29[36], stage0_29[37], stage0_29[38], stage0_29[39], stage0_29[40], stage0_29[41]},
      {stage1_31[6],stage1_30[18],stage1_29[89],stage1_28[162],stage1_27[166]}
   );
   gpc606_5 gpc1139 (
      {stage0_28[73], stage0_28[74], stage0_28[75], stage0_28[76], stage0_28[77], stage0_28[78]},
      {stage0_30[0], stage0_30[1], stage0_30[2], stage0_30[3], stage0_30[4], stage0_30[5]},
      {stage1_32[0],stage1_31[7],stage1_30[19],stage1_29[90],stage1_28[163]}
   );
   gpc606_5 gpc1140 (
      {stage0_28[79], stage0_28[80], stage0_28[81], stage0_28[82], stage0_28[83], stage0_28[84]},
      {stage0_30[6], stage0_30[7], stage0_30[8], stage0_30[9], stage0_30[10], stage0_30[11]},
      {stage1_32[1],stage1_31[8],stage1_30[20],stage1_29[91],stage1_28[164]}
   );
   gpc606_5 gpc1141 (
      {stage0_28[85], stage0_28[86], stage0_28[87], stage0_28[88], stage0_28[89], stage0_28[90]},
      {stage0_30[12], stage0_30[13], stage0_30[14], stage0_30[15], stage0_30[16], stage0_30[17]},
      {stage1_32[2],stage1_31[9],stage1_30[21],stage1_29[92],stage1_28[165]}
   );
   gpc606_5 gpc1142 (
      {stage0_28[91], stage0_28[92], stage0_28[93], stage0_28[94], stage0_28[95], stage0_28[96]},
      {stage0_30[18], stage0_30[19], stage0_30[20], stage0_30[21], stage0_30[22], stage0_30[23]},
      {stage1_32[3],stage1_31[10],stage1_30[22],stage1_29[93],stage1_28[166]}
   );
   gpc606_5 gpc1143 (
      {stage0_28[97], stage0_28[98], stage0_28[99], stage0_28[100], stage0_28[101], stage0_28[102]},
      {stage0_30[24], stage0_30[25], stage0_30[26], stage0_30[27], stage0_30[28], stage0_30[29]},
      {stage1_32[4],stage1_31[11],stage1_30[23],stage1_29[94],stage1_28[167]}
   );
   gpc606_5 gpc1144 (
      {stage0_28[103], stage0_28[104], stage0_28[105], stage0_28[106], stage0_28[107], stage0_28[108]},
      {stage0_30[30], stage0_30[31], stage0_30[32], stage0_30[33], stage0_30[34], stage0_30[35]},
      {stage1_32[5],stage1_31[12],stage1_30[24],stage1_29[95],stage1_28[168]}
   );
   gpc606_5 gpc1145 (
      {stage0_28[109], stage0_28[110], stage0_28[111], stage0_28[112], stage0_28[113], stage0_28[114]},
      {stage0_30[36], stage0_30[37], stage0_30[38], stage0_30[39], stage0_30[40], stage0_30[41]},
      {stage1_32[6],stage1_31[13],stage1_30[25],stage1_29[96],stage1_28[169]}
   );
   gpc606_5 gpc1146 (
      {stage0_28[115], stage0_28[116], stage0_28[117], stage0_28[118], stage0_28[119], stage0_28[120]},
      {stage0_30[42], stage0_30[43], stage0_30[44], stage0_30[45], stage0_30[46], stage0_30[47]},
      {stage1_32[7],stage1_31[14],stage1_30[26],stage1_29[97],stage1_28[170]}
   );
   gpc606_5 gpc1147 (
      {stage0_28[121], stage0_28[122], stage0_28[123], stage0_28[124], stage0_28[125], stage0_28[126]},
      {stage0_30[48], stage0_30[49], stage0_30[50], stage0_30[51], stage0_30[52], stage0_30[53]},
      {stage1_32[8],stage1_31[15],stage1_30[27],stage1_29[98],stage1_28[171]}
   );
   gpc606_5 gpc1148 (
      {stage0_28[127], stage0_28[128], stage0_28[129], stage0_28[130], stage0_28[131], stage0_28[132]},
      {stage0_30[54], stage0_30[55], stage0_30[56], stage0_30[57], stage0_30[58], stage0_30[59]},
      {stage1_32[9],stage1_31[16],stage1_30[28],stage1_29[99],stage1_28[172]}
   );
   gpc606_5 gpc1149 (
      {stage0_28[133], stage0_28[134], stage0_28[135], stage0_28[136], stage0_28[137], stage0_28[138]},
      {stage0_30[60], stage0_30[61], stage0_30[62], stage0_30[63], stage0_30[64], stage0_30[65]},
      {stage1_32[10],stage1_31[17],stage1_30[29],stage1_29[100],stage1_28[173]}
   );
   gpc606_5 gpc1150 (
      {stage0_28[139], stage0_28[140], stage0_28[141], stage0_28[142], stage0_28[143], stage0_28[144]},
      {stage0_30[66], stage0_30[67], stage0_30[68], stage0_30[69], stage0_30[70], stage0_30[71]},
      {stage1_32[11],stage1_31[18],stage1_30[30],stage1_29[101],stage1_28[174]}
   );
   gpc606_5 gpc1151 (
      {stage0_28[145], stage0_28[146], stage0_28[147], stage0_28[148], stage0_28[149], stage0_28[150]},
      {stage0_30[72], stage0_30[73], stage0_30[74], stage0_30[75], stage0_30[76], stage0_30[77]},
      {stage1_32[12],stage1_31[19],stage1_30[31],stage1_29[102],stage1_28[175]}
   );
   gpc606_5 gpc1152 (
      {stage0_28[151], stage0_28[152], stage0_28[153], stage0_28[154], stage0_28[155], stage0_28[156]},
      {stage0_30[78], stage0_30[79], stage0_30[80], stage0_30[81], stage0_30[82], stage0_30[83]},
      {stage1_32[13],stage1_31[20],stage1_30[32],stage1_29[103],stage1_28[176]}
   );
   gpc606_5 gpc1153 (
      {stage0_28[157], stage0_28[158], stage0_28[159], stage0_28[160], stage0_28[161], stage0_28[162]},
      {stage0_30[84], stage0_30[85], stage0_30[86], stage0_30[87], stage0_30[88], stage0_30[89]},
      {stage1_32[14],stage1_31[21],stage1_30[33],stage1_29[104],stage1_28[177]}
   );
   gpc606_5 gpc1154 (
      {stage0_28[163], stage0_28[164], stage0_28[165], stage0_28[166], stage0_28[167], stage0_28[168]},
      {stage0_30[90], stage0_30[91], stage0_30[92], stage0_30[93], stage0_30[94], stage0_30[95]},
      {stage1_32[15],stage1_31[22],stage1_30[34],stage1_29[105],stage1_28[178]}
   );
   gpc606_5 gpc1155 (
      {stage0_28[169], stage0_28[170], stage0_28[171], stage0_28[172], stage0_28[173], stage0_28[174]},
      {stage0_30[96], stage0_30[97], stage0_30[98], stage0_30[99], stage0_30[100], stage0_30[101]},
      {stage1_32[16],stage1_31[23],stage1_30[35],stage1_29[106],stage1_28[179]}
   );
   gpc606_5 gpc1156 (
      {stage0_28[175], stage0_28[176], stage0_28[177], stage0_28[178], stage0_28[179], stage0_28[180]},
      {stage0_30[102], stage0_30[103], stage0_30[104], stage0_30[105], stage0_30[106], stage0_30[107]},
      {stage1_32[17],stage1_31[24],stage1_30[36],stage1_29[107],stage1_28[180]}
   );
   gpc606_5 gpc1157 (
      {stage0_28[181], stage0_28[182], stage0_28[183], stage0_28[184], stage0_28[185], stage0_28[186]},
      {stage0_30[108], stage0_30[109], stage0_30[110], stage0_30[111], stage0_30[112], stage0_30[113]},
      {stage1_32[18],stage1_31[25],stage1_30[37],stage1_29[108],stage1_28[181]}
   );
   gpc606_5 gpc1158 (
      {stage0_28[187], stage0_28[188], stage0_28[189], stage0_28[190], stage0_28[191], stage0_28[192]},
      {stage0_30[114], stage0_30[115], stage0_30[116], stage0_30[117], stage0_30[118], stage0_30[119]},
      {stage1_32[19],stage1_31[26],stage1_30[38],stage1_29[109],stage1_28[182]}
   );
   gpc606_5 gpc1159 (
      {stage0_28[193], stage0_28[194], stage0_28[195], stage0_28[196], stage0_28[197], stage0_28[198]},
      {stage0_30[120], stage0_30[121], stage0_30[122], stage0_30[123], stage0_30[124], stage0_30[125]},
      {stage1_32[20],stage1_31[27],stage1_30[39],stage1_29[110],stage1_28[183]}
   );
   gpc606_5 gpc1160 (
      {stage0_28[199], stage0_28[200], stage0_28[201], stage0_28[202], stage0_28[203], stage0_28[204]},
      {stage0_30[126], stage0_30[127], stage0_30[128], stage0_30[129], stage0_30[130], stage0_30[131]},
      {stage1_32[21],stage1_31[28],stage1_30[40],stage1_29[111],stage1_28[184]}
   );
   gpc606_5 gpc1161 (
      {stage0_28[205], stage0_28[206], stage0_28[207], stage0_28[208], stage0_28[209], stage0_28[210]},
      {stage0_30[132], stage0_30[133], stage0_30[134], stage0_30[135], stage0_30[136], stage0_30[137]},
      {stage1_32[22],stage1_31[29],stage1_30[41],stage1_29[112],stage1_28[185]}
   );
   gpc606_5 gpc1162 (
      {stage0_28[211], stage0_28[212], stage0_28[213], stage0_28[214], stage0_28[215], stage0_28[216]},
      {stage0_30[138], stage0_30[139], stage0_30[140], stage0_30[141], stage0_30[142], stage0_30[143]},
      {stage1_32[23],stage1_31[30],stage1_30[42],stage1_29[113],stage1_28[186]}
   );
   gpc606_5 gpc1163 (
      {stage0_28[217], stage0_28[218], stage0_28[219], stage0_28[220], stage0_28[221], stage0_28[222]},
      {stage0_30[144], stage0_30[145], stage0_30[146], stage0_30[147], stage0_30[148], stage0_30[149]},
      {stage1_32[24],stage1_31[31],stage1_30[43],stage1_29[114],stage1_28[187]}
   );
   gpc606_5 gpc1164 (
      {stage0_28[223], stage0_28[224], stage0_28[225], stage0_28[226], stage0_28[227], stage0_28[228]},
      {stage0_30[150], stage0_30[151], stage0_30[152], stage0_30[153], stage0_30[154], stage0_30[155]},
      {stage1_32[25],stage1_31[32],stage1_30[44],stage1_29[115],stage1_28[188]}
   );
   gpc606_5 gpc1165 (
      {stage0_28[229], stage0_28[230], stage0_28[231], stage0_28[232], stage0_28[233], stage0_28[234]},
      {stage0_30[156], stage0_30[157], stage0_30[158], stage0_30[159], stage0_30[160], stage0_30[161]},
      {stage1_32[26],stage1_31[33],stage1_30[45],stage1_29[116],stage1_28[189]}
   );
   gpc606_5 gpc1166 (
      {stage0_28[235], stage0_28[236], stage0_28[237], stage0_28[238], stage0_28[239], stage0_28[240]},
      {stage0_30[162], stage0_30[163], stage0_30[164], stage0_30[165], stage0_30[166], stage0_30[167]},
      {stage1_32[27],stage1_31[34],stage1_30[46],stage1_29[117],stage1_28[190]}
   );
   gpc606_5 gpc1167 (
      {stage0_28[241], stage0_28[242], stage0_28[243], stage0_28[244], stage0_28[245], stage0_28[246]},
      {stage0_30[168], stage0_30[169], stage0_30[170], stage0_30[171], stage0_30[172], stage0_30[173]},
      {stage1_32[28],stage1_31[35],stage1_30[47],stage1_29[118],stage1_28[191]}
   );
   gpc606_5 gpc1168 (
      {stage0_28[247], stage0_28[248], stage0_28[249], stage0_28[250], stage0_28[251], stage0_28[252]},
      {stage0_30[174], stage0_30[175], stage0_30[176], stage0_30[177], stage0_30[178], stage0_30[179]},
      {stage1_32[29],stage1_31[36],stage1_30[48],stage1_29[119],stage1_28[192]}
   );
   gpc606_5 gpc1169 (
      {stage0_28[253], stage0_28[254], stage0_28[255], stage0_28[256], stage0_28[257], stage0_28[258]},
      {stage0_30[180], stage0_30[181], stage0_30[182], stage0_30[183], stage0_30[184], stage0_30[185]},
      {stage1_32[30],stage1_31[37],stage1_30[49],stage1_29[120],stage1_28[193]}
   );
   gpc606_5 gpc1170 (
      {stage0_28[259], stage0_28[260], stage0_28[261], stage0_28[262], stage0_28[263], stage0_28[264]},
      {stage0_30[186], stage0_30[187], stage0_30[188], stage0_30[189], stage0_30[190], stage0_30[191]},
      {stage1_32[31],stage1_31[38],stage1_30[50],stage1_29[121],stage1_28[194]}
   );
   gpc606_5 gpc1171 (
      {stage0_28[265], stage0_28[266], stage0_28[267], stage0_28[268], stage0_28[269], stage0_28[270]},
      {stage0_30[192], stage0_30[193], stage0_30[194], stage0_30[195], stage0_30[196], stage0_30[197]},
      {stage1_32[32],stage1_31[39],stage1_30[51],stage1_29[122],stage1_28[195]}
   );
   gpc606_5 gpc1172 (
      {stage0_28[271], stage0_28[272], stage0_28[273], stage0_28[274], stage0_28[275], stage0_28[276]},
      {stage0_30[198], stage0_30[199], stage0_30[200], stage0_30[201], stage0_30[202], stage0_30[203]},
      {stage1_32[33],stage1_31[40],stage1_30[52],stage1_29[123],stage1_28[196]}
   );
   gpc606_5 gpc1173 (
      {stage0_28[277], stage0_28[278], stage0_28[279], stage0_28[280], stage0_28[281], stage0_28[282]},
      {stage0_30[204], stage0_30[205], stage0_30[206], stage0_30[207], stage0_30[208], stage0_30[209]},
      {stage1_32[34],stage1_31[41],stage1_30[53],stage1_29[124],stage1_28[197]}
   );
   gpc606_5 gpc1174 (
      {stage0_28[283], stage0_28[284], stage0_28[285], stage0_28[286], stage0_28[287], stage0_28[288]},
      {stage0_30[210], stage0_30[211], stage0_30[212], stage0_30[213], stage0_30[214], stage0_30[215]},
      {stage1_32[35],stage1_31[42],stage1_30[54],stage1_29[125],stage1_28[198]}
   );
   gpc606_5 gpc1175 (
      {stage0_28[289], stage0_28[290], stage0_28[291], stage0_28[292], stage0_28[293], stage0_28[294]},
      {stage0_30[216], stage0_30[217], stage0_30[218], stage0_30[219], stage0_30[220], stage0_30[221]},
      {stage1_32[36],stage1_31[43],stage1_30[55],stage1_29[126],stage1_28[199]}
   );
   gpc606_5 gpc1176 (
      {stage0_28[295], stage0_28[296], stage0_28[297], stage0_28[298], stage0_28[299], stage0_28[300]},
      {stage0_30[222], stage0_30[223], stage0_30[224], stage0_30[225], stage0_30[226], stage0_30[227]},
      {stage1_32[37],stage1_31[44],stage1_30[56],stage1_29[127],stage1_28[200]}
   );
   gpc615_5 gpc1177 (
      {stage0_28[301], stage0_28[302], stage0_28[303], stage0_28[304], stage0_28[305]},
      {stage0_29[42]},
      {stage0_30[228], stage0_30[229], stage0_30[230], stage0_30[231], stage0_30[232], stage0_30[233]},
      {stage1_32[38],stage1_31[45],stage1_30[57],stage1_29[128],stage1_28[201]}
   );
   gpc615_5 gpc1178 (
      {stage0_28[306], stage0_28[307], stage0_28[308], stage0_28[309], stage0_28[310]},
      {stage0_29[43]},
      {stage0_30[234], stage0_30[235], stage0_30[236], stage0_30[237], stage0_30[238], stage0_30[239]},
      {stage1_32[39],stage1_31[46],stage1_30[58],stage1_29[129],stage1_28[202]}
   );
   gpc615_5 gpc1179 (
      {stage0_28[311], stage0_28[312], stage0_28[313], stage0_28[314], stage0_28[315]},
      {stage0_29[44]},
      {stage0_30[240], stage0_30[241], stage0_30[242], stage0_30[243], stage0_30[244], stage0_30[245]},
      {stage1_32[40],stage1_31[47],stage1_30[59],stage1_29[130],stage1_28[203]}
   );
   gpc615_5 gpc1180 (
      {stage0_28[316], stage0_28[317], stage0_28[318], stage0_28[319], stage0_28[320]},
      {stage0_29[45]},
      {stage0_30[246], stage0_30[247], stage0_30[248], stage0_30[249], stage0_30[250], stage0_30[251]},
      {stage1_32[41],stage1_31[48],stage1_30[60],stage1_29[131],stage1_28[204]}
   );
   gpc615_5 gpc1181 (
      {stage0_28[321], stage0_28[322], stage0_28[323], stage0_28[324], stage0_28[325]},
      {stage0_29[46]},
      {stage0_30[252], stage0_30[253], stage0_30[254], stage0_30[255], stage0_30[256], stage0_30[257]},
      {stage1_32[42],stage1_31[49],stage1_30[61],stage1_29[132],stage1_28[205]}
   );
   gpc615_5 gpc1182 (
      {stage0_28[326], stage0_28[327], stage0_28[328], stage0_28[329], stage0_28[330]},
      {stage0_29[47]},
      {stage0_30[258], stage0_30[259], stage0_30[260], stage0_30[261], stage0_30[262], stage0_30[263]},
      {stage1_32[43],stage1_31[50],stage1_30[62],stage1_29[133],stage1_28[206]}
   );
   gpc615_5 gpc1183 (
      {stage0_28[331], stage0_28[332], stage0_28[333], stage0_28[334], stage0_28[335]},
      {stage0_29[48]},
      {stage0_30[264], stage0_30[265], stage0_30[266], stage0_30[267], stage0_30[268], stage0_30[269]},
      {stage1_32[44],stage1_31[51],stage1_30[63],stage1_29[134],stage1_28[207]}
   );
   gpc615_5 gpc1184 (
      {stage0_28[336], stage0_28[337], stage0_28[338], stage0_28[339], stage0_28[340]},
      {stage0_29[49]},
      {stage0_30[270], stage0_30[271], stage0_30[272], stage0_30[273], stage0_30[274], stage0_30[275]},
      {stage1_32[45],stage1_31[52],stage1_30[64],stage1_29[135],stage1_28[208]}
   );
   gpc615_5 gpc1185 (
      {stage0_28[341], stage0_28[342], stage0_28[343], stage0_28[344], stage0_28[345]},
      {stage0_29[50]},
      {stage0_30[276], stage0_30[277], stage0_30[278], stage0_30[279], stage0_30[280], stage0_30[281]},
      {stage1_32[46],stage1_31[53],stage1_30[65],stage1_29[136],stage1_28[209]}
   );
   gpc615_5 gpc1186 (
      {stage0_28[346], stage0_28[347], stage0_28[348], stage0_28[349], stage0_28[350]},
      {stage0_29[51]},
      {stage0_30[282], stage0_30[283], stage0_30[284], stage0_30[285], stage0_30[286], stage0_30[287]},
      {stage1_32[47],stage1_31[54],stage1_30[66],stage1_29[137],stage1_28[210]}
   );
   gpc615_5 gpc1187 (
      {stage0_28[351], stage0_28[352], stage0_28[353], stage0_28[354], stage0_28[355]},
      {stage0_29[52]},
      {stage0_30[288], stage0_30[289], stage0_30[290], stage0_30[291], stage0_30[292], stage0_30[293]},
      {stage1_32[48],stage1_31[55],stage1_30[67],stage1_29[138],stage1_28[211]}
   );
   gpc615_5 gpc1188 (
      {stage0_28[356], stage0_28[357], stage0_28[358], stage0_28[359], stage0_28[360]},
      {stage0_29[53]},
      {stage0_30[294], stage0_30[295], stage0_30[296], stage0_30[297], stage0_30[298], stage0_30[299]},
      {stage1_32[49],stage1_31[56],stage1_30[68],stage1_29[139],stage1_28[212]}
   );
   gpc615_5 gpc1189 (
      {stage0_28[361], stage0_28[362], stage0_28[363], stage0_28[364], stage0_28[365]},
      {stage0_29[54]},
      {stage0_30[300], stage0_30[301], stage0_30[302], stage0_30[303], stage0_30[304], stage0_30[305]},
      {stage1_32[50],stage1_31[57],stage1_30[69],stage1_29[140],stage1_28[213]}
   );
   gpc615_5 gpc1190 (
      {stage0_28[366], stage0_28[367], stage0_28[368], stage0_28[369], stage0_28[370]},
      {stage0_29[55]},
      {stage0_30[306], stage0_30[307], stage0_30[308], stage0_30[309], stage0_30[310], stage0_30[311]},
      {stage1_32[51],stage1_31[58],stage1_30[70],stage1_29[141],stage1_28[214]}
   );
   gpc615_5 gpc1191 (
      {stage0_28[371], stage0_28[372], stage0_28[373], stage0_28[374], stage0_28[375]},
      {stage0_29[56]},
      {stage0_30[312], stage0_30[313], stage0_30[314], stage0_30[315], stage0_30[316], stage0_30[317]},
      {stage1_32[52],stage1_31[59],stage1_30[71],stage1_29[142],stage1_28[215]}
   );
   gpc615_5 gpc1192 (
      {stage0_28[376], stage0_28[377], stage0_28[378], stage0_28[379], stage0_28[380]},
      {stage0_29[57]},
      {stage0_30[318], stage0_30[319], stage0_30[320], stage0_30[321], stage0_30[322], stage0_30[323]},
      {stage1_32[53],stage1_31[60],stage1_30[72],stage1_29[143],stage1_28[216]}
   );
   gpc615_5 gpc1193 (
      {stage0_28[381], stage0_28[382], stage0_28[383], stage0_28[384], stage0_28[385]},
      {stage0_29[58]},
      {stage0_30[324], stage0_30[325], stage0_30[326], stage0_30[327], stage0_30[328], stage0_30[329]},
      {stage1_32[54],stage1_31[61],stage1_30[73],stage1_29[144],stage1_28[217]}
   );
   gpc615_5 gpc1194 (
      {stage0_28[386], stage0_28[387], stage0_28[388], stage0_28[389], stage0_28[390]},
      {stage0_29[59]},
      {stage0_30[330], stage0_30[331], stage0_30[332], stage0_30[333], stage0_30[334], stage0_30[335]},
      {stage1_32[55],stage1_31[62],stage1_30[74],stage1_29[145],stage1_28[218]}
   );
   gpc615_5 gpc1195 (
      {stage0_28[391], stage0_28[392], stage0_28[393], stage0_28[394], stage0_28[395]},
      {stage0_29[60]},
      {stage0_30[336], stage0_30[337], stage0_30[338], stage0_30[339], stage0_30[340], stage0_30[341]},
      {stage1_32[56],stage1_31[63],stage1_30[75],stage1_29[146],stage1_28[219]}
   );
   gpc615_5 gpc1196 (
      {stage0_28[396], stage0_28[397], stage0_28[398], stage0_28[399], stage0_28[400]},
      {stage0_29[61]},
      {stage0_30[342], stage0_30[343], stage0_30[344], stage0_30[345], stage0_30[346], stage0_30[347]},
      {stage1_32[57],stage1_31[64],stage1_30[76],stage1_29[147],stage1_28[220]}
   );
   gpc615_5 gpc1197 (
      {stage0_28[401], stage0_28[402], stage0_28[403], stage0_28[404], stage0_28[405]},
      {stage0_29[62]},
      {stage0_30[348], stage0_30[349], stage0_30[350], stage0_30[351], stage0_30[352], stage0_30[353]},
      {stage1_32[58],stage1_31[65],stage1_30[77],stage1_29[148],stage1_28[221]}
   );
   gpc615_5 gpc1198 (
      {stage0_28[406], stage0_28[407], stage0_28[408], stage0_28[409], stage0_28[410]},
      {stage0_29[63]},
      {stage0_30[354], stage0_30[355], stage0_30[356], stage0_30[357], stage0_30[358], stage0_30[359]},
      {stage1_32[59],stage1_31[66],stage1_30[78],stage1_29[149],stage1_28[222]}
   );
   gpc615_5 gpc1199 (
      {stage0_28[411], stage0_28[412], stage0_28[413], stage0_28[414], stage0_28[415]},
      {stage0_29[64]},
      {stage0_30[360], stage0_30[361], stage0_30[362], stage0_30[363], stage0_30[364], stage0_30[365]},
      {stage1_32[60],stage1_31[67],stage1_30[79],stage1_29[150],stage1_28[223]}
   );
   gpc615_5 gpc1200 (
      {stage0_28[416], stage0_28[417], stage0_28[418], stage0_28[419], stage0_28[420]},
      {stage0_29[65]},
      {stage0_30[366], stage0_30[367], stage0_30[368], stage0_30[369], stage0_30[370], stage0_30[371]},
      {stage1_32[61],stage1_31[68],stage1_30[80],stage1_29[151],stage1_28[224]}
   );
   gpc615_5 gpc1201 (
      {stage0_28[421], stage0_28[422], stage0_28[423], stage0_28[424], stage0_28[425]},
      {stage0_29[66]},
      {stage0_30[372], stage0_30[373], stage0_30[374], stage0_30[375], stage0_30[376], stage0_30[377]},
      {stage1_32[62],stage1_31[69],stage1_30[81],stage1_29[152],stage1_28[225]}
   );
   gpc615_5 gpc1202 (
      {stage0_28[426], stage0_28[427], stage0_28[428], stage0_28[429], stage0_28[430]},
      {stage0_29[67]},
      {stage0_30[378], stage0_30[379], stage0_30[380], stage0_30[381], stage0_30[382], stage0_30[383]},
      {stage1_32[63],stage1_31[70],stage1_30[82],stage1_29[153],stage1_28[226]}
   );
   gpc615_5 gpc1203 (
      {stage0_28[431], stage0_28[432], stage0_28[433], stage0_28[434], stage0_28[435]},
      {stage0_29[68]},
      {stage0_30[384], stage0_30[385], stage0_30[386], stage0_30[387], stage0_30[388], stage0_30[389]},
      {stage1_32[64],stage1_31[71],stage1_30[83],stage1_29[154],stage1_28[227]}
   );
   gpc615_5 gpc1204 (
      {stage0_28[436], stage0_28[437], stage0_28[438], stage0_28[439], stage0_28[440]},
      {stage0_29[69]},
      {stage0_30[390], stage0_30[391], stage0_30[392], stage0_30[393], stage0_30[394], stage0_30[395]},
      {stage1_32[65],stage1_31[72],stage1_30[84],stage1_29[155],stage1_28[228]}
   );
   gpc615_5 gpc1205 (
      {stage0_28[441], stage0_28[442], stage0_28[443], stage0_28[444], stage0_28[445]},
      {stage0_29[70]},
      {stage0_30[396], stage0_30[397], stage0_30[398], stage0_30[399], stage0_30[400], stage0_30[401]},
      {stage1_32[66],stage1_31[73],stage1_30[85],stage1_29[156],stage1_28[229]}
   );
   gpc615_5 gpc1206 (
      {stage0_28[446], stage0_28[447], stage0_28[448], stage0_28[449], stage0_28[450]},
      {stage0_29[71]},
      {stage0_30[402], stage0_30[403], stage0_30[404], stage0_30[405], stage0_30[406], stage0_30[407]},
      {stage1_32[67],stage1_31[74],stage1_30[86],stage1_29[157],stage1_28[230]}
   );
   gpc615_5 gpc1207 (
      {stage0_28[451], stage0_28[452], stage0_28[453], stage0_28[454], stage0_28[455]},
      {stage0_29[72]},
      {stage0_30[408], stage0_30[409], stage0_30[410], stage0_30[411], stage0_30[412], stage0_30[413]},
      {stage1_32[68],stage1_31[75],stage1_30[87],stage1_29[158],stage1_28[231]}
   );
   gpc615_5 gpc1208 (
      {stage0_28[456], stage0_28[457], stage0_28[458], stage0_28[459], stage0_28[460]},
      {stage0_29[73]},
      {stage0_30[414], stage0_30[415], stage0_30[416], stage0_30[417], stage0_30[418], stage0_30[419]},
      {stage1_32[69],stage1_31[76],stage1_30[88],stage1_29[159],stage1_28[232]}
   );
   gpc615_5 gpc1209 (
      {stage0_28[461], stage0_28[462], stage0_28[463], stage0_28[464], stage0_28[465]},
      {stage0_29[74]},
      {stage0_30[420], stage0_30[421], stage0_30[422], stage0_30[423], stage0_30[424], stage0_30[425]},
      {stage1_32[70],stage1_31[77],stage1_30[89],stage1_29[160],stage1_28[233]}
   );
   gpc615_5 gpc1210 (
      {stage0_28[466], stage0_28[467], stage0_28[468], stage0_28[469], stage0_28[470]},
      {stage0_29[75]},
      {stage0_30[426], stage0_30[427], stage0_30[428], stage0_30[429], stage0_30[430], stage0_30[431]},
      {stage1_32[71],stage1_31[78],stage1_30[90],stage1_29[161],stage1_28[234]}
   );
   gpc615_5 gpc1211 (
      {stage0_28[471], stage0_28[472], stage0_28[473], stage0_28[474], stage0_28[475]},
      {stage0_29[76]},
      {stage0_30[432], stage0_30[433], stage0_30[434], stage0_30[435], stage0_30[436], stage0_30[437]},
      {stage1_32[72],stage1_31[79],stage1_30[91],stage1_29[162],stage1_28[235]}
   );
   gpc615_5 gpc1212 (
      {stage0_28[476], stage0_28[477], stage0_28[478], stage0_28[479], stage0_28[480]},
      {stage0_29[77]},
      {stage0_30[438], stage0_30[439], stage0_30[440], stage0_30[441], stage0_30[442], stage0_30[443]},
      {stage1_32[73],stage1_31[80],stage1_30[92],stage1_29[163],stage1_28[236]}
   );
   gpc615_5 gpc1213 (
      {stage0_28[481], stage0_28[482], stage0_28[483], stage0_28[484], stage0_28[485]},
      {stage0_29[78]},
      {stage0_30[444], stage0_30[445], stage0_30[446], stage0_30[447], stage0_30[448], stage0_30[449]},
      {stage1_32[74],stage1_31[81],stage1_30[93],stage1_29[164],stage1_28[237]}
   );
   gpc615_5 gpc1214 (
      {stage0_28[486], stage0_28[487], stage0_28[488], stage0_28[489], stage0_28[490]},
      {stage0_29[79]},
      {stage0_30[450], stage0_30[451], stage0_30[452], stage0_30[453], stage0_30[454], stage0_30[455]},
      {stage1_32[75],stage1_31[82],stage1_30[94],stage1_29[165],stage1_28[238]}
   );
   gpc615_5 gpc1215 (
      {stage0_28[491], stage0_28[492], stage0_28[493], stage0_28[494], stage0_28[495]},
      {stage0_29[80]},
      {stage0_30[456], stage0_30[457], stage0_30[458], stage0_30[459], stage0_30[460], stage0_30[461]},
      {stage1_32[76],stage1_31[83],stage1_30[95],stage1_29[166],stage1_28[239]}
   );
   gpc615_5 gpc1216 (
      {stage0_28[496], stage0_28[497], stage0_28[498], stage0_28[499], stage0_28[500]},
      {stage0_29[81]},
      {stage0_30[462], stage0_30[463], stage0_30[464], stage0_30[465], stage0_30[466], stage0_30[467]},
      {stage1_32[77],stage1_31[84],stage1_30[96],stage1_29[167],stage1_28[240]}
   );
   gpc615_5 gpc1217 (
      {stage0_28[501], stage0_28[502], stage0_28[503], stage0_28[504], stage0_28[505]},
      {stage0_29[82]},
      {stage0_30[468], stage0_30[469], stage0_30[470], stage0_30[471], stage0_30[472], stage0_30[473]},
      {stage1_32[78],stage1_31[85],stage1_30[97],stage1_29[168],stage1_28[241]}
   );
   gpc606_5 gpc1218 (
      {stage0_29[83], stage0_29[84], stage0_29[85], stage0_29[86], stage0_29[87], stage0_29[88]},
      {stage0_31[0], stage0_31[1], stage0_31[2], stage0_31[3], stage0_31[4], stage0_31[5]},
      {stage1_33[0],stage1_32[79],stage1_31[86],stage1_30[98],stage1_29[169]}
   );
   gpc606_5 gpc1219 (
      {stage0_29[89], stage0_29[90], stage0_29[91], stage0_29[92], stage0_29[93], stage0_29[94]},
      {stage0_31[6], stage0_31[7], stage0_31[8], stage0_31[9], stage0_31[10], stage0_31[11]},
      {stage1_33[1],stage1_32[80],stage1_31[87],stage1_30[99],stage1_29[170]}
   );
   gpc606_5 gpc1220 (
      {stage0_29[95], stage0_29[96], stage0_29[97], stage0_29[98], stage0_29[99], stage0_29[100]},
      {stage0_31[12], stage0_31[13], stage0_31[14], stage0_31[15], stage0_31[16], stage0_31[17]},
      {stage1_33[2],stage1_32[81],stage1_31[88],stage1_30[100],stage1_29[171]}
   );
   gpc606_5 gpc1221 (
      {stage0_29[101], stage0_29[102], stage0_29[103], stage0_29[104], stage0_29[105], stage0_29[106]},
      {stage0_31[18], stage0_31[19], stage0_31[20], stage0_31[21], stage0_31[22], stage0_31[23]},
      {stage1_33[3],stage1_32[82],stage1_31[89],stage1_30[101],stage1_29[172]}
   );
   gpc606_5 gpc1222 (
      {stage0_29[107], stage0_29[108], stage0_29[109], stage0_29[110], stage0_29[111], stage0_29[112]},
      {stage0_31[24], stage0_31[25], stage0_31[26], stage0_31[27], stage0_31[28], stage0_31[29]},
      {stage1_33[4],stage1_32[83],stage1_31[90],stage1_30[102],stage1_29[173]}
   );
   gpc606_5 gpc1223 (
      {stage0_29[113], stage0_29[114], stage0_29[115], stage0_29[116], stage0_29[117], stage0_29[118]},
      {stage0_31[30], stage0_31[31], stage0_31[32], stage0_31[33], stage0_31[34], stage0_31[35]},
      {stage1_33[5],stage1_32[84],stage1_31[91],stage1_30[103],stage1_29[174]}
   );
   gpc606_5 gpc1224 (
      {stage0_29[119], stage0_29[120], stage0_29[121], stage0_29[122], stage0_29[123], stage0_29[124]},
      {stage0_31[36], stage0_31[37], stage0_31[38], stage0_31[39], stage0_31[40], stage0_31[41]},
      {stage1_33[6],stage1_32[85],stage1_31[92],stage1_30[104],stage1_29[175]}
   );
   gpc606_5 gpc1225 (
      {stage0_29[125], stage0_29[126], stage0_29[127], stage0_29[128], stage0_29[129], stage0_29[130]},
      {stage0_31[42], stage0_31[43], stage0_31[44], stage0_31[45], stage0_31[46], stage0_31[47]},
      {stage1_33[7],stage1_32[86],stage1_31[93],stage1_30[105],stage1_29[176]}
   );
   gpc606_5 gpc1226 (
      {stage0_29[131], stage0_29[132], stage0_29[133], stage0_29[134], stage0_29[135], stage0_29[136]},
      {stage0_31[48], stage0_31[49], stage0_31[50], stage0_31[51], stage0_31[52], stage0_31[53]},
      {stage1_33[8],stage1_32[87],stage1_31[94],stage1_30[106],stage1_29[177]}
   );
   gpc606_5 gpc1227 (
      {stage0_29[137], stage0_29[138], stage0_29[139], stage0_29[140], stage0_29[141], stage0_29[142]},
      {stage0_31[54], stage0_31[55], stage0_31[56], stage0_31[57], stage0_31[58], stage0_31[59]},
      {stage1_33[9],stage1_32[88],stage1_31[95],stage1_30[107],stage1_29[178]}
   );
   gpc606_5 gpc1228 (
      {stage0_29[143], stage0_29[144], stage0_29[145], stage0_29[146], stage0_29[147], stage0_29[148]},
      {stage0_31[60], stage0_31[61], stage0_31[62], stage0_31[63], stage0_31[64], stage0_31[65]},
      {stage1_33[10],stage1_32[89],stage1_31[96],stage1_30[108],stage1_29[179]}
   );
   gpc606_5 gpc1229 (
      {stage0_29[149], stage0_29[150], stage0_29[151], stage0_29[152], stage0_29[153], stage0_29[154]},
      {stage0_31[66], stage0_31[67], stage0_31[68], stage0_31[69], stage0_31[70], stage0_31[71]},
      {stage1_33[11],stage1_32[90],stage1_31[97],stage1_30[109],stage1_29[180]}
   );
   gpc606_5 gpc1230 (
      {stage0_29[155], stage0_29[156], stage0_29[157], stage0_29[158], stage0_29[159], stage0_29[160]},
      {stage0_31[72], stage0_31[73], stage0_31[74], stage0_31[75], stage0_31[76], stage0_31[77]},
      {stage1_33[12],stage1_32[91],stage1_31[98],stage1_30[110],stage1_29[181]}
   );
   gpc606_5 gpc1231 (
      {stage0_29[161], stage0_29[162], stage0_29[163], stage0_29[164], stage0_29[165], stage0_29[166]},
      {stage0_31[78], stage0_31[79], stage0_31[80], stage0_31[81], stage0_31[82], stage0_31[83]},
      {stage1_33[13],stage1_32[92],stage1_31[99],stage1_30[111],stage1_29[182]}
   );
   gpc606_5 gpc1232 (
      {stage0_29[167], stage0_29[168], stage0_29[169], stage0_29[170], stage0_29[171], stage0_29[172]},
      {stage0_31[84], stage0_31[85], stage0_31[86], stage0_31[87], stage0_31[88], stage0_31[89]},
      {stage1_33[14],stage1_32[93],stage1_31[100],stage1_30[112],stage1_29[183]}
   );
   gpc606_5 gpc1233 (
      {stage0_29[173], stage0_29[174], stage0_29[175], stage0_29[176], stage0_29[177], stage0_29[178]},
      {stage0_31[90], stage0_31[91], stage0_31[92], stage0_31[93], stage0_31[94], stage0_31[95]},
      {stage1_33[15],stage1_32[94],stage1_31[101],stage1_30[113],stage1_29[184]}
   );
   gpc606_5 gpc1234 (
      {stage0_29[179], stage0_29[180], stage0_29[181], stage0_29[182], stage0_29[183], stage0_29[184]},
      {stage0_31[96], stage0_31[97], stage0_31[98], stage0_31[99], stage0_31[100], stage0_31[101]},
      {stage1_33[16],stage1_32[95],stage1_31[102],stage1_30[114],stage1_29[185]}
   );
   gpc606_5 gpc1235 (
      {stage0_29[185], stage0_29[186], stage0_29[187], stage0_29[188], stage0_29[189], stage0_29[190]},
      {stage0_31[102], stage0_31[103], stage0_31[104], stage0_31[105], stage0_31[106], stage0_31[107]},
      {stage1_33[17],stage1_32[96],stage1_31[103],stage1_30[115],stage1_29[186]}
   );
   gpc606_5 gpc1236 (
      {stage0_29[191], stage0_29[192], stage0_29[193], stage0_29[194], stage0_29[195], stage0_29[196]},
      {stage0_31[108], stage0_31[109], stage0_31[110], stage0_31[111], stage0_31[112], stage0_31[113]},
      {stage1_33[18],stage1_32[97],stage1_31[104],stage1_30[116],stage1_29[187]}
   );
   gpc606_5 gpc1237 (
      {stage0_29[197], stage0_29[198], stage0_29[199], stage0_29[200], stage0_29[201], stage0_29[202]},
      {stage0_31[114], stage0_31[115], stage0_31[116], stage0_31[117], stage0_31[118], stage0_31[119]},
      {stage1_33[19],stage1_32[98],stage1_31[105],stage1_30[117],stage1_29[188]}
   );
   gpc606_5 gpc1238 (
      {stage0_29[203], stage0_29[204], stage0_29[205], stage0_29[206], stage0_29[207], stage0_29[208]},
      {stage0_31[120], stage0_31[121], stage0_31[122], stage0_31[123], stage0_31[124], stage0_31[125]},
      {stage1_33[20],stage1_32[99],stage1_31[106],stage1_30[118],stage1_29[189]}
   );
   gpc606_5 gpc1239 (
      {stage0_29[209], stage0_29[210], stage0_29[211], stage0_29[212], stage0_29[213], stage0_29[214]},
      {stage0_31[126], stage0_31[127], stage0_31[128], stage0_31[129], stage0_31[130], stage0_31[131]},
      {stage1_33[21],stage1_32[100],stage1_31[107],stage1_30[119],stage1_29[190]}
   );
   gpc606_5 gpc1240 (
      {stage0_29[215], stage0_29[216], stage0_29[217], stage0_29[218], stage0_29[219], stage0_29[220]},
      {stage0_31[132], stage0_31[133], stage0_31[134], stage0_31[135], stage0_31[136], stage0_31[137]},
      {stage1_33[22],stage1_32[101],stage1_31[108],stage1_30[120],stage1_29[191]}
   );
   gpc606_5 gpc1241 (
      {stage0_29[221], stage0_29[222], stage0_29[223], stage0_29[224], stage0_29[225], stage0_29[226]},
      {stage0_31[138], stage0_31[139], stage0_31[140], stage0_31[141], stage0_31[142], stage0_31[143]},
      {stage1_33[23],stage1_32[102],stage1_31[109],stage1_30[121],stage1_29[192]}
   );
   gpc606_5 gpc1242 (
      {stage0_29[227], stage0_29[228], stage0_29[229], stage0_29[230], stage0_29[231], stage0_29[232]},
      {stage0_31[144], stage0_31[145], stage0_31[146], stage0_31[147], stage0_31[148], stage0_31[149]},
      {stage1_33[24],stage1_32[103],stage1_31[110],stage1_30[122],stage1_29[193]}
   );
   gpc606_5 gpc1243 (
      {stage0_29[233], stage0_29[234], stage0_29[235], stage0_29[236], stage0_29[237], stage0_29[238]},
      {stage0_31[150], stage0_31[151], stage0_31[152], stage0_31[153], stage0_31[154], stage0_31[155]},
      {stage1_33[25],stage1_32[104],stage1_31[111],stage1_30[123],stage1_29[194]}
   );
   gpc606_5 gpc1244 (
      {stage0_29[239], stage0_29[240], stage0_29[241], stage0_29[242], stage0_29[243], stage0_29[244]},
      {stage0_31[156], stage0_31[157], stage0_31[158], stage0_31[159], stage0_31[160], stage0_31[161]},
      {stage1_33[26],stage1_32[105],stage1_31[112],stage1_30[124],stage1_29[195]}
   );
   gpc606_5 gpc1245 (
      {stage0_29[245], stage0_29[246], stage0_29[247], stage0_29[248], stage0_29[249], stage0_29[250]},
      {stage0_31[162], stage0_31[163], stage0_31[164], stage0_31[165], stage0_31[166], stage0_31[167]},
      {stage1_33[27],stage1_32[106],stage1_31[113],stage1_30[125],stage1_29[196]}
   );
   gpc606_5 gpc1246 (
      {stage0_29[251], stage0_29[252], stage0_29[253], stage0_29[254], stage0_29[255], stage0_29[256]},
      {stage0_31[168], stage0_31[169], stage0_31[170], stage0_31[171], stage0_31[172], stage0_31[173]},
      {stage1_33[28],stage1_32[107],stage1_31[114],stage1_30[126],stage1_29[197]}
   );
   gpc606_5 gpc1247 (
      {stage0_29[257], stage0_29[258], stage0_29[259], stage0_29[260], stage0_29[261], stage0_29[262]},
      {stage0_31[174], stage0_31[175], stage0_31[176], stage0_31[177], stage0_31[178], stage0_31[179]},
      {stage1_33[29],stage1_32[108],stage1_31[115],stage1_30[127],stage1_29[198]}
   );
   gpc606_5 gpc1248 (
      {stage0_29[263], stage0_29[264], stage0_29[265], stage0_29[266], stage0_29[267], stage0_29[268]},
      {stage0_31[180], stage0_31[181], stage0_31[182], stage0_31[183], stage0_31[184], stage0_31[185]},
      {stage1_33[30],stage1_32[109],stage1_31[116],stage1_30[128],stage1_29[199]}
   );
   gpc606_5 gpc1249 (
      {stage0_29[269], stage0_29[270], stage0_29[271], stage0_29[272], stage0_29[273], stage0_29[274]},
      {stage0_31[186], stage0_31[187], stage0_31[188], stage0_31[189], stage0_31[190], stage0_31[191]},
      {stage1_33[31],stage1_32[110],stage1_31[117],stage1_30[129],stage1_29[200]}
   );
   gpc606_5 gpc1250 (
      {stage0_29[275], stage0_29[276], stage0_29[277], stage0_29[278], stage0_29[279], stage0_29[280]},
      {stage0_31[192], stage0_31[193], stage0_31[194], stage0_31[195], stage0_31[196], stage0_31[197]},
      {stage1_33[32],stage1_32[111],stage1_31[118],stage1_30[130],stage1_29[201]}
   );
   gpc606_5 gpc1251 (
      {stage0_29[281], stage0_29[282], stage0_29[283], stage0_29[284], stage0_29[285], stage0_29[286]},
      {stage0_31[198], stage0_31[199], stage0_31[200], stage0_31[201], stage0_31[202], stage0_31[203]},
      {stage1_33[33],stage1_32[112],stage1_31[119],stage1_30[131],stage1_29[202]}
   );
   gpc606_5 gpc1252 (
      {stage0_29[287], stage0_29[288], stage0_29[289], stage0_29[290], stage0_29[291], stage0_29[292]},
      {stage0_31[204], stage0_31[205], stage0_31[206], stage0_31[207], stage0_31[208], stage0_31[209]},
      {stage1_33[34],stage1_32[113],stage1_31[120],stage1_30[132],stage1_29[203]}
   );
   gpc606_5 gpc1253 (
      {stage0_29[293], stage0_29[294], stage0_29[295], stage0_29[296], stage0_29[297], stage0_29[298]},
      {stage0_31[210], stage0_31[211], stage0_31[212], stage0_31[213], stage0_31[214], stage0_31[215]},
      {stage1_33[35],stage1_32[114],stage1_31[121],stage1_30[133],stage1_29[204]}
   );
   gpc606_5 gpc1254 (
      {stage0_29[299], stage0_29[300], stage0_29[301], stage0_29[302], stage0_29[303], stage0_29[304]},
      {stage0_31[216], stage0_31[217], stage0_31[218], stage0_31[219], stage0_31[220], stage0_31[221]},
      {stage1_33[36],stage1_32[115],stage1_31[122],stage1_30[134],stage1_29[205]}
   );
   gpc606_5 gpc1255 (
      {stage0_29[305], stage0_29[306], stage0_29[307], stage0_29[308], stage0_29[309], stage0_29[310]},
      {stage0_31[222], stage0_31[223], stage0_31[224], stage0_31[225], stage0_31[226], stage0_31[227]},
      {stage1_33[37],stage1_32[116],stage1_31[123],stage1_30[135],stage1_29[206]}
   );
   gpc606_5 gpc1256 (
      {stage0_29[311], stage0_29[312], stage0_29[313], stage0_29[314], stage0_29[315], stage0_29[316]},
      {stage0_31[228], stage0_31[229], stage0_31[230], stage0_31[231], stage0_31[232], stage0_31[233]},
      {stage1_33[38],stage1_32[117],stage1_31[124],stage1_30[136],stage1_29[207]}
   );
   gpc606_5 gpc1257 (
      {stage0_29[317], stage0_29[318], stage0_29[319], stage0_29[320], stage0_29[321], stage0_29[322]},
      {stage0_31[234], stage0_31[235], stage0_31[236], stage0_31[237], stage0_31[238], stage0_31[239]},
      {stage1_33[39],stage1_32[118],stage1_31[125],stage1_30[137],stage1_29[208]}
   );
   gpc606_5 gpc1258 (
      {stage0_29[323], stage0_29[324], stage0_29[325], stage0_29[326], stage0_29[327], stage0_29[328]},
      {stage0_31[240], stage0_31[241], stage0_31[242], stage0_31[243], stage0_31[244], stage0_31[245]},
      {stage1_33[40],stage1_32[119],stage1_31[126],stage1_30[138],stage1_29[209]}
   );
   gpc606_5 gpc1259 (
      {stage0_29[329], stage0_29[330], stage0_29[331], stage0_29[332], stage0_29[333], stage0_29[334]},
      {stage0_31[246], stage0_31[247], stage0_31[248], stage0_31[249], stage0_31[250], stage0_31[251]},
      {stage1_33[41],stage1_32[120],stage1_31[127],stage1_30[139],stage1_29[210]}
   );
   gpc606_5 gpc1260 (
      {stage0_29[335], stage0_29[336], stage0_29[337], stage0_29[338], stage0_29[339], stage0_29[340]},
      {stage0_31[252], stage0_31[253], stage0_31[254], stage0_31[255], stage0_31[256], stage0_31[257]},
      {stage1_33[42],stage1_32[121],stage1_31[128],stage1_30[140],stage1_29[211]}
   );
   gpc606_5 gpc1261 (
      {stage0_29[341], stage0_29[342], stage0_29[343], stage0_29[344], stage0_29[345], stage0_29[346]},
      {stage0_31[258], stage0_31[259], stage0_31[260], stage0_31[261], stage0_31[262], stage0_31[263]},
      {stage1_33[43],stage1_32[122],stage1_31[129],stage1_30[141],stage1_29[212]}
   );
   gpc606_5 gpc1262 (
      {stage0_29[347], stage0_29[348], stage0_29[349], stage0_29[350], stage0_29[351], stage0_29[352]},
      {stage0_31[264], stage0_31[265], stage0_31[266], stage0_31[267], stage0_31[268], stage0_31[269]},
      {stage1_33[44],stage1_32[123],stage1_31[130],stage1_30[142],stage1_29[213]}
   );
   gpc606_5 gpc1263 (
      {stage0_29[353], stage0_29[354], stage0_29[355], stage0_29[356], stage0_29[357], stage0_29[358]},
      {stage0_31[270], stage0_31[271], stage0_31[272], stage0_31[273], stage0_31[274], stage0_31[275]},
      {stage1_33[45],stage1_32[124],stage1_31[131],stage1_30[143],stage1_29[214]}
   );
   gpc606_5 gpc1264 (
      {stage0_29[359], stage0_29[360], stage0_29[361], stage0_29[362], stage0_29[363], stage0_29[364]},
      {stage0_31[276], stage0_31[277], stage0_31[278], stage0_31[279], stage0_31[280], stage0_31[281]},
      {stage1_33[46],stage1_32[125],stage1_31[132],stage1_30[144],stage1_29[215]}
   );
   gpc606_5 gpc1265 (
      {stage0_29[365], stage0_29[366], stage0_29[367], stage0_29[368], stage0_29[369], stage0_29[370]},
      {stage0_31[282], stage0_31[283], stage0_31[284], stage0_31[285], stage0_31[286], stage0_31[287]},
      {stage1_33[47],stage1_32[126],stage1_31[133],stage1_30[145],stage1_29[216]}
   );
   gpc606_5 gpc1266 (
      {stage0_29[371], stage0_29[372], stage0_29[373], stage0_29[374], stage0_29[375], stage0_29[376]},
      {stage0_31[288], stage0_31[289], stage0_31[290], stage0_31[291], stage0_31[292], stage0_31[293]},
      {stage1_33[48],stage1_32[127],stage1_31[134],stage1_30[146],stage1_29[217]}
   );
   gpc606_5 gpc1267 (
      {stage0_29[377], stage0_29[378], stage0_29[379], stage0_29[380], stage0_29[381], stage0_29[382]},
      {stage0_31[294], stage0_31[295], stage0_31[296], stage0_31[297], stage0_31[298], stage0_31[299]},
      {stage1_33[49],stage1_32[128],stage1_31[135],stage1_30[147],stage1_29[218]}
   );
   gpc606_5 gpc1268 (
      {stage0_29[383], stage0_29[384], stage0_29[385], stage0_29[386], stage0_29[387], stage0_29[388]},
      {stage0_31[300], stage0_31[301], stage0_31[302], stage0_31[303], stage0_31[304], stage0_31[305]},
      {stage1_33[50],stage1_32[129],stage1_31[136],stage1_30[148],stage1_29[219]}
   );
   gpc606_5 gpc1269 (
      {stage0_29[389], stage0_29[390], stage0_29[391], stage0_29[392], stage0_29[393], stage0_29[394]},
      {stage0_31[306], stage0_31[307], stage0_31[308], stage0_31[309], stage0_31[310], stage0_31[311]},
      {stage1_33[51],stage1_32[130],stage1_31[137],stage1_30[149],stage1_29[220]}
   );
   gpc606_5 gpc1270 (
      {stage0_29[395], stage0_29[396], stage0_29[397], stage0_29[398], stage0_29[399], stage0_29[400]},
      {stage0_31[312], stage0_31[313], stage0_31[314], stage0_31[315], stage0_31[316], stage0_31[317]},
      {stage1_33[52],stage1_32[131],stage1_31[138],stage1_30[150],stage1_29[221]}
   );
   gpc606_5 gpc1271 (
      {stage0_29[401], stage0_29[402], stage0_29[403], stage0_29[404], stage0_29[405], stage0_29[406]},
      {stage0_31[318], stage0_31[319], stage0_31[320], stage0_31[321], stage0_31[322], stage0_31[323]},
      {stage1_33[53],stage1_32[132],stage1_31[139],stage1_30[151],stage1_29[222]}
   );
   gpc606_5 gpc1272 (
      {stage0_29[407], stage0_29[408], stage0_29[409], stage0_29[410], stage0_29[411], stage0_29[412]},
      {stage0_31[324], stage0_31[325], stage0_31[326], stage0_31[327], stage0_31[328], stage0_31[329]},
      {stage1_33[54],stage1_32[133],stage1_31[140],stage1_30[152],stage1_29[223]}
   );
   gpc606_5 gpc1273 (
      {stage0_29[413], stage0_29[414], stage0_29[415], stage0_29[416], stage0_29[417], stage0_29[418]},
      {stage0_31[330], stage0_31[331], stage0_31[332], stage0_31[333], stage0_31[334], stage0_31[335]},
      {stage1_33[55],stage1_32[134],stage1_31[141],stage1_30[153],stage1_29[224]}
   );
   gpc606_5 gpc1274 (
      {stage0_29[419], stage0_29[420], stage0_29[421], stage0_29[422], stage0_29[423], stage0_29[424]},
      {stage0_31[336], stage0_31[337], stage0_31[338], stage0_31[339], stage0_31[340], stage0_31[341]},
      {stage1_33[56],stage1_32[135],stage1_31[142],stage1_30[154],stage1_29[225]}
   );
   gpc606_5 gpc1275 (
      {stage0_29[425], stage0_29[426], stage0_29[427], stage0_29[428], stage0_29[429], stage0_29[430]},
      {stage0_31[342], stage0_31[343], stage0_31[344], stage0_31[345], stage0_31[346], stage0_31[347]},
      {stage1_33[57],stage1_32[136],stage1_31[143],stage1_30[155],stage1_29[226]}
   );
   gpc606_5 gpc1276 (
      {stage0_29[431], stage0_29[432], stage0_29[433], stage0_29[434], stage0_29[435], stage0_29[436]},
      {stage0_31[348], stage0_31[349], stage0_31[350], stage0_31[351], stage0_31[352], stage0_31[353]},
      {stage1_33[58],stage1_32[137],stage1_31[144],stage1_30[156],stage1_29[227]}
   );
   gpc606_5 gpc1277 (
      {stage0_29[437], stage0_29[438], stage0_29[439], stage0_29[440], stage0_29[441], stage0_29[442]},
      {stage0_31[354], stage0_31[355], stage0_31[356], stage0_31[357], stage0_31[358], stage0_31[359]},
      {stage1_33[59],stage1_32[138],stage1_31[145],stage1_30[157],stage1_29[228]}
   );
   gpc606_5 gpc1278 (
      {stage0_29[443], stage0_29[444], stage0_29[445], stage0_29[446], stage0_29[447], stage0_29[448]},
      {stage0_31[360], stage0_31[361], stage0_31[362], stage0_31[363], stage0_31[364], stage0_31[365]},
      {stage1_33[60],stage1_32[139],stage1_31[146],stage1_30[158],stage1_29[229]}
   );
   gpc606_5 gpc1279 (
      {stage0_29[449], stage0_29[450], stage0_29[451], stage0_29[452], stage0_29[453], stage0_29[454]},
      {stage0_31[366], stage0_31[367], stage0_31[368], stage0_31[369], stage0_31[370], stage0_31[371]},
      {stage1_33[61],stage1_32[140],stage1_31[147],stage1_30[159],stage1_29[230]}
   );
   gpc606_5 gpc1280 (
      {stage0_29[455], stage0_29[456], stage0_29[457], stage0_29[458], stage0_29[459], stage0_29[460]},
      {stage0_31[372], stage0_31[373], stage0_31[374], stage0_31[375], stage0_31[376], stage0_31[377]},
      {stage1_33[62],stage1_32[141],stage1_31[148],stage1_30[160],stage1_29[231]}
   );
   gpc606_5 gpc1281 (
      {stage0_29[461], stage0_29[462], stage0_29[463], stage0_29[464], stage0_29[465], stage0_29[466]},
      {stage0_31[378], stage0_31[379], stage0_31[380], stage0_31[381], stage0_31[382], stage0_31[383]},
      {stage1_33[63],stage1_32[142],stage1_31[149],stage1_30[161],stage1_29[232]}
   );
   gpc606_5 gpc1282 (
      {stage0_29[467], stage0_29[468], stage0_29[469], stage0_29[470], stage0_29[471], stage0_29[472]},
      {stage0_31[384], stage0_31[385], stage0_31[386], stage0_31[387], stage0_31[388], stage0_31[389]},
      {stage1_33[64],stage1_32[143],stage1_31[150],stage1_30[162],stage1_29[233]}
   );
   gpc606_5 gpc1283 (
      {stage0_29[473], stage0_29[474], stage0_29[475], stage0_29[476], stage0_29[477], stage0_29[478]},
      {stage0_31[390], stage0_31[391], stage0_31[392], stage0_31[393], stage0_31[394], stage0_31[395]},
      {stage1_33[65],stage1_32[144],stage1_31[151],stage1_30[163],stage1_29[234]}
   );
   gpc606_5 gpc1284 (
      {stage0_29[479], stage0_29[480], stage0_29[481], stage0_29[482], stage0_29[483], stage0_29[484]},
      {stage0_31[396], stage0_31[397], stage0_31[398], stage0_31[399], stage0_31[400], stage0_31[401]},
      {stage1_33[66],stage1_32[145],stage1_31[152],stage1_30[164],stage1_29[235]}
   );
   gpc606_5 gpc1285 (
      {stage0_29[485], stage0_29[486], stage0_29[487], stage0_29[488], stage0_29[489], stage0_29[490]},
      {stage0_31[402], stage0_31[403], stage0_31[404], stage0_31[405], stage0_31[406], stage0_31[407]},
      {stage1_33[67],stage1_32[146],stage1_31[153],stage1_30[165],stage1_29[236]}
   );
   gpc606_5 gpc1286 (
      {stage0_29[491], stage0_29[492], stage0_29[493], stage0_29[494], stage0_29[495], stage0_29[496]},
      {stage0_31[408], stage0_31[409], stage0_31[410], stage0_31[411], stage0_31[412], stage0_31[413]},
      {stage1_33[68],stage1_32[147],stage1_31[154],stage1_30[166],stage1_29[237]}
   );
   gpc606_5 gpc1287 (
      {stage0_29[497], stage0_29[498], stage0_29[499], stage0_29[500], stage0_29[501], stage0_29[502]},
      {stage0_31[414], stage0_31[415], stage0_31[416], stage0_31[417], stage0_31[418], stage0_31[419]},
      {stage1_33[69],stage1_32[148],stage1_31[155],stage1_30[167],stage1_29[238]}
   );
   gpc606_5 gpc1288 (
      {stage0_29[503], stage0_29[504], stage0_29[505], stage0_29[506], stage0_29[507], stage0_29[508]},
      {stage0_31[420], stage0_31[421], stage0_31[422], stage0_31[423], stage0_31[424], stage0_31[425]},
      {stage1_33[70],stage1_32[149],stage1_31[156],stage1_30[168],stage1_29[239]}
   );
   gpc1_1 gpc1289 (
      {stage0_0[502]},
      {stage1_0[101]}
   );
   gpc1_1 gpc1290 (
      {stage0_0[503]},
      {stage1_0[102]}
   );
   gpc1_1 gpc1291 (
      {stage0_0[504]},
      {stage1_0[103]}
   );
   gpc1_1 gpc1292 (
      {stage0_0[505]},
      {stage1_0[104]}
   );
   gpc1_1 gpc1293 (
      {stage0_0[506]},
      {stage1_0[105]}
   );
   gpc1_1 gpc1294 (
      {stage0_0[507]},
      {stage1_0[106]}
   );
   gpc1_1 gpc1295 (
      {stage0_0[508]},
      {stage1_0[107]}
   );
   gpc1_1 gpc1296 (
      {stage0_0[509]},
      {stage1_0[108]}
   );
   gpc1_1 gpc1297 (
      {stage0_0[510]},
      {stage1_0[109]}
   );
   gpc1_1 gpc1298 (
      {stage0_0[511]},
      {stage1_0[110]}
   );
   gpc1_1 gpc1299 (
      {stage0_1[453]},
      {stage1_1[140]}
   );
   gpc1_1 gpc1300 (
      {stage0_1[454]},
      {stage1_1[141]}
   );
   gpc1_1 gpc1301 (
      {stage0_1[455]},
      {stage1_1[142]}
   );
   gpc1_1 gpc1302 (
      {stage0_1[456]},
      {stage1_1[143]}
   );
   gpc1_1 gpc1303 (
      {stage0_1[457]},
      {stage1_1[144]}
   );
   gpc1_1 gpc1304 (
      {stage0_1[458]},
      {stage1_1[145]}
   );
   gpc1_1 gpc1305 (
      {stage0_1[459]},
      {stage1_1[146]}
   );
   gpc1_1 gpc1306 (
      {stage0_1[460]},
      {stage1_1[147]}
   );
   gpc1_1 gpc1307 (
      {stage0_1[461]},
      {stage1_1[148]}
   );
   gpc1_1 gpc1308 (
      {stage0_1[462]},
      {stage1_1[149]}
   );
   gpc1_1 gpc1309 (
      {stage0_1[463]},
      {stage1_1[150]}
   );
   gpc1_1 gpc1310 (
      {stage0_1[464]},
      {stage1_1[151]}
   );
   gpc1_1 gpc1311 (
      {stage0_1[465]},
      {stage1_1[152]}
   );
   gpc1_1 gpc1312 (
      {stage0_1[466]},
      {stage1_1[153]}
   );
   gpc1_1 gpc1313 (
      {stage0_1[467]},
      {stage1_1[154]}
   );
   gpc1_1 gpc1314 (
      {stage0_1[468]},
      {stage1_1[155]}
   );
   gpc1_1 gpc1315 (
      {stage0_1[469]},
      {stage1_1[156]}
   );
   gpc1_1 gpc1316 (
      {stage0_1[470]},
      {stage1_1[157]}
   );
   gpc1_1 gpc1317 (
      {stage0_1[471]},
      {stage1_1[158]}
   );
   gpc1_1 gpc1318 (
      {stage0_1[472]},
      {stage1_1[159]}
   );
   gpc1_1 gpc1319 (
      {stage0_1[473]},
      {stage1_1[160]}
   );
   gpc1_1 gpc1320 (
      {stage0_1[474]},
      {stage1_1[161]}
   );
   gpc1_1 gpc1321 (
      {stage0_1[475]},
      {stage1_1[162]}
   );
   gpc1_1 gpc1322 (
      {stage0_1[476]},
      {stage1_1[163]}
   );
   gpc1_1 gpc1323 (
      {stage0_1[477]},
      {stage1_1[164]}
   );
   gpc1_1 gpc1324 (
      {stage0_1[478]},
      {stage1_1[165]}
   );
   gpc1_1 gpc1325 (
      {stage0_1[479]},
      {stage1_1[166]}
   );
   gpc1_1 gpc1326 (
      {stage0_1[480]},
      {stage1_1[167]}
   );
   gpc1_1 gpc1327 (
      {stage0_1[481]},
      {stage1_1[168]}
   );
   gpc1_1 gpc1328 (
      {stage0_1[482]},
      {stage1_1[169]}
   );
   gpc1_1 gpc1329 (
      {stage0_1[483]},
      {stage1_1[170]}
   );
   gpc1_1 gpc1330 (
      {stage0_1[484]},
      {stage1_1[171]}
   );
   gpc1_1 gpc1331 (
      {stage0_1[485]},
      {stage1_1[172]}
   );
   gpc1_1 gpc1332 (
      {stage0_1[486]},
      {stage1_1[173]}
   );
   gpc1_1 gpc1333 (
      {stage0_1[487]},
      {stage1_1[174]}
   );
   gpc1_1 gpc1334 (
      {stage0_1[488]},
      {stage1_1[175]}
   );
   gpc1_1 gpc1335 (
      {stage0_1[489]},
      {stage1_1[176]}
   );
   gpc1_1 gpc1336 (
      {stage0_1[490]},
      {stage1_1[177]}
   );
   gpc1_1 gpc1337 (
      {stage0_1[491]},
      {stage1_1[178]}
   );
   gpc1_1 gpc1338 (
      {stage0_1[492]},
      {stage1_1[179]}
   );
   gpc1_1 gpc1339 (
      {stage0_1[493]},
      {stage1_1[180]}
   );
   gpc1_1 gpc1340 (
      {stage0_1[494]},
      {stage1_1[181]}
   );
   gpc1_1 gpc1341 (
      {stage0_1[495]},
      {stage1_1[182]}
   );
   gpc1_1 gpc1342 (
      {stage0_1[496]},
      {stage1_1[183]}
   );
   gpc1_1 gpc1343 (
      {stage0_1[497]},
      {stage1_1[184]}
   );
   gpc1_1 gpc1344 (
      {stage0_1[498]},
      {stage1_1[185]}
   );
   gpc1_1 gpc1345 (
      {stage0_1[499]},
      {stage1_1[186]}
   );
   gpc1_1 gpc1346 (
      {stage0_1[500]},
      {stage1_1[187]}
   );
   gpc1_1 gpc1347 (
      {stage0_1[501]},
      {stage1_1[188]}
   );
   gpc1_1 gpc1348 (
      {stage0_1[502]},
      {stage1_1[189]}
   );
   gpc1_1 gpc1349 (
      {stage0_1[503]},
      {stage1_1[190]}
   );
   gpc1_1 gpc1350 (
      {stage0_1[504]},
      {stage1_1[191]}
   );
   gpc1_1 gpc1351 (
      {stage0_1[505]},
      {stage1_1[192]}
   );
   gpc1_1 gpc1352 (
      {stage0_1[506]},
      {stage1_1[193]}
   );
   gpc1_1 gpc1353 (
      {stage0_1[507]},
      {stage1_1[194]}
   );
   gpc1_1 gpc1354 (
      {stage0_1[508]},
      {stage1_1[195]}
   );
   gpc1_1 gpc1355 (
      {stage0_1[509]},
      {stage1_1[196]}
   );
   gpc1_1 gpc1356 (
      {stage0_1[510]},
      {stage1_1[197]}
   );
   gpc1_1 gpc1357 (
      {stage0_1[511]},
      {stage1_1[198]}
   );
   gpc1_1 gpc1358 (
      {stage0_2[481]},
      {stage1_2[157]}
   );
   gpc1_1 gpc1359 (
      {stage0_2[482]},
      {stage1_2[158]}
   );
   gpc1_1 gpc1360 (
      {stage0_2[483]},
      {stage1_2[159]}
   );
   gpc1_1 gpc1361 (
      {stage0_2[484]},
      {stage1_2[160]}
   );
   gpc1_1 gpc1362 (
      {stage0_2[485]},
      {stage1_2[161]}
   );
   gpc1_1 gpc1363 (
      {stage0_2[486]},
      {stage1_2[162]}
   );
   gpc1_1 gpc1364 (
      {stage0_2[487]},
      {stage1_2[163]}
   );
   gpc1_1 gpc1365 (
      {stage0_2[488]},
      {stage1_2[164]}
   );
   gpc1_1 gpc1366 (
      {stage0_2[489]},
      {stage1_2[165]}
   );
   gpc1_1 gpc1367 (
      {stage0_2[490]},
      {stage1_2[166]}
   );
   gpc1_1 gpc1368 (
      {stage0_2[491]},
      {stage1_2[167]}
   );
   gpc1_1 gpc1369 (
      {stage0_2[492]},
      {stage1_2[168]}
   );
   gpc1_1 gpc1370 (
      {stage0_2[493]},
      {stage1_2[169]}
   );
   gpc1_1 gpc1371 (
      {stage0_2[494]},
      {stage1_2[170]}
   );
   gpc1_1 gpc1372 (
      {stage0_2[495]},
      {stage1_2[171]}
   );
   gpc1_1 gpc1373 (
      {stage0_2[496]},
      {stage1_2[172]}
   );
   gpc1_1 gpc1374 (
      {stage0_2[497]},
      {stage1_2[173]}
   );
   gpc1_1 gpc1375 (
      {stage0_2[498]},
      {stage1_2[174]}
   );
   gpc1_1 gpc1376 (
      {stage0_2[499]},
      {stage1_2[175]}
   );
   gpc1_1 gpc1377 (
      {stage0_2[500]},
      {stage1_2[176]}
   );
   gpc1_1 gpc1378 (
      {stage0_2[501]},
      {stage1_2[177]}
   );
   gpc1_1 gpc1379 (
      {stage0_2[502]},
      {stage1_2[178]}
   );
   gpc1_1 gpc1380 (
      {stage0_2[503]},
      {stage1_2[179]}
   );
   gpc1_1 gpc1381 (
      {stage0_2[504]},
      {stage1_2[180]}
   );
   gpc1_1 gpc1382 (
      {stage0_2[505]},
      {stage1_2[181]}
   );
   gpc1_1 gpc1383 (
      {stage0_2[506]},
      {stage1_2[182]}
   );
   gpc1_1 gpc1384 (
      {stage0_2[507]},
      {stage1_2[183]}
   );
   gpc1_1 gpc1385 (
      {stage0_2[508]},
      {stage1_2[184]}
   );
   gpc1_1 gpc1386 (
      {stage0_2[509]},
      {stage1_2[185]}
   );
   gpc1_1 gpc1387 (
      {stage0_2[510]},
      {stage1_2[186]}
   );
   gpc1_1 gpc1388 (
      {stage0_2[511]},
      {stage1_2[187]}
   );
   gpc1_1 gpc1389 (
      {stage0_3[414]},
      {stage1_3[179]}
   );
   gpc1_1 gpc1390 (
      {stage0_3[415]},
      {stage1_3[180]}
   );
   gpc1_1 gpc1391 (
      {stage0_3[416]},
      {stage1_3[181]}
   );
   gpc1_1 gpc1392 (
      {stage0_3[417]},
      {stage1_3[182]}
   );
   gpc1_1 gpc1393 (
      {stage0_3[418]},
      {stage1_3[183]}
   );
   gpc1_1 gpc1394 (
      {stage0_3[419]},
      {stage1_3[184]}
   );
   gpc1_1 gpc1395 (
      {stage0_3[420]},
      {stage1_3[185]}
   );
   gpc1_1 gpc1396 (
      {stage0_3[421]},
      {stage1_3[186]}
   );
   gpc1_1 gpc1397 (
      {stage0_3[422]},
      {stage1_3[187]}
   );
   gpc1_1 gpc1398 (
      {stage0_3[423]},
      {stage1_3[188]}
   );
   gpc1_1 gpc1399 (
      {stage0_3[424]},
      {stage1_3[189]}
   );
   gpc1_1 gpc1400 (
      {stage0_3[425]},
      {stage1_3[190]}
   );
   gpc1_1 gpc1401 (
      {stage0_3[426]},
      {stage1_3[191]}
   );
   gpc1_1 gpc1402 (
      {stage0_3[427]},
      {stage1_3[192]}
   );
   gpc1_1 gpc1403 (
      {stage0_3[428]},
      {stage1_3[193]}
   );
   gpc1_1 gpc1404 (
      {stage0_3[429]},
      {stage1_3[194]}
   );
   gpc1_1 gpc1405 (
      {stage0_3[430]},
      {stage1_3[195]}
   );
   gpc1_1 gpc1406 (
      {stage0_3[431]},
      {stage1_3[196]}
   );
   gpc1_1 gpc1407 (
      {stage0_3[432]},
      {stage1_3[197]}
   );
   gpc1_1 gpc1408 (
      {stage0_3[433]},
      {stage1_3[198]}
   );
   gpc1_1 gpc1409 (
      {stage0_3[434]},
      {stage1_3[199]}
   );
   gpc1_1 gpc1410 (
      {stage0_3[435]},
      {stage1_3[200]}
   );
   gpc1_1 gpc1411 (
      {stage0_3[436]},
      {stage1_3[201]}
   );
   gpc1_1 gpc1412 (
      {stage0_3[437]},
      {stage1_3[202]}
   );
   gpc1_1 gpc1413 (
      {stage0_3[438]},
      {stage1_3[203]}
   );
   gpc1_1 gpc1414 (
      {stage0_3[439]},
      {stage1_3[204]}
   );
   gpc1_1 gpc1415 (
      {stage0_3[440]},
      {stage1_3[205]}
   );
   gpc1_1 gpc1416 (
      {stage0_3[441]},
      {stage1_3[206]}
   );
   gpc1_1 gpc1417 (
      {stage0_3[442]},
      {stage1_3[207]}
   );
   gpc1_1 gpc1418 (
      {stage0_3[443]},
      {stage1_3[208]}
   );
   gpc1_1 gpc1419 (
      {stage0_3[444]},
      {stage1_3[209]}
   );
   gpc1_1 gpc1420 (
      {stage0_3[445]},
      {stage1_3[210]}
   );
   gpc1_1 gpc1421 (
      {stage0_3[446]},
      {stage1_3[211]}
   );
   gpc1_1 gpc1422 (
      {stage0_3[447]},
      {stage1_3[212]}
   );
   gpc1_1 gpc1423 (
      {stage0_3[448]},
      {stage1_3[213]}
   );
   gpc1_1 gpc1424 (
      {stage0_3[449]},
      {stage1_3[214]}
   );
   gpc1_1 gpc1425 (
      {stage0_3[450]},
      {stage1_3[215]}
   );
   gpc1_1 gpc1426 (
      {stage0_3[451]},
      {stage1_3[216]}
   );
   gpc1_1 gpc1427 (
      {stage0_3[452]},
      {stage1_3[217]}
   );
   gpc1_1 gpc1428 (
      {stage0_3[453]},
      {stage1_3[218]}
   );
   gpc1_1 gpc1429 (
      {stage0_3[454]},
      {stage1_3[219]}
   );
   gpc1_1 gpc1430 (
      {stage0_3[455]},
      {stage1_3[220]}
   );
   gpc1_1 gpc1431 (
      {stage0_3[456]},
      {stage1_3[221]}
   );
   gpc1_1 gpc1432 (
      {stage0_3[457]},
      {stage1_3[222]}
   );
   gpc1_1 gpc1433 (
      {stage0_3[458]},
      {stage1_3[223]}
   );
   gpc1_1 gpc1434 (
      {stage0_3[459]},
      {stage1_3[224]}
   );
   gpc1_1 gpc1435 (
      {stage0_3[460]},
      {stage1_3[225]}
   );
   gpc1_1 gpc1436 (
      {stage0_3[461]},
      {stage1_3[226]}
   );
   gpc1_1 gpc1437 (
      {stage0_3[462]},
      {stage1_3[227]}
   );
   gpc1_1 gpc1438 (
      {stage0_3[463]},
      {stage1_3[228]}
   );
   gpc1_1 gpc1439 (
      {stage0_3[464]},
      {stage1_3[229]}
   );
   gpc1_1 gpc1440 (
      {stage0_3[465]},
      {stage1_3[230]}
   );
   gpc1_1 gpc1441 (
      {stage0_3[466]},
      {stage1_3[231]}
   );
   gpc1_1 gpc1442 (
      {stage0_3[467]},
      {stage1_3[232]}
   );
   gpc1_1 gpc1443 (
      {stage0_3[468]},
      {stage1_3[233]}
   );
   gpc1_1 gpc1444 (
      {stage0_3[469]},
      {stage1_3[234]}
   );
   gpc1_1 gpc1445 (
      {stage0_3[470]},
      {stage1_3[235]}
   );
   gpc1_1 gpc1446 (
      {stage0_3[471]},
      {stage1_3[236]}
   );
   gpc1_1 gpc1447 (
      {stage0_3[472]},
      {stage1_3[237]}
   );
   gpc1_1 gpc1448 (
      {stage0_3[473]},
      {stage1_3[238]}
   );
   gpc1_1 gpc1449 (
      {stage0_3[474]},
      {stage1_3[239]}
   );
   gpc1_1 gpc1450 (
      {stage0_3[475]},
      {stage1_3[240]}
   );
   gpc1_1 gpc1451 (
      {stage0_3[476]},
      {stage1_3[241]}
   );
   gpc1_1 gpc1452 (
      {stage0_3[477]},
      {stage1_3[242]}
   );
   gpc1_1 gpc1453 (
      {stage0_3[478]},
      {stage1_3[243]}
   );
   gpc1_1 gpc1454 (
      {stage0_3[479]},
      {stage1_3[244]}
   );
   gpc1_1 gpc1455 (
      {stage0_3[480]},
      {stage1_3[245]}
   );
   gpc1_1 gpc1456 (
      {stage0_3[481]},
      {stage1_3[246]}
   );
   gpc1_1 gpc1457 (
      {stage0_3[482]},
      {stage1_3[247]}
   );
   gpc1_1 gpc1458 (
      {stage0_3[483]},
      {stage1_3[248]}
   );
   gpc1_1 gpc1459 (
      {stage0_3[484]},
      {stage1_3[249]}
   );
   gpc1_1 gpc1460 (
      {stage0_3[485]},
      {stage1_3[250]}
   );
   gpc1_1 gpc1461 (
      {stage0_3[486]},
      {stage1_3[251]}
   );
   gpc1_1 gpc1462 (
      {stage0_3[487]},
      {stage1_3[252]}
   );
   gpc1_1 gpc1463 (
      {stage0_3[488]},
      {stage1_3[253]}
   );
   gpc1_1 gpc1464 (
      {stage0_3[489]},
      {stage1_3[254]}
   );
   gpc1_1 gpc1465 (
      {stage0_3[490]},
      {stage1_3[255]}
   );
   gpc1_1 gpc1466 (
      {stage0_3[491]},
      {stage1_3[256]}
   );
   gpc1_1 gpc1467 (
      {stage0_3[492]},
      {stage1_3[257]}
   );
   gpc1_1 gpc1468 (
      {stage0_3[493]},
      {stage1_3[258]}
   );
   gpc1_1 gpc1469 (
      {stage0_3[494]},
      {stage1_3[259]}
   );
   gpc1_1 gpc1470 (
      {stage0_3[495]},
      {stage1_3[260]}
   );
   gpc1_1 gpc1471 (
      {stage0_3[496]},
      {stage1_3[261]}
   );
   gpc1_1 gpc1472 (
      {stage0_3[497]},
      {stage1_3[262]}
   );
   gpc1_1 gpc1473 (
      {stage0_3[498]},
      {stage1_3[263]}
   );
   gpc1_1 gpc1474 (
      {stage0_3[499]},
      {stage1_3[264]}
   );
   gpc1_1 gpc1475 (
      {stage0_3[500]},
      {stage1_3[265]}
   );
   gpc1_1 gpc1476 (
      {stage0_3[501]},
      {stage1_3[266]}
   );
   gpc1_1 gpc1477 (
      {stage0_3[502]},
      {stage1_3[267]}
   );
   gpc1_1 gpc1478 (
      {stage0_3[503]},
      {stage1_3[268]}
   );
   gpc1_1 gpc1479 (
      {stage0_3[504]},
      {stage1_3[269]}
   );
   gpc1_1 gpc1480 (
      {stage0_3[505]},
      {stage1_3[270]}
   );
   gpc1_1 gpc1481 (
      {stage0_3[506]},
      {stage1_3[271]}
   );
   gpc1_1 gpc1482 (
      {stage0_3[507]},
      {stage1_3[272]}
   );
   gpc1_1 gpc1483 (
      {stage0_3[508]},
      {stage1_3[273]}
   );
   gpc1_1 gpc1484 (
      {stage0_3[509]},
      {stage1_3[274]}
   );
   gpc1_1 gpc1485 (
      {stage0_3[510]},
      {stage1_3[275]}
   );
   gpc1_1 gpc1486 (
      {stage0_3[511]},
      {stage1_3[276]}
   );
   gpc1_1 gpc1487 (
      {stage0_6[446]},
      {stage1_6[177]}
   );
   gpc1_1 gpc1488 (
      {stage0_6[447]},
      {stage1_6[178]}
   );
   gpc1_1 gpc1489 (
      {stage0_6[448]},
      {stage1_6[179]}
   );
   gpc1_1 gpc1490 (
      {stage0_6[449]},
      {stage1_6[180]}
   );
   gpc1_1 gpc1491 (
      {stage0_6[450]},
      {stage1_6[181]}
   );
   gpc1_1 gpc1492 (
      {stage0_6[451]},
      {stage1_6[182]}
   );
   gpc1_1 gpc1493 (
      {stage0_6[452]},
      {stage1_6[183]}
   );
   gpc1_1 gpc1494 (
      {stage0_6[453]},
      {stage1_6[184]}
   );
   gpc1_1 gpc1495 (
      {stage0_6[454]},
      {stage1_6[185]}
   );
   gpc1_1 gpc1496 (
      {stage0_6[455]},
      {stage1_6[186]}
   );
   gpc1_1 gpc1497 (
      {stage0_6[456]},
      {stage1_6[187]}
   );
   gpc1_1 gpc1498 (
      {stage0_6[457]},
      {stage1_6[188]}
   );
   gpc1_1 gpc1499 (
      {stage0_6[458]},
      {stage1_6[189]}
   );
   gpc1_1 gpc1500 (
      {stage0_6[459]},
      {stage1_6[190]}
   );
   gpc1_1 gpc1501 (
      {stage0_6[460]},
      {stage1_6[191]}
   );
   gpc1_1 gpc1502 (
      {stage0_6[461]},
      {stage1_6[192]}
   );
   gpc1_1 gpc1503 (
      {stage0_6[462]},
      {stage1_6[193]}
   );
   gpc1_1 gpc1504 (
      {stage0_6[463]},
      {stage1_6[194]}
   );
   gpc1_1 gpc1505 (
      {stage0_6[464]},
      {stage1_6[195]}
   );
   gpc1_1 gpc1506 (
      {stage0_6[465]},
      {stage1_6[196]}
   );
   gpc1_1 gpc1507 (
      {stage0_6[466]},
      {stage1_6[197]}
   );
   gpc1_1 gpc1508 (
      {stage0_6[467]},
      {stage1_6[198]}
   );
   gpc1_1 gpc1509 (
      {stage0_6[468]},
      {stage1_6[199]}
   );
   gpc1_1 gpc1510 (
      {stage0_6[469]},
      {stage1_6[200]}
   );
   gpc1_1 gpc1511 (
      {stage0_6[470]},
      {stage1_6[201]}
   );
   gpc1_1 gpc1512 (
      {stage0_6[471]},
      {stage1_6[202]}
   );
   gpc1_1 gpc1513 (
      {stage0_6[472]},
      {stage1_6[203]}
   );
   gpc1_1 gpc1514 (
      {stage0_6[473]},
      {stage1_6[204]}
   );
   gpc1_1 gpc1515 (
      {stage0_6[474]},
      {stage1_6[205]}
   );
   gpc1_1 gpc1516 (
      {stage0_6[475]},
      {stage1_6[206]}
   );
   gpc1_1 gpc1517 (
      {stage0_6[476]},
      {stage1_6[207]}
   );
   gpc1_1 gpc1518 (
      {stage0_6[477]},
      {stage1_6[208]}
   );
   gpc1_1 gpc1519 (
      {stage0_6[478]},
      {stage1_6[209]}
   );
   gpc1_1 gpc1520 (
      {stage0_6[479]},
      {stage1_6[210]}
   );
   gpc1_1 gpc1521 (
      {stage0_6[480]},
      {stage1_6[211]}
   );
   gpc1_1 gpc1522 (
      {stage0_6[481]},
      {stage1_6[212]}
   );
   gpc1_1 gpc1523 (
      {stage0_6[482]},
      {stage1_6[213]}
   );
   gpc1_1 gpc1524 (
      {stage0_6[483]},
      {stage1_6[214]}
   );
   gpc1_1 gpc1525 (
      {stage0_6[484]},
      {stage1_6[215]}
   );
   gpc1_1 gpc1526 (
      {stage0_6[485]},
      {stage1_6[216]}
   );
   gpc1_1 gpc1527 (
      {stage0_6[486]},
      {stage1_6[217]}
   );
   gpc1_1 gpc1528 (
      {stage0_6[487]},
      {stage1_6[218]}
   );
   gpc1_1 gpc1529 (
      {stage0_6[488]},
      {stage1_6[219]}
   );
   gpc1_1 gpc1530 (
      {stage0_6[489]},
      {stage1_6[220]}
   );
   gpc1_1 gpc1531 (
      {stage0_6[490]},
      {stage1_6[221]}
   );
   gpc1_1 gpc1532 (
      {stage0_6[491]},
      {stage1_6[222]}
   );
   gpc1_1 gpc1533 (
      {stage0_6[492]},
      {stage1_6[223]}
   );
   gpc1_1 gpc1534 (
      {stage0_6[493]},
      {stage1_6[224]}
   );
   gpc1_1 gpc1535 (
      {stage0_6[494]},
      {stage1_6[225]}
   );
   gpc1_1 gpc1536 (
      {stage0_6[495]},
      {stage1_6[226]}
   );
   gpc1_1 gpc1537 (
      {stage0_6[496]},
      {stage1_6[227]}
   );
   gpc1_1 gpc1538 (
      {stage0_6[497]},
      {stage1_6[228]}
   );
   gpc1_1 gpc1539 (
      {stage0_6[498]},
      {stage1_6[229]}
   );
   gpc1_1 gpc1540 (
      {stage0_6[499]},
      {stage1_6[230]}
   );
   gpc1_1 gpc1541 (
      {stage0_6[500]},
      {stage1_6[231]}
   );
   gpc1_1 gpc1542 (
      {stage0_6[501]},
      {stage1_6[232]}
   );
   gpc1_1 gpc1543 (
      {stage0_6[502]},
      {stage1_6[233]}
   );
   gpc1_1 gpc1544 (
      {stage0_6[503]},
      {stage1_6[234]}
   );
   gpc1_1 gpc1545 (
      {stage0_6[504]},
      {stage1_6[235]}
   );
   gpc1_1 gpc1546 (
      {stage0_6[505]},
      {stage1_6[236]}
   );
   gpc1_1 gpc1547 (
      {stage0_6[506]},
      {stage1_6[237]}
   );
   gpc1_1 gpc1548 (
      {stage0_6[507]},
      {stage1_6[238]}
   );
   gpc1_1 gpc1549 (
      {stage0_6[508]},
      {stage1_6[239]}
   );
   gpc1_1 gpc1550 (
      {stage0_6[509]},
      {stage1_6[240]}
   );
   gpc1_1 gpc1551 (
      {stage0_6[510]},
      {stage1_6[241]}
   );
   gpc1_1 gpc1552 (
      {stage0_6[511]},
      {stage1_6[242]}
   );
   gpc1_1 gpc1553 (
      {stage0_8[377]},
      {stage1_8[214]}
   );
   gpc1_1 gpc1554 (
      {stage0_8[378]},
      {stage1_8[215]}
   );
   gpc1_1 gpc1555 (
      {stage0_8[379]},
      {stage1_8[216]}
   );
   gpc1_1 gpc1556 (
      {stage0_8[380]},
      {stage1_8[217]}
   );
   gpc1_1 gpc1557 (
      {stage0_8[381]},
      {stage1_8[218]}
   );
   gpc1_1 gpc1558 (
      {stage0_8[382]},
      {stage1_8[219]}
   );
   gpc1_1 gpc1559 (
      {stage0_8[383]},
      {stage1_8[220]}
   );
   gpc1_1 gpc1560 (
      {stage0_8[384]},
      {stage1_8[221]}
   );
   gpc1_1 gpc1561 (
      {stage0_8[385]},
      {stage1_8[222]}
   );
   gpc1_1 gpc1562 (
      {stage0_8[386]},
      {stage1_8[223]}
   );
   gpc1_1 gpc1563 (
      {stage0_8[387]},
      {stage1_8[224]}
   );
   gpc1_1 gpc1564 (
      {stage0_8[388]},
      {stage1_8[225]}
   );
   gpc1_1 gpc1565 (
      {stage0_8[389]},
      {stage1_8[226]}
   );
   gpc1_1 gpc1566 (
      {stage0_8[390]},
      {stage1_8[227]}
   );
   gpc1_1 gpc1567 (
      {stage0_8[391]},
      {stage1_8[228]}
   );
   gpc1_1 gpc1568 (
      {stage0_8[392]},
      {stage1_8[229]}
   );
   gpc1_1 gpc1569 (
      {stage0_8[393]},
      {stage1_8[230]}
   );
   gpc1_1 gpc1570 (
      {stage0_8[394]},
      {stage1_8[231]}
   );
   gpc1_1 gpc1571 (
      {stage0_8[395]},
      {stage1_8[232]}
   );
   gpc1_1 gpc1572 (
      {stage0_8[396]},
      {stage1_8[233]}
   );
   gpc1_1 gpc1573 (
      {stage0_8[397]},
      {stage1_8[234]}
   );
   gpc1_1 gpc1574 (
      {stage0_8[398]},
      {stage1_8[235]}
   );
   gpc1_1 gpc1575 (
      {stage0_8[399]},
      {stage1_8[236]}
   );
   gpc1_1 gpc1576 (
      {stage0_8[400]},
      {stage1_8[237]}
   );
   gpc1_1 gpc1577 (
      {stage0_8[401]},
      {stage1_8[238]}
   );
   gpc1_1 gpc1578 (
      {stage0_8[402]},
      {stage1_8[239]}
   );
   gpc1_1 gpc1579 (
      {stage0_8[403]},
      {stage1_8[240]}
   );
   gpc1_1 gpc1580 (
      {stage0_8[404]},
      {stage1_8[241]}
   );
   gpc1_1 gpc1581 (
      {stage0_8[405]},
      {stage1_8[242]}
   );
   gpc1_1 gpc1582 (
      {stage0_8[406]},
      {stage1_8[243]}
   );
   gpc1_1 gpc1583 (
      {stage0_8[407]},
      {stage1_8[244]}
   );
   gpc1_1 gpc1584 (
      {stage0_8[408]},
      {stage1_8[245]}
   );
   gpc1_1 gpc1585 (
      {stage0_8[409]},
      {stage1_8[246]}
   );
   gpc1_1 gpc1586 (
      {stage0_8[410]},
      {stage1_8[247]}
   );
   gpc1_1 gpc1587 (
      {stage0_8[411]},
      {stage1_8[248]}
   );
   gpc1_1 gpc1588 (
      {stage0_8[412]},
      {stage1_8[249]}
   );
   gpc1_1 gpc1589 (
      {stage0_8[413]},
      {stage1_8[250]}
   );
   gpc1_1 gpc1590 (
      {stage0_8[414]},
      {stage1_8[251]}
   );
   gpc1_1 gpc1591 (
      {stage0_8[415]},
      {stage1_8[252]}
   );
   gpc1_1 gpc1592 (
      {stage0_8[416]},
      {stage1_8[253]}
   );
   gpc1_1 gpc1593 (
      {stage0_8[417]},
      {stage1_8[254]}
   );
   gpc1_1 gpc1594 (
      {stage0_8[418]},
      {stage1_8[255]}
   );
   gpc1_1 gpc1595 (
      {stage0_8[419]},
      {stage1_8[256]}
   );
   gpc1_1 gpc1596 (
      {stage0_8[420]},
      {stage1_8[257]}
   );
   gpc1_1 gpc1597 (
      {stage0_8[421]},
      {stage1_8[258]}
   );
   gpc1_1 gpc1598 (
      {stage0_8[422]},
      {stage1_8[259]}
   );
   gpc1_1 gpc1599 (
      {stage0_8[423]},
      {stage1_8[260]}
   );
   gpc1_1 gpc1600 (
      {stage0_8[424]},
      {stage1_8[261]}
   );
   gpc1_1 gpc1601 (
      {stage0_8[425]},
      {stage1_8[262]}
   );
   gpc1_1 gpc1602 (
      {stage0_8[426]},
      {stage1_8[263]}
   );
   gpc1_1 gpc1603 (
      {stage0_8[427]},
      {stage1_8[264]}
   );
   gpc1_1 gpc1604 (
      {stage0_8[428]},
      {stage1_8[265]}
   );
   gpc1_1 gpc1605 (
      {stage0_8[429]},
      {stage1_8[266]}
   );
   gpc1_1 gpc1606 (
      {stage0_8[430]},
      {stage1_8[267]}
   );
   gpc1_1 gpc1607 (
      {stage0_8[431]},
      {stage1_8[268]}
   );
   gpc1_1 gpc1608 (
      {stage0_8[432]},
      {stage1_8[269]}
   );
   gpc1_1 gpc1609 (
      {stage0_8[433]},
      {stage1_8[270]}
   );
   gpc1_1 gpc1610 (
      {stage0_8[434]},
      {stage1_8[271]}
   );
   gpc1_1 gpc1611 (
      {stage0_8[435]},
      {stage1_8[272]}
   );
   gpc1_1 gpc1612 (
      {stage0_8[436]},
      {stage1_8[273]}
   );
   gpc1_1 gpc1613 (
      {stage0_8[437]},
      {stage1_8[274]}
   );
   gpc1_1 gpc1614 (
      {stage0_8[438]},
      {stage1_8[275]}
   );
   gpc1_1 gpc1615 (
      {stage0_8[439]},
      {stage1_8[276]}
   );
   gpc1_1 gpc1616 (
      {stage0_8[440]},
      {stage1_8[277]}
   );
   gpc1_1 gpc1617 (
      {stage0_8[441]},
      {stage1_8[278]}
   );
   gpc1_1 gpc1618 (
      {stage0_8[442]},
      {stage1_8[279]}
   );
   gpc1_1 gpc1619 (
      {stage0_8[443]},
      {stage1_8[280]}
   );
   gpc1_1 gpc1620 (
      {stage0_8[444]},
      {stage1_8[281]}
   );
   gpc1_1 gpc1621 (
      {stage0_8[445]},
      {stage1_8[282]}
   );
   gpc1_1 gpc1622 (
      {stage0_8[446]},
      {stage1_8[283]}
   );
   gpc1_1 gpc1623 (
      {stage0_8[447]},
      {stage1_8[284]}
   );
   gpc1_1 gpc1624 (
      {stage0_8[448]},
      {stage1_8[285]}
   );
   gpc1_1 gpc1625 (
      {stage0_8[449]},
      {stage1_8[286]}
   );
   gpc1_1 gpc1626 (
      {stage0_8[450]},
      {stage1_8[287]}
   );
   gpc1_1 gpc1627 (
      {stage0_8[451]},
      {stage1_8[288]}
   );
   gpc1_1 gpc1628 (
      {stage0_8[452]},
      {stage1_8[289]}
   );
   gpc1_1 gpc1629 (
      {stage0_8[453]},
      {stage1_8[290]}
   );
   gpc1_1 gpc1630 (
      {stage0_8[454]},
      {stage1_8[291]}
   );
   gpc1_1 gpc1631 (
      {stage0_8[455]},
      {stage1_8[292]}
   );
   gpc1_1 gpc1632 (
      {stage0_8[456]},
      {stage1_8[293]}
   );
   gpc1_1 gpc1633 (
      {stage0_8[457]},
      {stage1_8[294]}
   );
   gpc1_1 gpc1634 (
      {stage0_8[458]},
      {stage1_8[295]}
   );
   gpc1_1 gpc1635 (
      {stage0_8[459]},
      {stage1_8[296]}
   );
   gpc1_1 gpc1636 (
      {stage0_8[460]},
      {stage1_8[297]}
   );
   gpc1_1 gpc1637 (
      {stage0_8[461]},
      {stage1_8[298]}
   );
   gpc1_1 gpc1638 (
      {stage0_8[462]},
      {stage1_8[299]}
   );
   gpc1_1 gpc1639 (
      {stage0_8[463]},
      {stage1_8[300]}
   );
   gpc1_1 gpc1640 (
      {stage0_8[464]},
      {stage1_8[301]}
   );
   gpc1_1 gpc1641 (
      {stage0_8[465]},
      {stage1_8[302]}
   );
   gpc1_1 gpc1642 (
      {stage0_8[466]},
      {stage1_8[303]}
   );
   gpc1_1 gpc1643 (
      {stage0_8[467]},
      {stage1_8[304]}
   );
   gpc1_1 gpc1644 (
      {stage0_8[468]},
      {stage1_8[305]}
   );
   gpc1_1 gpc1645 (
      {stage0_8[469]},
      {stage1_8[306]}
   );
   gpc1_1 gpc1646 (
      {stage0_8[470]},
      {stage1_8[307]}
   );
   gpc1_1 gpc1647 (
      {stage0_8[471]},
      {stage1_8[308]}
   );
   gpc1_1 gpc1648 (
      {stage0_8[472]},
      {stage1_8[309]}
   );
   gpc1_1 gpc1649 (
      {stage0_8[473]},
      {stage1_8[310]}
   );
   gpc1_1 gpc1650 (
      {stage0_8[474]},
      {stage1_8[311]}
   );
   gpc1_1 gpc1651 (
      {stage0_8[475]},
      {stage1_8[312]}
   );
   gpc1_1 gpc1652 (
      {stage0_8[476]},
      {stage1_8[313]}
   );
   gpc1_1 gpc1653 (
      {stage0_8[477]},
      {stage1_8[314]}
   );
   gpc1_1 gpc1654 (
      {stage0_8[478]},
      {stage1_8[315]}
   );
   gpc1_1 gpc1655 (
      {stage0_8[479]},
      {stage1_8[316]}
   );
   gpc1_1 gpc1656 (
      {stage0_8[480]},
      {stage1_8[317]}
   );
   gpc1_1 gpc1657 (
      {stage0_8[481]},
      {stage1_8[318]}
   );
   gpc1_1 gpc1658 (
      {stage0_8[482]},
      {stage1_8[319]}
   );
   gpc1_1 gpc1659 (
      {stage0_8[483]},
      {stage1_8[320]}
   );
   gpc1_1 gpc1660 (
      {stage0_8[484]},
      {stage1_8[321]}
   );
   gpc1_1 gpc1661 (
      {stage0_8[485]},
      {stage1_8[322]}
   );
   gpc1_1 gpc1662 (
      {stage0_8[486]},
      {stage1_8[323]}
   );
   gpc1_1 gpc1663 (
      {stage0_8[487]},
      {stage1_8[324]}
   );
   gpc1_1 gpc1664 (
      {stage0_8[488]},
      {stage1_8[325]}
   );
   gpc1_1 gpc1665 (
      {stage0_8[489]},
      {stage1_8[326]}
   );
   gpc1_1 gpc1666 (
      {stage0_8[490]},
      {stage1_8[327]}
   );
   gpc1_1 gpc1667 (
      {stage0_8[491]},
      {stage1_8[328]}
   );
   gpc1_1 gpc1668 (
      {stage0_8[492]},
      {stage1_8[329]}
   );
   gpc1_1 gpc1669 (
      {stage0_8[493]},
      {stage1_8[330]}
   );
   gpc1_1 gpc1670 (
      {stage0_8[494]},
      {stage1_8[331]}
   );
   gpc1_1 gpc1671 (
      {stage0_8[495]},
      {stage1_8[332]}
   );
   gpc1_1 gpc1672 (
      {stage0_8[496]},
      {stage1_8[333]}
   );
   gpc1_1 gpc1673 (
      {stage0_8[497]},
      {stage1_8[334]}
   );
   gpc1_1 gpc1674 (
      {stage0_8[498]},
      {stage1_8[335]}
   );
   gpc1_1 gpc1675 (
      {stage0_8[499]},
      {stage1_8[336]}
   );
   gpc1_1 gpc1676 (
      {stage0_8[500]},
      {stage1_8[337]}
   );
   gpc1_1 gpc1677 (
      {stage0_8[501]},
      {stage1_8[338]}
   );
   gpc1_1 gpc1678 (
      {stage0_8[502]},
      {stage1_8[339]}
   );
   gpc1_1 gpc1679 (
      {stage0_8[503]},
      {stage1_8[340]}
   );
   gpc1_1 gpc1680 (
      {stage0_8[504]},
      {stage1_8[341]}
   );
   gpc1_1 gpc1681 (
      {stage0_8[505]},
      {stage1_8[342]}
   );
   gpc1_1 gpc1682 (
      {stage0_8[506]},
      {stage1_8[343]}
   );
   gpc1_1 gpc1683 (
      {stage0_8[507]},
      {stage1_8[344]}
   );
   gpc1_1 gpc1684 (
      {stage0_8[508]},
      {stage1_8[345]}
   );
   gpc1_1 gpc1685 (
      {stage0_8[509]},
      {stage1_8[346]}
   );
   gpc1_1 gpc1686 (
      {stage0_8[510]},
      {stage1_8[347]}
   );
   gpc1_1 gpc1687 (
      {stage0_8[511]},
      {stage1_8[348]}
   );
   gpc1_1 gpc1688 (
      {stage0_9[509]},
      {stage1_9[209]}
   );
   gpc1_1 gpc1689 (
      {stage0_9[510]},
      {stage1_9[210]}
   );
   gpc1_1 gpc1690 (
      {stage0_9[511]},
      {stage1_9[211]}
   );
   gpc1_1 gpc1691 (
      {stage0_11[501]},
      {stage1_11[195]}
   );
   gpc1_1 gpc1692 (
      {stage0_11[502]},
      {stage1_11[196]}
   );
   gpc1_1 gpc1693 (
      {stage0_11[503]},
      {stage1_11[197]}
   );
   gpc1_1 gpc1694 (
      {stage0_11[504]},
      {stage1_11[198]}
   );
   gpc1_1 gpc1695 (
      {stage0_11[505]},
      {stage1_11[199]}
   );
   gpc1_1 gpc1696 (
      {stage0_11[506]},
      {stage1_11[200]}
   );
   gpc1_1 gpc1697 (
      {stage0_11[507]},
      {stage1_11[201]}
   );
   gpc1_1 gpc1698 (
      {stage0_11[508]},
      {stage1_11[202]}
   );
   gpc1_1 gpc1699 (
      {stage0_11[509]},
      {stage1_11[203]}
   );
   gpc1_1 gpc1700 (
      {stage0_11[510]},
      {stage1_11[204]}
   );
   gpc1_1 gpc1701 (
      {stage0_11[511]},
      {stage1_11[205]}
   );
   gpc1_1 gpc1702 (
      {stage0_13[507]},
      {stage1_13[227]}
   );
   gpc1_1 gpc1703 (
      {stage0_13[508]},
      {stage1_13[228]}
   );
   gpc1_1 gpc1704 (
      {stage0_13[509]},
      {stage1_13[229]}
   );
   gpc1_1 gpc1705 (
      {stage0_13[510]},
      {stage1_13[230]}
   );
   gpc1_1 gpc1706 (
      {stage0_13[511]},
      {stage1_13[231]}
   );
   gpc1_1 gpc1707 (
      {stage0_14[472]},
      {stage1_14[192]}
   );
   gpc1_1 gpc1708 (
      {stage0_14[473]},
      {stage1_14[193]}
   );
   gpc1_1 gpc1709 (
      {stage0_14[474]},
      {stage1_14[194]}
   );
   gpc1_1 gpc1710 (
      {stage0_14[475]},
      {stage1_14[195]}
   );
   gpc1_1 gpc1711 (
      {stage0_14[476]},
      {stage1_14[196]}
   );
   gpc1_1 gpc1712 (
      {stage0_14[477]},
      {stage1_14[197]}
   );
   gpc1_1 gpc1713 (
      {stage0_14[478]},
      {stage1_14[198]}
   );
   gpc1_1 gpc1714 (
      {stage0_14[479]},
      {stage1_14[199]}
   );
   gpc1_1 gpc1715 (
      {stage0_14[480]},
      {stage1_14[200]}
   );
   gpc1_1 gpc1716 (
      {stage0_14[481]},
      {stage1_14[201]}
   );
   gpc1_1 gpc1717 (
      {stage0_14[482]},
      {stage1_14[202]}
   );
   gpc1_1 gpc1718 (
      {stage0_14[483]},
      {stage1_14[203]}
   );
   gpc1_1 gpc1719 (
      {stage0_14[484]},
      {stage1_14[204]}
   );
   gpc1_1 gpc1720 (
      {stage0_14[485]},
      {stage1_14[205]}
   );
   gpc1_1 gpc1721 (
      {stage0_14[486]},
      {stage1_14[206]}
   );
   gpc1_1 gpc1722 (
      {stage0_14[487]},
      {stage1_14[207]}
   );
   gpc1_1 gpc1723 (
      {stage0_14[488]},
      {stage1_14[208]}
   );
   gpc1_1 gpc1724 (
      {stage0_14[489]},
      {stage1_14[209]}
   );
   gpc1_1 gpc1725 (
      {stage0_14[490]},
      {stage1_14[210]}
   );
   gpc1_1 gpc1726 (
      {stage0_14[491]},
      {stage1_14[211]}
   );
   gpc1_1 gpc1727 (
      {stage0_14[492]},
      {stage1_14[212]}
   );
   gpc1_1 gpc1728 (
      {stage0_14[493]},
      {stage1_14[213]}
   );
   gpc1_1 gpc1729 (
      {stage0_14[494]},
      {stage1_14[214]}
   );
   gpc1_1 gpc1730 (
      {stage0_14[495]},
      {stage1_14[215]}
   );
   gpc1_1 gpc1731 (
      {stage0_14[496]},
      {stage1_14[216]}
   );
   gpc1_1 gpc1732 (
      {stage0_14[497]},
      {stage1_14[217]}
   );
   gpc1_1 gpc1733 (
      {stage0_14[498]},
      {stage1_14[218]}
   );
   gpc1_1 gpc1734 (
      {stage0_14[499]},
      {stage1_14[219]}
   );
   gpc1_1 gpc1735 (
      {stage0_14[500]},
      {stage1_14[220]}
   );
   gpc1_1 gpc1736 (
      {stage0_14[501]},
      {stage1_14[221]}
   );
   gpc1_1 gpc1737 (
      {stage0_14[502]},
      {stage1_14[222]}
   );
   gpc1_1 gpc1738 (
      {stage0_14[503]},
      {stage1_14[223]}
   );
   gpc1_1 gpc1739 (
      {stage0_14[504]},
      {stage1_14[224]}
   );
   gpc1_1 gpc1740 (
      {stage0_14[505]},
      {stage1_14[225]}
   );
   gpc1_1 gpc1741 (
      {stage0_14[506]},
      {stage1_14[226]}
   );
   gpc1_1 gpc1742 (
      {stage0_14[507]},
      {stage1_14[227]}
   );
   gpc1_1 gpc1743 (
      {stage0_14[508]},
      {stage1_14[228]}
   );
   gpc1_1 gpc1744 (
      {stage0_14[509]},
      {stage1_14[229]}
   );
   gpc1_1 gpc1745 (
      {stage0_14[510]},
      {stage1_14[230]}
   );
   gpc1_1 gpc1746 (
      {stage0_14[511]},
      {stage1_14[231]}
   );
   gpc1_1 gpc1747 (
      {stage0_15[456]},
      {stage1_15[181]}
   );
   gpc1_1 gpc1748 (
      {stage0_15[457]},
      {stage1_15[182]}
   );
   gpc1_1 gpc1749 (
      {stage0_15[458]},
      {stage1_15[183]}
   );
   gpc1_1 gpc1750 (
      {stage0_15[459]},
      {stage1_15[184]}
   );
   gpc1_1 gpc1751 (
      {stage0_15[460]},
      {stage1_15[185]}
   );
   gpc1_1 gpc1752 (
      {stage0_15[461]},
      {stage1_15[186]}
   );
   gpc1_1 gpc1753 (
      {stage0_15[462]},
      {stage1_15[187]}
   );
   gpc1_1 gpc1754 (
      {stage0_15[463]},
      {stage1_15[188]}
   );
   gpc1_1 gpc1755 (
      {stage0_15[464]},
      {stage1_15[189]}
   );
   gpc1_1 gpc1756 (
      {stage0_15[465]},
      {stage1_15[190]}
   );
   gpc1_1 gpc1757 (
      {stage0_15[466]},
      {stage1_15[191]}
   );
   gpc1_1 gpc1758 (
      {stage0_15[467]},
      {stage1_15[192]}
   );
   gpc1_1 gpc1759 (
      {stage0_15[468]},
      {stage1_15[193]}
   );
   gpc1_1 gpc1760 (
      {stage0_15[469]},
      {stage1_15[194]}
   );
   gpc1_1 gpc1761 (
      {stage0_15[470]},
      {stage1_15[195]}
   );
   gpc1_1 gpc1762 (
      {stage0_15[471]},
      {stage1_15[196]}
   );
   gpc1_1 gpc1763 (
      {stage0_15[472]},
      {stage1_15[197]}
   );
   gpc1_1 gpc1764 (
      {stage0_15[473]},
      {stage1_15[198]}
   );
   gpc1_1 gpc1765 (
      {stage0_15[474]},
      {stage1_15[199]}
   );
   gpc1_1 gpc1766 (
      {stage0_15[475]},
      {stage1_15[200]}
   );
   gpc1_1 gpc1767 (
      {stage0_15[476]},
      {stage1_15[201]}
   );
   gpc1_1 gpc1768 (
      {stage0_15[477]},
      {stage1_15[202]}
   );
   gpc1_1 gpc1769 (
      {stage0_15[478]},
      {stage1_15[203]}
   );
   gpc1_1 gpc1770 (
      {stage0_15[479]},
      {stage1_15[204]}
   );
   gpc1_1 gpc1771 (
      {stage0_15[480]},
      {stage1_15[205]}
   );
   gpc1_1 gpc1772 (
      {stage0_15[481]},
      {stage1_15[206]}
   );
   gpc1_1 gpc1773 (
      {stage0_15[482]},
      {stage1_15[207]}
   );
   gpc1_1 gpc1774 (
      {stage0_15[483]},
      {stage1_15[208]}
   );
   gpc1_1 gpc1775 (
      {stage0_15[484]},
      {stage1_15[209]}
   );
   gpc1_1 gpc1776 (
      {stage0_15[485]},
      {stage1_15[210]}
   );
   gpc1_1 gpc1777 (
      {stage0_15[486]},
      {stage1_15[211]}
   );
   gpc1_1 gpc1778 (
      {stage0_15[487]},
      {stage1_15[212]}
   );
   gpc1_1 gpc1779 (
      {stage0_15[488]},
      {stage1_15[213]}
   );
   gpc1_1 gpc1780 (
      {stage0_15[489]},
      {stage1_15[214]}
   );
   gpc1_1 gpc1781 (
      {stage0_15[490]},
      {stage1_15[215]}
   );
   gpc1_1 gpc1782 (
      {stage0_15[491]},
      {stage1_15[216]}
   );
   gpc1_1 gpc1783 (
      {stage0_15[492]},
      {stage1_15[217]}
   );
   gpc1_1 gpc1784 (
      {stage0_15[493]},
      {stage1_15[218]}
   );
   gpc1_1 gpc1785 (
      {stage0_15[494]},
      {stage1_15[219]}
   );
   gpc1_1 gpc1786 (
      {stage0_15[495]},
      {stage1_15[220]}
   );
   gpc1_1 gpc1787 (
      {stage0_15[496]},
      {stage1_15[221]}
   );
   gpc1_1 gpc1788 (
      {stage0_15[497]},
      {stage1_15[222]}
   );
   gpc1_1 gpc1789 (
      {stage0_15[498]},
      {stage1_15[223]}
   );
   gpc1_1 gpc1790 (
      {stage0_15[499]},
      {stage1_15[224]}
   );
   gpc1_1 gpc1791 (
      {stage0_15[500]},
      {stage1_15[225]}
   );
   gpc1_1 gpc1792 (
      {stage0_15[501]},
      {stage1_15[226]}
   );
   gpc1_1 gpc1793 (
      {stage0_15[502]},
      {stage1_15[227]}
   );
   gpc1_1 gpc1794 (
      {stage0_15[503]},
      {stage1_15[228]}
   );
   gpc1_1 gpc1795 (
      {stage0_15[504]},
      {stage1_15[229]}
   );
   gpc1_1 gpc1796 (
      {stage0_15[505]},
      {stage1_15[230]}
   );
   gpc1_1 gpc1797 (
      {stage0_15[506]},
      {stage1_15[231]}
   );
   gpc1_1 gpc1798 (
      {stage0_15[507]},
      {stage1_15[232]}
   );
   gpc1_1 gpc1799 (
      {stage0_15[508]},
      {stage1_15[233]}
   );
   gpc1_1 gpc1800 (
      {stage0_15[509]},
      {stage1_15[234]}
   );
   gpc1_1 gpc1801 (
      {stage0_15[510]},
      {stage1_15[235]}
   );
   gpc1_1 gpc1802 (
      {stage0_15[511]},
      {stage1_15[236]}
   );
   gpc1_1 gpc1803 (
      {stage0_17[510]},
      {stage1_17[222]}
   );
   gpc1_1 gpc1804 (
      {stage0_17[511]},
      {stage1_17[223]}
   );
   gpc1_1 gpc1805 (
      {stage0_18[511]},
      {stage1_18[202]}
   );
   gpc1_1 gpc1806 (
      {stage0_19[431]},
      {stage1_19[182]}
   );
   gpc1_1 gpc1807 (
      {stage0_19[432]},
      {stage1_19[183]}
   );
   gpc1_1 gpc1808 (
      {stage0_19[433]},
      {stage1_19[184]}
   );
   gpc1_1 gpc1809 (
      {stage0_19[434]},
      {stage1_19[185]}
   );
   gpc1_1 gpc1810 (
      {stage0_19[435]},
      {stage1_19[186]}
   );
   gpc1_1 gpc1811 (
      {stage0_19[436]},
      {stage1_19[187]}
   );
   gpc1_1 gpc1812 (
      {stage0_19[437]},
      {stage1_19[188]}
   );
   gpc1_1 gpc1813 (
      {stage0_19[438]},
      {stage1_19[189]}
   );
   gpc1_1 gpc1814 (
      {stage0_19[439]},
      {stage1_19[190]}
   );
   gpc1_1 gpc1815 (
      {stage0_19[440]},
      {stage1_19[191]}
   );
   gpc1_1 gpc1816 (
      {stage0_19[441]},
      {stage1_19[192]}
   );
   gpc1_1 gpc1817 (
      {stage0_19[442]},
      {stage1_19[193]}
   );
   gpc1_1 gpc1818 (
      {stage0_19[443]},
      {stage1_19[194]}
   );
   gpc1_1 gpc1819 (
      {stage0_19[444]},
      {stage1_19[195]}
   );
   gpc1_1 gpc1820 (
      {stage0_19[445]},
      {stage1_19[196]}
   );
   gpc1_1 gpc1821 (
      {stage0_19[446]},
      {stage1_19[197]}
   );
   gpc1_1 gpc1822 (
      {stage0_19[447]},
      {stage1_19[198]}
   );
   gpc1_1 gpc1823 (
      {stage0_19[448]},
      {stage1_19[199]}
   );
   gpc1_1 gpc1824 (
      {stage0_19[449]},
      {stage1_19[200]}
   );
   gpc1_1 gpc1825 (
      {stage0_19[450]},
      {stage1_19[201]}
   );
   gpc1_1 gpc1826 (
      {stage0_19[451]},
      {stage1_19[202]}
   );
   gpc1_1 gpc1827 (
      {stage0_19[452]},
      {stage1_19[203]}
   );
   gpc1_1 gpc1828 (
      {stage0_19[453]},
      {stage1_19[204]}
   );
   gpc1_1 gpc1829 (
      {stage0_19[454]},
      {stage1_19[205]}
   );
   gpc1_1 gpc1830 (
      {stage0_19[455]},
      {stage1_19[206]}
   );
   gpc1_1 gpc1831 (
      {stage0_19[456]},
      {stage1_19[207]}
   );
   gpc1_1 gpc1832 (
      {stage0_19[457]},
      {stage1_19[208]}
   );
   gpc1_1 gpc1833 (
      {stage0_19[458]},
      {stage1_19[209]}
   );
   gpc1_1 gpc1834 (
      {stage0_19[459]},
      {stage1_19[210]}
   );
   gpc1_1 gpc1835 (
      {stage0_19[460]},
      {stage1_19[211]}
   );
   gpc1_1 gpc1836 (
      {stage0_19[461]},
      {stage1_19[212]}
   );
   gpc1_1 gpc1837 (
      {stage0_19[462]},
      {stage1_19[213]}
   );
   gpc1_1 gpc1838 (
      {stage0_19[463]},
      {stage1_19[214]}
   );
   gpc1_1 gpc1839 (
      {stage0_19[464]},
      {stage1_19[215]}
   );
   gpc1_1 gpc1840 (
      {stage0_19[465]},
      {stage1_19[216]}
   );
   gpc1_1 gpc1841 (
      {stage0_19[466]},
      {stage1_19[217]}
   );
   gpc1_1 gpc1842 (
      {stage0_19[467]},
      {stage1_19[218]}
   );
   gpc1_1 gpc1843 (
      {stage0_19[468]},
      {stage1_19[219]}
   );
   gpc1_1 gpc1844 (
      {stage0_19[469]},
      {stage1_19[220]}
   );
   gpc1_1 gpc1845 (
      {stage0_19[470]},
      {stage1_19[221]}
   );
   gpc1_1 gpc1846 (
      {stage0_19[471]},
      {stage1_19[222]}
   );
   gpc1_1 gpc1847 (
      {stage0_19[472]},
      {stage1_19[223]}
   );
   gpc1_1 gpc1848 (
      {stage0_19[473]},
      {stage1_19[224]}
   );
   gpc1_1 gpc1849 (
      {stage0_19[474]},
      {stage1_19[225]}
   );
   gpc1_1 gpc1850 (
      {stage0_19[475]},
      {stage1_19[226]}
   );
   gpc1_1 gpc1851 (
      {stage0_19[476]},
      {stage1_19[227]}
   );
   gpc1_1 gpc1852 (
      {stage0_19[477]},
      {stage1_19[228]}
   );
   gpc1_1 gpc1853 (
      {stage0_19[478]},
      {stage1_19[229]}
   );
   gpc1_1 gpc1854 (
      {stage0_19[479]},
      {stage1_19[230]}
   );
   gpc1_1 gpc1855 (
      {stage0_19[480]},
      {stage1_19[231]}
   );
   gpc1_1 gpc1856 (
      {stage0_19[481]},
      {stage1_19[232]}
   );
   gpc1_1 gpc1857 (
      {stage0_19[482]},
      {stage1_19[233]}
   );
   gpc1_1 gpc1858 (
      {stage0_19[483]},
      {stage1_19[234]}
   );
   gpc1_1 gpc1859 (
      {stage0_19[484]},
      {stage1_19[235]}
   );
   gpc1_1 gpc1860 (
      {stage0_19[485]},
      {stage1_19[236]}
   );
   gpc1_1 gpc1861 (
      {stage0_19[486]},
      {stage1_19[237]}
   );
   gpc1_1 gpc1862 (
      {stage0_19[487]},
      {stage1_19[238]}
   );
   gpc1_1 gpc1863 (
      {stage0_19[488]},
      {stage1_19[239]}
   );
   gpc1_1 gpc1864 (
      {stage0_19[489]},
      {stage1_19[240]}
   );
   gpc1_1 gpc1865 (
      {stage0_19[490]},
      {stage1_19[241]}
   );
   gpc1_1 gpc1866 (
      {stage0_19[491]},
      {stage1_19[242]}
   );
   gpc1_1 gpc1867 (
      {stage0_19[492]},
      {stage1_19[243]}
   );
   gpc1_1 gpc1868 (
      {stage0_19[493]},
      {stage1_19[244]}
   );
   gpc1_1 gpc1869 (
      {stage0_19[494]},
      {stage1_19[245]}
   );
   gpc1_1 gpc1870 (
      {stage0_19[495]},
      {stage1_19[246]}
   );
   gpc1_1 gpc1871 (
      {stage0_19[496]},
      {stage1_19[247]}
   );
   gpc1_1 gpc1872 (
      {stage0_19[497]},
      {stage1_19[248]}
   );
   gpc1_1 gpc1873 (
      {stage0_19[498]},
      {stage1_19[249]}
   );
   gpc1_1 gpc1874 (
      {stage0_19[499]},
      {stage1_19[250]}
   );
   gpc1_1 gpc1875 (
      {stage0_19[500]},
      {stage1_19[251]}
   );
   gpc1_1 gpc1876 (
      {stage0_19[501]},
      {stage1_19[252]}
   );
   gpc1_1 gpc1877 (
      {stage0_19[502]},
      {stage1_19[253]}
   );
   gpc1_1 gpc1878 (
      {stage0_19[503]},
      {stage1_19[254]}
   );
   gpc1_1 gpc1879 (
      {stage0_19[504]},
      {stage1_19[255]}
   );
   gpc1_1 gpc1880 (
      {stage0_19[505]},
      {stage1_19[256]}
   );
   gpc1_1 gpc1881 (
      {stage0_19[506]},
      {stage1_19[257]}
   );
   gpc1_1 gpc1882 (
      {stage0_19[507]},
      {stage1_19[258]}
   );
   gpc1_1 gpc1883 (
      {stage0_19[508]},
      {stage1_19[259]}
   );
   gpc1_1 gpc1884 (
      {stage0_19[509]},
      {stage1_19[260]}
   );
   gpc1_1 gpc1885 (
      {stage0_19[510]},
      {stage1_19[261]}
   );
   gpc1_1 gpc1886 (
      {stage0_19[511]},
      {stage1_19[262]}
   );
   gpc1_1 gpc1887 (
      {stage0_20[504]},
      {stage1_20[206]}
   );
   gpc1_1 gpc1888 (
      {stage0_20[505]},
      {stage1_20[207]}
   );
   gpc1_1 gpc1889 (
      {stage0_20[506]},
      {stage1_20[208]}
   );
   gpc1_1 gpc1890 (
      {stage0_20[507]},
      {stage1_20[209]}
   );
   gpc1_1 gpc1891 (
      {stage0_20[508]},
      {stage1_20[210]}
   );
   gpc1_1 gpc1892 (
      {stage0_20[509]},
      {stage1_20[211]}
   );
   gpc1_1 gpc1893 (
      {stage0_20[510]},
      {stage1_20[212]}
   );
   gpc1_1 gpc1894 (
      {stage0_20[511]},
      {stage1_20[213]}
   );
   gpc1_1 gpc1895 (
      {stage0_21[471]},
      {stage1_21[229]}
   );
   gpc1_1 gpc1896 (
      {stage0_21[472]},
      {stage1_21[230]}
   );
   gpc1_1 gpc1897 (
      {stage0_21[473]},
      {stage1_21[231]}
   );
   gpc1_1 gpc1898 (
      {stage0_21[474]},
      {stage1_21[232]}
   );
   gpc1_1 gpc1899 (
      {stage0_21[475]},
      {stage1_21[233]}
   );
   gpc1_1 gpc1900 (
      {stage0_21[476]},
      {stage1_21[234]}
   );
   gpc1_1 gpc1901 (
      {stage0_21[477]},
      {stage1_21[235]}
   );
   gpc1_1 gpc1902 (
      {stage0_21[478]},
      {stage1_21[236]}
   );
   gpc1_1 gpc1903 (
      {stage0_21[479]},
      {stage1_21[237]}
   );
   gpc1_1 gpc1904 (
      {stage0_21[480]},
      {stage1_21[238]}
   );
   gpc1_1 gpc1905 (
      {stage0_21[481]},
      {stage1_21[239]}
   );
   gpc1_1 gpc1906 (
      {stage0_21[482]},
      {stage1_21[240]}
   );
   gpc1_1 gpc1907 (
      {stage0_21[483]},
      {stage1_21[241]}
   );
   gpc1_1 gpc1908 (
      {stage0_21[484]},
      {stage1_21[242]}
   );
   gpc1_1 gpc1909 (
      {stage0_21[485]},
      {stage1_21[243]}
   );
   gpc1_1 gpc1910 (
      {stage0_21[486]},
      {stage1_21[244]}
   );
   gpc1_1 gpc1911 (
      {stage0_21[487]},
      {stage1_21[245]}
   );
   gpc1_1 gpc1912 (
      {stage0_21[488]},
      {stage1_21[246]}
   );
   gpc1_1 gpc1913 (
      {stage0_21[489]},
      {stage1_21[247]}
   );
   gpc1_1 gpc1914 (
      {stage0_21[490]},
      {stage1_21[248]}
   );
   gpc1_1 gpc1915 (
      {stage0_21[491]},
      {stage1_21[249]}
   );
   gpc1_1 gpc1916 (
      {stage0_21[492]},
      {stage1_21[250]}
   );
   gpc1_1 gpc1917 (
      {stage0_21[493]},
      {stage1_21[251]}
   );
   gpc1_1 gpc1918 (
      {stage0_21[494]},
      {stage1_21[252]}
   );
   gpc1_1 gpc1919 (
      {stage0_21[495]},
      {stage1_21[253]}
   );
   gpc1_1 gpc1920 (
      {stage0_21[496]},
      {stage1_21[254]}
   );
   gpc1_1 gpc1921 (
      {stage0_21[497]},
      {stage1_21[255]}
   );
   gpc1_1 gpc1922 (
      {stage0_21[498]},
      {stage1_21[256]}
   );
   gpc1_1 gpc1923 (
      {stage0_21[499]},
      {stage1_21[257]}
   );
   gpc1_1 gpc1924 (
      {stage0_21[500]},
      {stage1_21[258]}
   );
   gpc1_1 gpc1925 (
      {stage0_21[501]},
      {stage1_21[259]}
   );
   gpc1_1 gpc1926 (
      {stage0_21[502]},
      {stage1_21[260]}
   );
   gpc1_1 gpc1927 (
      {stage0_21[503]},
      {stage1_21[261]}
   );
   gpc1_1 gpc1928 (
      {stage0_21[504]},
      {stage1_21[262]}
   );
   gpc1_1 gpc1929 (
      {stage0_21[505]},
      {stage1_21[263]}
   );
   gpc1_1 gpc1930 (
      {stage0_21[506]},
      {stage1_21[264]}
   );
   gpc1_1 gpc1931 (
      {stage0_21[507]},
      {stage1_21[265]}
   );
   gpc1_1 gpc1932 (
      {stage0_21[508]},
      {stage1_21[266]}
   );
   gpc1_1 gpc1933 (
      {stage0_21[509]},
      {stage1_21[267]}
   );
   gpc1_1 gpc1934 (
      {stage0_21[510]},
      {stage1_21[268]}
   );
   gpc1_1 gpc1935 (
      {stage0_21[511]},
      {stage1_21[269]}
   );
   gpc1_1 gpc1936 (
      {stage0_22[423]},
      {stage1_22[185]}
   );
   gpc1_1 gpc1937 (
      {stage0_22[424]},
      {stage1_22[186]}
   );
   gpc1_1 gpc1938 (
      {stage0_22[425]},
      {stage1_22[187]}
   );
   gpc1_1 gpc1939 (
      {stage0_22[426]},
      {stage1_22[188]}
   );
   gpc1_1 gpc1940 (
      {stage0_22[427]},
      {stage1_22[189]}
   );
   gpc1_1 gpc1941 (
      {stage0_22[428]},
      {stage1_22[190]}
   );
   gpc1_1 gpc1942 (
      {stage0_22[429]},
      {stage1_22[191]}
   );
   gpc1_1 gpc1943 (
      {stage0_22[430]},
      {stage1_22[192]}
   );
   gpc1_1 gpc1944 (
      {stage0_22[431]},
      {stage1_22[193]}
   );
   gpc1_1 gpc1945 (
      {stage0_22[432]},
      {stage1_22[194]}
   );
   gpc1_1 gpc1946 (
      {stage0_22[433]},
      {stage1_22[195]}
   );
   gpc1_1 gpc1947 (
      {stage0_22[434]},
      {stage1_22[196]}
   );
   gpc1_1 gpc1948 (
      {stage0_22[435]},
      {stage1_22[197]}
   );
   gpc1_1 gpc1949 (
      {stage0_22[436]},
      {stage1_22[198]}
   );
   gpc1_1 gpc1950 (
      {stage0_22[437]},
      {stage1_22[199]}
   );
   gpc1_1 gpc1951 (
      {stage0_22[438]},
      {stage1_22[200]}
   );
   gpc1_1 gpc1952 (
      {stage0_22[439]},
      {stage1_22[201]}
   );
   gpc1_1 gpc1953 (
      {stage0_22[440]},
      {stage1_22[202]}
   );
   gpc1_1 gpc1954 (
      {stage0_22[441]},
      {stage1_22[203]}
   );
   gpc1_1 gpc1955 (
      {stage0_22[442]},
      {stage1_22[204]}
   );
   gpc1_1 gpc1956 (
      {stage0_22[443]},
      {stage1_22[205]}
   );
   gpc1_1 gpc1957 (
      {stage0_22[444]},
      {stage1_22[206]}
   );
   gpc1_1 gpc1958 (
      {stage0_22[445]},
      {stage1_22[207]}
   );
   gpc1_1 gpc1959 (
      {stage0_22[446]},
      {stage1_22[208]}
   );
   gpc1_1 gpc1960 (
      {stage0_22[447]},
      {stage1_22[209]}
   );
   gpc1_1 gpc1961 (
      {stage0_22[448]},
      {stage1_22[210]}
   );
   gpc1_1 gpc1962 (
      {stage0_22[449]},
      {stage1_22[211]}
   );
   gpc1_1 gpc1963 (
      {stage0_22[450]},
      {stage1_22[212]}
   );
   gpc1_1 gpc1964 (
      {stage0_22[451]},
      {stage1_22[213]}
   );
   gpc1_1 gpc1965 (
      {stage0_22[452]},
      {stage1_22[214]}
   );
   gpc1_1 gpc1966 (
      {stage0_22[453]},
      {stage1_22[215]}
   );
   gpc1_1 gpc1967 (
      {stage0_22[454]},
      {stage1_22[216]}
   );
   gpc1_1 gpc1968 (
      {stage0_22[455]},
      {stage1_22[217]}
   );
   gpc1_1 gpc1969 (
      {stage0_22[456]},
      {stage1_22[218]}
   );
   gpc1_1 gpc1970 (
      {stage0_22[457]},
      {stage1_22[219]}
   );
   gpc1_1 gpc1971 (
      {stage0_22[458]},
      {stage1_22[220]}
   );
   gpc1_1 gpc1972 (
      {stage0_22[459]},
      {stage1_22[221]}
   );
   gpc1_1 gpc1973 (
      {stage0_22[460]},
      {stage1_22[222]}
   );
   gpc1_1 gpc1974 (
      {stage0_22[461]},
      {stage1_22[223]}
   );
   gpc1_1 gpc1975 (
      {stage0_22[462]},
      {stage1_22[224]}
   );
   gpc1_1 gpc1976 (
      {stage0_22[463]},
      {stage1_22[225]}
   );
   gpc1_1 gpc1977 (
      {stage0_22[464]},
      {stage1_22[226]}
   );
   gpc1_1 gpc1978 (
      {stage0_22[465]},
      {stage1_22[227]}
   );
   gpc1_1 gpc1979 (
      {stage0_22[466]},
      {stage1_22[228]}
   );
   gpc1_1 gpc1980 (
      {stage0_22[467]},
      {stage1_22[229]}
   );
   gpc1_1 gpc1981 (
      {stage0_22[468]},
      {stage1_22[230]}
   );
   gpc1_1 gpc1982 (
      {stage0_22[469]},
      {stage1_22[231]}
   );
   gpc1_1 gpc1983 (
      {stage0_22[470]},
      {stage1_22[232]}
   );
   gpc1_1 gpc1984 (
      {stage0_22[471]},
      {stage1_22[233]}
   );
   gpc1_1 gpc1985 (
      {stage0_22[472]},
      {stage1_22[234]}
   );
   gpc1_1 gpc1986 (
      {stage0_22[473]},
      {stage1_22[235]}
   );
   gpc1_1 gpc1987 (
      {stage0_22[474]},
      {stage1_22[236]}
   );
   gpc1_1 gpc1988 (
      {stage0_22[475]},
      {stage1_22[237]}
   );
   gpc1_1 gpc1989 (
      {stage0_22[476]},
      {stage1_22[238]}
   );
   gpc1_1 gpc1990 (
      {stage0_22[477]},
      {stage1_22[239]}
   );
   gpc1_1 gpc1991 (
      {stage0_22[478]},
      {stage1_22[240]}
   );
   gpc1_1 gpc1992 (
      {stage0_22[479]},
      {stage1_22[241]}
   );
   gpc1_1 gpc1993 (
      {stage0_22[480]},
      {stage1_22[242]}
   );
   gpc1_1 gpc1994 (
      {stage0_22[481]},
      {stage1_22[243]}
   );
   gpc1_1 gpc1995 (
      {stage0_22[482]},
      {stage1_22[244]}
   );
   gpc1_1 gpc1996 (
      {stage0_22[483]},
      {stage1_22[245]}
   );
   gpc1_1 gpc1997 (
      {stage0_22[484]},
      {stage1_22[246]}
   );
   gpc1_1 gpc1998 (
      {stage0_22[485]},
      {stage1_22[247]}
   );
   gpc1_1 gpc1999 (
      {stage0_22[486]},
      {stage1_22[248]}
   );
   gpc1_1 gpc2000 (
      {stage0_22[487]},
      {stage1_22[249]}
   );
   gpc1_1 gpc2001 (
      {stage0_22[488]},
      {stage1_22[250]}
   );
   gpc1_1 gpc2002 (
      {stage0_22[489]},
      {stage1_22[251]}
   );
   gpc1_1 gpc2003 (
      {stage0_22[490]},
      {stage1_22[252]}
   );
   gpc1_1 gpc2004 (
      {stage0_22[491]},
      {stage1_22[253]}
   );
   gpc1_1 gpc2005 (
      {stage0_22[492]},
      {stage1_22[254]}
   );
   gpc1_1 gpc2006 (
      {stage0_22[493]},
      {stage1_22[255]}
   );
   gpc1_1 gpc2007 (
      {stage0_22[494]},
      {stage1_22[256]}
   );
   gpc1_1 gpc2008 (
      {stage0_22[495]},
      {stage1_22[257]}
   );
   gpc1_1 gpc2009 (
      {stage0_22[496]},
      {stage1_22[258]}
   );
   gpc1_1 gpc2010 (
      {stage0_22[497]},
      {stage1_22[259]}
   );
   gpc1_1 gpc2011 (
      {stage0_22[498]},
      {stage1_22[260]}
   );
   gpc1_1 gpc2012 (
      {stage0_22[499]},
      {stage1_22[261]}
   );
   gpc1_1 gpc2013 (
      {stage0_22[500]},
      {stage1_22[262]}
   );
   gpc1_1 gpc2014 (
      {stage0_22[501]},
      {stage1_22[263]}
   );
   gpc1_1 gpc2015 (
      {stage0_22[502]},
      {stage1_22[264]}
   );
   gpc1_1 gpc2016 (
      {stage0_22[503]},
      {stage1_22[265]}
   );
   gpc1_1 gpc2017 (
      {stage0_22[504]},
      {stage1_22[266]}
   );
   gpc1_1 gpc2018 (
      {stage0_22[505]},
      {stage1_22[267]}
   );
   gpc1_1 gpc2019 (
      {stage0_22[506]},
      {stage1_22[268]}
   );
   gpc1_1 gpc2020 (
      {stage0_22[507]},
      {stage1_22[269]}
   );
   gpc1_1 gpc2021 (
      {stage0_22[508]},
      {stage1_22[270]}
   );
   gpc1_1 gpc2022 (
      {stage0_22[509]},
      {stage1_22[271]}
   );
   gpc1_1 gpc2023 (
      {stage0_22[510]},
      {stage1_22[272]}
   );
   gpc1_1 gpc2024 (
      {stage0_22[511]},
      {stage1_22[273]}
   );
   gpc1_1 gpc2025 (
      {stage0_23[500]},
      {stage1_23[154]}
   );
   gpc1_1 gpc2026 (
      {stage0_23[501]},
      {stage1_23[155]}
   );
   gpc1_1 gpc2027 (
      {stage0_23[502]},
      {stage1_23[156]}
   );
   gpc1_1 gpc2028 (
      {stage0_23[503]},
      {stage1_23[157]}
   );
   gpc1_1 gpc2029 (
      {stage0_23[504]},
      {stage1_23[158]}
   );
   gpc1_1 gpc2030 (
      {stage0_23[505]},
      {stage1_23[159]}
   );
   gpc1_1 gpc2031 (
      {stage0_23[506]},
      {stage1_23[160]}
   );
   gpc1_1 gpc2032 (
      {stage0_23[507]},
      {stage1_23[161]}
   );
   gpc1_1 gpc2033 (
      {stage0_23[508]},
      {stage1_23[162]}
   );
   gpc1_1 gpc2034 (
      {stage0_23[509]},
      {stage1_23[163]}
   );
   gpc1_1 gpc2035 (
      {stage0_23[510]},
      {stage1_23[164]}
   );
   gpc1_1 gpc2036 (
      {stage0_23[511]},
      {stage1_23[165]}
   );
   gpc1_1 gpc2037 (
      {stage0_25[482]},
      {stage1_25[244]}
   );
   gpc1_1 gpc2038 (
      {stage0_25[483]},
      {stage1_25[245]}
   );
   gpc1_1 gpc2039 (
      {stage0_25[484]},
      {stage1_25[246]}
   );
   gpc1_1 gpc2040 (
      {stage0_25[485]},
      {stage1_25[247]}
   );
   gpc1_1 gpc2041 (
      {stage0_25[486]},
      {stage1_25[248]}
   );
   gpc1_1 gpc2042 (
      {stage0_25[487]},
      {stage1_25[249]}
   );
   gpc1_1 gpc2043 (
      {stage0_25[488]},
      {stage1_25[250]}
   );
   gpc1_1 gpc2044 (
      {stage0_25[489]},
      {stage1_25[251]}
   );
   gpc1_1 gpc2045 (
      {stage0_25[490]},
      {stage1_25[252]}
   );
   gpc1_1 gpc2046 (
      {stage0_25[491]},
      {stage1_25[253]}
   );
   gpc1_1 gpc2047 (
      {stage0_25[492]},
      {stage1_25[254]}
   );
   gpc1_1 gpc2048 (
      {stage0_25[493]},
      {stage1_25[255]}
   );
   gpc1_1 gpc2049 (
      {stage0_25[494]},
      {stage1_25[256]}
   );
   gpc1_1 gpc2050 (
      {stage0_25[495]},
      {stage1_25[257]}
   );
   gpc1_1 gpc2051 (
      {stage0_25[496]},
      {stage1_25[258]}
   );
   gpc1_1 gpc2052 (
      {stage0_25[497]},
      {stage1_25[259]}
   );
   gpc1_1 gpc2053 (
      {stage0_25[498]},
      {stage1_25[260]}
   );
   gpc1_1 gpc2054 (
      {stage0_25[499]},
      {stage1_25[261]}
   );
   gpc1_1 gpc2055 (
      {stage0_25[500]},
      {stage1_25[262]}
   );
   gpc1_1 gpc2056 (
      {stage0_25[501]},
      {stage1_25[263]}
   );
   gpc1_1 gpc2057 (
      {stage0_25[502]},
      {stage1_25[264]}
   );
   gpc1_1 gpc2058 (
      {stage0_25[503]},
      {stage1_25[265]}
   );
   gpc1_1 gpc2059 (
      {stage0_25[504]},
      {stage1_25[266]}
   );
   gpc1_1 gpc2060 (
      {stage0_25[505]},
      {stage1_25[267]}
   );
   gpc1_1 gpc2061 (
      {stage0_25[506]},
      {stage1_25[268]}
   );
   gpc1_1 gpc2062 (
      {stage0_25[507]},
      {stage1_25[269]}
   );
   gpc1_1 gpc2063 (
      {stage0_25[508]},
      {stage1_25[270]}
   );
   gpc1_1 gpc2064 (
      {stage0_25[509]},
      {stage1_25[271]}
   );
   gpc1_1 gpc2065 (
      {stage0_25[510]},
      {stage1_25[272]}
   );
   gpc1_1 gpc2066 (
      {stage0_25[511]},
      {stage1_25[273]}
   );
   gpc1_1 gpc2067 (
      {stage0_26[498]},
      {stage1_26[177]}
   );
   gpc1_1 gpc2068 (
      {stage0_26[499]},
      {stage1_26[178]}
   );
   gpc1_1 gpc2069 (
      {stage0_26[500]},
      {stage1_26[179]}
   );
   gpc1_1 gpc2070 (
      {stage0_26[501]},
      {stage1_26[180]}
   );
   gpc1_1 gpc2071 (
      {stage0_26[502]},
      {stage1_26[181]}
   );
   gpc1_1 gpc2072 (
      {stage0_26[503]},
      {stage1_26[182]}
   );
   gpc1_1 gpc2073 (
      {stage0_26[504]},
      {stage1_26[183]}
   );
   gpc1_1 gpc2074 (
      {stage0_26[505]},
      {stage1_26[184]}
   );
   gpc1_1 gpc2075 (
      {stage0_26[506]},
      {stage1_26[185]}
   );
   gpc1_1 gpc2076 (
      {stage0_26[507]},
      {stage1_26[186]}
   );
   gpc1_1 gpc2077 (
      {stage0_26[508]},
      {stage1_26[187]}
   );
   gpc1_1 gpc2078 (
      {stage0_26[509]},
      {stage1_26[188]}
   );
   gpc1_1 gpc2079 (
      {stage0_26[510]},
      {stage1_26[189]}
   );
   gpc1_1 gpc2080 (
      {stage0_26[511]},
      {stage1_26[190]}
   );
   gpc1_1 gpc2081 (
      {stage0_27[479]},
      {stage1_27[167]}
   );
   gpc1_1 gpc2082 (
      {stage0_27[480]},
      {stage1_27[168]}
   );
   gpc1_1 gpc2083 (
      {stage0_27[481]},
      {stage1_27[169]}
   );
   gpc1_1 gpc2084 (
      {stage0_27[482]},
      {stage1_27[170]}
   );
   gpc1_1 gpc2085 (
      {stage0_27[483]},
      {stage1_27[171]}
   );
   gpc1_1 gpc2086 (
      {stage0_27[484]},
      {stage1_27[172]}
   );
   gpc1_1 gpc2087 (
      {stage0_27[485]},
      {stage1_27[173]}
   );
   gpc1_1 gpc2088 (
      {stage0_27[486]},
      {stage1_27[174]}
   );
   gpc1_1 gpc2089 (
      {stage0_27[487]},
      {stage1_27[175]}
   );
   gpc1_1 gpc2090 (
      {stage0_27[488]},
      {stage1_27[176]}
   );
   gpc1_1 gpc2091 (
      {stage0_27[489]},
      {stage1_27[177]}
   );
   gpc1_1 gpc2092 (
      {stage0_27[490]},
      {stage1_27[178]}
   );
   gpc1_1 gpc2093 (
      {stage0_27[491]},
      {stage1_27[179]}
   );
   gpc1_1 gpc2094 (
      {stage0_27[492]},
      {stage1_27[180]}
   );
   gpc1_1 gpc2095 (
      {stage0_27[493]},
      {stage1_27[181]}
   );
   gpc1_1 gpc2096 (
      {stage0_27[494]},
      {stage1_27[182]}
   );
   gpc1_1 gpc2097 (
      {stage0_27[495]},
      {stage1_27[183]}
   );
   gpc1_1 gpc2098 (
      {stage0_27[496]},
      {stage1_27[184]}
   );
   gpc1_1 gpc2099 (
      {stage0_27[497]},
      {stage1_27[185]}
   );
   gpc1_1 gpc2100 (
      {stage0_27[498]},
      {stage1_27[186]}
   );
   gpc1_1 gpc2101 (
      {stage0_27[499]},
      {stage1_27[187]}
   );
   gpc1_1 gpc2102 (
      {stage0_27[500]},
      {stage1_27[188]}
   );
   gpc1_1 gpc2103 (
      {stage0_27[501]},
      {stage1_27[189]}
   );
   gpc1_1 gpc2104 (
      {stage0_27[502]},
      {stage1_27[190]}
   );
   gpc1_1 gpc2105 (
      {stage0_27[503]},
      {stage1_27[191]}
   );
   gpc1_1 gpc2106 (
      {stage0_27[504]},
      {stage1_27[192]}
   );
   gpc1_1 gpc2107 (
      {stage0_27[505]},
      {stage1_27[193]}
   );
   gpc1_1 gpc2108 (
      {stage0_27[506]},
      {stage1_27[194]}
   );
   gpc1_1 gpc2109 (
      {stage0_27[507]},
      {stage1_27[195]}
   );
   gpc1_1 gpc2110 (
      {stage0_27[508]},
      {stage1_27[196]}
   );
   gpc1_1 gpc2111 (
      {stage0_27[509]},
      {stage1_27[197]}
   );
   gpc1_1 gpc2112 (
      {stage0_27[510]},
      {stage1_27[198]}
   );
   gpc1_1 gpc2113 (
      {stage0_27[511]},
      {stage1_27[199]}
   );
   gpc1_1 gpc2114 (
      {stage0_28[506]},
      {stage1_28[242]}
   );
   gpc1_1 gpc2115 (
      {stage0_28[507]},
      {stage1_28[243]}
   );
   gpc1_1 gpc2116 (
      {stage0_28[508]},
      {stage1_28[244]}
   );
   gpc1_1 gpc2117 (
      {stage0_28[509]},
      {stage1_28[245]}
   );
   gpc1_1 gpc2118 (
      {stage0_28[510]},
      {stage1_28[246]}
   );
   gpc1_1 gpc2119 (
      {stage0_28[511]},
      {stage1_28[247]}
   );
   gpc1_1 gpc2120 (
      {stage0_29[509]},
      {stage1_29[240]}
   );
   gpc1_1 gpc2121 (
      {stage0_29[510]},
      {stage1_29[241]}
   );
   gpc1_1 gpc2122 (
      {stage0_29[511]},
      {stage1_29[242]}
   );
   gpc1_1 gpc2123 (
      {stage0_30[474]},
      {stage1_30[169]}
   );
   gpc1_1 gpc2124 (
      {stage0_30[475]},
      {stage1_30[170]}
   );
   gpc1_1 gpc2125 (
      {stage0_30[476]},
      {stage1_30[171]}
   );
   gpc1_1 gpc2126 (
      {stage0_30[477]},
      {stage1_30[172]}
   );
   gpc1_1 gpc2127 (
      {stage0_30[478]},
      {stage1_30[173]}
   );
   gpc1_1 gpc2128 (
      {stage0_30[479]},
      {stage1_30[174]}
   );
   gpc1_1 gpc2129 (
      {stage0_30[480]},
      {stage1_30[175]}
   );
   gpc1_1 gpc2130 (
      {stage0_30[481]},
      {stage1_30[176]}
   );
   gpc1_1 gpc2131 (
      {stage0_30[482]},
      {stage1_30[177]}
   );
   gpc1_1 gpc2132 (
      {stage0_30[483]},
      {stage1_30[178]}
   );
   gpc1_1 gpc2133 (
      {stage0_30[484]},
      {stage1_30[179]}
   );
   gpc1_1 gpc2134 (
      {stage0_30[485]},
      {stage1_30[180]}
   );
   gpc1_1 gpc2135 (
      {stage0_30[486]},
      {stage1_30[181]}
   );
   gpc1_1 gpc2136 (
      {stage0_30[487]},
      {stage1_30[182]}
   );
   gpc1_1 gpc2137 (
      {stage0_30[488]},
      {stage1_30[183]}
   );
   gpc1_1 gpc2138 (
      {stage0_30[489]},
      {stage1_30[184]}
   );
   gpc1_1 gpc2139 (
      {stage0_30[490]},
      {stage1_30[185]}
   );
   gpc1_1 gpc2140 (
      {stage0_30[491]},
      {stage1_30[186]}
   );
   gpc1_1 gpc2141 (
      {stage0_30[492]},
      {stage1_30[187]}
   );
   gpc1_1 gpc2142 (
      {stage0_30[493]},
      {stage1_30[188]}
   );
   gpc1_1 gpc2143 (
      {stage0_30[494]},
      {stage1_30[189]}
   );
   gpc1_1 gpc2144 (
      {stage0_30[495]},
      {stage1_30[190]}
   );
   gpc1_1 gpc2145 (
      {stage0_30[496]},
      {stage1_30[191]}
   );
   gpc1_1 gpc2146 (
      {stage0_30[497]},
      {stage1_30[192]}
   );
   gpc1_1 gpc2147 (
      {stage0_30[498]},
      {stage1_30[193]}
   );
   gpc1_1 gpc2148 (
      {stage0_30[499]},
      {stage1_30[194]}
   );
   gpc1_1 gpc2149 (
      {stage0_30[500]},
      {stage1_30[195]}
   );
   gpc1_1 gpc2150 (
      {stage0_30[501]},
      {stage1_30[196]}
   );
   gpc1_1 gpc2151 (
      {stage0_30[502]},
      {stage1_30[197]}
   );
   gpc1_1 gpc2152 (
      {stage0_30[503]},
      {stage1_30[198]}
   );
   gpc1_1 gpc2153 (
      {stage0_30[504]},
      {stage1_30[199]}
   );
   gpc1_1 gpc2154 (
      {stage0_30[505]},
      {stage1_30[200]}
   );
   gpc1_1 gpc2155 (
      {stage0_30[506]},
      {stage1_30[201]}
   );
   gpc1_1 gpc2156 (
      {stage0_30[507]},
      {stage1_30[202]}
   );
   gpc1_1 gpc2157 (
      {stage0_30[508]},
      {stage1_30[203]}
   );
   gpc1_1 gpc2158 (
      {stage0_30[509]},
      {stage1_30[204]}
   );
   gpc1_1 gpc2159 (
      {stage0_30[510]},
      {stage1_30[205]}
   );
   gpc1_1 gpc2160 (
      {stage0_30[511]},
      {stage1_30[206]}
   );
   gpc1_1 gpc2161 (
      {stage0_31[426]},
      {stage1_31[157]}
   );
   gpc1_1 gpc2162 (
      {stage0_31[427]},
      {stage1_31[158]}
   );
   gpc1_1 gpc2163 (
      {stage0_31[428]},
      {stage1_31[159]}
   );
   gpc1_1 gpc2164 (
      {stage0_31[429]},
      {stage1_31[160]}
   );
   gpc1_1 gpc2165 (
      {stage0_31[430]},
      {stage1_31[161]}
   );
   gpc1_1 gpc2166 (
      {stage0_31[431]},
      {stage1_31[162]}
   );
   gpc1_1 gpc2167 (
      {stage0_31[432]},
      {stage1_31[163]}
   );
   gpc1_1 gpc2168 (
      {stage0_31[433]},
      {stage1_31[164]}
   );
   gpc1_1 gpc2169 (
      {stage0_31[434]},
      {stage1_31[165]}
   );
   gpc1_1 gpc2170 (
      {stage0_31[435]},
      {stage1_31[166]}
   );
   gpc1_1 gpc2171 (
      {stage0_31[436]},
      {stage1_31[167]}
   );
   gpc1_1 gpc2172 (
      {stage0_31[437]},
      {stage1_31[168]}
   );
   gpc1_1 gpc2173 (
      {stage0_31[438]},
      {stage1_31[169]}
   );
   gpc1_1 gpc2174 (
      {stage0_31[439]},
      {stage1_31[170]}
   );
   gpc1_1 gpc2175 (
      {stage0_31[440]},
      {stage1_31[171]}
   );
   gpc1_1 gpc2176 (
      {stage0_31[441]},
      {stage1_31[172]}
   );
   gpc1_1 gpc2177 (
      {stage0_31[442]},
      {stage1_31[173]}
   );
   gpc1_1 gpc2178 (
      {stage0_31[443]},
      {stage1_31[174]}
   );
   gpc1_1 gpc2179 (
      {stage0_31[444]},
      {stage1_31[175]}
   );
   gpc1_1 gpc2180 (
      {stage0_31[445]},
      {stage1_31[176]}
   );
   gpc1_1 gpc2181 (
      {stage0_31[446]},
      {stage1_31[177]}
   );
   gpc1_1 gpc2182 (
      {stage0_31[447]},
      {stage1_31[178]}
   );
   gpc1_1 gpc2183 (
      {stage0_31[448]},
      {stage1_31[179]}
   );
   gpc1_1 gpc2184 (
      {stage0_31[449]},
      {stage1_31[180]}
   );
   gpc1_1 gpc2185 (
      {stage0_31[450]},
      {stage1_31[181]}
   );
   gpc1_1 gpc2186 (
      {stage0_31[451]},
      {stage1_31[182]}
   );
   gpc1_1 gpc2187 (
      {stage0_31[452]},
      {stage1_31[183]}
   );
   gpc1_1 gpc2188 (
      {stage0_31[453]},
      {stage1_31[184]}
   );
   gpc1_1 gpc2189 (
      {stage0_31[454]},
      {stage1_31[185]}
   );
   gpc1_1 gpc2190 (
      {stage0_31[455]},
      {stage1_31[186]}
   );
   gpc1_1 gpc2191 (
      {stage0_31[456]},
      {stage1_31[187]}
   );
   gpc1_1 gpc2192 (
      {stage0_31[457]},
      {stage1_31[188]}
   );
   gpc1_1 gpc2193 (
      {stage0_31[458]},
      {stage1_31[189]}
   );
   gpc1_1 gpc2194 (
      {stage0_31[459]},
      {stage1_31[190]}
   );
   gpc1_1 gpc2195 (
      {stage0_31[460]},
      {stage1_31[191]}
   );
   gpc1_1 gpc2196 (
      {stage0_31[461]},
      {stage1_31[192]}
   );
   gpc1_1 gpc2197 (
      {stage0_31[462]},
      {stage1_31[193]}
   );
   gpc1_1 gpc2198 (
      {stage0_31[463]},
      {stage1_31[194]}
   );
   gpc1_1 gpc2199 (
      {stage0_31[464]},
      {stage1_31[195]}
   );
   gpc1_1 gpc2200 (
      {stage0_31[465]},
      {stage1_31[196]}
   );
   gpc1_1 gpc2201 (
      {stage0_31[466]},
      {stage1_31[197]}
   );
   gpc1_1 gpc2202 (
      {stage0_31[467]},
      {stage1_31[198]}
   );
   gpc1_1 gpc2203 (
      {stage0_31[468]},
      {stage1_31[199]}
   );
   gpc1_1 gpc2204 (
      {stage0_31[469]},
      {stage1_31[200]}
   );
   gpc1_1 gpc2205 (
      {stage0_31[470]},
      {stage1_31[201]}
   );
   gpc1_1 gpc2206 (
      {stage0_31[471]},
      {stage1_31[202]}
   );
   gpc1_1 gpc2207 (
      {stage0_31[472]},
      {stage1_31[203]}
   );
   gpc1_1 gpc2208 (
      {stage0_31[473]},
      {stage1_31[204]}
   );
   gpc1_1 gpc2209 (
      {stage0_31[474]},
      {stage1_31[205]}
   );
   gpc1_1 gpc2210 (
      {stage0_31[475]},
      {stage1_31[206]}
   );
   gpc1_1 gpc2211 (
      {stage0_31[476]},
      {stage1_31[207]}
   );
   gpc1_1 gpc2212 (
      {stage0_31[477]},
      {stage1_31[208]}
   );
   gpc1_1 gpc2213 (
      {stage0_31[478]},
      {stage1_31[209]}
   );
   gpc1_1 gpc2214 (
      {stage0_31[479]},
      {stage1_31[210]}
   );
   gpc1_1 gpc2215 (
      {stage0_31[480]},
      {stage1_31[211]}
   );
   gpc1_1 gpc2216 (
      {stage0_31[481]},
      {stage1_31[212]}
   );
   gpc1_1 gpc2217 (
      {stage0_31[482]},
      {stage1_31[213]}
   );
   gpc1_1 gpc2218 (
      {stage0_31[483]},
      {stage1_31[214]}
   );
   gpc1_1 gpc2219 (
      {stage0_31[484]},
      {stage1_31[215]}
   );
   gpc1_1 gpc2220 (
      {stage0_31[485]},
      {stage1_31[216]}
   );
   gpc1_1 gpc2221 (
      {stage0_31[486]},
      {stage1_31[217]}
   );
   gpc1_1 gpc2222 (
      {stage0_31[487]},
      {stage1_31[218]}
   );
   gpc1_1 gpc2223 (
      {stage0_31[488]},
      {stage1_31[219]}
   );
   gpc1_1 gpc2224 (
      {stage0_31[489]},
      {stage1_31[220]}
   );
   gpc1_1 gpc2225 (
      {stage0_31[490]},
      {stage1_31[221]}
   );
   gpc1_1 gpc2226 (
      {stage0_31[491]},
      {stage1_31[222]}
   );
   gpc1_1 gpc2227 (
      {stage0_31[492]},
      {stage1_31[223]}
   );
   gpc1_1 gpc2228 (
      {stage0_31[493]},
      {stage1_31[224]}
   );
   gpc1_1 gpc2229 (
      {stage0_31[494]},
      {stage1_31[225]}
   );
   gpc1_1 gpc2230 (
      {stage0_31[495]},
      {stage1_31[226]}
   );
   gpc1_1 gpc2231 (
      {stage0_31[496]},
      {stage1_31[227]}
   );
   gpc1_1 gpc2232 (
      {stage0_31[497]},
      {stage1_31[228]}
   );
   gpc1_1 gpc2233 (
      {stage0_31[498]},
      {stage1_31[229]}
   );
   gpc1_1 gpc2234 (
      {stage0_31[499]},
      {stage1_31[230]}
   );
   gpc1_1 gpc2235 (
      {stage0_31[500]},
      {stage1_31[231]}
   );
   gpc1_1 gpc2236 (
      {stage0_31[501]},
      {stage1_31[232]}
   );
   gpc1_1 gpc2237 (
      {stage0_31[502]},
      {stage1_31[233]}
   );
   gpc1_1 gpc2238 (
      {stage0_31[503]},
      {stage1_31[234]}
   );
   gpc1_1 gpc2239 (
      {stage0_31[504]},
      {stage1_31[235]}
   );
   gpc1_1 gpc2240 (
      {stage0_31[505]},
      {stage1_31[236]}
   );
   gpc1_1 gpc2241 (
      {stage0_31[506]},
      {stage1_31[237]}
   );
   gpc1_1 gpc2242 (
      {stage0_31[507]},
      {stage1_31[238]}
   );
   gpc1_1 gpc2243 (
      {stage0_31[508]},
      {stage1_31[239]}
   );
   gpc1_1 gpc2244 (
      {stage0_31[509]},
      {stage1_31[240]}
   );
   gpc1_1 gpc2245 (
      {stage0_31[510]},
      {stage1_31[241]}
   );
   gpc1_1 gpc2246 (
      {stage0_31[511]},
      {stage1_31[242]}
   );
   gpc2135_5 gpc2247 (
      {stage1_0[0], stage1_0[1], stage1_0[2], stage1_0[3], stage1_0[4]},
      {stage1_1[0], stage1_1[1], stage1_1[2]},
      {stage1_2[0]},
      {stage1_3[0], stage1_3[1]},
      {stage2_4[0],stage2_3[0],stage2_2[0],stage2_1[0],stage2_0[0]}
   );
   gpc2135_5 gpc2248 (
      {stage1_0[5], stage1_0[6], stage1_0[7], stage1_0[8], stage1_0[9]},
      {stage1_1[3], stage1_1[4], stage1_1[5]},
      {stage1_2[1]},
      {stage1_3[2], stage1_3[3]},
      {stage2_4[1],stage2_3[1],stage2_2[1],stage2_1[1],stage2_0[1]}
   );
   gpc2135_5 gpc2249 (
      {stage1_0[10], stage1_0[11], stage1_0[12], stage1_0[13], stage1_0[14]},
      {stage1_1[6], stage1_1[7], stage1_1[8]},
      {stage1_2[2]},
      {stage1_3[4], stage1_3[5]},
      {stage2_4[2],stage2_3[2],stage2_2[2],stage2_1[2],stage2_0[2]}
   );
   gpc2135_5 gpc2250 (
      {stage1_0[15], stage1_0[16], stage1_0[17], stage1_0[18], stage1_0[19]},
      {stage1_1[9], stage1_1[10], stage1_1[11]},
      {stage1_2[3]},
      {stage1_3[6], stage1_3[7]},
      {stage2_4[3],stage2_3[3],stage2_2[3],stage2_1[3],stage2_0[3]}
   );
   gpc615_5 gpc2251 (
      {stage1_0[20], stage1_0[21], stage1_0[22], stage1_0[23], stage1_0[24]},
      {stage1_1[12]},
      {stage1_2[4], stage1_2[5], stage1_2[6], stage1_2[7], stage1_2[8], stage1_2[9]},
      {stage2_4[4],stage2_3[4],stage2_2[4],stage2_1[4],stage2_0[4]}
   );
   gpc615_5 gpc2252 (
      {stage1_0[25], stage1_0[26], stage1_0[27], stage1_0[28], stage1_0[29]},
      {stage1_1[13]},
      {stage1_2[10], stage1_2[11], stage1_2[12], stage1_2[13], stage1_2[14], stage1_2[15]},
      {stage2_4[5],stage2_3[5],stage2_2[5],stage2_1[5],stage2_0[5]}
   );
   gpc615_5 gpc2253 (
      {stage1_0[30], stage1_0[31], stage1_0[32], stage1_0[33], stage1_0[34]},
      {stage1_1[14]},
      {stage1_2[16], stage1_2[17], stage1_2[18], stage1_2[19], stage1_2[20], stage1_2[21]},
      {stage2_4[6],stage2_3[6],stage2_2[6],stage2_1[6],stage2_0[6]}
   );
   gpc615_5 gpc2254 (
      {stage1_0[35], stage1_0[36], stage1_0[37], stage1_0[38], stage1_0[39]},
      {stage1_1[15]},
      {stage1_2[22], stage1_2[23], stage1_2[24], stage1_2[25], stage1_2[26], stage1_2[27]},
      {stage2_4[7],stage2_3[7],stage2_2[7],stage2_1[7],stage2_0[7]}
   );
   gpc615_5 gpc2255 (
      {stage1_0[40], stage1_0[41], stage1_0[42], stage1_0[43], stage1_0[44]},
      {stage1_1[16]},
      {stage1_2[28], stage1_2[29], stage1_2[30], stage1_2[31], stage1_2[32], stage1_2[33]},
      {stage2_4[8],stage2_3[8],stage2_2[8],stage2_1[8],stage2_0[8]}
   );
   gpc615_5 gpc2256 (
      {stage1_0[45], stage1_0[46], stage1_0[47], stage1_0[48], stage1_0[49]},
      {stage1_1[17]},
      {stage1_2[34], stage1_2[35], stage1_2[36], stage1_2[37], stage1_2[38], stage1_2[39]},
      {stage2_4[9],stage2_3[9],stage2_2[9],stage2_1[9],stage2_0[9]}
   );
   gpc615_5 gpc2257 (
      {stage1_0[50], stage1_0[51], stage1_0[52], stage1_0[53], stage1_0[54]},
      {stage1_1[18]},
      {stage1_2[40], stage1_2[41], stage1_2[42], stage1_2[43], stage1_2[44], stage1_2[45]},
      {stage2_4[10],stage2_3[10],stage2_2[10],stage2_1[10],stage2_0[10]}
   );
   gpc615_5 gpc2258 (
      {stage1_0[55], stage1_0[56], stage1_0[57], stage1_0[58], stage1_0[59]},
      {stage1_1[19]},
      {stage1_2[46], stage1_2[47], stage1_2[48], stage1_2[49], stage1_2[50], stage1_2[51]},
      {stage2_4[11],stage2_3[11],stage2_2[11],stage2_1[11],stage2_0[11]}
   );
   gpc606_5 gpc2259 (
      {stage1_1[20], stage1_1[21], stage1_1[22], stage1_1[23], stage1_1[24], stage1_1[25]},
      {stage1_3[8], stage1_3[9], stage1_3[10], stage1_3[11], stage1_3[12], stage1_3[13]},
      {stage2_5[0],stage2_4[12],stage2_3[12],stage2_2[12],stage2_1[12]}
   );
   gpc606_5 gpc2260 (
      {stage1_1[26], stage1_1[27], stage1_1[28], stage1_1[29], stage1_1[30], stage1_1[31]},
      {stage1_3[14], stage1_3[15], stage1_3[16], stage1_3[17], stage1_3[18], stage1_3[19]},
      {stage2_5[1],stage2_4[13],stage2_3[13],stage2_2[13],stage2_1[13]}
   );
   gpc606_5 gpc2261 (
      {stage1_1[32], stage1_1[33], stage1_1[34], stage1_1[35], stage1_1[36], stage1_1[37]},
      {stage1_3[20], stage1_3[21], stage1_3[22], stage1_3[23], stage1_3[24], stage1_3[25]},
      {stage2_5[2],stage2_4[14],stage2_3[14],stage2_2[14],stage2_1[14]}
   );
   gpc606_5 gpc2262 (
      {stage1_1[38], stage1_1[39], stage1_1[40], stage1_1[41], stage1_1[42], stage1_1[43]},
      {stage1_3[26], stage1_3[27], stage1_3[28], stage1_3[29], stage1_3[30], stage1_3[31]},
      {stage2_5[3],stage2_4[15],stage2_3[15],stage2_2[15],stage2_1[15]}
   );
   gpc606_5 gpc2263 (
      {stage1_1[44], stage1_1[45], stage1_1[46], stage1_1[47], stage1_1[48], stage1_1[49]},
      {stage1_3[32], stage1_3[33], stage1_3[34], stage1_3[35], stage1_3[36], stage1_3[37]},
      {stage2_5[4],stage2_4[16],stage2_3[16],stage2_2[16],stage2_1[16]}
   );
   gpc606_5 gpc2264 (
      {stage1_1[50], stage1_1[51], stage1_1[52], stage1_1[53], stage1_1[54], stage1_1[55]},
      {stage1_3[38], stage1_3[39], stage1_3[40], stage1_3[41], stage1_3[42], stage1_3[43]},
      {stage2_5[5],stage2_4[17],stage2_3[17],stage2_2[17],stage2_1[17]}
   );
   gpc606_5 gpc2265 (
      {stage1_1[56], stage1_1[57], stage1_1[58], stage1_1[59], stage1_1[60], stage1_1[61]},
      {stage1_3[44], stage1_3[45], stage1_3[46], stage1_3[47], stage1_3[48], stage1_3[49]},
      {stage2_5[6],stage2_4[18],stage2_3[18],stage2_2[18],stage2_1[18]}
   );
   gpc606_5 gpc2266 (
      {stage1_1[62], stage1_1[63], stage1_1[64], stage1_1[65], stage1_1[66], stage1_1[67]},
      {stage1_3[50], stage1_3[51], stage1_3[52], stage1_3[53], stage1_3[54], stage1_3[55]},
      {stage2_5[7],stage2_4[19],stage2_3[19],stage2_2[19],stage2_1[19]}
   );
   gpc606_5 gpc2267 (
      {stage1_1[68], stage1_1[69], stage1_1[70], stage1_1[71], stage1_1[72], stage1_1[73]},
      {stage1_3[56], stage1_3[57], stage1_3[58], stage1_3[59], stage1_3[60], stage1_3[61]},
      {stage2_5[8],stage2_4[20],stage2_3[20],stage2_2[20],stage2_1[20]}
   );
   gpc606_5 gpc2268 (
      {stage1_1[74], stage1_1[75], stage1_1[76], stage1_1[77], stage1_1[78], stage1_1[79]},
      {stage1_3[62], stage1_3[63], stage1_3[64], stage1_3[65], stage1_3[66], stage1_3[67]},
      {stage2_5[9],stage2_4[21],stage2_3[21],stage2_2[21],stage2_1[21]}
   );
   gpc606_5 gpc2269 (
      {stage1_1[80], stage1_1[81], stage1_1[82], stage1_1[83], stage1_1[84], stage1_1[85]},
      {stage1_3[68], stage1_3[69], stage1_3[70], stage1_3[71], stage1_3[72], stage1_3[73]},
      {stage2_5[10],stage2_4[22],stage2_3[22],stage2_2[22],stage2_1[22]}
   );
   gpc606_5 gpc2270 (
      {stage1_1[86], stage1_1[87], stage1_1[88], stage1_1[89], stage1_1[90], stage1_1[91]},
      {stage1_3[74], stage1_3[75], stage1_3[76], stage1_3[77], stage1_3[78], stage1_3[79]},
      {stage2_5[11],stage2_4[23],stage2_3[23],stage2_2[23],stage2_1[23]}
   );
   gpc606_5 gpc2271 (
      {stage1_1[92], stage1_1[93], stage1_1[94], stage1_1[95], stage1_1[96], stage1_1[97]},
      {stage1_3[80], stage1_3[81], stage1_3[82], stage1_3[83], stage1_3[84], stage1_3[85]},
      {stage2_5[12],stage2_4[24],stage2_3[24],stage2_2[24],stage2_1[24]}
   );
   gpc606_5 gpc2272 (
      {stage1_1[98], stage1_1[99], stage1_1[100], stage1_1[101], stage1_1[102], stage1_1[103]},
      {stage1_3[86], stage1_3[87], stage1_3[88], stage1_3[89], stage1_3[90], stage1_3[91]},
      {stage2_5[13],stage2_4[25],stage2_3[25],stage2_2[25],stage2_1[25]}
   );
   gpc606_5 gpc2273 (
      {stage1_1[104], stage1_1[105], stage1_1[106], stage1_1[107], stage1_1[108], stage1_1[109]},
      {stage1_3[92], stage1_3[93], stage1_3[94], stage1_3[95], stage1_3[96], stage1_3[97]},
      {stage2_5[14],stage2_4[26],stage2_3[26],stage2_2[26],stage2_1[26]}
   );
   gpc606_5 gpc2274 (
      {stage1_1[110], stage1_1[111], stage1_1[112], stage1_1[113], stage1_1[114], stage1_1[115]},
      {stage1_3[98], stage1_3[99], stage1_3[100], stage1_3[101], stage1_3[102], stage1_3[103]},
      {stage2_5[15],stage2_4[27],stage2_3[27],stage2_2[27],stage2_1[27]}
   );
   gpc606_5 gpc2275 (
      {stage1_1[116], stage1_1[117], stage1_1[118], stage1_1[119], stage1_1[120], stage1_1[121]},
      {stage1_3[104], stage1_3[105], stage1_3[106], stage1_3[107], stage1_3[108], stage1_3[109]},
      {stage2_5[16],stage2_4[28],stage2_3[28],stage2_2[28],stage2_1[28]}
   );
   gpc606_5 gpc2276 (
      {stage1_1[122], stage1_1[123], stage1_1[124], stage1_1[125], stage1_1[126], stage1_1[127]},
      {stage1_3[110], stage1_3[111], stage1_3[112], stage1_3[113], stage1_3[114], stage1_3[115]},
      {stage2_5[17],stage2_4[29],stage2_3[29],stage2_2[29],stage2_1[29]}
   );
   gpc606_5 gpc2277 (
      {stage1_1[128], stage1_1[129], stage1_1[130], stage1_1[131], stage1_1[132], stage1_1[133]},
      {stage1_3[116], stage1_3[117], stage1_3[118], stage1_3[119], stage1_3[120], stage1_3[121]},
      {stage2_5[18],stage2_4[30],stage2_3[30],stage2_2[30],stage2_1[30]}
   );
   gpc606_5 gpc2278 (
      {stage1_1[134], stage1_1[135], stage1_1[136], stage1_1[137], stage1_1[138], stage1_1[139]},
      {stage1_3[122], stage1_3[123], stage1_3[124], stage1_3[125], stage1_3[126], stage1_3[127]},
      {stage2_5[19],stage2_4[31],stage2_3[31],stage2_2[31],stage2_1[31]}
   );
   gpc606_5 gpc2279 (
      {stage1_1[140], stage1_1[141], stage1_1[142], stage1_1[143], stage1_1[144], stage1_1[145]},
      {stage1_3[128], stage1_3[129], stage1_3[130], stage1_3[131], stage1_3[132], stage1_3[133]},
      {stage2_5[20],stage2_4[32],stage2_3[32],stage2_2[32],stage2_1[32]}
   );
   gpc606_5 gpc2280 (
      {stage1_1[146], stage1_1[147], stage1_1[148], stage1_1[149], stage1_1[150], stage1_1[151]},
      {stage1_3[134], stage1_3[135], stage1_3[136], stage1_3[137], stage1_3[138], stage1_3[139]},
      {stage2_5[21],stage2_4[33],stage2_3[33],stage2_2[33],stage2_1[33]}
   );
   gpc606_5 gpc2281 (
      {stage1_1[152], stage1_1[153], stage1_1[154], stage1_1[155], stage1_1[156], stage1_1[157]},
      {stage1_3[140], stage1_3[141], stage1_3[142], stage1_3[143], stage1_3[144], stage1_3[145]},
      {stage2_5[22],stage2_4[34],stage2_3[34],stage2_2[34],stage2_1[34]}
   );
   gpc606_5 gpc2282 (
      {stage1_1[158], stage1_1[159], stage1_1[160], stage1_1[161], stage1_1[162], stage1_1[163]},
      {stage1_3[146], stage1_3[147], stage1_3[148], stage1_3[149], stage1_3[150], stage1_3[151]},
      {stage2_5[23],stage2_4[35],stage2_3[35],stage2_2[35],stage2_1[35]}
   );
   gpc606_5 gpc2283 (
      {stage1_1[164], stage1_1[165], stage1_1[166], stage1_1[167], stage1_1[168], stage1_1[169]},
      {stage1_3[152], stage1_3[153], stage1_3[154], stage1_3[155], stage1_3[156], stage1_3[157]},
      {stage2_5[24],stage2_4[36],stage2_3[36],stage2_2[36],stage2_1[36]}
   );
   gpc606_5 gpc2284 (
      {stage1_1[170], stage1_1[171], stage1_1[172], stage1_1[173], stage1_1[174], stage1_1[175]},
      {stage1_3[158], stage1_3[159], stage1_3[160], stage1_3[161], stage1_3[162], stage1_3[163]},
      {stage2_5[25],stage2_4[37],stage2_3[37],stage2_2[37],stage2_1[37]}
   );
   gpc606_5 gpc2285 (
      {stage1_1[176], stage1_1[177], stage1_1[178], stage1_1[179], stage1_1[180], stage1_1[181]},
      {stage1_3[164], stage1_3[165], stage1_3[166], stage1_3[167], stage1_3[168], stage1_3[169]},
      {stage2_5[26],stage2_4[38],stage2_3[38],stage2_2[38],stage2_1[38]}
   );
   gpc615_5 gpc2286 (
      {stage1_2[52], stage1_2[53], stage1_2[54], stage1_2[55], stage1_2[56]},
      {stage1_3[170]},
      {stage1_4[0], stage1_4[1], stage1_4[2], stage1_4[3], stage1_4[4], stage1_4[5]},
      {stage2_6[0],stage2_5[27],stage2_4[39],stage2_3[39],stage2_2[39]}
   );
   gpc615_5 gpc2287 (
      {stage1_2[57], stage1_2[58], stage1_2[59], stage1_2[60], stage1_2[61]},
      {stage1_3[171]},
      {stage1_4[6], stage1_4[7], stage1_4[8], stage1_4[9], stage1_4[10], stage1_4[11]},
      {stage2_6[1],stage2_5[28],stage2_4[40],stage2_3[40],stage2_2[40]}
   );
   gpc615_5 gpc2288 (
      {stage1_2[62], stage1_2[63], stage1_2[64], stage1_2[65], stage1_2[66]},
      {stage1_3[172]},
      {stage1_4[12], stage1_4[13], stage1_4[14], stage1_4[15], stage1_4[16], stage1_4[17]},
      {stage2_6[2],stage2_5[29],stage2_4[41],stage2_3[41],stage2_2[41]}
   );
   gpc615_5 gpc2289 (
      {stage1_2[67], stage1_2[68], stage1_2[69], stage1_2[70], stage1_2[71]},
      {stage1_3[173]},
      {stage1_4[18], stage1_4[19], stage1_4[20], stage1_4[21], stage1_4[22], stage1_4[23]},
      {stage2_6[3],stage2_5[30],stage2_4[42],stage2_3[42],stage2_2[42]}
   );
   gpc615_5 gpc2290 (
      {stage1_2[72], stage1_2[73], stage1_2[74], stage1_2[75], stage1_2[76]},
      {stage1_3[174]},
      {stage1_4[24], stage1_4[25], stage1_4[26], stage1_4[27], stage1_4[28], stage1_4[29]},
      {stage2_6[4],stage2_5[31],stage2_4[43],stage2_3[43],stage2_2[43]}
   );
   gpc615_5 gpc2291 (
      {stage1_2[77], stage1_2[78], stage1_2[79], stage1_2[80], stage1_2[81]},
      {stage1_3[175]},
      {stage1_4[30], stage1_4[31], stage1_4[32], stage1_4[33], stage1_4[34], stage1_4[35]},
      {stage2_6[5],stage2_5[32],stage2_4[44],stage2_3[44],stage2_2[44]}
   );
   gpc615_5 gpc2292 (
      {stage1_2[82], stage1_2[83], stage1_2[84], stage1_2[85], stage1_2[86]},
      {stage1_3[176]},
      {stage1_4[36], stage1_4[37], stage1_4[38], stage1_4[39], stage1_4[40], stage1_4[41]},
      {stage2_6[6],stage2_5[33],stage2_4[45],stage2_3[45],stage2_2[45]}
   );
   gpc615_5 gpc2293 (
      {stage1_2[87], stage1_2[88], stage1_2[89], stage1_2[90], stage1_2[91]},
      {stage1_3[177]},
      {stage1_4[42], stage1_4[43], stage1_4[44], stage1_4[45], stage1_4[46], stage1_4[47]},
      {stage2_6[7],stage2_5[34],stage2_4[46],stage2_3[46],stage2_2[46]}
   );
   gpc615_5 gpc2294 (
      {stage1_2[92], stage1_2[93], stage1_2[94], stage1_2[95], stage1_2[96]},
      {stage1_3[178]},
      {stage1_4[48], stage1_4[49], stage1_4[50], stage1_4[51], stage1_4[52], stage1_4[53]},
      {stage2_6[8],stage2_5[35],stage2_4[47],stage2_3[47],stage2_2[47]}
   );
   gpc615_5 gpc2295 (
      {stage1_2[97], stage1_2[98], stage1_2[99], stage1_2[100], stage1_2[101]},
      {stage1_3[179]},
      {stage1_4[54], stage1_4[55], stage1_4[56], stage1_4[57], stage1_4[58], stage1_4[59]},
      {stage2_6[9],stage2_5[36],stage2_4[48],stage2_3[48],stage2_2[48]}
   );
   gpc615_5 gpc2296 (
      {stage1_2[102], stage1_2[103], stage1_2[104], stage1_2[105], stage1_2[106]},
      {stage1_3[180]},
      {stage1_4[60], stage1_4[61], stage1_4[62], stage1_4[63], stage1_4[64], stage1_4[65]},
      {stage2_6[10],stage2_5[37],stage2_4[49],stage2_3[49],stage2_2[49]}
   );
   gpc615_5 gpc2297 (
      {stage1_2[107], stage1_2[108], stage1_2[109], stage1_2[110], stage1_2[111]},
      {stage1_3[181]},
      {stage1_4[66], stage1_4[67], stage1_4[68], stage1_4[69], stage1_4[70], stage1_4[71]},
      {stage2_6[11],stage2_5[38],stage2_4[50],stage2_3[50],stage2_2[50]}
   );
   gpc615_5 gpc2298 (
      {stage1_2[112], stage1_2[113], stage1_2[114], stage1_2[115], stage1_2[116]},
      {stage1_3[182]},
      {stage1_4[72], stage1_4[73], stage1_4[74], stage1_4[75], stage1_4[76], stage1_4[77]},
      {stage2_6[12],stage2_5[39],stage2_4[51],stage2_3[51],stage2_2[51]}
   );
   gpc615_5 gpc2299 (
      {stage1_2[117], stage1_2[118], stage1_2[119], stage1_2[120], stage1_2[121]},
      {stage1_3[183]},
      {stage1_4[78], stage1_4[79], stage1_4[80], stage1_4[81], stage1_4[82], stage1_4[83]},
      {stage2_6[13],stage2_5[40],stage2_4[52],stage2_3[52],stage2_2[52]}
   );
   gpc615_5 gpc2300 (
      {stage1_2[122], stage1_2[123], stage1_2[124], stage1_2[125], stage1_2[126]},
      {stage1_3[184]},
      {stage1_4[84], stage1_4[85], stage1_4[86], stage1_4[87], stage1_4[88], stage1_4[89]},
      {stage2_6[14],stage2_5[41],stage2_4[53],stage2_3[53],stage2_2[53]}
   );
   gpc615_5 gpc2301 (
      {stage1_2[127], stage1_2[128], stage1_2[129], stage1_2[130], stage1_2[131]},
      {stage1_3[185]},
      {stage1_4[90], stage1_4[91], stage1_4[92], stage1_4[93], stage1_4[94], stage1_4[95]},
      {stage2_6[15],stage2_5[42],stage2_4[54],stage2_3[54],stage2_2[54]}
   );
   gpc615_5 gpc2302 (
      {stage1_2[132], stage1_2[133], stage1_2[134], stage1_2[135], stage1_2[136]},
      {stage1_3[186]},
      {stage1_4[96], stage1_4[97], stage1_4[98], stage1_4[99], stage1_4[100], stage1_4[101]},
      {stage2_6[16],stage2_5[43],stage2_4[55],stage2_3[55],stage2_2[55]}
   );
   gpc615_5 gpc2303 (
      {stage1_2[137], stage1_2[138], stage1_2[139], stage1_2[140], stage1_2[141]},
      {stage1_3[187]},
      {stage1_4[102], stage1_4[103], stage1_4[104], stage1_4[105], stage1_4[106], stage1_4[107]},
      {stage2_6[17],stage2_5[44],stage2_4[56],stage2_3[56],stage2_2[56]}
   );
   gpc615_5 gpc2304 (
      {stage1_2[142], stage1_2[143], stage1_2[144], stage1_2[145], stage1_2[146]},
      {stage1_3[188]},
      {stage1_4[108], stage1_4[109], stage1_4[110], stage1_4[111], stage1_4[112], stage1_4[113]},
      {stage2_6[18],stage2_5[45],stage2_4[57],stage2_3[57],stage2_2[57]}
   );
   gpc615_5 gpc2305 (
      {stage1_2[147], stage1_2[148], stage1_2[149], stage1_2[150], stage1_2[151]},
      {stage1_3[189]},
      {stage1_4[114], stage1_4[115], stage1_4[116], stage1_4[117], stage1_4[118], stage1_4[119]},
      {stage2_6[19],stage2_5[46],stage2_4[58],stage2_3[58],stage2_2[58]}
   );
   gpc615_5 gpc2306 (
      {stage1_3[190], stage1_3[191], stage1_3[192], stage1_3[193], stage1_3[194]},
      {stage1_4[120]},
      {stage1_5[0], stage1_5[1], stage1_5[2], stage1_5[3], stage1_5[4], stage1_5[5]},
      {stage2_7[0],stage2_6[20],stage2_5[47],stage2_4[59],stage2_3[59]}
   );
   gpc615_5 gpc2307 (
      {stage1_3[195], stage1_3[196], stage1_3[197], stage1_3[198], stage1_3[199]},
      {stage1_4[121]},
      {stage1_5[6], stage1_5[7], stage1_5[8], stage1_5[9], stage1_5[10], stage1_5[11]},
      {stage2_7[1],stage2_6[21],stage2_5[48],stage2_4[60],stage2_3[60]}
   );
   gpc615_5 gpc2308 (
      {stage1_3[200], stage1_3[201], stage1_3[202], stage1_3[203], stage1_3[204]},
      {stage1_4[122]},
      {stage1_5[12], stage1_5[13], stage1_5[14], stage1_5[15], stage1_5[16], stage1_5[17]},
      {stage2_7[2],stage2_6[22],stage2_5[49],stage2_4[61],stage2_3[61]}
   );
   gpc615_5 gpc2309 (
      {stage1_3[205], stage1_3[206], stage1_3[207], stage1_3[208], stage1_3[209]},
      {stage1_4[123]},
      {stage1_5[18], stage1_5[19], stage1_5[20], stage1_5[21], stage1_5[22], stage1_5[23]},
      {stage2_7[3],stage2_6[23],stage2_5[50],stage2_4[62],stage2_3[62]}
   );
   gpc615_5 gpc2310 (
      {stage1_3[210], stage1_3[211], stage1_3[212], stage1_3[213], stage1_3[214]},
      {stage1_4[124]},
      {stage1_5[24], stage1_5[25], stage1_5[26], stage1_5[27], stage1_5[28], stage1_5[29]},
      {stage2_7[4],stage2_6[24],stage2_5[51],stage2_4[63],stage2_3[63]}
   );
   gpc615_5 gpc2311 (
      {stage1_3[215], stage1_3[216], stage1_3[217], stage1_3[218], stage1_3[219]},
      {stage1_4[125]},
      {stage1_5[30], stage1_5[31], stage1_5[32], stage1_5[33], stage1_5[34], stage1_5[35]},
      {stage2_7[5],stage2_6[25],stage2_5[52],stage2_4[64],stage2_3[64]}
   );
   gpc615_5 gpc2312 (
      {stage1_3[220], stage1_3[221], stage1_3[222], stage1_3[223], stage1_3[224]},
      {stage1_4[126]},
      {stage1_5[36], stage1_5[37], stage1_5[38], stage1_5[39], stage1_5[40], stage1_5[41]},
      {stage2_7[6],stage2_6[26],stage2_5[53],stage2_4[65],stage2_3[65]}
   );
   gpc615_5 gpc2313 (
      {stage1_3[225], stage1_3[226], stage1_3[227], stage1_3[228], stage1_3[229]},
      {stage1_4[127]},
      {stage1_5[42], stage1_5[43], stage1_5[44], stage1_5[45], stage1_5[46], stage1_5[47]},
      {stage2_7[7],stage2_6[27],stage2_5[54],stage2_4[66],stage2_3[66]}
   );
   gpc615_5 gpc2314 (
      {stage1_3[230], stage1_3[231], stage1_3[232], stage1_3[233], stage1_3[234]},
      {stage1_4[128]},
      {stage1_5[48], stage1_5[49], stage1_5[50], stage1_5[51], stage1_5[52], stage1_5[53]},
      {stage2_7[8],stage2_6[28],stage2_5[55],stage2_4[67],stage2_3[67]}
   );
   gpc615_5 gpc2315 (
      {stage1_3[235], stage1_3[236], stage1_3[237], stage1_3[238], stage1_3[239]},
      {stage1_4[129]},
      {stage1_5[54], stage1_5[55], stage1_5[56], stage1_5[57], stage1_5[58], stage1_5[59]},
      {stage2_7[9],stage2_6[29],stage2_5[56],stage2_4[68],stage2_3[68]}
   );
   gpc615_5 gpc2316 (
      {stage1_3[240], stage1_3[241], stage1_3[242], stage1_3[243], stage1_3[244]},
      {stage1_4[130]},
      {stage1_5[60], stage1_5[61], stage1_5[62], stage1_5[63], stage1_5[64], stage1_5[65]},
      {stage2_7[10],stage2_6[30],stage2_5[57],stage2_4[69],stage2_3[69]}
   );
   gpc615_5 gpc2317 (
      {stage1_3[245], stage1_3[246], stage1_3[247], stage1_3[248], stage1_3[249]},
      {stage1_4[131]},
      {stage1_5[66], stage1_5[67], stage1_5[68], stage1_5[69], stage1_5[70], stage1_5[71]},
      {stage2_7[11],stage2_6[31],stage2_5[58],stage2_4[70],stage2_3[70]}
   );
   gpc615_5 gpc2318 (
      {stage1_3[250], stage1_3[251], stage1_3[252], stage1_3[253], stage1_3[254]},
      {stage1_4[132]},
      {stage1_5[72], stage1_5[73], stage1_5[74], stage1_5[75], stage1_5[76], stage1_5[77]},
      {stage2_7[12],stage2_6[32],stage2_5[59],stage2_4[71],stage2_3[71]}
   );
   gpc615_5 gpc2319 (
      {stage1_3[255], stage1_3[256], stage1_3[257], stage1_3[258], stage1_3[259]},
      {stage1_4[133]},
      {stage1_5[78], stage1_5[79], stage1_5[80], stage1_5[81], stage1_5[82], stage1_5[83]},
      {stage2_7[13],stage2_6[33],stage2_5[60],stage2_4[72],stage2_3[72]}
   );
   gpc615_5 gpc2320 (
      {stage1_3[260], stage1_3[261], stage1_3[262], stage1_3[263], stage1_3[264]},
      {stage1_4[134]},
      {stage1_5[84], stage1_5[85], stage1_5[86], stage1_5[87], stage1_5[88], stage1_5[89]},
      {stage2_7[14],stage2_6[34],stage2_5[61],stage2_4[73],stage2_3[73]}
   );
   gpc615_5 gpc2321 (
      {stage1_3[265], stage1_3[266], stage1_3[267], stage1_3[268], stage1_3[269]},
      {stage1_4[135]},
      {stage1_5[90], stage1_5[91], stage1_5[92], stage1_5[93], stage1_5[94], stage1_5[95]},
      {stage2_7[15],stage2_6[35],stage2_5[62],stage2_4[74],stage2_3[74]}
   );
   gpc615_5 gpc2322 (
      {stage1_3[270], stage1_3[271], stage1_3[272], stage1_3[273], stage1_3[274]},
      {stage1_4[136]},
      {stage1_5[96], stage1_5[97], stage1_5[98], stage1_5[99], stage1_5[100], stage1_5[101]},
      {stage2_7[16],stage2_6[36],stage2_5[63],stage2_4[75],stage2_3[75]}
   );
   gpc615_5 gpc2323 (
      {stage1_3[275], stage1_3[276], 1'b0, 1'b0, 1'b0},
      {stage1_4[137]},
      {stage1_5[102], stage1_5[103], stage1_5[104], stage1_5[105], stage1_5[106], stage1_5[107]},
      {stage2_7[17],stage2_6[37],stage2_5[64],stage2_4[76],stage2_3[76]}
   );
   gpc1163_5 gpc2324 (
      {stage1_4[138], stage1_4[139], stage1_4[140]},
      {stage1_5[108], stage1_5[109], stage1_5[110], stage1_5[111], stage1_5[112], stage1_5[113]},
      {stage1_6[0]},
      {stage1_7[0]},
      {stage2_8[0],stage2_7[18],stage2_6[38],stage2_5[65],stage2_4[77]}
   );
   gpc606_5 gpc2325 (
      {stage1_4[141], stage1_4[142], stage1_4[143], stage1_4[144], stage1_4[145], stage1_4[146]},
      {stage1_6[1], stage1_6[2], stage1_6[3], stage1_6[4], stage1_6[5], stage1_6[6]},
      {stage2_8[1],stage2_7[19],stage2_6[39],stage2_5[66],stage2_4[78]}
   );
   gpc606_5 gpc2326 (
      {stage1_4[147], stage1_4[148], stage1_4[149], stage1_4[150], stage1_4[151], stage1_4[152]},
      {stage1_6[7], stage1_6[8], stage1_6[9], stage1_6[10], stage1_6[11], stage1_6[12]},
      {stage2_8[2],stage2_7[20],stage2_6[40],stage2_5[67],stage2_4[79]}
   );
   gpc606_5 gpc2327 (
      {stage1_4[153], stage1_4[154], stage1_4[155], stage1_4[156], stage1_4[157], stage1_4[158]},
      {stage1_6[13], stage1_6[14], stage1_6[15], stage1_6[16], stage1_6[17], stage1_6[18]},
      {stage2_8[3],stage2_7[21],stage2_6[41],stage2_5[68],stage2_4[80]}
   );
   gpc606_5 gpc2328 (
      {stage1_4[159], stage1_4[160], stage1_4[161], stage1_4[162], stage1_4[163], stage1_4[164]},
      {stage1_6[19], stage1_6[20], stage1_6[21], stage1_6[22], stage1_6[23], stage1_6[24]},
      {stage2_8[4],stage2_7[22],stage2_6[42],stage2_5[69],stage2_4[81]}
   );
   gpc606_5 gpc2329 (
      {stage1_4[165], stage1_4[166], stage1_4[167], stage1_4[168], stage1_4[169], stage1_4[170]},
      {stage1_6[25], stage1_6[26], stage1_6[27], stage1_6[28], stage1_6[29], stage1_6[30]},
      {stage2_8[5],stage2_7[23],stage2_6[43],stage2_5[70],stage2_4[82]}
   );
   gpc606_5 gpc2330 (
      {stage1_4[171], stage1_4[172], stage1_4[173], stage1_4[174], stage1_4[175], stage1_4[176]},
      {stage1_6[31], stage1_6[32], stage1_6[33], stage1_6[34], stage1_6[35], stage1_6[36]},
      {stage2_8[6],stage2_7[24],stage2_6[44],stage2_5[71],stage2_4[83]}
   );
   gpc606_5 gpc2331 (
      {stage1_4[177], stage1_4[178], stage1_4[179], stage1_4[180], stage1_4[181], stage1_4[182]},
      {stage1_6[37], stage1_6[38], stage1_6[39], stage1_6[40], stage1_6[41], stage1_6[42]},
      {stage2_8[7],stage2_7[25],stage2_6[45],stage2_5[72],stage2_4[84]}
   );
   gpc606_5 gpc2332 (
      {stage1_4[183], stage1_4[184], stage1_4[185], stage1_4[186], stage1_4[187], stage1_4[188]},
      {stage1_6[43], stage1_6[44], stage1_6[45], stage1_6[46], stage1_6[47], stage1_6[48]},
      {stage2_8[8],stage2_7[26],stage2_6[46],stage2_5[73],stage2_4[85]}
   );
   gpc606_5 gpc2333 (
      {stage1_4[189], stage1_4[190], stage1_4[191], stage1_4[192], stage1_4[193], stage1_4[194]},
      {stage1_6[49], stage1_6[50], stage1_6[51], stage1_6[52], stage1_6[53], stage1_6[54]},
      {stage2_8[9],stage2_7[27],stage2_6[47],stage2_5[74],stage2_4[86]}
   );
   gpc606_5 gpc2334 (
      {stage1_4[195], stage1_4[196], stage1_4[197], stage1_4[198], stage1_4[199], stage1_4[200]},
      {stage1_6[55], stage1_6[56], stage1_6[57], stage1_6[58], stage1_6[59], stage1_6[60]},
      {stage2_8[10],stage2_7[28],stage2_6[48],stage2_5[75],stage2_4[87]}
   );
   gpc606_5 gpc2335 (
      {stage1_4[201], stage1_4[202], stage1_4[203], stage1_4[204], stage1_4[205], stage1_4[206]},
      {stage1_6[61], stage1_6[62], stage1_6[63], stage1_6[64], stage1_6[65], stage1_6[66]},
      {stage2_8[11],stage2_7[29],stage2_6[49],stage2_5[76],stage2_4[88]}
   );
   gpc615_5 gpc2336 (
      {stage1_4[207], stage1_4[208], stage1_4[209], stage1_4[210], stage1_4[211]},
      {stage1_5[114]},
      {stage1_6[67], stage1_6[68], stage1_6[69], stage1_6[70], stage1_6[71], stage1_6[72]},
      {stage2_8[12],stage2_7[30],stage2_6[50],stage2_5[77],stage2_4[89]}
   );
   gpc615_5 gpc2337 (
      {stage1_4[212], stage1_4[213], stage1_4[214], stage1_4[215], stage1_4[216]},
      {stage1_5[115]},
      {stage1_6[73], stage1_6[74], stage1_6[75], stage1_6[76], stage1_6[77], stage1_6[78]},
      {stage2_8[13],stage2_7[31],stage2_6[51],stage2_5[78],stage2_4[90]}
   );
   gpc606_5 gpc2338 (
      {stage1_5[116], stage1_5[117], stage1_5[118], stage1_5[119], stage1_5[120], stage1_5[121]},
      {stage1_7[1], stage1_7[2], stage1_7[3], stage1_7[4], stage1_7[5], stage1_7[6]},
      {stage2_9[0],stage2_8[14],stage2_7[32],stage2_6[52],stage2_5[79]}
   );
   gpc606_5 gpc2339 (
      {stage1_5[122], stage1_5[123], stage1_5[124], stage1_5[125], stage1_5[126], stage1_5[127]},
      {stage1_7[7], stage1_7[8], stage1_7[9], stage1_7[10], stage1_7[11], stage1_7[12]},
      {stage2_9[1],stage2_8[15],stage2_7[33],stage2_6[53],stage2_5[80]}
   );
   gpc606_5 gpc2340 (
      {stage1_5[128], stage1_5[129], stage1_5[130], stage1_5[131], stage1_5[132], stage1_5[133]},
      {stage1_7[13], stage1_7[14], stage1_7[15], stage1_7[16], stage1_7[17], stage1_7[18]},
      {stage2_9[2],stage2_8[16],stage2_7[34],stage2_6[54],stage2_5[81]}
   );
   gpc606_5 gpc2341 (
      {stage1_5[134], stage1_5[135], stage1_5[136], stage1_5[137], stage1_5[138], stage1_5[139]},
      {stage1_7[19], stage1_7[20], stage1_7[21], stage1_7[22], stage1_7[23], stage1_7[24]},
      {stage2_9[3],stage2_8[17],stage2_7[35],stage2_6[55],stage2_5[82]}
   );
   gpc606_5 gpc2342 (
      {stage1_5[140], stage1_5[141], stage1_5[142], stage1_5[143], stage1_5[144], stage1_5[145]},
      {stage1_7[25], stage1_7[26], stage1_7[27], stage1_7[28], stage1_7[29], stage1_7[30]},
      {stage2_9[4],stage2_8[18],stage2_7[36],stage2_6[56],stage2_5[83]}
   );
   gpc606_5 gpc2343 (
      {stage1_5[146], stage1_5[147], stage1_5[148], stage1_5[149], stage1_5[150], stage1_5[151]},
      {stage1_7[31], stage1_7[32], stage1_7[33], stage1_7[34], stage1_7[35], stage1_7[36]},
      {stage2_9[5],stage2_8[19],stage2_7[37],stage2_6[57],stage2_5[84]}
   );
   gpc606_5 gpc2344 (
      {stage1_5[152], stage1_5[153], stage1_5[154], stage1_5[155], stage1_5[156], stage1_5[157]},
      {stage1_7[37], stage1_7[38], stage1_7[39], stage1_7[40], stage1_7[41], stage1_7[42]},
      {stage2_9[6],stage2_8[20],stage2_7[38],stage2_6[58],stage2_5[85]}
   );
   gpc606_5 gpc2345 (
      {stage1_5[158], stage1_5[159], stage1_5[160], stage1_5[161], stage1_5[162], stage1_5[163]},
      {stage1_7[43], stage1_7[44], stage1_7[45], stage1_7[46], stage1_7[47], stage1_7[48]},
      {stage2_9[7],stage2_8[21],stage2_7[39],stage2_6[59],stage2_5[86]}
   );
   gpc606_5 gpc2346 (
      {stage1_5[164], stage1_5[165], stage1_5[166], stage1_5[167], stage1_5[168], stage1_5[169]},
      {stage1_7[49], stage1_7[50], stage1_7[51], stage1_7[52], stage1_7[53], stage1_7[54]},
      {stage2_9[8],stage2_8[22],stage2_7[40],stage2_6[60],stage2_5[87]}
   );
   gpc606_5 gpc2347 (
      {stage1_5[170], stage1_5[171], stage1_5[172], stage1_5[173], stage1_5[174], stage1_5[175]},
      {stage1_7[55], stage1_7[56], stage1_7[57], stage1_7[58], stage1_7[59], stage1_7[60]},
      {stage2_9[9],stage2_8[23],stage2_7[41],stage2_6[61],stage2_5[88]}
   );
   gpc606_5 gpc2348 (
      {stage1_5[176], stage1_5[177], stage1_5[178], stage1_5[179], stage1_5[180], stage1_5[181]},
      {stage1_7[61], stage1_7[62], stage1_7[63], stage1_7[64], stage1_7[65], stage1_7[66]},
      {stage2_9[10],stage2_8[24],stage2_7[42],stage2_6[62],stage2_5[89]}
   );
   gpc606_5 gpc2349 (
      {stage1_5[182], stage1_5[183], stage1_5[184], stage1_5[185], stage1_5[186], stage1_5[187]},
      {stage1_7[67], stage1_7[68], stage1_7[69], stage1_7[70], stage1_7[71], stage1_7[72]},
      {stage2_9[11],stage2_8[25],stage2_7[43],stage2_6[63],stage2_5[90]}
   );
   gpc606_5 gpc2350 (
      {stage1_5[188], stage1_5[189], stage1_5[190], stage1_5[191], stage1_5[192], stage1_5[193]},
      {stage1_7[73], stage1_7[74], stage1_7[75], stage1_7[76], stage1_7[77], stage1_7[78]},
      {stage2_9[12],stage2_8[26],stage2_7[44],stage2_6[64],stage2_5[91]}
   );
   gpc606_5 gpc2351 (
      {stage1_5[194], stage1_5[195], stage1_5[196], stage1_5[197], stage1_5[198], stage1_5[199]},
      {stage1_7[79], stage1_7[80], stage1_7[81], stage1_7[82], stage1_7[83], stage1_7[84]},
      {stage2_9[13],stage2_8[27],stage2_7[45],stage2_6[65],stage2_5[92]}
   );
   gpc606_5 gpc2352 (
      {stage1_5[200], stage1_5[201], stage1_5[202], stage1_5[203], stage1_5[204], stage1_5[205]},
      {stage1_7[85], stage1_7[86], stage1_7[87], stage1_7[88], stage1_7[89], stage1_7[90]},
      {stage2_9[14],stage2_8[28],stage2_7[46],stage2_6[66],stage2_5[93]}
   );
   gpc606_5 gpc2353 (
      {stage1_6[79], stage1_6[80], stage1_6[81], stage1_6[82], stage1_6[83], stage1_6[84]},
      {stage1_8[0], stage1_8[1], stage1_8[2], stage1_8[3], stage1_8[4], stage1_8[5]},
      {stage2_10[0],stage2_9[15],stage2_8[29],stage2_7[47],stage2_6[67]}
   );
   gpc606_5 gpc2354 (
      {stage1_6[85], stage1_6[86], stage1_6[87], stage1_6[88], stage1_6[89], stage1_6[90]},
      {stage1_8[6], stage1_8[7], stage1_8[8], stage1_8[9], stage1_8[10], stage1_8[11]},
      {stage2_10[1],stage2_9[16],stage2_8[30],stage2_7[48],stage2_6[68]}
   );
   gpc606_5 gpc2355 (
      {stage1_6[91], stage1_6[92], stage1_6[93], stage1_6[94], stage1_6[95], stage1_6[96]},
      {stage1_8[12], stage1_8[13], stage1_8[14], stage1_8[15], stage1_8[16], stage1_8[17]},
      {stage2_10[2],stage2_9[17],stage2_8[31],stage2_7[49],stage2_6[69]}
   );
   gpc606_5 gpc2356 (
      {stage1_6[97], stage1_6[98], stage1_6[99], stage1_6[100], stage1_6[101], stage1_6[102]},
      {stage1_8[18], stage1_8[19], stage1_8[20], stage1_8[21], stage1_8[22], stage1_8[23]},
      {stage2_10[3],stage2_9[18],stage2_8[32],stage2_7[50],stage2_6[70]}
   );
   gpc606_5 gpc2357 (
      {stage1_6[103], stage1_6[104], stage1_6[105], stage1_6[106], stage1_6[107], stage1_6[108]},
      {stage1_8[24], stage1_8[25], stage1_8[26], stage1_8[27], stage1_8[28], stage1_8[29]},
      {stage2_10[4],stage2_9[19],stage2_8[33],stage2_7[51],stage2_6[71]}
   );
   gpc606_5 gpc2358 (
      {stage1_6[109], stage1_6[110], stage1_6[111], stage1_6[112], stage1_6[113], stage1_6[114]},
      {stage1_8[30], stage1_8[31], stage1_8[32], stage1_8[33], stage1_8[34], stage1_8[35]},
      {stage2_10[5],stage2_9[20],stage2_8[34],stage2_7[52],stage2_6[72]}
   );
   gpc606_5 gpc2359 (
      {stage1_6[115], stage1_6[116], stage1_6[117], stage1_6[118], stage1_6[119], stage1_6[120]},
      {stage1_8[36], stage1_8[37], stage1_8[38], stage1_8[39], stage1_8[40], stage1_8[41]},
      {stage2_10[6],stage2_9[21],stage2_8[35],stage2_7[53],stage2_6[73]}
   );
   gpc606_5 gpc2360 (
      {stage1_6[121], stage1_6[122], stage1_6[123], stage1_6[124], stage1_6[125], stage1_6[126]},
      {stage1_8[42], stage1_8[43], stage1_8[44], stage1_8[45], stage1_8[46], stage1_8[47]},
      {stage2_10[7],stage2_9[22],stage2_8[36],stage2_7[54],stage2_6[74]}
   );
   gpc606_5 gpc2361 (
      {stage1_6[127], stage1_6[128], stage1_6[129], stage1_6[130], stage1_6[131], stage1_6[132]},
      {stage1_8[48], stage1_8[49], stage1_8[50], stage1_8[51], stage1_8[52], stage1_8[53]},
      {stage2_10[8],stage2_9[23],stage2_8[37],stage2_7[55],stage2_6[75]}
   );
   gpc606_5 gpc2362 (
      {stage1_6[133], stage1_6[134], stage1_6[135], stage1_6[136], stage1_6[137], stage1_6[138]},
      {stage1_8[54], stage1_8[55], stage1_8[56], stage1_8[57], stage1_8[58], stage1_8[59]},
      {stage2_10[9],stage2_9[24],stage2_8[38],stage2_7[56],stage2_6[76]}
   );
   gpc606_5 gpc2363 (
      {stage1_6[139], stage1_6[140], stage1_6[141], stage1_6[142], stage1_6[143], stage1_6[144]},
      {stage1_8[60], stage1_8[61], stage1_8[62], stage1_8[63], stage1_8[64], stage1_8[65]},
      {stage2_10[10],stage2_9[25],stage2_8[39],stage2_7[57],stage2_6[77]}
   );
   gpc606_5 gpc2364 (
      {stage1_6[145], stage1_6[146], stage1_6[147], stage1_6[148], stage1_6[149], stage1_6[150]},
      {stage1_8[66], stage1_8[67], stage1_8[68], stage1_8[69], stage1_8[70], stage1_8[71]},
      {stage2_10[11],stage2_9[26],stage2_8[40],stage2_7[58],stage2_6[78]}
   );
   gpc606_5 gpc2365 (
      {stage1_6[151], stage1_6[152], stage1_6[153], stage1_6[154], stage1_6[155], stage1_6[156]},
      {stage1_8[72], stage1_8[73], stage1_8[74], stage1_8[75], stage1_8[76], stage1_8[77]},
      {stage2_10[12],stage2_9[27],stage2_8[41],stage2_7[59],stage2_6[79]}
   );
   gpc606_5 gpc2366 (
      {stage1_6[157], stage1_6[158], stage1_6[159], stage1_6[160], stage1_6[161], stage1_6[162]},
      {stage1_8[78], stage1_8[79], stage1_8[80], stage1_8[81], stage1_8[82], stage1_8[83]},
      {stage2_10[13],stage2_9[28],stage2_8[42],stage2_7[60],stage2_6[80]}
   );
   gpc606_5 gpc2367 (
      {stage1_6[163], stage1_6[164], stage1_6[165], stage1_6[166], stage1_6[167], stage1_6[168]},
      {stage1_8[84], stage1_8[85], stage1_8[86], stage1_8[87], stage1_8[88], stage1_8[89]},
      {stage2_10[14],stage2_9[29],stage2_8[43],stage2_7[61],stage2_6[81]}
   );
   gpc606_5 gpc2368 (
      {stage1_6[169], stage1_6[170], stage1_6[171], stage1_6[172], stage1_6[173], stage1_6[174]},
      {stage1_8[90], stage1_8[91], stage1_8[92], stage1_8[93], stage1_8[94], stage1_8[95]},
      {stage2_10[15],stage2_9[30],stage2_8[44],stage2_7[62],stage2_6[82]}
   );
   gpc606_5 gpc2369 (
      {stage1_6[175], stage1_6[176], stage1_6[177], stage1_6[178], stage1_6[179], stage1_6[180]},
      {stage1_8[96], stage1_8[97], stage1_8[98], stage1_8[99], stage1_8[100], stage1_8[101]},
      {stage2_10[16],stage2_9[31],stage2_8[45],stage2_7[63],stage2_6[83]}
   );
   gpc606_5 gpc2370 (
      {stage1_6[181], stage1_6[182], stage1_6[183], stage1_6[184], stage1_6[185], stage1_6[186]},
      {stage1_8[102], stage1_8[103], stage1_8[104], stage1_8[105], stage1_8[106], stage1_8[107]},
      {stage2_10[17],stage2_9[32],stage2_8[46],stage2_7[64],stage2_6[84]}
   );
   gpc606_5 gpc2371 (
      {stage1_6[187], stage1_6[188], stage1_6[189], stage1_6[190], stage1_6[191], stage1_6[192]},
      {stage1_8[108], stage1_8[109], stage1_8[110], stage1_8[111], stage1_8[112], stage1_8[113]},
      {stage2_10[18],stage2_9[33],stage2_8[47],stage2_7[65],stage2_6[85]}
   );
   gpc615_5 gpc2372 (
      {stage1_6[193], stage1_6[194], stage1_6[195], stage1_6[196], stage1_6[197]},
      {stage1_7[91]},
      {stage1_8[114], stage1_8[115], stage1_8[116], stage1_8[117], stage1_8[118], stage1_8[119]},
      {stage2_10[19],stage2_9[34],stage2_8[48],stage2_7[66],stage2_6[86]}
   );
   gpc615_5 gpc2373 (
      {stage1_6[198], stage1_6[199], stage1_6[200], stage1_6[201], stage1_6[202]},
      {stage1_7[92]},
      {stage1_8[120], stage1_8[121], stage1_8[122], stage1_8[123], stage1_8[124], stage1_8[125]},
      {stage2_10[20],stage2_9[35],stage2_8[49],stage2_7[67],stage2_6[87]}
   );
   gpc615_5 gpc2374 (
      {stage1_6[203], stage1_6[204], stage1_6[205], stage1_6[206], stage1_6[207]},
      {stage1_7[93]},
      {stage1_8[126], stage1_8[127], stage1_8[128], stage1_8[129], stage1_8[130], stage1_8[131]},
      {stage2_10[21],stage2_9[36],stage2_8[50],stage2_7[68],stage2_6[88]}
   );
   gpc615_5 gpc2375 (
      {stage1_6[208], stage1_6[209], stage1_6[210], stage1_6[211], stage1_6[212]},
      {stage1_7[94]},
      {stage1_8[132], stage1_8[133], stage1_8[134], stage1_8[135], stage1_8[136], stage1_8[137]},
      {stage2_10[22],stage2_9[37],stage2_8[51],stage2_7[69],stage2_6[89]}
   );
   gpc615_5 gpc2376 (
      {stage1_6[213], stage1_6[214], stage1_6[215], stage1_6[216], stage1_6[217]},
      {stage1_7[95]},
      {stage1_8[138], stage1_8[139], stage1_8[140], stage1_8[141], stage1_8[142], stage1_8[143]},
      {stage2_10[23],stage2_9[38],stage2_8[52],stage2_7[70],stage2_6[90]}
   );
   gpc615_5 gpc2377 (
      {stage1_6[218], stage1_6[219], stage1_6[220], stage1_6[221], stage1_6[222]},
      {stage1_7[96]},
      {stage1_8[144], stage1_8[145], stage1_8[146], stage1_8[147], stage1_8[148], stage1_8[149]},
      {stage2_10[24],stage2_9[39],stage2_8[53],stage2_7[71],stage2_6[91]}
   );
   gpc615_5 gpc2378 (
      {stage1_6[223], stage1_6[224], stage1_6[225], stage1_6[226], stage1_6[227]},
      {stage1_7[97]},
      {stage1_8[150], stage1_8[151], stage1_8[152], stage1_8[153], stage1_8[154], stage1_8[155]},
      {stage2_10[25],stage2_9[40],stage2_8[54],stage2_7[72],stage2_6[92]}
   );
   gpc615_5 gpc2379 (
      {stage1_6[228], stage1_6[229], stage1_6[230], stage1_6[231], stage1_6[232]},
      {stage1_7[98]},
      {stage1_8[156], stage1_8[157], stage1_8[158], stage1_8[159], stage1_8[160], stage1_8[161]},
      {stage2_10[26],stage2_9[41],stage2_8[55],stage2_7[73],stage2_6[93]}
   );
   gpc615_5 gpc2380 (
      {stage1_6[233], stage1_6[234], stage1_6[235], stage1_6[236], stage1_6[237]},
      {stage1_7[99]},
      {stage1_8[162], stage1_8[163], stage1_8[164], stage1_8[165], stage1_8[166], stage1_8[167]},
      {stage2_10[27],stage2_9[42],stage2_8[56],stage2_7[74],stage2_6[94]}
   );
   gpc615_5 gpc2381 (
      {stage1_6[238], stage1_6[239], stage1_6[240], stage1_6[241], stage1_6[242]},
      {stage1_7[100]},
      {stage1_8[168], stage1_8[169], stage1_8[170], stage1_8[171], stage1_8[172], stage1_8[173]},
      {stage2_10[28],stage2_9[43],stage2_8[57],stage2_7[75],stage2_6[95]}
   );
   gpc615_5 gpc2382 (
      {stage1_7[101], stage1_7[102], stage1_7[103], stage1_7[104], stage1_7[105]},
      {stage1_8[174]},
      {stage1_9[0], stage1_9[1], stage1_9[2], stage1_9[3], stage1_9[4], stage1_9[5]},
      {stage2_11[0],stage2_10[29],stage2_9[44],stage2_8[58],stage2_7[76]}
   );
   gpc615_5 gpc2383 (
      {stage1_7[106], stage1_7[107], stage1_7[108], stage1_7[109], stage1_7[110]},
      {stage1_8[175]},
      {stage1_9[6], stage1_9[7], stage1_9[8], stage1_9[9], stage1_9[10], stage1_9[11]},
      {stage2_11[1],stage2_10[30],stage2_9[45],stage2_8[59],stage2_7[77]}
   );
   gpc615_5 gpc2384 (
      {stage1_7[111], stage1_7[112], stage1_7[113], stage1_7[114], stage1_7[115]},
      {stage1_8[176]},
      {stage1_9[12], stage1_9[13], stage1_9[14], stage1_9[15], stage1_9[16], stage1_9[17]},
      {stage2_11[2],stage2_10[31],stage2_9[46],stage2_8[60],stage2_7[78]}
   );
   gpc615_5 gpc2385 (
      {stage1_7[116], stage1_7[117], stage1_7[118], stage1_7[119], stage1_7[120]},
      {stage1_8[177]},
      {stage1_9[18], stage1_9[19], stage1_9[20], stage1_9[21], stage1_9[22], stage1_9[23]},
      {stage2_11[3],stage2_10[32],stage2_9[47],stage2_8[61],stage2_7[79]}
   );
   gpc615_5 gpc2386 (
      {stage1_7[121], stage1_7[122], stage1_7[123], stage1_7[124], stage1_7[125]},
      {stage1_8[178]},
      {stage1_9[24], stage1_9[25], stage1_9[26], stage1_9[27], stage1_9[28], stage1_9[29]},
      {stage2_11[4],stage2_10[33],stage2_9[48],stage2_8[62],stage2_7[80]}
   );
   gpc615_5 gpc2387 (
      {stage1_7[126], stage1_7[127], stage1_7[128], stage1_7[129], stage1_7[130]},
      {stage1_8[179]},
      {stage1_9[30], stage1_9[31], stage1_9[32], stage1_9[33], stage1_9[34], stage1_9[35]},
      {stage2_11[5],stage2_10[34],stage2_9[49],stage2_8[63],stage2_7[81]}
   );
   gpc615_5 gpc2388 (
      {stage1_7[131], stage1_7[132], stage1_7[133], stage1_7[134], stage1_7[135]},
      {stage1_8[180]},
      {stage1_9[36], stage1_9[37], stage1_9[38], stage1_9[39], stage1_9[40], stage1_9[41]},
      {stage2_11[6],stage2_10[35],stage2_9[50],stage2_8[64],stage2_7[82]}
   );
   gpc615_5 gpc2389 (
      {stage1_7[136], stage1_7[137], stage1_7[138], stage1_7[139], stage1_7[140]},
      {stage1_8[181]},
      {stage1_9[42], stage1_9[43], stage1_9[44], stage1_9[45], stage1_9[46], stage1_9[47]},
      {stage2_11[7],stage2_10[36],stage2_9[51],stage2_8[65],stage2_7[83]}
   );
   gpc615_5 gpc2390 (
      {stage1_7[141], stage1_7[142], stage1_7[143], stage1_7[144], stage1_7[145]},
      {stage1_8[182]},
      {stage1_9[48], stage1_9[49], stage1_9[50], stage1_9[51], stage1_9[52], stage1_9[53]},
      {stage2_11[8],stage2_10[37],stage2_9[52],stage2_8[66],stage2_7[84]}
   );
   gpc615_5 gpc2391 (
      {stage1_7[146], stage1_7[147], stage1_7[148], stage1_7[149], stage1_7[150]},
      {stage1_8[183]},
      {stage1_9[54], stage1_9[55], stage1_9[56], stage1_9[57], stage1_9[58], stage1_9[59]},
      {stage2_11[9],stage2_10[38],stage2_9[53],stage2_8[67],stage2_7[85]}
   );
   gpc615_5 gpc2392 (
      {stage1_7[151], stage1_7[152], stage1_7[153], stage1_7[154], stage1_7[155]},
      {stage1_8[184]},
      {stage1_9[60], stage1_9[61], stage1_9[62], stage1_9[63], stage1_9[64], stage1_9[65]},
      {stage2_11[10],stage2_10[39],stage2_9[54],stage2_8[68],stage2_7[86]}
   );
   gpc615_5 gpc2393 (
      {stage1_7[156], stage1_7[157], stage1_7[158], stage1_7[159], stage1_7[160]},
      {stage1_8[185]},
      {stage1_9[66], stage1_9[67], stage1_9[68], stage1_9[69], stage1_9[70], stage1_9[71]},
      {stage2_11[11],stage2_10[40],stage2_9[55],stage2_8[69],stage2_7[87]}
   );
   gpc615_5 gpc2394 (
      {stage1_7[161], stage1_7[162], stage1_7[163], stage1_7[164], stage1_7[165]},
      {stage1_8[186]},
      {stage1_9[72], stage1_9[73], stage1_9[74], stage1_9[75], stage1_9[76], stage1_9[77]},
      {stage2_11[12],stage2_10[41],stage2_9[56],stage2_8[70],stage2_7[88]}
   );
   gpc606_5 gpc2395 (
      {stage1_8[187], stage1_8[188], stage1_8[189], stage1_8[190], stage1_8[191], stage1_8[192]},
      {stage1_10[0], stage1_10[1], stage1_10[2], stage1_10[3], stage1_10[4], stage1_10[5]},
      {stage2_12[0],stage2_11[13],stage2_10[42],stage2_9[57],stage2_8[71]}
   );
   gpc606_5 gpc2396 (
      {stage1_8[193], stage1_8[194], stage1_8[195], stage1_8[196], stage1_8[197], stage1_8[198]},
      {stage1_10[6], stage1_10[7], stage1_10[8], stage1_10[9], stage1_10[10], stage1_10[11]},
      {stage2_12[1],stage2_11[14],stage2_10[43],stage2_9[58],stage2_8[72]}
   );
   gpc606_5 gpc2397 (
      {stage1_8[199], stage1_8[200], stage1_8[201], stage1_8[202], stage1_8[203], stage1_8[204]},
      {stage1_10[12], stage1_10[13], stage1_10[14], stage1_10[15], stage1_10[16], stage1_10[17]},
      {stage2_12[2],stage2_11[15],stage2_10[44],stage2_9[59],stage2_8[73]}
   );
   gpc606_5 gpc2398 (
      {stage1_8[205], stage1_8[206], stage1_8[207], stage1_8[208], stage1_8[209], stage1_8[210]},
      {stage1_10[18], stage1_10[19], stage1_10[20], stage1_10[21], stage1_10[22], stage1_10[23]},
      {stage2_12[3],stage2_11[16],stage2_10[45],stage2_9[60],stage2_8[74]}
   );
   gpc606_5 gpc2399 (
      {stage1_8[211], stage1_8[212], stage1_8[213], stage1_8[214], stage1_8[215], stage1_8[216]},
      {stage1_10[24], stage1_10[25], stage1_10[26], stage1_10[27], stage1_10[28], stage1_10[29]},
      {stage2_12[4],stage2_11[17],stage2_10[46],stage2_9[61],stage2_8[75]}
   );
   gpc606_5 gpc2400 (
      {stage1_8[217], stage1_8[218], stage1_8[219], stage1_8[220], stage1_8[221], stage1_8[222]},
      {stage1_10[30], stage1_10[31], stage1_10[32], stage1_10[33], stage1_10[34], stage1_10[35]},
      {stage2_12[5],stage2_11[18],stage2_10[47],stage2_9[62],stage2_8[76]}
   );
   gpc606_5 gpc2401 (
      {stage1_8[223], stage1_8[224], stage1_8[225], stage1_8[226], stage1_8[227], stage1_8[228]},
      {stage1_10[36], stage1_10[37], stage1_10[38], stage1_10[39], stage1_10[40], stage1_10[41]},
      {stage2_12[6],stage2_11[19],stage2_10[48],stage2_9[63],stage2_8[77]}
   );
   gpc606_5 gpc2402 (
      {stage1_8[229], stage1_8[230], stage1_8[231], stage1_8[232], stage1_8[233], stage1_8[234]},
      {stage1_10[42], stage1_10[43], stage1_10[44], stage1_10[45], stage1_10[46], stage1_10[47]},
      {stage2_12[7],stage2_11[20],stage2_10[49],stage2_9[64],stage2_8[78]}
   );
   gpc606_5 gpc2403 (
      {stage1_8[235], stage1_8[236], stage1_8[237], stage1_8[238], stage1_8[239], stage1_8[240]},
      {stage1_10[48], stage1_10[49], stage1_10[50], stage1_10[51], stage1_10[52], stage1_10[53]},
      {stage2_12[8],stage2_11[21],stage2_10[50],stage2_9[65],stage2_8[79]}
   );
   gpc606_5 gpc2404 (
      {stage1_8[241], stage1_8[242], stage1_8[243], stage1_8[244], stage1_8[245], stage1_8[246]},
      {stage1_10[54], stage1_10[55], stage1_10[56], stage1_10[57], stage1_10[58], stage1_10[59]},
      {stage2_12[9],stage2_11[22],stage2_10[51],stage2_9[66],stage2_8[80]}
   );
   gpc606_5 gpc2405 (
      {stage1_8[247], stage1_8[248], stage1_8[249], stage1_8[250], stage1_8[251], stage1_8[252]},
      {stage1_10[60], stage1_10[61], stage1_10[62], stage1_10[63], stage1_10[64], stage1_10[65]},
      {stage2_12[10],stage2_11[23],stage2_10[52],stage2_9[67],stage2_8[81]}
   );
   gpc606_5 gpc2406 (
      {stage1_8[253], stage1_8[254], stage1_8[255], stage1_8[256], stage1_8[257], stage1_8[258]},
      {stage1_10[66], stage1_10[67], stage1_10[68], stage1_10[69], stage1_10[70], stage1_10[71]},
      {stage2_12[11],stage2_11[24],stage2_10[53],stage2_9[68],stage2_8[82]}
   );
   gpc606_5 gpc2407 (
      {stage1_8[259], stage1_8[260], stage1_8[261], stage1_8[262], stage1_8[263], stage1_8[264]},
      {stage1_10[72], stage1_10[73], stage1_10[74], stage1_10[75], stage1_10[76], stage1_10[77]},
      {stage2_12[12],stage2_11[25],stage2_10[54],stage2_9[69],stage2_8[83]}
   );
   gpc606_5 gpc2408 (
      {stage1_8[265], stage1_8[266], stage1_8[267], stage1_8[268], stage1_8[269], stage1_8[270]},
      {stage1_10[78], stage1_10[79], stage1_10[80], stage1_10[81], stage1_10[82], stage1_10[83]},
      {stage2_12[13],stage2_11[26],stage2_10[55],stage2_9[70],stage2_8[84]}
   );
   gpc606_5 gpc2409 (
      {stage1_8[271], stage1_8[272], stage1_8[273], stage1_8[274], stage1_8[275], stage1_8[276]},
      {stage1_10[84], stage1_10[85], stage1_10[86], stage1_10[87], stage1_10[88], stage1_10[89]},
      {stage2_12[14],stage2_11[27],stage2_10[56],stage2_9[71],stage2_8[85]}
   );
   gpc606_5 gpc2410 (
      {stage1_8[277], stage1_8[278], stage1_8[279], stage1_8[280], stage1_8[281], stage1_8[282]},
      {stage1_10[90], stage1_10[91], stage1_10[92], stage1_10[93], stage1_10[94], stage1_10[95]},
      {stage2_12[15],stage2_11[28],stage2_10[57],stage2_9[72],stage2_8[86]}
   );
   gpc606_5 gpc2411 (
      {stage1_8[283], stage1_8[284], stage1_8[285], stage1_8[286], stage1_8[287], stage1_8[288]},
      {stage1_10[96], stage1_10[97], stage1_10[98], stage1_10[99], stage1_10[100], stage1_10[101]},
      {stage2_12[16],stage2_11[29],stage2_10[58],stage2_9[73],stage2_8[87]}
   );
   gpc606_5 gpc2412 (
      {stage1_8[289], stage1_8[290], stage1_8[291], stage1_8[292], stage1_8[293], stage1_8[294]},
      {stage1_10[102], stage1_10[103], stage1_10[104], stage1_10[105], stage1_10[106], stage1_10[107]},
      {stage2_12[17],stage2_11[30],stage2_10[59],stage2_9[74],stage2_8[88]}
   );
   gpc606_5 gpc2413 (
      {stage1_8[295], stage1_8[296], stage1_8[297], stage1_8[298], stage1_8[299], stage1_8[300]},
      {stage1_10[108], stage1_10[109], stage1_10[110], stage1_10[111], stage1_10[112], stage1_10[113]},
      {stage2_12[18],stage2_11[31],stage2_10[60],stage2_9[75],stage2_8[89]}
   );
   gpc606_5 gpc2414 (
      {stage1_8[301], stage1_8[302], stage1_8[303], stage1_8[304], stage1_8[305], stage1_8[306]},
      {stage1_10[114], stage1_10[115], stage1_10[116], stage1_10[117], stage1_10[118], stage1_10[119]},
      {stage2_12[19],stage2_11[32],stage2_10[61],stage2_9[76],stage2_8[90]}
   );
   gpc606_5 gpc2415 (
      {stage1_8[307], stage1_8[308], stage1_8[309], stage1_8[310], stage1_8[311], stage1_8[312]},
      {stage1_10[120], stage1_10[121], stage1_10[122], stage1_10[123], stage1_10[124], stage1_10[125]},
      {stage2_12[20],stage2_11[33],stage2_10[62],stage2_9[77],stage2_8[91]}
   );
   gpc606_5 gpc2416 (
      {stage1_8[313], stage1_8[314], stage1_8[315], stage1_8[316], stage1_8[317], stage1_8[318]},
      {stage1_10[126], stage1_10[127], stage1_10[128], stage1_10[129], stage1_10[130], stage1_10[131]},
      {stage2_12[21],stage2_11[34],stage2_10[63],stage2_9[78],stage2_8[92]}
   );
   gpc606_5 gpc2417 (
      {stage1_8[319], stage1_8[320], stage1_8[321], stage1_8[322], stage1_8[323], stage1_8[324]},
      {stage1_10[132], stage1_10[133], stage1_10[134], stage1_10[135], stage1_10[136], stage1_10[137]},
      {stage2_12[22],stage2_11[35],stage2_10[64],stage2_9[79],stage2_8[93]}
   );
   gpc606_5 gpc2418 (
      {stage1_8[325], stage1_8[326], stage1_8[327], stage1_8[328], stage1_8[329], stage1_8[330]},
      {stage1_10[138], stage1_10[139], stage1_10[140], stage1_10[141], stage1_10[142], stage1_10[143]},
      {stage2_12[23],stage2_11[36],stage2_10[65],stage2_9[80],stage2_8[94]}
   );
   gpc606_5 gpc2419 (
      {stage1_8[331], stage1_8[332], stage1_8[333], stage1_8[334], stage1_8[335], stage1_8[336]},
      {stage1_10[144], stage1_10[145], stage1_10[146], stage1_10[147], stage1_10[148], stage1_10[149]},
      {stage2_12[24],stage2_11[37],stage2_10[66],stage2_9[81],stage2_8[95]}
   );
   gpc606_5 gpc2420 (
      {stage1_8[337], stage1_8[338], stage1_8[339], stage1_8[340], stage1_8[341], stage1_8[342]},
      {stage1_10[150], stage1_10[151], stage1_10[152], stage1_10[153], stage1_10[154], stage1_10[155]},
      {stage2_12[25],stage2_11[38],stage2_10[67],stage2_9[82],stage2_8[96]}
   );
   gpc606_5 gpc2421 (
      {stage1_8[343], stage1_8[344], stage1_8[345], stage1_8[346], stage1_8[347], stage1_8[348]},
      {stage1_10[156], stage1_10[157], stage1_10[158], stage1_10[159], stage1_10[160], stage1_10[161]},
      {stage2_12[26],stage2_11[39],stage2_10[68],stage2_9[83],stage2_8[97]}
   );
   gpc606_5 gpc2422 (
      {stage1_9[78], stage1_9[79], stage1_9[80], stage1_9[81], stage1_9[82], stage1_9[83]},
      {stage1_11[0], stage1_11[1], stage1_11[2], stage1_11[3], stage1_11[4], stage1_11[5]},
      {stage2_13[0],stage2_12[27],stage2_11[40],stage2_10[69],stage2_9[84]}
   );
   gpc606_5 gpc2423 (
      {stage1_9[84], stage1_9[85], stage1_9[86], stage1_9[87], stage1_9[88], stage1_9[89]},
      {stage1_11[6], stage1_11[7], stage1_11[8], stage1_11[9], stage1_11[10], stage1_11[11]},
      {stage2_13[1],stage2_12[28],stage2_11[41],stage2_10[70],stage2_9[85]}
   );
   gpc606_5 gpc2424 (
      {stage1_9[90], stage1_9[91], stage1_9[92], stage1_9[93], stage1_9[94], stage1_9[95]},
      {stage1_11[12], stage1_11[13], stage1_11[14], stage1_11[15], stage1_11[16], stage1_11[17]},
      {stage2_13[2],stage2_12[29],stage2_11[42],stage2_10[71],stage2_9[86]}
   );
   gpc606_5 gpc2425 (
      {stage1_9[96], stage1_9[97], stage1_9[98], stage1_9[99], stage1_9[100], stage1_9[101]},
      {stage1_11[18], stage1_11[19], stage1_11[20], stage1_11[21], stage1_11[22], stage1_11[23]},
      {stage2_13[3],stage2_12[30],stage2_11[43],stage2_10[72],stage2_9[87]}
   );
   gpc606_5 gpc2426 (
      {stage1_9[102], stage1_9[103], stage1_9[104], stage1_9[105], stage1_9[106], stage1_9[107]},
      {stage1_11[24], stage1_11[25], stage1_11[26], stage1_11[27], stage1_11[28], stage1_11[29]},
      {stage2_13[4],stage2_12[31],stage2_11[44],stage2_10[73],stage2_9[88]}
   );
   gpc606_5 gpc2427 (
      {stage1_9[108], stage1_9[109], stage1_9[110], stage1_9[111], stage1_9[112], stage1_9[113]},
      {stage1_11[30], stage1_11[31], stage1_11[32], stage1_11[33], stage1_11[34], stage1_11[35]},
      {stage2_13[5],stage2_12[32],stage2_11[45],stage2_10[74],stage2_9[89]}
   );
   gpc606_5 gpc2428 (
      {stage1_9[114], stage1_9[115], stage1_9[116], stage1_9[117], stage1_9[118], stage1_9[119]},
      {stage1_11[36], stage1_11[37], stage1_11[38], stage1_11[39], stage1_11[40], stage1_11[41]},
      {stage2_13[6],stage2_12[33],stage2_11[46],stage2_10[75],stage2_9[90]}
   );
   gpc606_5 gpc2429 (
      {stage1_9[120], stage1_9[121], stage1_9[122], stage1_9[123], stage1_9[124], stage1_9[125]},
      {stage1_11[42], stage1_11[43], stage1_11[44], stage1_11[45], stage1_11[46], stage1_11[47]},
      {stage2_13[7],stage2_12[34],stage2_11[47],stage2_10[76],stage2_9[91]}
   );
   gpc606_5 gpc2430 (
      {stage1_9[126], stage1_9[127], stage1_9[128], stage1_9[129], stage1_9[130], stage1_9[131]},
      {stage1_11[48], stage1_11[49], stage1_11[50], stage1_11[51], stage1_11[52], stage1_11[53]},
      {stage2_13[8],stage2_12[35],stage2_11[48],stage2_10[77],stage2_9[92]}
   );
   gpc606_5 gpc2431 (
      {stage1_9[132], stage1_9[133], stage1_9[134], stage1_9[135], stage1_9[136], stage1_9[137]},
      {stage1_11[54], stage1_11[55], stage1_11[56], stage1_11[57], stage1_11[58], stage1_11[59]},
      {stage2_13[9],stage2_12[36],stage2_11[49],stage2_10[78],stage2_9[93]}
   );
   gpc606_5 gpc2432 (
      {stage1_9[138], stage1_9[139], stage1_9[140], stage1_9[141], stage1_9[142], stage1_9[143]},
      {stage1_11[60], stage1_11[61], stage1_11[62], stage1_11[63], stage1_11[64], stage1_11[65]},
      {stage2_13[10],stage2_12[37],stage2_11[50],stage2_10[79],stage2_9[94]}
   );
   gpc606_5 gpc2433 (
      {stage1_9[144], stage1_9[145], stage1_9[146], stage1_9[147], stage1_9[148], stage1_9[149]},
      {stage1_11[66], stage1_11[67], stage1_11[68], stage1_11[69], stage1_11[70], stage1_11[71]},
      {stage2_13[11],stage2_12[38],stage2_11[51],stage2_10[80],stage2_9[95]}
   );
   gpc606_5 gpc2434 (
      {stage1_9[150], stage1_9[151], stage1_9[152], stage1_9[153], stage1_9[154], stage1_9[155]},
      {stage1_11[72], stage1_11[73], stage1_11[74], stage1_11[75], stage1_11[76], stage1_11[77]},
      {stage2_13[12],stage2_12[39],stage2_11[52],stage2_10[81],stage2_9[96]}
   );
   gpc606_5 gpc2435 (
      {stage1_9[156], stage1_9[157], stage1_9[158], stage1_9[159], stage1_9[160], stage1_9[161]},
      {stage1_11[78], stage1_11[79], stage1_11[80], stage1_11[81], stage1_11[82], stage1_11[83]},
      {stage2_13[13],stage2_12[40],stage2_11[53],stage2_10[82],stage2_9[97]}
   );
   gpc606_5 gpc2436 (
      {stage1_9[162], stage1_9[163], stage1_9[164], stage1_9[165], stage1_9[166], stage1_9[167]},
      {stage1_11[84], stage1_11[85], stage1_11[86], stage1_11[87], stage1_11[88], stage1_11[89]},
      {stage2_13[14],stage2_12[41],stage2_11[54],stage2_10[83],stage2_9[98]}
   );
   gpc606_5 gpc2437 (
      {stage1_9[168], stage1_9[169], stage1_9[170], stage1_9[171], stage1_9[172], stage1_9[173]},
      {stage1_11[90], stage1_11[91], stage1_11[92], stage1_11[93], stage1_11[94], stage1_11[95]},
      {stage2_13[15],stage2_12[42],stage2_11[55],stage2_10[84],stage2_9[99]}
   );
   gpc606_5 gpc2438 (
      {stage1_9[174], stage1_9[175], stage1_9[176], stage1_9[177], stage1_9[178], stage1_9[179]},
      {stage1_11[96], stage1_11[97], stage1_11[98], stage1_11[99], stage1_11[100], stage1_11[101]},
      {stage2_13[16],stage2_12[43],stage2_11[56],stage2_10[85],stage2_9[100]}
   );
   gpc606_5 gpc2439 (
      {stage1_9[180], stage1_9[181], stage1_9[182], stage1_9[183], stage1_9[184], stage1_9[185]},
      {stage1_11[102], stage1_11[103], stage1_11[104], stage1_11[105], stage1_11[106], stage1_11[107]},
      {stage2_13[17],stage2_12[44],stage2_11[57],stage2_10[86],stage2_9[101]}
   );
   gpc606_5 gpc2440 (
      {stage1_9[186], stage1_9[187], stage1_9[188], stage1_9[189], stage1_9[190], stage1_9[191]},
      {stage1_11[108], stage1_11[109], stage1_11[110], stage1_11[111], stage1_11[112], stage1_11[113]},
      {stage2_13[18],stage2_12[45],stage2_11[58],stage2_10[87],stage2_9[102]}
   );
   gpc606_5 gpc2441 (
      {stage1_9[192], stage1_9[193], stage1_9[194], stage1_9[195], stage1_9[196], stage1_9[197]},
      {stage1_11[114], stage1_11[115], stage1_11[116], stage1_11[117], stage1_11[118], stage1_11[119]},
      {stage2_13[19],stage2_12[46],stage2_11[59],stage2_10[88],stage2_9[103]}
   );
   gpc606_5 gpc2442 (
      {stage1_9[198], stage1_9[199], stage1_9[200], stage1_9[201], stage1_9[202], stage1_9[203]},
      {stage1_11[120], stage1_11[121], stage1_11[122], stage1_11[123], stage1_11[124], stage1_11[125]},
      {stage2_13[20],stage2_12[47],stage2_11[60],stage2_10[89],stage2_9[104]}
   );
   gpc606_5 gpc2443 (
      {stage1_9[204], stage1_9[205], stage1_9[206], stage1_9[207], stage1_9[208], stage1_9[209]},
      {stage1_11[126], stage1_11[127], stage1_11[128], stage1_11[129], stage1_11[130], stage1_11[131]},
      {stage2_13[21],stage2_12[48],stage2_11[61],stage2_10[90],stage2_9[105]}
   );
   gpc615_5 gpc2444 (
      {stage1_10[162], stage1_10[163], stage1_10[164], stage1_10[165], stage1_10[166]},
      {stage1_11[132]},
      {stage1_12[0], stage1_12[1], stage1_12[2], stage1_12[3], stage1_12[4], stage1_12[5]},
      {stage2_14[0],stage2_13[22],stage2_12[49],stage2_11[62],stage2_10[91]}
   );
   gpc615_5 gpc2445 (
      {stage1_10[167], stage1_10[168], stage1_10[169], stage1_10[170], stage1_10[171]},
      {stage1_11[133]},
      {stage1_12[6], stage1_12[7], stage1_12[8], stage1_12[9], stage1_12[10], stage1_12[11]},
      {stage2_14[1],stage2_13[23],stage2_12[50],stage2_11[63],stage2_10[92]}
   );
   gpc615_5 gpc2446 (
      {stage1_10[172], stage1_10[173], stage1_10[174], stage1_10[175], stage1_10[176]},
      {stage1_11[134]},
      {stage1_12[12], stage1_12[13], stage1_12[14], stage1_12[15], stage1_12[16], stage1_12[17]},
      {stage2_14[2],stage2_13[24],stage2_12[51],stage2_11[64],stage2_10[93]}
   );
   gpc615_5 gpc2447 (
      {stage1_10[177], stage1_10[178], stage1_10[179], stage1_10[180], stage1_10[181]},
      {stage1_11[135]},
      {stage1_12[18], stage1_12[19], stage1_12[20], stage1_12[21], stage1_12[22], stage1_12[23]},
      {stage2_14[3],stage2_13[25],stage2_12[52],stage2_11[65],stage2_10[94]}
   );
   gpc615_5 gpc2448 (
      {stage1_11[136], stage1_11[137], stage1_11[138], stage1_11[139], stage1_11[140]},
      {stage1_12[24]},
      {stage1_13[0], stage1_13[1], stage1_13[2], stage1_13[3], stage1_13[4], stage1_13[5]},
      {stage2_15[0],stage2_14[4],stage2_13[26],stage2_12[53],stage2_11[66]}
   );
   gpc615_5 gpc2449 (
      {stage1_11[141], stage1_11[142], stage1_11[143], stage1_11[144], stage1_11[145]},
      {stage1_12[25]},
      {stage1_13[6], stage1_13[7], stage1_13[8], stage1_13[9], stage1_13[10], stage1_13[11]},
      {stage2_15[1],stage2_14[5],stage2_13[27],stage2_12[54],stage2_11[67]}
   );
   gpc615_5 gpc2450 (
      {stage1_11[146], stage1_11[147], stage1_11[148], stage1_11[149], stage1_11[150]},
      {stage1_12[26]},
      {stage1_13[12], stage1_13[13], stage1_13[14], stage1_13[15], stage1_13[16], stage1_13[17]},
      {stage2_15[2],stage2_14[6],stage2_13[28],stage2_12[55],stage2_11[68]}
   );
   gpc615_5 gpc2451 (
      {stage1_11[151], stage1_11[152], stage1_11[153], stage1_11[154], stage1_11[155]},
      {stage1_12[27]},
      {stage1_13[18], stage1_13[19], stage1_13[20], stage1_13[21], stage1_13[22], stage1_13[23]},
      {stage2_15[3],stage2_14[7],stage2_13[29],stage2_12[56],stage2_11[69]}
   );
   gpc615_5 gpc2452 (
      {stage1_11[156], stage1_11[157], stage1_11[158], stage1_11[159], stage1_11[160]},
      {stage1_12[28]},
      {stage1_13[24], stage1_13[25], stage1_13[26], stage1_13[27], stage1_13[28], stage1_13[29]},
      {stage2_15[4],stage2_14[8],stage2_13[30],stage2_12[57],stage2_11[70]}
   );
   gpc606_5 gpc2453 (
      {stage1_12[29], stage1_12[30], stage1_12[31], stage1_12[32], stage1_12[33], stage1_12[34]},
      {stage1_14[0], stage1_14[1], stage1_14[2], stage1_14[3], stage1_14[4], stage1_14[5]},
      {stage2_16[0],stage2_15[5],stage2_14[9],stage2_13[31],stage2_12[58]}
   );
   gpc615_5 gpc2454 (
      {stage1_12[35], stage1_12[36], stage1_12[37], stage1_12[38], stage1_12[39]},
      {stage1_13[30]},
      {stage1_14[6], stage1_14[7], stage1_14[8], stage1_14[9], stage1_14[10], stage1_14[11]},
      {stage2_16[1],stage2_15[6],stage2_14[10],stage2_13[32],stage2_12[59]}
   );
   gpc615_5 gpc2455 (
      {stage1_12[40], stage1_12[41], stage1_12[42], stage1_12[43], stage1_12[44]},
      {stage1_13[31]},
      {stage1_14[12], stage1_14[13], stage1_14[14], stage1_14[15], stage1_14[16], stage1_14[17]},
      {stage2_16[2],stage2_15[7],stage2_14[11],stage2_13[33],stage2_12[60]}
   );
   gpc615_5 gpc2456 (
      {stage1_12[45], stage1_12[46], stage1_12[47], stage1_12[48], stage1_12[49]},
      {stage1_13[32]},
      {stage1_14[18], stage1_14[19], stage1_14[20], stage1_14[21], stage1_14[22], stage1_14[23]},
      {stage2_16[3],stage2_15[8],stage2_14[12],stage2_13[34],stage2_12[61]}
   );
   gpc615_5 gpc2457 (
      {stage1_12[50], stage1_12[51], stage1_12[52], stage1_12[53], stage1_12[54]},
      {stage1_13[33]},
      {stage1_14[24], stage1_14[25], stage1_14[26], stage1_14[27], stage1_14[28], stage1_14[29]},
      {stage2_16[4],stage2_15[9],stage2_14[13],stage2_13[35],stage2_12[62]}
   );
   gpc615_5 gpc2458 (
      {stage1_12[55], stage1_12[56], stage1_12[57], stage1_12[58], stage1_12[59]},
      {stage1_13[34]},
      {stage1_14[30], stage1_14[31], stage1_14[32], stage1_14[33], stage1_14[34], stage1_14[35]},
      {stage2_16[5],stage2_15[10],stage2_14[14],stage2_13[36],stage2_12[63]}
   );
   gpc615_5 gpc2459 (
      {stage1_12[60], stage1_12[61], stage1_12[62], stage1_12[63], stage1_12[64]},
      {stage1_13[35]},
      {stage1_14[36], stage1_14[37], stage1_14[38], stage1_14[39], stage1_14[40], stage1_14[41]},
      {stage2_16[6],stage2_15[11],stage2_14[15],stage2_13[37],stage2_12[64]}
   );
   gpc615_5 gpc2460 (
      {stage1_12[65], stage1_12[66], stage1_12[67], stage1_12[68], stage1_12[69]},
      {stage1_13[36]},
      {stage1_14[42], stage1_14[43], stage1_14[44], stage1_14[45], stage1_14[46], stage1_14[47]},
      {stage2_16[7],stage2_15[12],stage2_14[16],stage2_13[38],stage2_12[65]}
   );
   gpc615_5 gpc2461 (
      {stage1_12[70], stage1_12[71], stage1_12[72], stage1_12[73], stage1_12[74]},
      {stage1_13[37]},
      {stage1_14[48], stage1_14[49], stage1_14[50], stage1_14[51], stage1_14[52], stage1_14[53]},
      {stage2_16[8],stage2_15[13],stage2_14[17],stage2_13[39],stage2_12[66]}
   );
   gpc615_5 gpc2462 (
      {stage1_12[75], stage1_12[76], stage1_12[77], stage1_12[78], stage1_12[79]},
      {stage1_13[38]},
      {stage1_14[54], stage1_14[55], stage1_14[56], stage1_14[57], stage1_14[58], stage1_14[59]},
      {stage2_16[9],stage2_15[14],stage2_14[18],stage2_13[40],stage2_12[67]}
   );
   gpc615_5 gpc2463 (
      {stage1_12[80], stage1_12[81], stage1_12[82], stage1_12[83], stage1_12[84]},
      {stage1_13[39]},
      {stage1_14[60], stage1_14[61], stage1_14[62], stage1_14[63], stage1_14[64], stage1_14[65]},
      {stage2_16[10],stage2_15[15],stage2_14[19],stage2_13[41],stage2_12[68]}
   );
   gpc615_5 gpc2464 (
      {stage1_12[85], stage1_12[86], stage1_12[87], stage1_12[88], stage1_12[89]},
      {stage1_13[40]},
      {stage1_14[66], stage1_14[67], stage1_14[68], stage1_14[69], stage1_14[70], stage1_14[71]},
      {stage2_16[11],stage2_15[16],stage2_14[20],stage2_13[42],stage2_12[69]}
   );
   gpc615_5 gpc2465 (
      {stage1_12[90], stage1_12[91], stage1_12[92], stage1_12[93], stage1_12[94]},
      {stage1_13[41]},
      {stage1_14[72], stage1_14[73], stage1_14[74], stage1_14[75], stage1_14[76], stage1_14[77]},
      {stage2_16[12],stage2_15[17],stage2_14[21],stage2_13[43],stage2_12[70]}
   );
   gpc615_5 gpc2466 (
      {stage1_12[95], stage1_12[96], stage1_12[97], stage1_12[98], stage1_12[99]},
      {stage1_13[42]},
      {stage1_14[78], stage1_14[79], stage1_14[80], stage1_14[81], stage1_14[82], stage1_14[83]},
      {stage2_16[13],stage2_15[18],stage2_14[22],stage2_13[44],stage2_12[71]}
   );
   gpc615_5 gpc2467 (
      {stage1_12[100], stage1_12[101], stage1_12[102], stage1_12[103], stage1_12[104]},
      {stage1_13[43]},
      {stage1_14[84], stage1_14[85], stage1_14[86], stage1_14[87], stage1_14[88], stage1_14[89]},
      {stage2_16[14],stage2_15[19],stage2_14[23],stage2_13[45],stage2_12[72]}
   );
   gpc615_5 gpc2468 (
      {stage1_12[105], stage1_12[106], stage1_12[107], stage1_12[108], stage1_12[109]},
      {stage1_13[44]},
      {stage1_14[90], stage1_14[91], stage1_14[92], stage1_14[93], stage1_14[94], stage1_14[95]},
      {stage2_16[15],stage2_15[20],stage2_14[24],stage2_13[46],stage2_12[73]}
   );
   gpc615_5 gpc2469 (
      {stage1_12[110], stage1_12[111], stage1_12[112], stage1_12[113], stage1_12[114]},
      {stage1_13[45]},
      {stage1_14[96], stage1_14[97], stage1_14[98], stage1_14[99], stage1_14[100], stage1_14[101]},
      {stage2_16[16],stage2_15[21],stage2_14[25],stage2_13[47],stage2_12[74]}
   );
   gpc615_5 gpc2470 (
      {stage1_12[115], stage1_12[116], stage1_12[117], stage1_12[118], stage1_12[119]},
      {stage1_13[46]},
      {stage1_14[102], stage1_14[103], stage1_14[104], stage1_14[105], stage1_14[106], stage1_14[107]},
      {stage2_16[17],stage2_15[22],stage2_14[26],stage2_13[48],stage2_12[75]}
   );
   gpc615_5 gpc2471 (
      {stage1_12[120], stage1_12[121], stage1_12[122], stage1_12[123], stage1_12[124]},
      {stage1_13[47]},
      {stage1_14[108], stage1_14[109], stage1_14[110], stage1_14[111], stage1_14[112], stage1_14[113]},
      {stage2_16[18],stage2_15[23],stage2_14[27],stage2_13[49],stage2_12[76]}
   );
   gpc615_5 gpc2472 (
      {stage1_12[125], stage1_12[126], stage1_12[127], stage1_12[128], stage1_12[129]},
      {stage1_13[48]},
      {stage1_14[114], stage1_14[115], stage1_14[116], stage1_14[117], stage1_14[118], stage1_14[119]},
      {stage2_16[19],stage2_15[24],stage2_14[28],stage2_13[50],stage2_12[77]}
   );
   gpc615_5 gpc2473 (
      {stage1_12[130], stage1_12[131], stage1_12[132], stage1_12[133], stage1_12[134]},
      {stage1_13[49]},
      {stage1_14[120], stage1_14[121], stage1_14[122], stage1_14[123], stage1_14[124], stage1_14[125]},
      {stage2_16[20],stage2_15[25],stage2_14[29],stage2_13[51],stage2_12[78]}
   );
   gpc615_5 gpc2474 (
      {stage1_12[135], stage1_12[136], stage1_12[137], stage1_12[138], stage1_12[139]},
      {stage1_13[50]},
      {stage1_14[126], stage1_14[127], stage1_14[128], stage1_14[129], stage1_14[130], stage1_14[131]},
      {stage2_16[21],stage2_15[26],stage2_14[30],stage2_13[52],stage2_12[79]}
   );
   gpc615_5 gpc2475 (
      {stage1_12[140], stage1_12[141], stage1_12[142], stage1_12[143], stage1_12[144]},
      {stage1_13[51]},
      {stage1_14[132], stage1_14[133], stage1_14[134], stage1_14[135], stage1_14[136], stage1_14[137]},
      {stage2_16[22],stage2_15[27],stage2_14[31],stage2_13[53],stage2_12[80]}
   );
   gpc615_5 gpc2476 (
      {stage1_12[145], stage1_12[146], stage1_12[147], stage1_12[148], stage1_12[149]},
      {stage1_13[52]},
      {stage1_14[138], stage1_14[139], stage1_14[140], stage1_14[141], stage1_14[142], stage1_14[143]},
      {stage2_16[23],stage2_15[28],stage2_14[32],stage2_13[54],stage2_12[81]}
   );
   gpc615_5 gpc2477 (
      {stage1_12[150], stage1_12[151], stage1_12[152], stage1_12[153], stage1_12[154]},
      {stage1_13[53]},
      {stage1_14[144], stage1_14[145], stage1_14[146], stage1_14[147], stage1_14[148], stage1_14[149]},
      {stage2_16[24],stage2_15[29],stage2_14[33],stage2_13[55],stage2_12[82]}
   );
   gpc615_5 gpc2478 (
      {stage1_12[155], stage1_12[156], stage1_12[157], stage1_12[158], stage1_12[159]},
      {stage1_13[54]},
      {stage1_14[150], stage1_14[151], stage1_14[152], stage1_14[153], stage1_14[154], stage1_14[155]},
      {stage2_16[25],stage2_15[30],stage2_14[34],stage2_13[56],stage2_12[83]}
   );
   gpc615_5 gpc2479 (
      {stage1_12[160], stage1_12[161], stage1_12[162], stage1_12[163], stage1_12[164]},
      {stage1_13[55]},
      {stage1_14[156], stage1_14[157], stage1_14[158], stage1_14[159], stage1_14[160], stage1_14[161]},
      {stage2_16[26],stage2_15[31],stage2_14[35],stage2_13[57],stage2_12[84]}
   );
   gpc615_5 gpc2480 (
      {stage1_12[165], stage1_12[166], stage1_12[167], stage1_12[168], stage1_12[169]},
      {stage1_13[56]},
      {stage1_14[162], stage1_14[163], stage1_14[164], stage1_14[165], stage1_14[166], stage1_14[167]},
      {stage2_16[27],stage2_15[32],stage2_14[36],stage2_13[58],stage2_12[85]}
   );
   gpc615_5 gpc2481 (
      {stage1_12[170], stage1_12[171], stage1_12[172], stage1_12[173], stage1_12[174]},
      {stage1_13[57]},
      {stage1_14[168], stage1_14[169], stage1_14[170], stage1_14[171], stage1_14[172], stage1_14[173]},
      {stage2_16[28],stage2_15[33],stage2_14[37],stage2_13[59],stage2_12[86]}
   );
   gpc615_5 gpc2482 (
      {stage1_12[175], stage1_12[176], stage1_12[177], stage1_12[178], stage1_12[179]},
      {stage1_13[58]},
      {stage1_14[174], stage1_14[175], stage1_14[176], stage1_14[177], stage1_14[178], stage1_14[179]},
      {stage2_16[29],stage2_15[34],stage2_14[38],stage2_13[60],stage2_12[87]}
   );
   gpc615_5 gpc2483 (
      {stage1_12[180], stage1_12[181], stage1_12[182], stage1_12[183], stage1_12[184]},
      {stage1_13[59]},
      {stage1_14[180], stage1_14[181], stage1_14[182], stage1_14[183], stage1_14[184], stage1_14[185]},
      {stage2_16[30],stage2_15[35],stage2_14[39],stage2_13[61],stage2_12[88]}
   );
   gpc615_5 gpc2484 (
      {stage1_12[185], stage1_12[186], stage1_12[187], stage1_12[188], stage1_12[189]},
      {stage1_13[60]},
      {stage1_14[186], stage1_14[187], stage1_14[188], stage1_14[189], stage1_14[190], stage1_14[191]},
      {stage2_16[31],stage2_15[36],stage2_14[40],stage2_13[62],stage2_12[89]}
   );
   gpc615_5 gpc2485 (
      {stage1_12[190], stage1_12[191], stage1_12[192], stage1_12[193], stage1_12[194]},
      {stage1_13[61]},
      {stage1_14[192], stage1_14[193], stage1_14[194], stage1_14[195], stage1_14[196], stage1_14[197]},
      {stage2_16[32],stage2_15[37],stage2_14[41],stage2_13[63],stage2_12[90]}
   );
   gpc615_5 gpc2486 (
      {stage1_12[195], stage1_12[196], stage1_12[197], stage1_12[198], stage1_12[199]},
      {stage1_13[62]},
      {stage1_14[198], stage1_14[199], stage1_14[200], stage1_14[201], stage1_14[202], stage1_14[203]},
      {stage2_16[33],stage2_15[38],stage2_14[42],stage2_13[64],stage2_12[91]}
   );
   gpc615_5 gpc2487 (
      {stage1_12[200], stage1_12[201], stage1_12[202], stage1_12[203], stage1_12[204]},
      {stage1_13[63]},
      {stage1_14[204], stage1_14[205], stage1_14[206], stage1_14[207], stage1_14[208], stage1_14[209]},
      {stage2_16[34],stage2_15[39],stage2_14[43],stage2_13[65],stage2_12[92]}
   );
   gpc615_5 gpc2488 (
      {stage1_12[205], stage1_12[206], stage1_12[207], stage1_12[208], stage1_12[209]},
      {stage1_13[64]},
      {stage1_14[210], stage1_14[211], stage1_14[212], stage1_14[213], stage1_14[214], stage1_14[215]},
      {stage2_16[35],stage2_15[40],stage2_14[44],stage2_13[66],stage2_12[93]}
   );
   gpc615_5 gpc2489 (
      {stage1_12[210], stage1_12[211], stage1_12[212], stage1_12[213], stage1_12[214]},
      {stage1_13[65]},
      {stage1_14[216], stage1_14[217], stage1_14[218], stage1_14[219], stage1_14[220], stage1_14[221]},
      {stage2_16[36],stage2_15[41],stage2_14[45],stage2_13[67],stage2_12[94]}
   );
   gpc606_5 gpc2490 (
      {stage1_13[66], stage1_13[67], stage1_13[68], stage1_13[69], stage1_13[70], stage1_13[71]},
      {stage1_15[0], stage1_15[1], stage1_15[2], stage1_15[3], stage1_15[4], stage1_15[5]},
      {stage2_17[0],stage2_16[37],stage2_15[42],stage2_14[46],stage2_13[68]}
   );
   gpc606_5 gpc2491 (
      {stage1_13[72], stage1_13[73], stage1_13[74], stage1_13[75], stage1_13[76], stage1_13[77]},
      {stage1_15[6], stage1_15[7], stage1_15[8], stage1_15[9], stage1_15[10], stage1_15[11]},
      {stage2_17[1],stage2_16[38],stage2_15[43],stage2_14[47],stage2_13[69]}
   );
   gpc606_5 gpc2492 (
      {stage1_13[78], stage1_13[79], stage1_13[80], stage1_13[81], stage1_13[82], stage1_13[83]},
      {stage1_15[12], stage1_15[13], stage1_15[14], stage1_15[15], stage1_15[16], stage1_15[17]},
      {stage2_17[2],stage2_16[39],stage2_15[44],stage2_14[48],stage2_13[70]}
   );
   gpc606_5 gpc2493 (
      {stage1_13[84], stage1_13[85], stage1_13[86], stage1_13[87], stage1_13[88], stage1_13[89]},
      {stage1_15[18], stage1_15[19], stage1_15[20], stage1_15[21], stage1_15[22], stage1_15[23]},
      {stage2_17[3],stage2_16[40],stage2_15[45],stage2_14[49],stage2_13[71]}
   );
   gpc606_5 gpc2494 (
      {stage1_13[90], stage1_13[91], stage1_13[92], stage1_13[93], stage1_13[94], stage1_13[95]},
      {stage1_15[24], stage1_15[25], stage1_15[26], stage1_15[27], stage1_15[28], stage1_15[29]},
      {stage2_17[4],stage2_16[41],stage2_15[46],stage2_14[50],stage2_13[72]}
   );
   gpc606_5 gpc2495 (
      {stage1_13[96], stage1_13[97], stage1_13[98], stage1_13[99], stage1_13[100], stage1_13[101]},
      {stage1_15[30], stage1_15[31], stage1_15[32], stage1_15[33], stage1_15[34], stage1_15[35]},
      {stage2_17[5],stage2_16[42],stage2_15[47],stage2_14[51],stage2_13[73]}
   );
   gpc606_5 gpc2496 (
      {stage1_13[102], stage1_13[103], stage1_13[104], stage1_13[105], stage1_13[106], stage1_13[107]},
      {stage1_15[36], stage1_15[37], stage1_15[38], stage1_15[39], stage1_15[40], stage1_15[41]},
      {stage2_17[6],stage2_16[43],stage2_15[48],stage2_14[52],stage2_13[74]}
   );
   gpc606_5 gpc2497 (
      {stage1_13[108], stage1_13[109], stage1_13[110], stage1_13[111], stage1_13[112], stage1_13[113]},
      {stage1_15[42], stage1_15[43], stage1_15[44], stage1_15[45], stage1_15[46], stage1_15[47]},
      {stage2_17[7],stage2_16[44],stage2_15[49],stage2_14[53],stage2_13[75]}
   );
   gpc606_5 gpc2498 (
      {stage1_13[114], stage1_13[115], stage1_13[116], stage1_13[117], stage1_13[118], stage1_13[119]},
      {stage1_15[48], stage1_15[49], stage1_15[50], stage1_15[51], stage1_15[52], stage1_15[53]},
      {stage2_17[8],stage2_16[45],stage2_15[50],stage2_14[54],stage2_13[76]}
   );
   gpc606_5 gpc2499 (
      {stage1_13[120], stage1_13[121], stage1_13[122], stage1_13[123], stage1_13[124], stage1_13[125]},
      {stage1_15[54], stage1_15[55], stage1_15[56], stage1_15[57], stage1_15[58], stage1_15[59]},
      {stage2_17[9],stage2_16[46],stage2_15[51],stage2_14[55],stage2_13[77]}
   );
   gpc606_5 gpc2500 (
      {stage1_13[126], stage1_13[127], stage1_13[128], stage1_13[129], stage1_13[130], stage1_13[131]},
      {stage1_15[60], stage1_15[61], stage1_15[62], stage1_15[63], stage1_15[64], stage1_15[65]},
      {stage2_17[10],stage2_16[47],stage2_15[52],stage2_14[56],stage2_13[78]}
   );
   gpc606_5 gpc2501 (
      {stage1_13[132], stage1_13[133], stage1_13[134], stage1_13[135], stage1_13[136], stage1_13[137]},
      {stage1_15[66], stage1_15[67], stage1_15[68], stage1_15[69], stage1_15[70], stage1_15[71]},
      {stage2_17[11],stage2_16[48],stage2_15[53],stage2_14[57],stage2_13[79]}
   );
   gpc606_5 gpc2502 (
      {stage1_13[138], stage1_13[139], stage1_13[140], stage1_13[141], stage1_13[142], stage1_13[143]},
      {stage1_15[72], stage1_15[73], stage1_15[74], stage1_15[75], stage1_15[76], stage1_15[77]},
      {stage2_17[12],stage2_16[49],stage2_15[54],stage2_14[58],stage2_13[80]}
   );
   gpc606_5 gpc2503 (
      {stage1_13[144], stage1_13[145], stage1_13[146], stage1_13[147], stage1_13[148], stage1_13[149]},
      {stage1_15[78], stage1_15[79], stage1_15[80], stage1_15[81], stage1_15[82], stage1_15[83]},
      {stage2_17[13],stage2_16[50],stage2_15[55],stage2_14[59],stage2_13[81]}
   );
   gpc606_5 gpc2504 (
      {stage1_13[150], stage1_13[151], stage1_13[152], stage1_13[153], stage1_13[154], stage1_13[155]},
      {stage1_15[84], stage1_15[85], stage1_15[86], stage1_15[87], stage1_15[88], stage1_15[89]},
      {stage2_17[14],stage2_16[51],stage2_15[56],stage2_14[60],stage2_13[82]}
   );
   gpc606_5 gpc2505 (
      {stage1_13[156], stage1_13[157], stage1_13[158], stage1_13[159], stage1_13[160], stage1_13[161]},
      {stage1_15[90], stage1_15[91], stage1_15[92], stage1_15[93], stage1_15[94], stage1_15[95]},
      {stage2_17[15],stage2_16[52],stage2_15[57],stage2_14[61],stage2_13[83]}
   );
   gpc606_5 gpc2506 (
      {stage1_13[162], stage1_13[163], stage1_13[164], stage1_13[165], stage1_13[166], stage1_13[167]},
      {stage1_15[96], stage1_15[97], stage1_15[98], stage1_15[99], stage1_15[100], stage1_15[101]},
      {stage2_17[16],stage2_16[53],stage2_15[58],stage2_14[62],stage2_13[84]}
   );
   gpc606_5 gpc2507 (
      {stage1_13[168], stage1_13[169], stage1_13[170], stage1_13[171], stage1_13[172], stage1_13[173]},
      {stage1_15[102], stage1_15[103], stage1_15[104], stage1_15[105], stage1_15[106], stage1_15[107]},
      {stage2_17[17],stage2_16[54],stage2_15[59],stage2_14[63],stage2_13[85]}
   );
   gpc606_5 gpc2508 (
      {stage1_13[174], stage1_13[175], stage1_13[176], stage1_13[177], stage1_13[178], stage1_13[179]},
      {stage1_15[108], stage1_15[109], stage1_15[110], stage1_15[111], stage1_15[112], stage1_15[113]},
      {stage2_17[18],stage2_16[55],stage2_15[60],stage2_14[64],stage2_13[86]}
   );
   gpc606_5 gpc2509 (
      {stage1_13[180], stage1_13[181], stage1_13[182], stage1_13[183], stage1_13[184], stage1_13[185]},
      {stage1_15[114], stage1_15[115], stage1_15[116], stage1_15[117], stage1_15[118], stage1_15[119]},
      {stage2_17[19],stage2_16[56],stage2_15[61],stage2_14[65],stage2_13[87]}
   );
   gpc606_5 gpc2510 (
      {stage1_13[186], stage1_13[187], stage1_13[188], stage1_13[189], stage1_13[190], stage1_13[191]},
      {stage1_15[120], stage1_15[121], stage1_15[122], stage1_15[123], stage1_15[124], stage1_15[125]},
      {stage2_17[20],stage2_16[57],stage2_15[62],stage2_14[66],stage2_13[88]}
   );
   gpc606_5 gpc2511 (
      {stage1_13[192], stage1_13[193], stage1_13[194], stage1_13[195], stage1_13[196], stage1_13[197]},
      {stage1_15[126], stage1_15[127], stage1_15[128], stage1_15[129], stage1_15[130], stage1_15[131]},
      {stage2_17[21],stage2_16[58],stage2_15[63],stage2_14[67],stage2_13[89]}
   );
   gpc615_5 gpc2512 (
      {stage1_14[222], stage1_14[223], stage1_14[224], stage1_14[225], stage1_14[226]},
      {stage1_15[132]},
      {stage1_16[0], stage1_16[1], stage1_16[2], stage1_16[3], stage1_16[4], stage1_16[5]},
      {stage2_18[0],stage2_17[22],stage2_16[59],stage2_15[64],stage2_14[68]}
   );
   gpc615_5 gpc2513 (
      {stage1_14[227], stage1_14[228], stage1_14[229], stage1_14[230], stage1_14[231]},
      {stage1_15[133]},
      {stage1_16[6], stage1_16[7], stage1_16[8], stage1_16[9], stage1_16[10], stage1_16[11]},
      {stage2_18[1],stage2_17[23],stage2_16[60],stage2_15[65],stage2_14[69]}
   );
   gpc606_5 gpc2514 (
      {stage1_15[134], stage1_15[135], stage1_15[136], stage1_15[137], stage1_15[138], stage1_15[139]},
      {stage1_17[0], stage1_17[1], stage1_17[2], stage1_17[3], stage1_17[4], stage1_17[5]},
      {stage2_19[0],stage2_18[2],stage2_17[24],stage2_16[61],stage2_15[66]}
   );
   gpc606_5 gpc2515 (
      {stage1_15[140], stage1_15[141], stage1_15[142], stage1_15[143], stage1_15[144], stage1_15[145]},
      {stage1_17[6], stage1_17[7], stage1_17[8], stage1_17[9], stage1_17[10], stage1_17[11]},
      {stage2_19[1],stage2_18[3],stage2_17[25],stage2_16[62],stage2_15[67]}
   );
   gpc606_5 gpc2516 (
      {stage1_15[146], stage1_15[147], stage1_15[148], stage1_15[149], stage1_15[150], stage1_15[151]},
      {stage1_17[12], stage1_17[13], stage1_17[14], stage1_17[15], stage1_17[16], stage1_17[17]},
      {stage2_19[2],stage2_18[4],stage2_17[26],stage2_16[63],stage2_15[68]}
   );
   gpc615_5 gpc2517 (
      {stage1_15[152], stage1_15[153], stage1_15[154], stage1_15[155], stage1_15[156]},
      {stage1_16[12]},
      {stage1_17[18], stage1_17[19], stage1_17[20], stage1_17[21], stage1_17[22], stage1_17[23]},
      {stage2_19[3],stage2_18[5],stage2_17[27],stage2_16[64],stage2_15[69]}
   );
   gpc615_5 gpc2518 (
      {stage1_15[157], stage1_15[158], stage1_15[159], stage1_15[160], stage1_15[161]},
      {stage1_16[13]},
      {stage1_17[24], stage1_17[25], stage1_17[26], stage1_17[27], stage1_17[28], stage1_17[29]},
      {stage2_19[4],stage2_18[6],stage2_17[28],stage2_16[65],stage2_15[70]}
   );
   gpc615_5 gpc2519 (
      {stage1_15[162], stage1_15[163], stage1_15[164], stage1_15[165], stage1_15[166]},
      {stage1_16[14]},
      {stage1_17[30], stage1_17[31], stage1_17[32], stage1_17[33], stage1_17[34], stage1_17[35]},
      {stage2_19[5],stage2_18[7],stage2_17[29],stage2_16[66],stage2_15[71]}
   );
   gpc615_5 gpc2520 (
      {stage1_15[167], stage1_15[168], stage1_15[169], stage1_15[170], stage1_15[171]},
      {stage1_16[15]},
      {stage1_17[36], stage1_17[37], stage1_17[38], stage1_17[39], stage1_17[40], stage1_17[41]},
      {stage2_19[6],stage2_18[8],stage2_17[30],stage2_16[67],stage2_15[72]}
   );
   gpc615_5 gpc2521 (
      {stage1_15[172], stage1_15[173], stage1_15[174], stage1_15[175], stage1_15[176]},
      {stage1_16[16]},
      {stage1_17[42], stage1_17[43], stage1_17[44], stage1_17[45], stage1_17[46], stage1_17[47]},
      {stage2_19[7],stage2_18[9],stage2_17[31],stage2_16[68],stage2_15[73]}
   );
   gpc615_5 gpc2522 (
      {stage1_15[177], stage1_15[178], stage1_15[179], stage1_15[180], stage1_15[181]},
      {stage1_16[17]},
      {stage1_17[48], stage1_17[49], stage1_17[50], stage1_17[51], stage1_17[52], stage1_17[53]},
      {stage2_19[8],stage2_18[10],stage2_17[32],stage2_16[69],stage2_15[74]}
   );
   gpc615_5 gpc2523 (
      {stage1_15[182], stage1_15[183], stage1_15[184], stage1_15[185], stage1_15[186]},
      {stage1_16[18]},
      {stage1_17[54], stage1_17[55], stage1_17[56], stage1_17[57], stage1_17[58], stage1_17[59]},
      {stage2_19[9],stage2_18[11],stage2_17[33],stage2_16[70],stage2_15[75]}
   );
   gpc615_5 gpc2524 (
      {stage1_15[187], stage1_15[188], stage1_15[189], stage1_15[190], stage1_15[191]},
      {stage1_16[19]},
      {stage1_17[60], stage1_17[61], stage1_17[62], stage1_17[63], stage1_17[64], stage1_17[65]},
      {stage2_19[10],stage2_18[12],stage2_17[34],stage2_16[71],stage2_15[76]}
   );
   gpc615_5 gpc2525 (
      {stage1_15[192], stage1_15[193], stage1_15[194], stage1_15[195], stage1_15[196]},
      {stage1_16[20]},
      {stage1_17[66], stage1_17[67], stage1_17[68], stage1_17[69], stage1_17[70], stage1_17[71]},
      {stage2_19[11],stage2_18[13],stage2_17[35],stage2_16[72],stage2_15[77]}
   );
   gpc615_5 gpc2526 (
      {stage1_15[197], stage1_15[198], stage1_15[199], stage1_15[200], stage1_15[201]},
      {stage1_16[21]},
      {stage1_17[72], stage1_17[73], stage1_17[74], stage1_17[75], stage1_17[76], stage1_17[77]},
      {stage2_19[12],stage2_18[14],stage2_17[36],stage2_16[73],stage2_15[78]}
   );
   gpc615_5 gpc2527 (
      {stage1_15[202], stage1_15[203], stage1_15[204], stage1_15[205], stage1_15[206]},
      {stage1_16[22]},
      {stage1_17[78], stage1_17[79], stage1_17[80], stage1_17[81], stage1_17[82], stage1_17[83]},
      {stage2_19[13],stage2_18[15],stage2_17[37],stage2_16[74],stage2_15[79]}
   );
   gpc615_5 gpc2528 (
      {stage1_15[207], stage1_15[208], stage1_15[209], stage1_15[210], stage1_15[211]},
      {stage1_16[23]},
      {stage1_17[84], stage1_17[85], stage1_17[86], stage1_17[87], stage1_17[88], stage1_17[89]},
      {stage2_19[14],stage2_18[16],stage2_17[38],stage2_16[75],stage2_15[80]}
   );
   gpc615_5 gpc2529 (
      {stage1_15[212], stage1_15[213], stage1_15[214], stage1_15[215], stage1_15[216]},
      {stage1_16[24]},
      {stage1_17[90], stage1_17[91], stage1_17[92], stage1_17[93], stage1_17[94], stage1_17[95]},
      {stage2_19[15],stage2_18[17],stage2_17[39],stage2_16[76],stage2_15[81]}
   );
   gpc615_5 gpc2530 (
      {stage1_15[217], stage1_15[218], stage1_15[219], stage1_15[220], stage1_15[221]},
      {stage1_16[25]},
      {stage1_17[96], stage1_17[97], stage1_17[98], stage1_17[99], stage1_17[100], stage1_17[101]},
      {stage2_19[16],stage2_18[18],stage2_17[40],stage2_16[77],stage2_15[82]}
   );
   gpc606_5 gpc2531 (
      {stage1_16[26], stage1_16[27], stage1_16[28], stage1_16[29], stage1_16[30], stage1_16[31]},
      {stage1_18[0], stage1_18[1], stage1_18[2], stage1_18[3], stage1_18[4], stage1_18[5]},
      {stage2_20[0],stage2_19[17],stage2_18[19],stage2_17[41],stage2_16[78]}
   );
   gpc606_5 gpc2532 (
      {stage1_16[32], stage1_16[33], stage1_16[34], stage1_16[35], stage1_16[36], stage1_16[37]},
      {stage1_18[6], stage1_18[7], stage1_18[8], stage1_18[9], stage1_18[10], stage1_18[11]},
      {stage2_20[1],stage2_19[18],stage2_18[20],stage2_17[42],stage2_16[79]}
   );
   gpc606_5 gpc2533 (
      {stage1_16[38], stage1_16[39], stage1_16[40], stage1_16[41], stage1_16[42], stage1_16[43]},
      {stage1_18[12], stage1_18[13], stage1_18[14], stage1_18[15], stage1_18[16], stage1_18[17]},
      {stage2_20[2],stage2_19[19],stage2_18[21],stage2_17[43],stage2_16[80]}
   );
   gpc606_5 gpc2534 (
      {stage1_16[44], stage1_16[45], stage1_16[46], stage1_16[47], stage1_16[48], stage1_16[49]},
      {stage1_18[18], stage1_18[19], stage1_18[20], stage1_18[21], stage1_18[22], stage1_18[23]},
      {stage2_20[3],stage2_19[20],stage2_18[22],stage2_17[44],stage2_16[81]}
   );
   gpc606_5 gpc2535 (
      {stage1_16[50], stage1_16[51], stage1_16[52], stage1_16[53], stage1_16[54], stage1_16[55]},
      {stage1_18[24], stage1_18[25], stage1_18[26], stage1_18[27], stage1_18[28], stage1_18[29]},
      {stage2_20[4],stage2_19[21],stage2_18[23],stage2_17[45],stage2_16[82]}
   );
   gpc606_5 gpc2536 (
      {stage1_16[56], stage1_16[57], stage1_16[58], stage1_16[59], stage1_16[60], stage1_16[61]},
      {stage1_18[30], stage1_18[31], stage1_18[32], stage1_18[33], stage1_18[34], stage1_18[35]},
      {stage2_20[5],stage2_19[22],stage2_18[24],stage2_17[46],stage2_16[83]}
   );
   gpc606_5 gpc2537 (
      {stage1_16[62], stage1_16[63], stage1_16[64], stage1_16[65], stage1_16[66], stage1_16[67]},
      {stage1_18[36], stage1_18[37], stage1_18[38], stage1_18[39], stage1_18[40], stage1_18[41]},
      {stage2_20[6],stage2_19[23],stage2_18[25],stage2_17[47],stage2_16[84]}
   );
   gpc606_5 gpc2538 (
      {stage1_16[68], stage1_16[69], stage1_16[70], stage1_16[71], stage1_16[72], stage1_16[73]},
      {stage1_18[42], stage1_18[43], stage1_18[44], stage1_18[45], stage1_18[46], stage1_18[47]},
      {stage2_20[7],stage2_19[24],stage2_18[26],stage2_17[48],stage2_16[85]}
   );
   gpc606_5 gpc2539 (
      {stage1_16[74], stage1_16[75], stage1_16[76], stage1_16[77], stage1_16[78], stage1_16[79]},
      {stage1_18[48], stage1_18[49], stage1_18[50], stage1_18[51], stage1_18[52], stage1_18[53]},
      {stage2_20[8],stage2_19[25],stage2_18[27],stage2_17[49],stage2_16[86]}
   );
   gpc606_5 gpc2540 (
      {stage1_16[80], stage1_16[81], stage1_16[82], stage1_16[83], stage1_16[84], stage1_16[85]},
      {stage1_18[54], stage1_18[55], stage1_18[56], stage1_18[57], stage1_18[58], stage1_18[59]},
      {stage2_20[9],stage2_19[26],stage2_18[28],stage2_17[50],stage2_16[87]}
   );
   gpc606_5 gpc2541 (
      {stage1_16[86], stage1_16[87], stage1_16[88], stage1_16[89], stage1_16[90], stage1_16[91]},
      {stage1_18[60], stage1_18[61], stage1_18[62], stage1_18[63], stage1_18[64], stage1_18[65]},
      {stage2_20[10],stage2_19[27],stage2_18[29],stage2_17[51],stage2_16[88]}
   );
   gpc606_5 gpc2542 (
      {stage1_16[92], stage1_16[93], stage1_16[94], stage1_16[95], stage1_16[96], stage1_16[97]},
      {stage1_18[66], stage1_18[67], stage1_18[68], stage1_18[69], stage1_18[70], stage1_18[71]},
      {stage2_20[11],stage2_19[28],stage2_18[30],stage2_17[52],stage2_16[89]}
   );
   gpc606_5 gpc2543 (
      {stage1_16[98], stage1_16[99], stage1_16[100], stage1_16[101], stage1_16[102], stage1_16[103]},
      {stage1_18[72], stage1_18[73], stage1_18[74], stage1_18[75], stage1_18[76], stage1_18[77]},
      {stage2_20[12],stage2_19[29],stage2_18[31],stage2_17[53],stage2_16[90]}
   );
   gpc606_5 gpc2544 (
      {stage1_16[104], stage1_16[105], stage1_16[106], stage1_16[107], stage1_16[108], stage1_16[109]},
      {stage1_18[78], stage1_18[79], stage1_18[80], stage1_18[81], stage1_18[82], stage1_18[83]},
      {stage2_20[13],stage2_19[30],stage2_18[32],stage2_17[54],stage2_16[91]}
   );
   gpc606_5 gpc2545 (
      {stage1_16[110], stage1_16[111], stage1_16[112], stage1_16[113], stage1_16[114], stage1_16[115]},
      {stage1_18[84], stage1_18[85], stage1_18[86], stage1_18[87], stage1_18[88], stage1_18[89]},
      {stage2_20[14],stage2_19[31],stage2_18[33],stage2_17[55],stage2_16[92]}
   );
   gpc606_5 gpc2546 (
      {stage1_16[116], stage1_16[117], stage1_16[118], stage1_16[119], stage1_16[120], stage1_16[121]},
      {stage1_18[90], stage1_18[91], stage1_18[92], stage1_18[93], stage1_18[94], stage1_18[95]},
      {stage2_20[15],stage2_19[32],stage2_18[34],stage2_17[56],stage2_16[93]}
   );
   gpc606_5 gpc2547 (
      {stage1_16[122], stage1_16[123], stage1_16[124], stage1_16[125], stage1_16[126], stage1_16[127]},
      {stage1_18[96], stage1_18[97], stage1_18[98], stage1_18[99], stage1_18[100], stage1_18[101]},
      {stage2_20[16],stage2_19[33],stage2_18[35],stage2_17[57],stage2_16[94]}
   );
   gpc606_5 gpc2548 (
      {stage1_16[128], stage1_16[129], stage1_16[130], stage1_16[131], stage1_16[132], stage1_16[133]},
      {stage1_18[102], stage1_18[103], stage1_18[104], stage1_18[105], stage1_18[106], stage1_18[107]},
      {stage2_20[17],stage2_19[34],stage2_18[36],stage2_17[58],stage2_16[95]}
   );
   gpc606_5 gpc2549 (
      {stage1_16[134], stage1_16[135], stage1_16[136], stage1_16[137], stage1_16[138], stage1_16[139]},
      {stage1_18[108], stage1_18[109], stage1_18[110], stage1_18[111], stage1_18[112], stage1_18[113]},
      {stage2_20[18],stage2_19[35],stage2_18[37],stage2_17[59],stage2_16[96]}
   );
   gpc606_5 gpc2550 (
      {stage1_16[140], stage1_16[141], stage1_16[142], stage1_16[143], stage1_16[144], stage1_16[145]},
      {stage1_18[114], stage1_18[115], stage1_18[116], stage1_18[117], stage1_18[118], stage1_18[119]},
      {stage2_20[19],stage2_19[36],stage2_18[38],stage2_17[60],stage2_16[97]}
   );
   gpc606_5 gpc2551 (
      {stage1_16[146], stage1_16[147], stage1_16[148], stage1_16[149], stage1_16[150], stage1_16[151]},
      {stage1_18[120], stage1_18[121], stage1_18[122], stage1_18[123], stage1_18[124], stage1_18[125]},
      {stage2_20[20],stage2_19[37],stage2_18[39],stage2_17[61],stage2_16[98]}
   );
   gpc606_5 gpc2552 (
      {stage1_16[152], stage1_16[153], stage1_16[154], stage1_16[155], stage1_16[156], stage1_16[157]},
      {stage1_18[126], stage1_18[127], stage1_18[128], stage1_18[129], stage1_18[130], stage1_18[131]},
      {stage2_20[21],stage2_19[38],stage2_18[40],stage2_17[62],stage2_16[99]}
   );
   gpc606_5 gpc2553 (
      {stage1_16[158], stage1_16[159], stage1_16[160], stage1_16[161], stage1_16[162], stage1_16[163]},
      {stage1_18[132], stage1_18[133], stage1_18[134], stage1_18[135], stage1_18[136], stage1_18[137]},
      {stage2_20[22],stage2_19[39],stage2_18[41],stage2_17[63],stage2_16[100]}
   );
   gpc606_5 gpc2554 (
      {stage1_16[164], stage1_16[165], stage1_16[166], stage1_16[167], stage1_16[168], stage1_16[169]},
      {stage1_18[138], stage1_18[139], stage1_18[140], stage1_18[141], stage1_18[142], stage1_18[143]},
      {stage2_20[23],stage2_19[40],stage2_18[42],stage2_17[64],stage2_16[101]}
   );
   gpc606_5 gpc2555 (
      {stage1_16[170], stage1_16[171], stage1_16[172], stage1_16[173], stage1_16[174], stage1_16[175]},
      {stage1_18[144], stage1_18[145], stage1_18[146], stage1_18[147], stage1_18[148], stage1_18[149]},
      {stage2_20[24],stage2_19[41],stage2_18[43],stage2_17[65],stage2_16[102]}
   );
   gpc615_5 gpc2556 (
      {stage1_16[176], stage1_16[177], stage1_16[178], stage1_16[179], stage1_16[180]},
      {stage1_17[102]},
      {stage1_18[150], stage1_18[151], stage1_18[152], stage1_18[153], stage1_18[154], stage1_18[155]},
      {stage2_20[25],stage2_19[42],stage2_18[44],stage2_17[66],stage2_16[103]}
   );
   gpc615_5 gpc2557 (
      {stage1_16[181], stage1_16[182], stage1_16[183], stage1_16[184], stage1_16[185]},
      {stage1_17[103]},
      {stage1_18[156], stage1_18[157], stage1_18[158], stage1_18[159], stage1_18[160], stage1_18[161]},
      {stage2_20[26],stage2_19[43],stage2_18[45],stage2_17[67],stage2_16[104]}
   );
   gpc615_5 gpc2558 (
      {stage1_16[186], stage1_16[187], stage1_16[188], stage1_16[189], stage1_16[190]},
      {stage1_17[104]},
      {stage1_18[162], stage1_18[163], stage1_18[164], stage1_18[165], stage1_18[166], stage1_18[167]},
      {stage2_20[27],stage2_19[44],stage2_18[46],stage2_17[68],stage2_16[105]}
   );
   gpc615_5 gpc2559 (
      {stage1_16[191], stage1_16[192], stage1_16[193], stage1_16[194], stage1_16[195]},
      {stage1_17[105]},
      {stage1_18[168], stage1_18[169], stage1_18[170], stage1_18[171], stage1_18[172], stage1_18[173]},
      {stage2_20[28],stage2_19[45],stage2_18[47],stage2_17[69],stage2_16[106]}
   );
   gpc606_5 gpc2560 (
      {stage1_17[106], stage1_17[107], stage1_17[108], stage1_17[109], stage1_17[110], stage1_17[111]},
      {stage1_19[0], stage1_19[1], stage1_19[2], stage1_19[3], stage1_19[4], stage1_19[5]},
      {stage2_21[0],stage2_20[29],stage2_19[46],stage2_18[48],stage2_17[70]}
   );
   gpc606_5 gpc2561 (
      {stage1_17[112], stage1_17[113], stage1_17[114], stage1_17[115], stage1_17[116], stage1_17[117]},
      {stage1_19[6], stage1_19[7], stage1_19[8], stage1_19[9], stage1_19[10], stage1_19[11]},
      {stage2_21[1],stage2_20[30],stage2_19[47],stage2_18[49],stage2_17[71]}
   );
   gpc606_5 gpc2562 (
      {stage1_17[118], stage1_17[119], stage1_17[120], stage1_17[121], stage1_17[122], stage1_17[123]},
      {stage1_19[12], stage1_19[13], stage1_19[14], stage1_19[15], stage1_19[16], stage1_19[17]},
      {stage2_21[2],stage2_20[31],stage2_19[48],stage2_18[50],stage2_17[72]}
   );
   gpc606_5 gpc2563 (
      {stage1_17[124], stage1_17[125], stage1_17[126], stage1_17[127], stage1_17[128], stage1_17[129]},
      {stage1_19[18], stage1_19[19], stage1_19[20], stage1_19[21], stage1_19[22], stage1_19[23]},
      {stage2_21[3],stage2_20[32],stage2_19[49],stage2_18[51],stage2_17[73]}
   );
   gpc606_5 gpc2564 (
      {stage1_17[130], stage1_17[131], stage1_17[132], stage1_17[133], stage1_17[134], stage1_17[135]},
      {stage1_19[24], stage1_19[25], stage1_19[26], stage1_19[27], stage1_19[28], stage1_19[29]},
      {stage2_21[4],stage2_20[33],stage2_19[50],stage2_18[52],stage2_17[74]}
   );
   gpc606_5 gpc2565 (
      {stage1_17[136], stage1_17[137], stage1_17[138], stage1_17[139], stage1_17[140], stage1_17[141]},
      {stage1_19[30], stage1_19[31], stage1_19[32], stage1_19[33], stage1_19[34], stage1_19[35]},
      {stage2_21[5],stage2_20[34],stage2_19[51],stage2_18[53],stage2_17[75]}
   );
   gpc606_5 gpc2566 (
      {stage1_17[142], stage1_17[143], stage1_17[144], stage1_17[145], stage1_17[146], stage1_17[147]},
      {stage1_19[36], stage1_19[37], stage1_19[38], stage1_19[39], stage1_19[40], stage1_19[41]},
      {stage2_21[6],stage2_20[35],stage2_19[52],stage2_18[54],stage2_17[76]}
   );
   gpc606_5 gpc2567 (
      {stage1_17[148], stage1_17[149], stage1_17[150], stage1_17[151], stage1_17[152], stage1_17[153]},
      {stage1_19[42], stage1_19[43], stage1_19[44], stage1_19[45], stage1_19[46], stage1_19[47]},
      {stage2_21[7],stage2_20[36],stage2_19[53],stage2_18[55],stage2_17[77]}
   );
   gpc606_5 gpc2568 (
      {stage1_17[154], stage1_17[155], stage1_17[156], stage1_17[157], stage1_17[158], stage1_17[159]},
      {stage1_19[48], stage1_19[49], stage1_19[50], stage1_19[51], stage1_19[52], stage1_19[53]},
      {stage2_21[8],stage2_20[37],stage2_19[54],stage2_18[56],stage2_17[78]}
   );
   gpc606_5 gpc2569 (
      {stage1_17[160], stage1_17[161], stage1_17[162], stage1_17[163], stage1_17[164], stage1_17[165]},
      {stage1_19[54], stage1_19[55], stage1_19[56], stage1_19[57], stage1_19[58], stage1_19[59]},
      {stage2_21[9],stage2_20[38],stage2_19[55],stage2_18[57],stage2_17[79]}
   );
   gpc606_5 gpc2570 (
      {stage1_17[166], stage1_17[167], stage1_17[168], stage1_17[169], stage1_17[170], stage1_17[171]},
      {stage1_19[60], stage1_19[61], stage1_19[62], stage1_19[63], stage1_19[64], stage1_19[65]},
      {stage2_21[10],stage2_20[39],stage2_19[56],stage2_18[58],stage2_17[80]}
   );
   gpc606_5 gpc2571 (
      {stage1_17[172], stage1_17[173], stage1_17[174], stage1_17[175], stage1_17[176], stage1_17[177]},
      {stage1_19[66], stage1_19[67], stage1_19[68], stage1_19[69], stage1_19[70], stage1_19[71]},
      {stage2_21[11],stage2_20[40],stage2_19[57],stage2_18[59],stage2_17[81]}
   );
   gpc615_5 gpc2572 (
      {stage1_18[174], stage1_18[175], stage1_18[176], stage1_18[177], stage1_18[178]},
      {stage1_19[72]},
      {stage1_20[0], stage1_20[1], stage1_20[2], stage1_20[3], stage1_20[4], stage1_20[5]},
      {stage2_22[0],stage2_21[12],stage2_20[41],stage2_19[58],stage2_18[60]}
   );
   gpc615_5 gpc2573 (
      {stage1_18[179], stage1_18[180], stage1_18[181], stage1_18[182], stage1_18[183]},
      {stage1_19[73]},
      {stage1_20[6], stage1_20[7], stage1_20[8], stage1_20[9], stage1_20[10], stage1_20[11]},
      {stage2_22[1],stage2_21[13],stage2_20[42],stage2_19[59],stage2_18[61]}
   );
   gpc615_5 gpc2574 (
      {stage1_18[184], stage1_18[185], stage1_18[186], stage1_18[187], stage1_18[188]},
      {stage1_19[74]},
      {stage1_20[12], stage1_20[13], stage1_20[14], stage1_20[15], stage1_20[16], stage1_20[17]},
      {stage2_22[2],stage2_21[14],stage2_20[43],stage2_19[60],stage2_18[62]}
   );
   gpc615_5 gpc2575 (
      {stage1_18[189], stage1_18[190], stage1_18[191], stage1_18[192], stage1_18[193]},
      {stage1_19[75]},
      {stage1_20[18], stage1_20[19], stage1_20[20], stage1_20[21], stage1_20[22], stage1_20[23]},
      {stage2_22[3],stage2_21[15],stage2_20[44],stage2_19[61],stage2_18[63]}
   );
   gpc606_5 gpc2576 (
      {stage1_19[76], stage1_19[77], stage1_19[78], stage1_19[79], stage1_19[80], stage1_19[81]},
      {stage1_21[0], stage1_21[1], stage1_21[2], stage1_21[3], stage1_21[4], stage1_21[5]},
      {stage2_23[0],stage2_22[4],stage2_21[16],stage2_20[45],stage2_19[62]}
   );
   gpc606_5 gpc2577 (
      {stage1_19[82], stage1_19[83], stage1_19[84], stage1_19[85], stage1_19[86], stage1_19[87]},
      {stage1_21[6], stage1_21[7], stage1_21[8], stage1_21[9], stage1_21[10], stage1_21[11]},
      {stage2_23[1],stage2_22[5],stage2_21[17],stage2_20[46],stage2_19[63]}
   );
   gpc606_5 gpc2578 (
      {stage1_19[88], stage1_19[89], stage1_19[90], stage1_19[91], stage1_19[92], stage1_19[93]},
      {stage1_21[12], stage1_21[13], stage1_21[14], stage1_21[15], stage1_21[16], stage1_21[17]},
      {stage2_23[2],stage2_22[6],stage2_21[18],stage2_20[47],stage2_19[64]}
   );
   gpc606_5 gpc2579 (
      {stage1_19[94], stage1_19[95], stage1_19[96], stage1_19[97], stage1_19[98], stage1_19[99]},
      {stage1_21[18], stage1_21[19], stage1_21[20], stage1_21[21], stage1_21[22], stage1_21[23]},
      {stage2_23[3],stage2_22[7],stage2_21[19],stage2_20[48],stage2_19[65]}
   );
   gpc606_5 gpc2580 (
      {stage1_19[100], stage1_19[101], stage1_19[102], stage1_19[103], stage1_19[104], stage1_19[105]},
      {stage1_21[24], stage1_21[25], stage1_21[26], stage1_21[27], stage1_21[28], stage1_21[29]},
      {stage2_23[4],stage2_22[8],stage2_21[20],stage2_20[49],stage2_19[66]}
   );
   gpc606_5 gpc2581 (
      {stage1_19[106], stage1_19[107], stage1_19[108], stage1_19[109], stage1_19[110], stage1_19[111]},
      {stage1_21[30], stage1_21[31], stage1_21[32], stage1_21[33], stage1_21[34], stage1_21[35]},
      {stage2_23[5],stage2_22[9],stage2_21[21],stage2_20[50],stage2_19[67]}
   );
   gpc606_5 gpc2582 (
      {stage1_19[112], stage1_19[113], stage1_19[114], stage1_19[115], stage1_19[116], stage1_19[117]},
      {stage1_21[36], stage1_21[37], stage1_21[38], stage1_21[39], stage1_21[40], stage1_21[41]},
      {stage2_23[6],stage2_22[10],stage2_21[22],stage2_20[51],stage2_19[68]}
   );
   gpc606_5 gpc2583 (
      {stage1_19[118], stage1_19[119], stage1_19[120], stage1_19[121], stage1_19[122], stage1_19[123]},
      {stage1_21[42], stage1_21[43], stage1_21[44], stage1_21[45], stage1_21[46], stage1_21[47]},
      {stage2_23[7],stage2_22[11],stage2_21[23],stage2_20[52],stage2_19[69]}
   );
   gpc606_5 gpc2584 (
      {stage1_19[124], stage1_19[125], stage1_19[126], stage1_19[127], stage1_19[128], stage1_19[129]},
      {stage1_21[48], stage1_21[49], stage1_21[50], stage1_21[51], stage1_21[52], stage1_21[53]},
      {stage2_23[8],stage2_22[12],stage2_21[24],stage2_20[53],stage2_19[70]}
   );
   gpc606_5 gpc2585 (
      {stage1_19[130], stage1_19[131], stage1_19[132], stage1_19[133], stage1_19[134], stage1_19[135]},
      {stage1_21[54], stage1_21[55], stage1_21[56], stage1_21[57], stage1_21[58], stage1_21[59]},
      {stage2_23[9],stage2_22[13],stage2_21[25],stage2_20[54],stage2_19[71]}
   );
   gpc606_5 gpc2586 (
      {stage1_19[136], stage1_19[137], stage1_19[138], stage1_19[139], stage1_19[140], stage1_19[141]},
      {stage1_21[60], stage1_21[61], stage1_21[62], stage1_21[63], stage1_21[64], stage1_21[65]},
      {stage2_23[10],stage2_22[14],stage2_21[26],stage2_20[55],stage2_19[72]}
   );
   gpc606_5 gpc2587 (
      {stage1_19[142], stage1_19[143], stage1_19[144], stage1_19[145], stage1_19[146], stage1_19[147]},
      {stage1_21[66], stage1_21[67], stage1_21[68], stage1_21[69], stage1_21[70], stage1_21[71]},
      {stage2_23[11],stage2_22[15],stage2_21[27],stage2_20[56],stage2_19[73]}
   );
   gpc606_5 gpc2588 (
      {stage1_19[148], stage1_19[149], stage1_19[150], stage1_19[151], stage1_19[152], stage1_19[153]},
      {stage1_21[72], stage1_21[73], stage1_21[74], stage1_21[75], stage1_21[76], stage1_21[77]},
      {stage2_23[12],stage2_22[16],stage2_21[28],stage2_20[57],stage2_19[74]}
   );
   gpc606_5 gpc2589 (
      {stage1_19[154], stage1_19[155], stage1_19[156], stage1_19[157], stage1_19[158], stage1_19[159]},
      {stage1_21[78], stage1_21[79], stage1_21[80], stage1_21[81], stage1_21[82], stage1_21[83]},
      {stage2_23[13],stage2_22[17],stage2_21[29],stage2_20[58],stage2_19[75]}
   );
   gpc606_5 gpc2590 (
      {stage1_19[160], stage1_19[161], stage1_19[162], stage1_19[163], stage1_19[164], stage1_19[165]},
      {stage1_21[84], stage1_21[85], stage1_21[86], stage1_21[87], stage1_21[88], stage1_21[89]},
      {stage2_23[14],stage2_22[18],stage2_21[30],stage2_20[59],stage2_19[76]}
   );
   gpc615_5 gpc2591 (
      {stage1_19[166], stage1_19[167], stage1_19[168], stage1_19[169], stage1_19[170]},
      {stage1_20[24]},
      {stage1_21[90], stage1_21[91], stage1_21[92], stage1_21[93], stage1_21[94], stage1_21[95]},
      {stage2_23[15],stage2_22[19],stage2_21[31],stage2_20[60],stage2_19[77]}
   );
   gpc615_5 gpc2592 (
      {stage1_19[171], stage1_19[172], stage1_19[173], stage1_19[174], stage1_19[175]},
      {stage1_20[25]},
      {stage1_21[96], stage1_21[97], stage1_21[98], stage1_21[99], stage1_21[100], stage1_21[101]},
      {stage2_23[16],stage2_22[20],stage2_21[32],stage2_20[61],stage2_19[78]}
   );
   gpc615_5 gpc2593 (
      {stage1_19[176], stage1_19[177], stage1_19[178], stage1_19[179], stage1_19[180]},
      {stage1_20[26]},
      {stage1_21[102], stage1_21[103], stage1_21[104], stage1_21[105], stage1_21[106], stage1_21[107]},
      {stage2_23[17],stage2_22[21],stage2_21[33],stage2_20[62],stage2_19[79]}
   );
   gpc615_5 gpc2594 (
      {stage1_19[181], stage1_19[182], stage1_19[183], stage1_19[184], stage1_19[185]},
      {stage1_20[27]},
      {stage1_21[108], stage1_21[109], stage1_21[110], stage1_21[111], stage1_21[112], stage1_21[113]},
      {stage2_23[18],stage2_22[22],stage2_21[34],stage2_20[63],stage2_19[80]}
   );
   gpc615_5 gpc2595 (
      {stage1_19[186], stage1_19[187], stage1_19[188], stage1_19[189], stage1_19[190]},
      {stage1_20[28]},
      {stage1_21[114], stage1_21[115], stage1_21[116], stage1_21[117], stage1_21[118], stage1_21[119]},
      {stage2_23[19],stage2_22[23],stage2_21[35],stage2_20[64],stage2_19[81]}
   );
   gpc615_5 gpc2596 (
      {stage1_19[191], stage1_19[192], stage1_19[193], stage1_19[194], stage1_19[195]},
      {stage1_20[29]},
      {stage1_21[120], stage1_21[121], stage1_21[122], stage1_21[123], stage1_21[124], stage1_21[125]},
      {stage2_23[20],stage2_22[24],stage2_21[36],stage2_20[65],stage2_19[82]}
   );
   gpc615_5 gpc2597 (
      {stage1_19[196], stage1_19[197], stage1_19[198], stage1_19[199], stage1_19[200]},
      {stage1_20[30]},
      {stage1_21[126], stage1_21[127], stage1_21[128], stage1_21[129], stage1_21[130], stage1_21[131]},
      {stage2_23[21],stage2_22[25],stage2_21[37],stage2_20[66],stage2_19[83]}
   );
   gpc615_5 gpc2598 (
      {stage1_19[201], stage1_19[202], stage1_19[203], stage1_19[204], stage1_19[205]},
      {stage1_20[31]},
      {stage1_21[132], stage1_21[133], stage1_21[134], stage1_21[135], stage1_21[136], stage1_21[137]},
      {stage2_23[22],stage2_22[26],stage2_21[38],stage2_20[67],stage2_19[84]}
   );
   gpc615_5 gpc2599 (
      {stage1_19[206], stage1_19[207], stage1_19[208], stage1_19[209], stage1_19[210]},
      {stage1_20[32]},
      {stage1_21[138], stage1_21[139], stage1_21[140], stage1_21[141], stage1_21[142], stage1_21[143]},
      {stage2_23[23],stage2_22[27],stage2_21[39],stage2_20[68],stage2_19[85]}
   );
   gpc615_5 gpc2600 (
      {stage1_19[211], stage1_19[212], stage1_19[213], stage1_19[214], stage1_19[215]},
      {stage1_20[33]},
      {stage1_21[144], stage1_21[145], stage1_21[146], stage1_21[147], stage1_21[148], stage1_21[149]},
      {stage2_23[24],stage2_22[28],stage2_21[40],stage2_20[69],stage2_19[86]}
   );
   gpc615_5 gpc2601 (
      {stage1_19[216], stage1_19[217], stage1_19[218], stage1_19[219], stage1_19[220]},
      {stage1_20[34]},
      {stage1_21[150], stage1_21[151], stage1_21[152], stage1_21[153], stage1_21[154], stage1_21[155]},
      {stage2_23[25],stage2_22[29],stage2_21[41],stage2_20[70],stage2_19[87]}
   );
   gpc615_5 gpc2602 (
      {stage1_19[221], stage1_19[222], stage1_19[223], stage1_19[224], stage1_19[225]},
      {stage1_20[35]},
      {stage1_21[156], stage1_21[157], stage1_21[158], stage1_21[159], stage1_21[160], stage1_21[161]},
      {stage2_23[26],stage2_22[30],stage2_21[42],stage2_20[71],stage2_19[88]}
   );
   gpc615_5 gpc2603 (
      {stage1_19[226], stage1_19[227], stage1_19[228], stage1_19[229], stage1_19[230]},
      {stage1_20[36]},
      {stage1_21[162], stage1_21[163], stage1_21[164], stage1_21[165], stage1_21[166], stage1_21[167]},
      {stage2_23[27],stage2_22[31],stage2_21[43],stage2_20[72],stage2_19[89]}
   );
   gpc615_5 gpc2604 (
      {stage1_19[231], stage1_19[232], stage1_19[233], stage1_19[234], stage1_19[235]},
      {stage1_20[37]},
      {stage1_21[168], stage1_21[169], stage1_21[170], stage1_21[171], stage1_21[172], stage1_21[173]},
      {stage2_23[28],stage2_22[32],stage2_21[44],stage2_20[73],stage2_19[90]}
   );
   gpc615_5 gpc2605 (
      {stage1_19[236], stage1_19[237], stage1_19[238], stage1_19[239], stage1_19[240]},
      {stage1_20[38]},
      {stage1_21[174], stage1_21[175], stage1_21[176], stage1_21[177], stage1_21[178], stage1_21[179]},
      {stage2_23[29],stage2_22[33],stage2_21[45],stage2_20[74],stage2_19[91]}
   );
   gpc615_5 gpc2606 (
      {stage1_19[241], stage1_19[242], stage1_19[243], stage1_19[244], stage1_19[245]},
      {stage1_20[39]},
      {stage1_21[180], stage1_21[181], stage1_21[182], stage1_21[183], stage1_21[184], stage1_21[185]},
      {stage2_23[30],stage2_22[34],stage2_21[46],stage2_20[75],stage2_19[92]}
   );
   gpc615_5 gpc2607 (
      {stage1_19[246], stage1_19[247], stage1_19[248], stage1_19[249], stage1_19[250]},
      {stage1_20[40]},
      {stage1_21[186], stage1_21[187], stage1_21[188], stage1_21[189], stage1_21[190], stage1_21[191]},
      {stage2_23[31],stage2_22[35],stage2_21[47],stage2_20[76],stage2_19[93]}
   );
   gpc615_5 gpc2608 (
      {stage1_19[251], stage1_19[252], stage1_19[253], stage1_19[254], stage1_19[255]},
      {stage1_20[41]},
      {stage1_21[192], stage1_21[193], stage1_21[194], stage1_21[195], stage1_21[196], stage1_21[197]},
      {stage2_23[32],stage2_22[36],stage2_21[48],stage2_20[77],stage2_19[94]}
   );
   gpc615_5 gpc2609 (
      {stage1_19[256], stage1_19[257], stage1_19[258], stage1_19[259], stage1_19[260]},
      {stage1_20[42]},
      {stage1_21[198], stage1_21[199], stage1_21[200], stage1_21[201], stage1_21[202], stage1_21[203]},
      {stage2_23[33],stage2_22[37],stage2_21[49],stage2_20[78],stage2_19[95]}
   );
   gpc606_5 gpc2610 (
      {stage1_20[43], stage1_20[44], stage1_20[45], stage1_20[46], stage1_20[47], stage1_20[48]},
      {stage1_22[0], stage1_22[1], stage1_22[2], stage1_22[3], stage1_22[4], stage1_22[5]},
      {stage2_24[0],stage2_23[34],stage2_22[38],stage2_21[50],stage2_20[79]}
   );
   gpc606_5 gpc2611 (
      {stage1_20[49], stage1_20[50], stage1_20[51], stage1_20[52], stage1_20[53], stage1_20[54]},
      {stage1_22[6], stage1_22[7], stage1_22[8], stage1_22[9], stage1_22[10], stage1_22[11]},
      {stage2_24[1],stage2_23[35],stage2_22[39],stage2_21[51],stage2_20[80]}
   );
   gpc606_5 gpc2612 (
      {stage1_20[55], stage1_20[56], stage1_20[57], stage1_20[58], stage1_20[59], stage1_20[60]},
      {stage1_22[12], stage1_22[13], stage1_22[14], stage1_22[15], stage1_22[16], stage1_22[17]},
      {stage2_24[2],stage2_23[36],stage2_22[40],stage2_21[52],stage2_20[81]}
   );
   gpc606_5 gpc2613 (
      {stage1_20[61], stage1_20[62], stage1_20[63], stage1_20[64], stage1_20[65], stage1_20[66]},
      {stage1_22[18], stage1_22[19], stage1_22[20], stage1_22[21], stage1_22[22], stage1_22[23]},
      {stage2_24[3],stage2_23[37],stage2_22[41],stage2_21[53],stage2_20[82]}
   );
   gpc606_5 gpc2614 (
      {stage1_20[67], stage1_20[68], stage1_20[69], stage1_20[70], stage1_20[71], stage1_20[72]},
      {stage1_22[24], stage1_22[25], stage1_22[26], stage1_22[27], stage1_22[28], stage1_22[29]},
      {stage2_24[4],stage2_23[38],stage2_22[42],stage2_21[54],stage2_20[83]}
   );
   gpc606_5 gpc2615 (
      {stage1_20[73], stage1_20[74], stage1_20[75], stage1_20[76], stage1_20[77], stage1_20[78]},
      {stage1_22[30], stage1_22[31], stage1_22[32], stage1_22[33], stage1_22[34], stage1_22[35]},
      {stage2_24[5],stage2_23[39],stage2_22[43],stage2_21[55],stage2_20[84]}
   );
   gpc606_5 gpc2616 (
      {stage1_20[79], stage1_20[80], stage1_20[81], stage1_20[82], stage1_20[83], stage1_20[84]},
      {stage1_22[36], stage1_22[37], stage1_22[38], stage1_22[39], stage1_22[40], stage1_22[41]},
      {stage2_24[6],stage2_23[40],stage2_22[44],stage2_21[56],stage2_20[85]}
   );
   gpc606_5 gpc2617 (
      {stage1_20[85], stage1_20[86], stage1_20[87], stage1_20[88], stage1_20[89], stage1_20[90]},
      {stage1_22[42], stage1_22[43], stage1_22[44], stage1_22[45], stage1_22[46], stage1_22[47]},
      {stage2_24[7],stage2_23[41],stage2_22[45],stage2_21[57],stage2_20[86]}
   );
   gpc606_5 gpc2618 (
      {stage1_20[91], stage1_20[92], stage1_20[93], stage1_20[94], stage1_20[95], stage1_20[96]},
      {stage1_22[48], stage1_22[49], stage1_22[50], stage1_22[51], stage1_22[52], stage1_22[53]},
      {stage2_24[8],stage2_23[42],stage2_22[46],stage2_21[58],stage2_20[87]}
   );
   gpc606_5 gpc2619 (
      {stage1_20[97], stage1_20[98], stage1_20[99], stage1_20[100], stage1_20[101], stage1_20[102]},
      {stage1_22[54], stage1_22[55], stage1_22[56], stage1_22[57], stage1_22[58], stage1_22[59]},
      {stage2_24[9],stage2_23[43],stage2_22[47],stage2_21[59],stage2_20[88]}
   );
   gpc606_5 gpc2620 (
      {stage1_20[103], stage1_20[104], stage1_20[105], stage1_20[106], stage1_20[107], stage1_20[108]},
      {stage1_22[60], stage1_22[61], stage1_22[62], stage1_22[63], stage1_22[64], stage1_22[65]},
      {stage2_24[10],stage2_23[44],stage2_22[48],stage2_21[60],stage2_20[89]}
   );
   gpc606_5 gpc2621 (
      {stage1_20[109], stage1_20[110], stage1_20[111], stage1_20[112], stage1_20[113], stage1_20[114]},
      {stage1_22[66], stage1_22[67], stage1_22[68], stage1_22[69], stage1_22[70], stage1_22[71]},
      {stage2_24[11],stage2_23[45],stage2_22[49],stage2_21[61],stage2_20[90]}
   );
   gpc606_5 gpc2622 (
      {stage1_20[115], stage1_20[116], stage1_20[117], stage1_20[118], stage1_20[119], stage1_20[120]},
      {stage1_22[72], stage1_22[73], stage1_22[74], stage1_22[75], stage1_22[76], stage1_22[77]},
      {stage2_24[12],stage2_23[46],stage2_22[50],stage2_21[62],stage2_20[91]}
   );
   gpc606_5 gpc2623 (
      {stage1_20[121], stage1_20[122], stage1_20[123], stage1_20[124], stage1_20[125], stage1_20[126]},
      {stage1_22[78], stage1_22[79], stage1_22[80], stage1_22[81], stage1_22[82], stage1_22[83]},
      {stage2_24[13],stage2_23[47],stage2_22[51],stage2_21[63],stage2_20[92]}
   );
   gpc606_5 gpc2624 (
      {stage1_20[127], stage1_20[128], stage1_20[129], stage1_20[130], stage1_20[131], stage1_20[132]},
      {stage1_22[84], stage1_22[85], stage1_22[86], stage1_22[87], stage1_22[88], stage1_22[89]},
      {stage2_24[14],stage2_23[48],stage2_22[52],stage2_21[64],stage2_20[93]}
   );
   gpc606_5 gpc2625 (
      {stage1_20[133], stage1_20[134], stage1_20[135], stage1_20[136], stage1_20[137], stage1_20[138]},
      {stage1_22[90], stage1_22[91], stage1_22[92], stage1_22[93], stage1_22[94], stage1_22[95]},
      {stage2_24[15],stage2_23[49],stage2_22[53],stage2_21[65],stage2_20[94]}
   );
   gpc606_5 gpc2626 (
      {stage1_20[139], stage1_20[140], stage1_20[141], stage1_20[142], stage1_20[143], stage1_20[144]},
      {stage1_22[96], stage1_22[97], stage1_22[98], stage1_22[99], stage1_22[100], stage1_22[101]},
      {stage2_24[16],stage2_23[50],stage2_22[54],stage2_21[66],stage2_20[95]}
   );
   gpc606_5 gpc2627 (
      {stage1_20[145], stage1_20[146], stage1_20[147], stage1_20[148], stage1_20[149], stage1_20[150]},
      {stage1_22[102], stage1_22[103], stage1_22[104], stage1_22[105], stage1_22[106], stage1_22[107]},
      {stage2_24[17],stage2_23[51],stage2_22[55],stage2_21[67],stage2_20[96]}
   );
   gpc606_5 gpc2628 (
      {stage1_20[151], stage1_20[152], stage1_20[153], stage1_20[154], stage1_20[155], stage1_20[156]},
      {stage1_22[108], stage1_22[109], stage1_22[110], stage1_22[111], stage1_22[112], stage1_22[113]},
      {stage2_24[18],stage2_23[52],stage2_22[56],stage2_21[68],stage2_20[97]}
   );
   gpc606_5 gpc2629 (
      {stage1_20[157], stage1_20[158], stage1_20[159], stage1_20[160], stage1_20[161], stage1_20[162]},
      {stage1_22[114], stage1_22[115], stage1_22[116], stage1_22[117], stage1_22[118], stage1_22[119]},
      {stage2_24[19],stage2_23[53],stage2_22[57],stage2_21[69],stage2_20[98]}
   );
   gpc606_5 gpc2630 (
      {stage1_20[163], stage1_20[164], stage1_20[165], stage1_20[166], stage1_20[167], stage1_20[168]},
      {stage1_22[120], stage1_22[121], stage1_22[122], stage1_22[123], stage1_22[124], stage1_22[125]},
      {stage2_24[20],stage2_23[54],stage2_22[58],stage2_21[70],stage2_20[99]}
   );
   gpc606_5 gpc2631 (
      {stage1_20[169], stage1_20[170], stage1_20[171], stage1_20[172], stage1_20[173], stage1_20[174]},
      {stage1_22[126], stage1_22[127], stage1_22[128], stage1_22[129], stage1_22[130], stage1_22[131]},
      {stage2_24[21],stage2_23[55],stage2_22[59],stage2_21[71],stage2_20[100]}
   );
   gpc606_5 gpc2632 (
      {stage1_20[175], stage1_20[176], stage1_20[177], stage1_20[178], stage1_20[179], stage1_20[180]},
      {stage1_22[132], stage1_22[133], stage1_22[134], stage1_22[135], stage1_22[136], stage1_22[137]},
      {stage2_24[22],stage2_23[56],stage2_22[60],stage2_21[72],stage2_20[101]}
   );
   gpc606_5 gpc2633 (
      {stage1_20[181], stage1_20[182], stage1_20[183], stage1_20[184], stage1_20[185], stage1_20[186]},
      {stage1_22[138], stage1_22[139], stage1_22[140], stage1_22[141], stage1_22[142], stage1_22[143]},
      {stage2_24[23],stage2_23[57],stage2_22[61],stage2_21[73],stage2_20[102]}
   );
   gpc606_5 gpc2634 (
      {stage1_20[187], stage1_20[188], stage1_20[189], stage1_20[190], stage1_20[191], stage1_20[192]},
      {stage1_22[144], stage1_22[145], stage1_22[146], stage1_22[147], stage1_22[148], stage1_22[149]},
      {stage2_24[24],stage2_23[58],stage2_22[62],stage2_21[74],stage2_20[103]}
   );
   gpc606_5 gpc2635 (
      {stage1_20[193], stage1_20[194], stage1_20[195], stage1_20[196], stage1_20[197], stage1_20[198]},
      {stage1_22[150], stage1_22[151], stage1_22[152], stage1_22[153], stage1_22[154], stage1_22[155]},
      {stage2_24[25],stage2_23[59],stage2_22[63],stage2_21[75],stage2_20[104]}
   );
   gpc606_5 gpc2636 (
      {stage1_20[199], stage1_20[200], stage1_20[201], stage1_20[202], stage1_20[203], stage1_20[204]},
      {stage1_22[156], stage1_22[157], stage1_22[158], stage1_22[159], stage1_22[160], stage1_22[161]},
      {stage2_24[26],stage2_23[60],stage2_22[64],stage2_21[76],stage2_20[105]}
   );
   gpc606_5 gpc2637 (
      {stage1_20[205], stage1_20[206], stage1_20[207], stage1_20[208], stage1_20[209], stage1_20[210]},
      {stage1_22[162], stage1_22[163], stage1_22[164], stage1_22[165], stage1_22[166], stage1_22[167]},
      {stage2_24[27],stage2_23[61],stage2_22[65],stage2_21[77],stage2_20[106]}
   );
   gpc606_5 gpc2638 (
      {stage1_21[204], stage1_21[205], stage1_21[206], stage1_21[207], stage1_21[208], stage1_21[209]},
      {stage1_23[0], stage1_23[1], stage1_23[2], stage1_23[3], stage1_23[4], stage1_23[5]},
      {stage2_25[0],stage2_24[28],stage2_23[62],stage2_22[66],stage2_21[78]}
   );
   gpc606_5 gpc2639 (
      {stage1_21[210], stage1_21[211], stage1_21[212], stage1_21[213], stage1_21[214], stage1_21[215]},
      {stage1_23[6], stage1_23[7], stage1_23[8], stage1_23[9], stage1_23[10], stage1_23[11]},
      {stage2_25[1],stage2_24[29],stage2_23[63],stage2_22[67],stage2_21[79]}
   );
   gpc606_5 gpc2640 (
      {stage1_21[216], stage1_21[217], stage1_21[218], stage1_21[219], stage1_21[220], stage1_21[221]},
      {stage1_23[12], stage1_23[13], stage1_23[14], stage1_23[15], stage1_23[16], stage1_23[17]},
      {stage2_25[2],stage2_24[30],stage2_23[64],stage2_22[68],stage2_21[80]}
   );
   gpc615_5 gpc2641 (
      {stage1_21[222], stage1_21[223], stage1_21[224], stage1_21[225], stage1_21[226]},
      {stage1_22[168]},
      {stage1_23[18], stage1_23[19], stage1_23[20], stage1_23[21], stage1_23[22], stage1_23[23]},
      {stage2_25[3],stage2_24[31],stage2_23[65],stage2_22[69],stage2_21[81]}
   );
   gpc606_5 gpc2642 (
      {stage1_22[169], stage1_22[170], stage1_22[171], stage1_22[172], stage1_22[173], stage1_22[174]},
      {stage1_24[0], stage1_24[1], stage1_24[2], stage1_24[3], stage1_24[4], stage1_24[5]},
      {stage2_26[0],stage2_25[4],stage2_24[32],stage2_23[66],stage2_22[70]}
   );
   gpc606_5 gpc2643 (
      {stage1_22[175], stage1_22[176], stage1_22[177], stage1_22[178], stage1_22[179], stage1_22[180]},
      {stage1_24[6], stage1_24[7], stage1_24[8], stage1_24[9], stage1_24[10], stage1_24[11]},
      {stage2_26[1],stage2_25[5],stage2_24[33],stage2_23[67],stage2_22[71]}
   );
   gpc606_5 gpc2644 (
      {stage1_22[181], stage1_22[182], stage1_22[183], stage1_22[184], stage1_22[185], stage1_22[186]},
      {stage1_24[12], stage1_24[13], stage1_24[14], stage1_24[15], stage1_24[16], stage1_24[17]},
      {stage2_26[2],stage2_25[6],stage2_24[34],stage2_23[68],stage2_22[72]}
   );
   gpc606_5 gpc2645 (
      {stage1_22[187], stage1_22[188], stage1_22[189], stage1_22[190], stage1_22[191], stage1_22[192]},
      {stage1_24[18], stage1_24[19], stage1_24[20], stage1_24[21], stage1_24[22], stage1_24[23]},
      {stage2_26[3],stage2_25[7],stage2_24[35],stage2_23[69],stage2_22[73]}
   );
   gpc615_5 gpc2646 (
      {stage1_22[193], stage1_22[194], stage1_22[195], stage1_22[196], stage1_22[197]},
      {stage1_23[24]},
      {stage1_24[24], stage1_24[25], stage1_24[26], stage1_24[27], stage1_24[28], stage1_24[29]},
      {stage2_26[4],stage2_25[8],stage2_24[36],stage2_23[70],stage2_22[74]}
   );
   gpc615_5 gpc2647 (
      {stage1_22[198], stage1_22[199], stage1_22[200], stage1_22[201], stage1_22[202]},
      {stage1_23[25]},
      {stage1_24[30], stage1_24[31], stage1_24[32], stage1_24[33], stage1_24[34], stage1_24[35]},
      {stage2_26[5],stage2_25[9],stage2_24[37],stage2_23[71],stage2_22[75]}
   );
   gpc615_5 gpc2648 (
      {stage1_22[203], stage1_22[204], stage1_22[205], stage1_22[206], stage1_22[207]},
      {stage1_23[26]},
      {stage1_24[36], stage1_24[37], stage1_24[38], stage1_24[39], stage1_24[40], stage1_24[41]},
      {stage2_26[6],stage2_25[10],stage2_24[38],stage2_23[72],stage2_22[76]}
   );
   gpc615_5 gpc2649 (
      {stage1_22[208], stage1_22[209], stage1_22[210], stage1_22[211], stage1_22[212]},
      {stage1_23[27]},
      {stage1_24[42], stage1_24[43], stage1_24[44], stage1_24[45], stage1_24[46], stage1_24[47]},
      {stage2_26[7],stage2_25[11],stage2_24[39],stage2_23[73],stage2_22[77]}
   );
   gpc615_5 gpc2650 (
      {stage1_22[213], stage1_22[214], stage1_22[215], stage1_22[216], stage1_22[217]},
      {stage1_23[28]},
      {stage1_24[48], stage1_24[49], stage1_24[50], stage1_24[51], stage1_24[52], stage1_24[53]},
      {stage2_26[8],stage2_25[12],stage2_24[40],stage2_23[74],stage2_22[78]}
   );
   gpc615_5 gpc2651 (
      {stage1_22[218], stage1_22[219], stage1_22[220], stage1_22[221], stage1_22[222]},
      {stage1_23[29]},
      {stage1_24[54], stage1_24[55], stage1_24[56], stage1_24[57], stage1_24[58], stage1_24[59]},
      {stage2_26[9],stage2_25[13],stage2_24[41],stage2_23[75],stage2_22[79]}
   );
   gpc615_5 gpc2652 (
      {stage1_22[223], stage1_22[224], stage1_22[225], stage1_22[226], stage1_22[227]},
      {stage1_23[30]},
      {stage1_24[60], stage1_24[61], stage1_24[62], stage1_24[63], stage1_24[64], stage1_24[65]},
      {stage2_26[10],stage2_25[14],stage2_24[42],stage2_23[76],stage2_22[80]}
   );
   gpc615_5 gpc2653 (
      {stage1_22[228], stage1_22[229], stage1_22[230], stage1_22[231], stage1_22[232]},
      {stage1_23[31]},
      {stage1_24[66], stage1_24[67], stage1_24[68], stage1_24[69], stage1_24[70], stage1_24[71]},
      {stage2_26[11],stage2_25[15],stage2_24[43],stage2_23[77],stage2_22[81]}
   );
   gpc615_5 gpc2654 (
      {stage1_22[233], stage1_22[234], stage1_22[235], stage1_22[236], stage1_22[237]},
      {stage1_23[32]},
      {stage1_24[72], stage1_24[73], stage1_24[74], stage1_24[75], stage1_24[76], stage1_24[77]},
      {stage2_26[12],stage2_25[16],stage2_24[44],stage2_23[78],stage2_22[82]}
   );
   gpc615_5 gpc2655 (
      {stage1_22[238], stage1_22[239], stage1_22[240], stage1_22[241], stage1_22[242]},
      {stage1_23[33]},
      {stage1_24[78], stage1_24[79], stage1_24[80], stage1_24[81], stage1_24[82], stage1_24[83]},
      {stage2_26[13],stage2_25[17],stage2_24[45],stage2_23[79],stage2_22[83]}
   );
   gpc615_5 gpc2656 (
      {stage1_22[243], stage1_22[244], stage1_22[245], stage1_22[246], stage1_22[247]},
      {stage1_23[34]},
      {stage1_24[84], stage1_24[85], stage1_24[86], stage1_24[87], stage1_24[88], stage1_24[89]},
      {stage2_26[14],stage2_25[18],stage2_24[46],stage2_23[80],stage2_22[84]}
   );
   gpc615_5 gpc2657 (
      {stage1_22[248], stage1_22[249], stage1_22[250], stage1_22[251], stage1_22[252]},
      {stage1_23[35]},
      {stage1_24[90], stage1_24[91], stage1_24[92], stage1_24[93], stage1_24[94], stage1_24[95]},
      {stage2_26[15],stage2_25[19],stage2_24[47],stage2_23[81],stage2_22[85]}
   );
   gpc615_5 gpc2658 (
      {stage1_22[253], stage1_22[254], stage1_22[255], stage1_22[256], stage1_22[257]},
      {stage1_23[36]},
      {stage1_24[96], stage1_24[97], stage1_24[98], stage1_24[99], stage1_24[100], stage1_24[101]},
      {stage2_26[16],stage2_25[20],stage2_24[48],stage2_23[82],stage2_22[86]}
   );
   gpc615_5 gpc2659 (
      {stage1_22[258], stage1_22[259], stage1_22[260], stage1_22[261], stage1_22[262]},
      {stage1_23[37]},
      {stage1_24[102], stage1_24[103], stage1_24[104], stage1_24[105], stage1_24[106], stage1_24[107]},
      {stage2_26[17],stage2_25[21],stage2_24[49],stage2_23[83],stage2_22[87]}
   );
   gpc615_5 gpc2660 (
      {stage1_22[263], stage1_22[264], stage1_22[265], stage1_22[266], stage1_22[267]},
      {stage1_23[38]},
      {stage1_24[108], stage1_24[109], stage1_24[110], stage1_24[111], stage1_24[112], stage1_24[113]},
      {stage2_26[18],stage2_25[22],stage2_24[50],stage2_23[84],stage2_22[88]}
   );
   gpc606_5 gpc2661 (
      {stage1_23[39], stage1_23[40], stage1_23[41], stage1_23[42], stage1_23[43], stage1_23[44]},
      {stage1_25[0], stage1_25[1], stage1_25[2], stage1_25[3], stage1_25[4], stage1_25[5]},
      {stage2_27[0],stage2_26[19],stage2_25[23],stage2_24[51],stage2_23[85]}
   );
   gpc606_5 gpc2662 (
      {stage1_23[45], stage1_23[46], stage1_23[47], stage1_23[48], stage1_23[49], stage1_23[50]},
      {stage1_25[6], stage1_25[7], stage1_25[8], stage1_25[9], stage1_25[10], stage1_25[11]},
      {stage2_27[1],stage2_26[20],stage2_25[24],stage2_24[52],stage2_23[86]}
   );
   gpc606_5 gpc2663 (
      {stage1_23[51], stage1_23[52], stage1_23[53], stage1_23[54], stage1_23[55], stage1_23[56]},
      {stage1_25[12], stage1_25[13], stage1_25[14], stage1_25[15], stage1_25[16], stage1_25[17]},
      {stage2_27[2],stage2_26[21],stage2_25[25],stage2_24[53],stage2_23[87]}
   );
   gpc606_5 gpc2664 (
      {stage1_23[57], stage1_23[58], stage1_23[59], stage1_23[60], stage1_23[61], stage1_23[62]},
      {stage1_25[18], stage1_25[19], stage1_25[20], stage1_25[21], stage1_25[22], stage1_25[23]},
      {stage2_27[3],stage2_26[22],stage2_25[26],stage2_24[54],stage2_23[88]}
   );
   gpc606_5 gpc2665 (
      {stage1_23[63], stage1_23[64], stage1_23[65], stage1_23[66], stage1_23[67], stage1_23[68]},
      {stage1_25[24], stage1_25[25], stage1_25[26], stage1_25[27], stage1_25[28], stage1_25[29]},
      {stage2_27[4],stage2_26[23],stage2_25[27],stage2_24[55],stage2_23[89]}
   );
   gpc606_5 gpc2666 (
      {stage1_23[69], stage1_23[70], stage1_23[71], stage1_23[72], stage1_23[73], stage1_23[74]},
      {stage1_25[30], stage1_25[31], stage1_25[32], stage1_25[33], stage1_25[34], stage1_25[35]},
      {stage2_27[5],stage2_26[24],stage2_25[28],stage2_24[56],stage2_23[90]}
   );
   gpc606_5 gpc2667 (
      {stage1_23[75], stage1_23[76], stage1_23[77], stage1_23[78], stage1_23[79], stage1_23[80]},
      {stage1_25[36], stage1_25[37], stage1_25[38], stage1_25[39], stage1_25[40], stage1_25[41]},
      {stage2_27[6],stage2_26[25],stage2_25[29],stage2_24[57],stage2_23[91]}
   );
   gpc606_5 gpc2668 (
      {stage1_23[81], stage1_23[82], stage1_23[83], stage1_23[84], stage1_23[85], stage1_23[86]},
      {stage1_25[42], stage1_25[43], stage1_25[44], stage1_25[45], stage1_25[46], stage1_25[47]},
      {stage2_27[7],stage2_26[26],stage2_25[30],stage2_24[58],stage2_23[92]}
   );
   gpc606_5 gpc2669 (
      {stage1_23[87], stage1_23[88], stage1_23[89], stage1_23[90], stage1_23[91], stage1_23[92]},
      {stage1_25[48], stage1_25[49], stage1_25[50], stage1_25[51], stage1_25[52], stage1_25[53]},
      {stage2_27[8],stage2_26[27],stage2_25[31],stage2_24[59],stage2_23[93]}
   );
   gpc606_5 gpc2670 (
      {stage1_23[93], stage1_23[94], stage1_23[95], stage1_23[96], stage1_23[97], stage1_23[98]},
      {stage1_25[54], stage1_25[55], stage1_25[56], stage1_25[57], stage1_25[58], stage1_25[59]},
      {stage2_27[9],stage2_26[28],stage2_25[32],stage2_24[60],stage2_23[94]}
   );
   gpc606_5 gpc2671 (
      {stage1_23[99], stage1_23[100], stage1_23[101], stage1_23[102], stage1_23[103], stage1_23[104]},
      {stage1_25[60], stage1_25[61], stage1_25[62], stage1_25[63], stage1_25[64], stage1_25[65]},
      {stage2_27[10],stage2_26[29],stage2_25[33],stage2_24[61],stage2_23[95]}
   );
   gpc606_5 gpc2672 (
      {stage1_23[105], stage1_23[106], stage1_23[107], stage1_23[108], stage1_23[109], stage1_23[110]},
      {stage1_25[66], stage1_25[67], stage1_25[68], stage1_25[69], stage1_25[70], stage1_25[71]},
      {stage2_27[11],stage2_26[30],stage2_25[34],stage2_24[62],stage2_23[96]}
   );
   gpc606_5 gpc2673 (
      {stage1_23[111], stage1_23[112], stage1_23[113], stage1_23[114], stage1_23[115], stage1_23[116]},
      {stage1_25[72], stage1_25[73], stage1_25[74], stage1_25[75], stage1_25[76], stage1_25[77]},
      {stage2_27[12],stage2_26[31],stage2_25[35],stage2_24[63],stage2_23[97]}
   );
   gpc606_5 gpc2674 (
      {stage1_23[117], stage1_23[118], stage1_23[119], stage1_23[120], stage1_23[121], stage1_23[122]},
      {stage1_25[78], stage1_25[79], stage1_25[80], stage1_25[81], stage1_25[82], stage1_25[83]},
      {stage2_27[13],stage2_26[32],stage2_25[36],stage2_24[64],stage2_23[98]}
   );
   gpc606_5 gpc2675 (
      {stage1_23[123], stage1_23[124], stage1_23[125], stage1_23[126], stage1_23[127], stage1_23[128]},
      {stage1_25[84], stage1_25[85], stage1_25[86], stage1_25[87], stage1_25[88], stage1_25[89]},
      {stage2_27[14],stage2_26[33],stage2_25[37],stage2_24[65],stage2_23[99]}
   );
   gpc606_5 gpc2676 (
      {stage1_23[129], stage1_23[130], stage1_23[131], stage1_23[132], stage1_23[133], stage1_23[134]},
      {stage1_25[90], stage1_25[91], stage1_25[92], stage1_25[93], stage1_25[94], stage1_25[95]},
      {stage2_27[15],stage2_26[34],stage2_25[38],stage2_24[66],stage2_23[100]}
   );
   gpc606_5 gpc2677 (
      {stage1_23[135], stage1_23[136], stage1_23[137], stage1_23[138], stage1_23[139], stage1_23[140]},
      {stage1_25[96], stage1_25[97], stage1_25[98], stage1_25[99], stage1_25[100], stage1_25[101]},
      {stage2_27[16],stage2_26[35],stage2_25[39],stage2_24[67],stage2_23[101]}
   );
   gpc615_5 gpc2678 (
      {stage1_23[141], stage1_23[142], stage1_23[143], stage1_23[144], stage1_23[145]},
      {stage1_24[114]},
      {stage1_25[102], stage1_25[103], stage1_25[104], stage1_25[105], stage1_25[106], stage1_25[107]},
      {stage2_27[17],stage2_26[36],stage2_25[40],stage2_24[68],stage2_23[102]}
   );
   gpc606_5 gpc2679 (
      {stage1_24[115], stage1_24[116], stage1_24[117], stage1_24[118], stage1_24[119], stage1_24[120]},
      {stage1_26[0], stage1_26[1], stage1_26[2], stage1_26[3], stage1_26[4], stage1_26[5]},
      {stage2_28[0],stage2_27[18],stage2_26[37],stage2_25[41],stage2_24[69]}
   );
   gpc606_5 gpc2680 (
      {stage1_24[121], stage1_24[122], stage1_24[123], stage1_24[124], stage1_24[125], stage1_24[126]},
      {stage1_26[6], stage1_26[7], stage1_26[8], stage1_26[9], stage1_26[10], stage1_26[11]},
      {stage2_28[1],stage2_27[19],stage2_26[38],stage2_25[42],stage2_24[70]}
   );
   gpc606_5 gpc2681 (
      {stage1_24[127], stage1_24[128], stage1_24[129], stage1_24[130], stage1_24[131], stage1_24[132]},
      {stage1_26[12], stage1_26[13], stage1_26[14], stage1_26[15], stage1_26[16], stage1_26[17]},
      {stage2_28[2],stage2_27[20],stage2_26[39],stage2_25[43],stage2_24[71]}
   );
   gpc606_5 gpc2682 (
      {stage1_24[133], stage1_24[134], stage1_24[135], stage1_24[136], stage1_24[137], stage1_24[138]},
      {stage1_26[18], stage1_26[19], stage1_26[20], stage1_26[21], stage1_26[22], stage1_26[23]},
      {stage2_28[3],stage2_27[21],stage2_26[40],stage2_25[44],stage2_24[72]}
   );
   gpc606_5 gpc2683 (
      {stage1_24[139], stage1_24[140], stage1_24[141], stage1_24[142], stage1_24[143], stage1_24[144]},
      {stage1_26[24], stage1_26[25], stage1_26[26], stage1_26[27], stage1_26[28], stage1_26[29]},
      {stage2_28[4],stage2_27[22],stage2_26[41],stage2_25[45],stage2_24[73]}
   );
   gpc606_5 gpc2684 (
      {stage1_24[145], stage1_24[146], stage1_24[147], stage1_24[148], stage1_24[149], stage1_24[150]},
      {stage1_26[30], stage1_26[31], stage1_26[32], stage1_26[33], stage1_26[34], stage1_26[35]},
      {stage2_28[5],stage2_27[23],stage2_26[42],stage2_25[46],stage2_24[74]}
   );
   gpc606_5 gpc2685 (
      {stage1_24[151], stage1_24[152], stage1_24[153], stage1_24[154], stage1_24[155], stage1_24[156]},
      {stage1_26[36], stage1_26[37], stage1_26[38], stage1_26[39], stage1_26[40], stage1_26[41]},
      {stage2_28[6],stage2_27[24],stage2_26[43],stage2_25[47],stage2_24[75]}
   );
   gpc606_5 gpc2686 (
      {stage1_24[157], stage1_24[158], stage1_24[159], stage1_24[160], stage1_24[161], stage1_24[162]},
      {stage1_26[42], stage1_26[43], stage1_26[44], stage1_26[45], stage1_26[46], stage1_26[47]},
      {stage2_28[7],stage2_27[25],stage2_26[44],stage2_25[48],stage2_24[76]}
   );
   gpc606_5 gpc2687 (
      {stage1_24[163], stage1_24[164], stage1_24[165], stage1_24[166], stage1_24[167], stage1_24[168]},
      {stage1_26[48], stage1_26[49], stage1_26[50], stage1_26[51], stage1_26[52], stage1_26[53]},
      {stage2_28[8],stage2_27[26],stage2_26[45],stage2_25[49],stage2_24[77]}
   );
   gpc606_5 gpc2688 (
      {stage1_24[169], stage1_24[170], stage1_24[171], stage1_24[172], stage1_24[173], stage1_24[174]},
      {stage1_26[54], stage1_26[55], stage1_26[56], stage1_26[57], stage1_26[58], stage1_26[59]},
      {stage2_28[9],stage2_27[27],stage2_26[46],stage2_25[50],stage2_24[78]}
   );
   gpc606_5 gpc2689 (
      {stage1_24[175], stage1_24[176], stage1_24[177], stage1_24[178], stage1_24[179], stage1_24[180]},
      {stage1_26[60], stage1_26[61], stage1_26[62], stage1_26[63], stage1_26[64], stage1_26[65]},
      {stage2_28[10],stage2_27[28],stage2_26[47],stage2_25[51],stage2_24[79]}
   );
   gpc606_5 gpc2690 (
      {stage1_24[181], stage1_24[182], stage1_24[183], stage1_24[184], stage1_24[185], stage1_24[186]},
      {stage1_26[66], stage1_26[67], stage1_26[68], stage1_26[69], stage1_26[70], stage1_26[71]},
      {stage2_28[11],stage2_27[29],stage2_26[48],stage2_25[52],stage2_24[80]}
   );
   gpc606_5 gpc2691 (
      {stage1_24[187], stage1_24[188], stage1_24[189], stage1_24[190], stage1_24[191], stage1_24[192]},
      {stage1_26[72], stage1_26[73], stage1_26[74], stage1_26[75], stage1_26[76], stage1_26[77]},
      {stage2_28[12],stage2_27[30],stage2_26[49],stage2_25[53],stage2_24[81]}
   );
   gpc606_5 gpc2692 (
      {stage1_24[193], stage1_24[194], stage1_24[195], stage1_24[196], stage1_24[197], stage1_24[198]},
      {stage1_26[78], stage1_26[79], stage1_26[80], stage1_26[81], stage1_26[82], stage1_26[83]},
      {stage2_28[13],stage2_27[31],stage2_26[50],stage2_25[54],stage2_24[82]}
   );
   gpc606_5 gpc2693 (
      {stage1_24[199], stage1_24[200], stage1_24[201], stage1_24[202], stage1_24[203], stage1_24[204]},
      {stage1_26[84], stage1_26[85], stage1_26[86], stage1_26[87], stage1_26[88], stage1_26[89]},
      {stage2_28[14],stage2_27[32],stage2_26[51],stage2_25[55],stage2_24[83]}
   );
   gpc606_5 gpc2694 (
      {stage1_24[205], stage1_24[206], stage1_24[207], stage1_24[208], stage1_24[209], stage1_24[210]},
      {stage1_26[90], stage1_26[91], stage1_26[92], stage1_26[93], stage1_26[94], stage1_26[95]},
      {stage2_28[15],stage2_27[33],stage2_26[52],stage2_25[56],stage2_24[84]}
   );
   gpc606_5 gpc2695 (
      {stage1_24[211], stage1_24[212], stage1_24[213], stage1_24[214], stage1_24[215], stage1_24[216]},
      {stage1_26[96], stage1_26[97], stage1_26[98], stage1_26[99], stage1_26[100], stage1_26[101]},
      {stage2_28[16],stage2_27[34],stage2_26[53],stage2_25[57],stage2_24[85]}
   );
   gpc606_5 gpc2696 (
      {stage1_25[108], stage1_25[109], stage1_25[110], stage1_25[111], stage1_25[112], stage1_25[113]},
      {stage1_27[0], stage1_27[1], stage1_27[2], stage1_27[3], stage1_27[4], stage1_27[5]},
      {stage2_29[0],stage2_28[17],stage2_27[35],stage2_26[54],stage2_25[58]}
   );
   gpc606_5 gpc2697 (
      {stage1_25[114], stage1_25[115], stage1_25[116], stage1_25[117], stage1_25[118], stage1_25[119]},
      {stage1_27[6], stage1_27[7], stage1_27[8], stage1_27[9], stage1_27[10], stage1_27[11]},
      {stage2_29[1],stage2_28[18],stage2_27[36],stage2_26[55],stage2_25[59]}
   );
   gpc606_5 gpc2698 (
      {stage1_25[120], stage1_25[121], stage1_25[122], stage1_25[123], stage1_25[124], stage1_25[125]},
      {stage1_27[12], stage1_27[13], stage1_27[14], stage1_27[15], stage1_27[16], stage1_27[17]},
      {stage2_29[2],stage2_28[19],stage2_27[37],stage2_26[56],stage2_25[60]}
   );
   gpc606_5 gpc2699 (
      {stage1_25[126], stage1_25[127], stage1_25[128], stage1_25[129], stage1_25[130], stage1_25[131]},
      {stage1_27[18], stage1_27[19], stage1_27[20], stage1_27[21], stage1_27[22], stage1_27[23]},
      {stage2_29[3],stage2_28[20],stage2_27[38],stage2_26[57],stage2_25[61]}
   );
   gpc606_5 gpc2700 (
      {stage1_25[132], stage1_25[133], stage1_25[134], stage1_25[135], stage1_25[136], stage1_25[137]},
      {stage1_27[24], stage1_27[25], stage1_27[26], stage1_27[27], stage1_27[28], stage1_27[29]},
      {stage2_29[4],stage2_28[21],stage2_27[39],stage2_26[58],stage2_25[62]}
   );
   gpc606_5 gpc2701 (
      {stage1_25[138], stage1_25[139], stage1_25[140], stage1_25[141], stage1_25[142], stage1_25[143]},
      {stage1_27[30], stage1_27[31], stage1_27[32], stage1_27[33], stage1_27[34], stage1_27[35]},
      {stage2_29[5],stage2_28[22],stage2_27[40],stage2_26[59],stage2_25[63]}
   );
   gpc606_5 gpc2702 (
      {stage1_25[144], stage1_25[145], stage1_25[146], stage1_25[147], stage1_25[148], stage1_25[149]},
      {stage1_27[36], stage1_27[37], stage1_27[38], stage1_27[39], stage1_27[40], stage1_27[41]},
      {stage2_29[6],stage2_28[23],stage2_27[41],stage2_26[60],stage2_25[64]}
   );
   gpc606_5 gpc2703 (
      {stage1_25[150], stage1_25[151], stage1_25[152], stage1_25[153], stage1_25[154], stage1_25[155]},
      {stage1_27[42], stage1_27[43], stage1_27[44], stage1_27[45], stage1_27[46], stage1_27[47]},
      {stage2_29[7],stage2_28[24],stage2_27[42],stage2_26[61],stage2_25[65]}
   );
   gpc606_5 gpc2704 (
      {stage1_25[156], stage1_25[157], stage1_25[158], stage1_25[159], stage1_25[160], stage1_25[161]},
      {stage1_27[48], stage1_27[49], stage1_27[50], stage1_27[51], stage1_27[52], stage1_27[53]},
      {stage2_29[8],stage2_28[25],stage2_27[43],stage2_26[62],stage2_25[66]}
   );
   gpc606_5 gpc2705 (
      {stage1_25[162], stage1_25[163], stage1_25[164], stage1_25[165], stage1_25[166], stage1_25[167]},
      {stage1_27[54], stage1_27[55], stage1_27[56], stage1_27[57], stage1_27[58], stage1_27[59]},
      {stage2_29[9],stage2_28[26],stage2_27[44],stage2_26[63],stage2_25[67]}
   );
   gpc606_5 gpc2706 (
      {stage1_25[168], stage1_25[169], stage1_25[170], stage1_25[171], stage1_25[172], stage1_25[173]},
      {stage1_27[60], stage1_27[61], stage1_27[62], stage1_27[63], stage1_27[64], stage1_27[65]},
      {stage2_29[10],stage2_28[27],stage2_27[45],stage2_26[64],stage2_25[68]}
   );
   gpc606_5 gpc2707 (
      {stage1_25[174], stage1_25[175], stage1_25[176], stage1_25[177], stage1_25[178], stage1_25[179]},
      {stage1_27[66], stage1_27[67], stage1_27[68], stage1_27[69], stage1_27[70], stage1_27[71]},
      {stage2_29[11],stage2_28[28],stage2_27[46],stage2_26[65],stage2_25[69]}
   );
   gpc606_5 gpc2708 (
      {stage1_25[180], stage1_25[181], stage1_25[182], stage1_25[183], stage1_25[184], stage1_25[185]},
      {stage1_27[72], stage1_27[73], stage1_27[74], stage1_27[75], stage1_27[76], stage1_27[77]},
      {stage2_29[12],stage2_28[29],stage2_27[47],stage2_26[66],stage2_25[70]}
   );
   gpc606_5 gpc2709 (
      {stage1_25[186], stage1_25[187], stage1_25[188], stage1_25[189], stage1_25[190], stage1_25[191]},
      {stage1_27[78], stage1_27[79], stage1_27[80], stage1_27[81], stage1_27[82], stage1_27[83]},
      {stage2_29[13],stage2_28[30],stage2_27[48],stage2_26[67],stage2_25[71]}
   );
   gpc606_5 gpc2710 (
      {stage1_25[192], stage1_25[193], stage1_25[194], stage1_25[195], stage1_25[196], stage1_25[197]},
      {stage1_27[84], stage1_27[85], stage1_27[86], stage1_27[87], stage1_27[88], stage1_27[89]},
      {stage2_29[14],stage2_28[31],stage2_27[49],stage2_26[68],stage2_25[72]}
   );
   gpc606_5 gpc2711 (
      {stage1_25[198], stage1_25[199], stage1_25[200], stage1_25[201], stage1_25[202], stage1_25[203]},
      {stage1_27[90], stage1_27[91], stage1_27[92], stage1_27[93], stage1_27[94], stage1_27[95]},
      {stage2_29[15],stage2_28[32],stage2_27[50],stage2_26[69],stage2_25[73]}
   );
   gpc606_5 gpc2712 (
      {stage1_25[204], stage1_25[205], stage1_25[206], stage1_25[207], stage1_25[208], stage1_25[209]},
      {stage1_27[96], stage1_27[97], stage1_27[98], stage1_27[99], stage1_27[100], stage1_27[101]},
      {stage2_29[16],stage2_28[33],stage2_27[51],stage2_26[70],stage2_25[74]}
   );
   gpc615_5 gpc2713 (
      {stage1_25[210], stage1_25[211], stage1_25[212], stage1_25[213], stage1_25[214]},
      {stage1_26[102]},
      {stage1_27[102], stage1_27[103], stage1_27[104], stage1_27[105], stage1_27[106], stage1_27[107]},
      {stage2_29[17],stage2_28[34],stage2_27[52],stage2_26[71],stage2_25[75]}
   );
   gpc615_5 gpc2714 (
      {stage1_25[215], stage1_25[216], stage1_25[217], stage1_25[218], stage1_25[219]},
      {stage1_26[103]},
      {stage1_27[108], stage1_27[109], stage1_27[110], stage1_27[111], stage1_27[112], stage1_27[113]},
      {stage2_29[18],stage2_28[35],stage2_27[53],stage2_26[72],stage2_25[76]}
   );
   gpc615_5 gpc2715 (
      {stage1_25[220], stage1_25[221], stage1_25[222], stage1_25[223], stage1_25[224]},
      {stage1_26[104]},
      {stage1_27[114], stage1_27[115], stage1_27[116], stage1_27[117], stage1_27[118], stage1_27[119]},
      {stage2_29[19],stage2_28[36],stage2_27[54],stage2_26[73],stage2_25[77]}
   );
   gpc615_5 gpc2716 (
      {stage1_25[225], stage1_25[226], stage1_25[227], stage1_25[228], stage1_25[229]},
      {stage1_26[105]},
      {stage1_27[120], stage1_27[121], stage1_27[122], stage1_27[123], stage1_27[124], stage1_27[125]},
      {stage2_29[20],stage2_28[37],stage2_27[55],stage2_26[74],stage2_25[78]}
   );
   gpc615_5 gpc2717 (
      {stage1_25[230], stage1_25[231], stage1_25[232], stage1_25[233], stage1_25[234]},
      {stage1_26[106]},
      {stage1_27[126], stage1_27[127], stage1_27[128], stage1_27[129], stage1_27[130], stage1_27[131]},
      {stage2_29[21],stage2_28[38],stage2_27[56],stage2_26[75],stage2_25[79]}
   );
   gpc615_5 gpc2718 (
      {stage1_25[235], stage1_25[236], stage1_25[237], stage1_25[238], stage1_25[239]},
      {stage1_26[107]},
      {stage1_27[132], stage1_27[133], stage1_27[134], stage1_27[135], stage1_27[136], stage1_27[137]},
      {stage2_29[22],stage2_28[39],stage2_27[57],stage2_26[76],stage2_25[80]}
   );
   gpc615_5 gpc2719 (
      {stage1_25[240], stage1_25[241], stage1_25[242], stage1_25[243], stage1_25[244]},
      {stage1_26[108]},
      {stage1_27[138], stage1_27[139], stage1_27[140], stage1_27[141], stage1_27[142], stage1_27[143]},
      {stage2_29[23],stage2_28[40],stage2_27[58],stage2_26[77],stage2_25[81]}
   );
   gpc615_5 gpc2720 (
      {stage1_25[245], stage1_25[246], stage1_25[247], stage1_25[248], stage1_25[249]},
      {stage1_26[109]},
      {stage1_27[144], stage1_27[145], stage1_27[146], stage1_27[147], stage1_27[148], stage1_27[149]},
      {stage2_29[24],stage2_28[41],stage2_27[59],stage2_26[78],stage2_25[82]}
   );
   gpc615_5 gpc2721 (
      {stage1_25[250], stage1_25[251], stage1_25[252], stage1_25[253], stage1_25[254]},
      {stage1_26[110]},
      {stage1_27[150], stage1_27[151], stage1_27[152], stage1_27[153], stage1_27[154], stage1_27[155]},
      {stage2_29[25],stage2_28[42],stage2_27[60],stage2_26[79],stage2_25[83]}
   );
   gpc615_5 gpc2722 (
      {stage1_26[111], stage1_26[112], stage1_26[113], stage1_26[114], stage1_26[115]},
      {stage1_27[156]},
      {stage1_28[0], stage1_28[1], stage1_28[2], stage1_28[3], stage1_28[4], stage1_28[5]},
      {stage2_30[0],stage2_29[26],stage2_28[43],stage2_27[61],stage2_26[80]}
   );
   gpc615_5 gpc2723 (
      {stage1_26[116], stage1_26[117], stage1_26[118], stage1_26[119], stage1_26[120]},
      {stage1_27[157]},
      {stage1_28[6], stage1_28[7], stage1_28[8], stage1_28[9], stage1_28[10], stage1_28[11]},
      {stage2_30[1],stage2_29[27],stage2_28[44],stage2_27[62],stage2_26[81]}
   );
   gpc615_5 gpc2724 (
      {stage1_26[121], stage1_26[122], stage1_26[123], stage1_26[124], stage1_26[125]},
      {stage1_27[158]},
      {stage1_28[12], stage1_28[13], stage1_28[14], stage1_28[15], stage1_28[16], stage1_28[17]},
      {stage2_30[2],stage2_29[28],stage2_28[45],stage2_27[63],stage2_26[82]}
   );
   gpc615_5 gpc2725 (
      {stage1_26[126], stage1_26[127], stage1_26[128], stage1_26[129], stage1_26[130]},
      {stage1_27[159]},
      {stage1_28[18], stage1_28[19], stage1_28[20], stage1_28[21], stage1_28[22], stage1_28[23]},
      {stage2_30[3],stage2_29[29],stage2_28[46],stage2_27[64],stage2_26[83]}
   );
   gpc615_5 gpc2726 (
      {stage1_26[131], stage1_26[132], stage1_26[133], stage1_26[134], stage1_26[135]},
      {stage1_27[160]},
      {stage1_28[24], stage1_28[25], stage1_28[26], stage1_28[27], stage1_28[28], stage1_28[29]},
      {stage2_30[4],stage2_29[30],stage2_28[47],stage2_27[65],stage2_26[84]}
   );
   gpc615_5 gpc2727 (
      {stage1_26[136], stage1_26[137], stage1_26[138], stage1_26[139], stage1_26[140]},
      {stage1_27[161]},
      {stage1_28[30], stage1_28[31], stage1_28[32], stage1_28[33], stage1_28[34], stage1_28[35]},
      {stage2_30[5],stage2_29[31],stage2_28[48],stage2_27[66],stage2_26[85]}
   );
   gpc615_5 gpc2728 (
      {stage1_26[141], stage1_26[142], stage1_26[143], stage1_26[144], stage1_26[145]},
      {stage1_27[162]},
      {stage1_28[36], stage1_28[37], stage1_28[38], stage1_28[39], stage1_28[40], stage1_28[41]},
      {stage2_30[6],stage2_29[32],stage2_28[49],stage2_27[67],stage2_26[86]}
   );
   gpc615_5 gpc2729 (
      {stage1_26[146], stage1_26[147], stage1_26[148], stage1_26[149], stage1_26[150]},
      {stage1_27[163]},
      {stage1_28[42], stage1_28[43], stage1_28[44], stage1_28[45], stage1_28[46], stage1_28[47]},
      {stage2_30[7],stage2_29[33],stage2_28[50],stage2_27[68],stage2_26[87]}
   );
   gpc615_5 gpc2730 (
      {stage1_26[151], stage1_26[152], stage1_26[153], stage1_26[154], stage1_26[155]},
      {stage1_27[164]},
      {stage1_28[48], stage1_28[49], stage1_28[50], stage1_28[51], stage1_28[52], stage1_28[53]},
      {stage2_30[8],stage2_29[34],stage2_28[51],stage2_27[69],stage2_26[88]}
   );
   gpc615_5 gpc2731 (
      {stage1_26[156], stage1_26[157], stage1_26[158], stage1_26[159], stage1_26[160]},
      {stage1_27[165]},
      {stage1_28[54], stage1_28[55], stage1_28[56], stage1_28[57], stage1_28[58], stage1_28[59]},
      {stage2_30[9],stage2_29[35],stage2_28[52],stage2_27[70],stage2_26[89]}
   );
   gpc615_5 gpc2732 (
      {stage1_26[161], stage1_26[162], stage1_26[163], stage1_26[164], stage1_26[165]},
      {stage1_27[166]},
      {stage1_28[60], stage1_28[61], stage1_28[62], stage1_28[63], stage1_28[64], stage1_28[65]},
      {stage2_30[10],stage2_29[36],stage2_28[53],stage2_27[71],stage2_26[90]}
   );
   gpc615_5 gpc2733 (
      {stage1_26[166], stage1_26[167], stage1_26[168], stage1_26[169], stage1_26[170]},
      {stage1_27[167]},
      {stage1_28[66], stage1_28[67], stage1_28[68], stage1_28[69], stage1_28[70], stage1_28[71]},
      {stage2_30[11],stage2_29[37],stage2_28[54],stage2_27[72],stage2_26[91]}
   );
   gpc615_5 gpc2734 (
      {stage1_26[171], stage1_26[172], stage1_26[173], stage1_26[174], stage1_26[175]},
      {stage1_27[168]},
      {stage1_28[72], stage1_28[73], stage1_28[74], stage1_28[75], stage1_28[76], stage1_28[77]},
      {stage2_30[12],stage2_29[38],stage2_28[55],stage2_27[73],stage2_26[92]}
   );
   gpc615_5 gpc2735 (
      {stage1_26[176], stage1_26[177], stage1_26[178], stage1_26[179], stage1_26[180]},
      {stage1_27[169]},
      {stage1_28[78], stage1_28[79], stage1_28[80], stage1_28[81], stage1_28[82], stage1_28[83]},
      {stage2_30[13],stage2_29[39],stage2_28[56],stage2_27[74],stage2_26[93]}
   );
   gpc615_5 gpc2736 (
      {stage1_26[181], stage1_26[182], stage1_26[183], stage1_26[184], stage1_26[185]},
      {stage1_27[170]},
      {stage1_28[84], stage1_28[85], stage1_28[86], stage1_28[87], stage1_28[88], stage1_28[89]},
      {stage2_30[14],stage2_29[40],stage2_28[57],stage2_27[75],stage2_26[94]}
   );
   gpc615_5 gpc2737 (
      {stage1_27[171], stage1_27[172], stage1_27[173], stage1_27[174], stage1_27[175]},
      {stage1_28[90]},
      {stage1_29[0], stage1_29[1], stage1_29[2], stage1_29[3], stage1_29[4], stage1_29[5]},
      {stage2_31[0],stage2_30[15],stage2_29[41],stage2_28[58],stage2_27[76]}
   );
   gpc615_5 gpc2738 (
      {stage1_27[176], stage1_27[177], stage1_27[178], stage1_27[179], stage1_27[180]},
      {stage1_28[91]},
      {stage1_29[6], stage1_29[7], stage1_29[8], stage1_29[9], stage1_29[10], stage1_29[11]},
      {stage2_31[1],stage2_30[16],stage2_29[42],stage2_28[59],stage2_27[77]}
   );
   gpc615_5 gpc2739 (
      {stage1_27[181], stage1_27[182], stage1_27[183], stage1_27[184], stage1_27[185]},
      {stage1_28[92]},
      {stage1_29[12], stage1_29[13], stage1_29[14], stage1_29[15], stage1_29[16], stage1_29[17]},
      {stage2_31[2],stage2_30[17],stage2_29[43],stage2_28[60],stage2_27[78]}
   );
   gpc615_5 gpc2740 (
      {stage1_27[186], stage1_27[187], stage1_27[188], stage1_27[189], stage1_27[190]},
      {stage1_28[93]},
      {stage1_29[18], stage1_29[19], stage1_29[20], stage1_29[21], stage1_29[22], stage1_29[23]},
      {stage2_31[3],stage2_30[18],stage2_29[44],stage2_28[61],stage2_27[79]}
   );
   gpc615_5 gpc2741 (
      {stage1_27[191], stage1_27[192], stage1_27[193], stage1_27[194], stage1_27[195]},
      {stage1_28[94]},
      {stage1_29[24], stage1_29[25], stage1_29[26], stage1_29[27], stage1_29[28], stage1_29[29]},
      {stage2_31[4],stage2_30[19],stage2_29[45],stage2_28[62],stage2_27[80]}
   );
   gpc606_5 gpc2742 (
      {stage1_28[95], stage1_28[96], stage1_28[97], stage1_28[98], stage1_28[99], stage1_28[100]},
      {stage1_30[0], stage1_30[1], stage1_30[2], stage1_30[3], stage1_30[4], stage1_30[5]},
      {stage2_32[0],stage2_31[5],stage2_30[20],stage2_29[46],stage2_28[63]}
   );
   gpc606_5 gpc2743 (
      {stage1_28[101], stage1_28[102], stage1_28[103], stage1_28[104], stage1_28[105], stage1_28[106]},
      {stage1_30[6], stage1_30[7], stage1_30[8], stage1_30[9], stage1_30[10], stage1_30[11]},
      {stage2_32[1],stage2_31[6],stage2_30[21],stage2_29[47],stage2_28[64]}
   );
   gpc606_5 gpc2744 (
      {stage1_28[107], stage1_28[108], stage1_28[109], stage1_28[110], stage1_28[111], stage1_28[112]},
      {stage1_30[12], stage1_30[13], stage1_30[14], stage1_30[15], stage1_30[16], stage1_30[17]},
      {stage2_32[2],stage2_31[7],stage2_30[22],stage2_29[48],stage2_28[65]}
   );
   gpc606_5 gpc2745 (
      {stage1_28[113], stage1_28[114], stage1_28[115], stage1_28[116], stage1_28[117], stage1_28[118]},
      {stage1_30[18], stage1_30[19], stage1_30[20], stage1_30[21], stage1_30[22], stage1_30[23]},
      {stage2_32[3],stage2_31[8],stage2_30[23],stage2_29[49],stage2_28[66]}
   );
   gpc606_5 gpc2746 (
      {stage1_28[119], stage1_28[120], stage1_28[121], stage1_28[122], stage1_28[123], stage1_28[124]},
      {stage1_30[24], stage1_30[25], stage1_30[26], stage1_30[27], stage1_30[28], stage1_30[29]},
      {stage2_32[4],stage2_31[9],stage2_30[24],stage2_29[50],stage2_28[67]}
   );
   gpc606_5 gpc2747 (
      {stage1_28[125], stage1_28[126], stage1_28[127], stage1_28[128], stage1_28[129], stage1_28[130]},
      {stage1_30[30], stage1_30[31], stage1_30[32], stage1_30[33], stage1_30[34], stage1_30[35]},
      {stage2_32[5],stage2_31[10],stage2_30[25],stage2_29[51],stage2_28[68]}
   );
   gpc606_5 gpc2748 (
      {stage1_28[131], stage1_28[132], stage1_28[133], stage1_28[134], stage1_28[135], stage1_28[136]},
      {stage1_30[36], stage1_30[37], stage1_30[38], stage1_30[39], stage1_30[40], stage1_30[41]},
      {stage2_32[6],stage2_31[11],stage2_30[26],stage2_29[52],stage2_28[69]}
   );
   gpc606_5 gpc2749 (
      {stage1_28[137], stage1_28[138], stage1_28[139], stage1_28[140], stage1_28[141], stage1_28[142]},
      {stage1_30[42], stage1_30[43], stage1_30[44], stage1_30[45], stage1_30[46], stage1_30[47]},
      {stage2_32[7],stage2_31[12],stage2_30[27],stage2_29[53],stage2_28[70]}
   );
   gpc606_5 gpc2750 (
      {stage1_28[143], stage1_28[144], stage1_28[145], stage1_28[146], stage1_28[147], stage1_28[148]},
      {stage1_30[48], stage1_30[49], stage1_30[50], stage1_30[51], stage1_30[52], stage1_30[53]},
      {stage2_32[8],stage2_31[13],stage2_30[28],stage2_29[54],stage2_28[71]}
   );
   gpc606_5 gpc2751 (
      {stage1_29[30], stage1_29[31], stage1_29[32], stage1_29[33], stage1_29[34], stage1_29[35]},
      {stage1_31[0], stage1_31[1], stage1_31[2], stage1_31[3], stage1_31[4], stage1_31[5]},
      {stage2_33[0],stage2_32[9],stage2_31[14],stage2_30[29],stage2_29[55]}
   );
   gpc606_5 gpc2752 (
      {stage1_29[36], stage1_29[37], stage1_29[38], stage1_29[39], stage1_29[40], stage1_29[41]},
      {stage1_31[6], stage1_31[7], stage1_31[8], stage1_31[9], stage1_31[10], stage1_31[11]},
      {stage2_33[1],stage2_32[10],stage2_31[15],stage2_30[30],stage2_29[56]}
   );
   gpc606_5 gpc2753 (
      {stage1_29[42], stage1_29[43], stage1_29[44], stage1_29[45], stage1_29[46], stage1_29[47]},
      {stage1_31[12], stage1_31[13], stage1_31[14], stage1_31[15], stage1_31[16], stage1_31[17]},
      {stage2_33[2],stage2_32[11],stage2_31[16],stage2_30[31],stage2_29[57]}
   );
   gpc606_5 gpc2754 (
      {stage1_29[48], stage1_29[49], stage1_29[50], stage1_29[51], stage1_29[52], stage1_29[53]},
      {stage1_31[18], stage1_31[19], stage1_31[20], stage1_31[21], stage1_31[22], stage1_31[23]},
      {stage2_33[3],stage2_32[12],stage2_31[17],stage2_30[32],stage2_29[58]}
   );
   gpc606_5 gpc2755 (
      {stage1_29[54], stage1_29[55], stage1_29[56], stage1_29[57], stage1_29[58], stage1_29[59]},
      {stage1_31[24], stage1_31[25], stage1_31[26], stage1_31[27], stage1_31[28], stage1_31[29]},
      {stage2_33[4],stage2_32[13],stage2_31[18],stage2_30[33],stage2_29[59]}
   );
   gpc606_5 gpc2756 (
      {stage1_29[60], stage1_29[61], stage1_29[62], stage1_29[63], stage1_29[64], stage1_29[65]},
      {stage1_31[30], stage1_31[31], stage1_31[32], stage1_31[33], stage1_31[34], stage1_31[35]},
      {stage2_33[5],stage2_32[14],stage2_31[19],stage2_30[34],stage2_29[60]}
   );
   gpc606_5 gpc2757 (
      {stage1_29[66], stage1_29[67], stage1_29[68], stage1_29[69], stage1_29[70], stage1_29[71]},
      {stage1_31[36], stage1_31[37], stage1_31[38], stage1_31[39], stage1_31[40], stage1_31[41]},
      {stage2_33[6],stage2_32[15],stage2_31[20],stage2_30[35],stage2_29[61]}
   );
   gpc606_5 gpc2758 (
      {stage1_29[72], stage1_29[73], stage1_29[74], stage1_29[75], stage1_29[76], stage1_29[77]},
      {stage1_31[42], stage1_31[43], stage1_31[44], stage1_31[45], stage1_31[46], stage1_31[47]},
      {stage2_33[7],stage2_32[16],stage2_31[21],stage2_30[36],stage2_29[62]}
   );
   gpc606_5 gpc2759 (
      {stage1_29[78], stage1_29[79], stage1_29[80], stage1_29[81], stage1_29[82], stage1_29[83]},
      {stage1_31[48], stage1_31[49], stage1_31[50], stage1_31[51], stage1_31[52], stage1_31[53]},
      {stage2_33[8],stage2_32[17],stage2_31[22],stage2_30[37],stage2_29[63]}
   );
   gpc606_5 gpc2760 (
      {stage1_29[84], stage1_29[85], stage1_29[86], stage1_29[87], stage1_29[88], stage1_29[89]},
      {stage1_31[54], stage1_31[55], stage1_31[56], stage1_31[57], stage1_31[58], stage1_31[59]},
      {stage2_33[9],stage2_32[18],stage2_31[23],stage2_30[38],stage2_29[64]}
   );
   gpc606_5 gpc2761 (
      {stage1_29[90], stage1_29[91], stage1_29[92], stage1_29[93], stage1_29[94], stage1_29[95]},
      {stage1_31[60], stage1_31[61], stage1_31[62], stage1_31[63], stage1_31[64], stage1_31[65]},
      {stage2_33[10],stage2_32[19],stage2_31[24],stage2_30[39],stage2_29[65]}
   );
   gpc606_5 gpc2762 (
      {stage1_29[96], stage1_29[97], stage1_29[98], stage1_29[99], stage1_29[100], stage1_29[101]},
      {stage1_31[66], stage1_31[67], stage1_31[68], stage1_31[69], stage1_31[70], stage1_31[71]},
      {stage2_33[11],stage2_32[20],stage2_31[25],stage2_30[40],stage2_29[66]}
   );
   gpc606_5 gpc2763 (
      {stage1_29[102], stage1_29[103], stage1_29[104], stage1_29[105], stage1_29[106], stage1_29[107]},
      {stage1_31[72], stage1_31[73], stage1_31[74], stage1_31[75], stage1_31[76], stage1_31[77]},
      {stage2_33[12],stage2_32[21],stage2_31[26],stage2_30[41],stage2_29[67]}
   );
   gpc606_5 gpc2764 (
      {stage1_29[108], stage1_29[109], stage1_29[110], stage1_29[111], stage1_29[112], stage1_29[113]},
      {stage1_31[78], stage1_31[79], stage1_31[80], stage1_31[81], stage1_31[82], stage1_31[83]},
      {stage2_33[13],stage2_32[22],stage2_31[27],stage2_30[42],stage2_29[68]}
   );
   gpc606_5 gpc2765 (
      {stage1_29[114], stage1_29[115], stage1_29[116], stage1_29[117], stage1_29[118], stage1_29[119]},
      {stage1_31[84], stage1_31[85], stage1_31[86], stage1_31[87], stage1_31[88], stage1_31[89]},
      {stage2_33[14],stage2_32[23],stage2_31[28],stage2_30[43],stage2_29[69]}
   );
   gpc606_5 gpc2766 (
      {stage1_29[120], stage1_29[121], stage1_29[122], stage1_29[123], stage1_29[124], stage1_29[125]},
      {stage1_31[90], stage1_31[91], stage1_31[92], stage1_31[93], stage1_31[94], stage1_31[95]},
      {stage2_33[15],stage2_32[24],stage2_31[29],stage2_30[44],stage2_29[70]}
   );
   gpc606_5 gpc2767 (
      {stage1_29[126], stage1_29[127], stage1_29[128], stage1_29[129], stage1_29[130], stage1_29[131]},
      {stage1_31[96], stage1_31[97], stage1_31[98], stage1_31[99], stage1_31[100], stage1_31[101]},
      {stage2_33[16],stage2_32[25],stage2_31[30],stage2_30[45],stage2_29[71]}
   );
   gpc606_5 gpc2768 (
      {stage1_29[132], stage1_29[133], stage1_29[134], stage1_29[135], stage1_29[136], stage1_29[137]},
      {stage1_31[102], stage1_31[103], stage1_31[104], stage1_31[105], stage1_31[106], stage1_31[107]},
      {stage2_33[17],stage2_32[26],stage2_31[31],stage2_30[46],stage2_29[72]}
   );
   gpc606_5 gpc2769 (
      {stage1_29[138], stage1_29[139], stage1_29[140], stage1_29[141], stage1_29[142], stage1_29[143]},
      {stage1_31[108], stage1_31[109], stage1_31[110], stage1_31[111], stage1_31[112], stage1_31[113]},
      {stage2_33[18],stage2_32[27],stage2_31[32],stage2_30[47],stage2_29[73]}
   );
   gpc606_5 gpc2770 (
      {stage1_29[144], stage1_29[145], stage1_29[146], stage1_29[147], stage1_29[148], stage1_29[149]},
      {stage1_31[114], stage1_31[115], stage1_31[116], stage1_31[117], stage1_31[118], stage1_31[119]},
      {stage2_33[19],stage2_32[28],stage2_31[33],stage2_30[48],stage2_29[74]}
   );
   gpc606_5 gpc2771 (
      {stage1_29[150], stage1_29[151], stage1_29[152], stage1_29[153], stage1_29[154], stage1_29[155]},
      {stage1_31[120], stage1_31[121], stage1_31[122], stage1_31[123], stage1_31[124], stage1_31[125]},
      {stage2_33[20],stage2_32[29],stage2_31[34],stage2_30[49],stage2_29[75]}
   );
   gpc606_5 gpc2772 (
      {stage1_29[156], stage1_29[157], stage1_29[158], stage1_29[159], stage1_29[160], stage1_29[161]},
      {stage1_31[126], stage1_31[127], stage1_31[128], stage1_31[129], stage1_31[130], stage1_31[131]},
      {stage2_33[21],stage2_32[30],stage2_31[35],stage2_30[50],stage2_29[76]}
   );
   gpc606_5 gpc2773 (
      {stage1_29[162], stage1_29[163], stage1_29[164], stage1_29[165], stage1_29[166], stage1_29[167]},
      {stage1_31[132], stage1_31[133], stage1_31[134], stage1_31[135], stage1_31[136], stage1_31[137]},
      {stage2_33[22],stage2_32[31],stage2_31[36],stage2_30[51],stage2_29[77]}
   );
   gpc606_5 gpc2774 (
      {stage1_29[168], stage1_29[169], stage1_29[170], stage1_29[171], stage1_29[172], stage1_29[173]},
      {stage1_31[138], stage1_31[139], stage1_31[140], stage1_31[141], stage1_31[142], stage1_31[143]},
      {stage2_33[23],stage2_32[32],stage2_31[37],stage2_30[52],stage2_29[78]}
   );
   gpc606_5 gpc2775 (
      {stage1_29[174], stage1_29[175], stage1_29[176], stage1_29[177], stage1_29[178], stage1_29[179]},
      {stage1_31[144], stage1_31[145], stage1_31[146], stage1_31[147], stage1_31[148], stage1_31[149]},
      {stage2_33[24],stage2_32[33],stage2_31[38],stage2_30[53],stage2_29[79]}
   );
   gpc606_5 gpc2776 (
      {stage1_30[54], stage1_30[55], stage1_30[56], stage1_30[57], stage1_30[58], stage1_30[59]},
      {stage1_32[0], stage1_32[1], stage1_32[2], stage1_32[3], stage1_32[4], stage1_32[5]},
      {stage2_34[0],stage2_33[25],stage2_32[34],stage2_31[39],stage2_30[54]}
   );
   gpc606_5 gpc2777 (
      {stage1_30[60], stage1_30[61], stage1_30[62], stage1_30[63], stage1_30[64], stage1_30[65]},
      {stage1_32[6], stage1_32[7], stage1_32[8], stage1_32[9], stage1_32[10], stage1_32[11]},
      {stage2_34[1],stage2_33[26],stage2_32[35],stage2_31[40],stage2_30[55]}
   );
   gpc606_5 gpc2778 (
      {stage1_30[66], stage1_30[67], stage1_30[68], stage1_30[69], stage1_30[70], stage1_30[71]},
      {stage1_32[12], stage1_32[13], stage1_32[14], stage1_32[15], stage1_32[16], stage1_32[17]},
      {stage2_34[2],stage2_33[27],stage2_32[36],stage2_31[41],stage2_30[56]}
   );
   gpc606_5 gpc2779 (
      {stage1_30[72], stage1_30[73], stage1_30[74], stage1_30[75], stage1_30[76], stage1_30[77]},
      {stage1_32[18], stage1_32[19], stage1_32[20], stage1_32[21], stage1_32[22], stage1_32[23]},
      {stage2_34[3],stage2_33[28],stage2_32[37],stage2_31[42],stage2_30[57]}
   );
   gpc606_5 gpc2780 (
      {stage1_30[78], stage1_30[79], stage1_30[80], stage1_30[81], stage1_30[82], stage1_30[83]},
      {stage1_32[24], stage1_32[25], stage1_32[26], stage1_32[27], stage1_32[28], stage1_32[29]},
      {stage2_34[4],stage2_33[29],stage2_32[38],stage2_31[43],stage2_30[58]}
   );
   gpc606_5 gpc2781 (
      {stage1_30[84], stage1_30[85], stage1_30[86], stage1_30[87], stage1_30[88], stage1_30[89]},
      {stage1_32[30], stage1_32[31], stage1_32[32], stage1_32[33], stage1_32[34], stage1_32[35]},
      {stage2_34[5],stage2_33[30],stage2_32[39],stage2_31[44],stage2_30[59]}
   );
   gpc606_5 gpc2782 (
      {stage1_30[90], stage1_30[91], stage1_30[92], stage1_30[93], stage1_30[94], stage1_30[95]},
      {stage1_32[36], stage1_32[37], stage1_32[38], stage1_32[39], stage1_32[40], stage1_32[41]},
      {stage2_34[6],stage2_33[31],stage2_32[40],stage2_31[45],stage2_30[60]}
   );
   gpc606_5 gpc2783 (
      {stage1_30[96], stage1_30[97], stage1_30[98], stage1_30[99], stage1_30[100], stage1_30[101]},
      {stage1_32[42], stage1_32[43], stage1_32[44], stage1_32[45], stage1_32[46], stage1_32[47]},
      {stage2_34[7],stage2_33[32],stage2_32[41],stage2_31[46],stage2_30[61]}
   );
   gpc606_5 gpc2784 (
      {stage1_30[102], stage1_30[103], stage1_30[104], stage1_30[105], stage1_30[106], stage1_30[107]},
      {stage1_32[48], stage1_32[49], stage1_32[50], stage1_32[51], stage1_32[52], stage1_32[53]},
      {stage2_34[8],stage2_33[33],stage2_32[42],stage2_31[47],stage2_30[62]}
   );
   gpc606_5 gpc2785 (
      {stage1_30[108], stage1_30[109], stage1_30[110], stage1_30[111], stage1_30[112], stage1_30[113]},
      {stage1_32[54], stage1_32[55], stage1_32[56], stage1_32[57], stage1_32[58], stage1_32[59]},
      {stage2_34[9],stage2_33[34],stage2_32[43],stage2_31[48],stage2_30[63]}
   );
   gpc606_5 gpc2786 (
      {stage1_30[114], stage1_30[115], stage1_30[116], stage1_30[117], stage1_30[118], stage1_30[119]},
      {stage1_32[60], stage1_32[61], stage1_32[62], stage1_32[63], stage1_32[64], stage1_32[65]},
      {stage2_34[10],stage2_33[35],stage2_32[44],stage2_31[49],stage2_30[64]}
   );
   gpc606_5 gpc2787 (
      {stage1_30[120], stage1_30[121], stage1_30[122], stage1_30[123], stage1_30[124], stage1_30[125]},
      {stage1_32[66], stage1_32[67], stage1_32[68], stage1_32[69], stage1_32[70], stage1_32[71]},
      {stage2_34[11],stage2_33[36],stage2_32[45],stage2_31[50],stage2_30[65]}
   );
   gpc606_5 gpc2788 (
      {stage1_30[126], stage1_30[127], stage1_30[128], stage1_30[129], stage1_30[130], stage1_30[131]},
      {stage1_32[72], stage1_32[73], stage1_32[74], stage1_32[75], stage1_32[76], stage1_32[77]},
      {stage2_34[12],stage2_33[37],stage2_32[46],stage2_31[51],stage2_30[66]}
   );
   gpc606_5 gpc2789 (
      {stage1_30[132], stage1_30[133], stage1_30[134], stage1_30[135], stage1_30[136], stage1_30[137]},
      {stage1_32[78], stage1_32[79], stage1_32[80], stage1_32[81], stage1_32[82], stage1_32[83]},
      {stage2_34[13],stage2_33[38],stage2_32[47],stage2_31[52],stage2_30[67]}
   );
   gpc606_5 gpc2790 (
      {stage1_30[138], stage1_30[139], stage1_30[140], stage1_30[141], stage1_30[142], stage1_30[143]},
      {stage1_32[84], stage1_32[85], stage1_32[86], stage1_32[87], stage1_32[88], stage1_32[89]},
      {stage2_34[14],stage2_33[39],stage2_32[48],stage2_31[53],stage2_30[68]}
   );
   gpc606_5 gpc2791 (
      {stage1_30[144], stage1_30[145], stage1_30[146], stage1_30[147], stage1_30[148], stage1_30[149]},
      {stage1_32[90], stage1_32[91], stage1_32[92], stage1_32[93], stage1_32[94], stage1_32[95]},
      {stage2_34[15],stage2_33[40],stage2_32[49],stage2_31[54],stage2_30[69]}
   );
   gpc606_5 gpc2792 (
      {stage1_30[150], stage1_30[151], stage1_30[152], stage1_30[153], stage1_30[154], stage1_30[155]},
      {stage1_32[96], stage1_32[97], stage1_32[98], stage1_32[99], stage1_32[100], stage1_32[101]},
      {stage2_34[16],stage2_33[41],stage2_32[50],stage2_31[55],stage2_30[70]}
   );
   gpc606_5 gpc2793 (
      {stage1_30[156], stage1_30[157], stage1_30[158], stage1_30[159], stage1_30[160], stage1_30[161]},
      {stage1_32[102], stage1_32[103], stage1_32[104], stage1_32[105], stage1_32[106], stage1_32[107]},
      {stage2_34[17],stage2_33[42],stage2_32[51],stage2_31[56],stage2_30[71]}
   );
   gpc606_5 gpc2794 (
      {stage1_30[162], stage1_30[163], stage1_30[164], stage1_30[165], stage1_30[166], stage1_30[167]},
      {stage1_32[108], stage1_32[109], stage1_32[110], stage1_32[111], stage1_32[112], stage1_32[113]},
      {stage2_34[18],stage2_33[43],stage2_32[52],stage2_31[57],stage2_30[72]}
   );
   gpc606_5 gpc2795 (
      {stage1_30[168], stage1_30[169], stage1_30[170], stage1_30[171], stage1_30[172], stage1_30[173]},
      {stage1_32[114], stage1_32[115], stage1_32[116], stage1_32[117], stage1_32[118], stage1_32[119]},
      {stage2_34[19],stage2_33[44],stage2_32[53],stage2_31[58],stage2_30[73]}
   );
   gpc606_5 gpc2796 (
      {stage1_30[174], stage1_30[175], stage1_30[176], stage1_30[177], stage1_30[178], stage1_30[179]},
      {stage1_32[120], stage1_32[121], stage1_32[122], stage1_32[123], stage1_32[124], stage1_32[125]},
      {stage2_34[20],stage2_33[45],stage2_32[54],stage2_31[59],stage2_30[74]}
   );
   gpc606_5 gpc2797 (
      {stage1_30[180], stage1_30[181], stage1_30[182], stage1_30[183], stage1_30[184], stage1_30[185]},
      {stage1_32[126], stage1_32[127], stage1_32[128], stage1_32[129], stage1_32[130], stage1_32[131]},
      {stage2_34[21],stage2_33[46],stage2_32[55],stage2_31[60],stage2_30[75]}
   );
   gpc606_5 gpc2798 (
      {stage1_30[186], stage1_30[187], stage1_30[188], stage1_30[189], stage1_30[190], stage1_30[191]},
      {stage1_32[132], stage1_32[133], stage1_32[134], stage1_32[135], stage1_32[136], stage1_32[137]},
      {stage2_34[22],stage2_33[47],stage2_32[56],stage2_31[61],stage2_30[76]}
   );
   gpc606_5 gpc2799 (
      {stage1_31[150], stage1_31[151], stage1_31[152], stage1_31[153], stage1_31[154], stage1_31[155]},
      {stage1_33[0], stage1_33[1], stage1_33[2], stage1_33[3], stage1_33[4], stage1_33[5]},
      {stage2_35[0],stage2_34[23],stage2_33[48],stage2_32[57],stage2_31[62]}
   );
   gpc606_5 gpc2800 (
      {stage1_31[156], stage1_31[157], stage1_31[158], stage1_31[159], stage1_31[160], stage1_31[161]},
      {stage1_33[6], stage1_33[7], stage1_33[8], stage1_33[9], stage1_33[10], stage1_33[11]},
      {stage2_35[1],stage2_34[24],stage2_33[49],stage2_32[58],stage2_31[63]}
   );
   gpc606_5 gpc2801 (
      {stage1_31[162], stage1_31[163], stage1_31[164], stage1_31[165], stage1_31[166], stage1_31[167]},
      {stage1_33[12], stage1_33[13], stage1_33[14], stage1_33[15], stage1_33[16], stage1_33[17]},
      {stage2_35[2],stage2_34[25],stage2_33[50],stage2_32[59],stage2_31[64]}
   );
   gpc606_5 gpc2802 (
      {stage1_31[168], stage1_31[169], stage1_31[170], stage1_31[171], stage1_31[172], stage1_31[173]},
      {stage1_33[18], stage1_33[19], stage1_33[20], stage1_33[21], stage1_33[22], stage1_33[23]},
      {stage2_35[3],stage2_34[26],stage2_33[51],stage2_32[60],stage2_31[65]}
   );
   gpc606_5 gpc2803 (
      {stage1_31[174], stage1_31[175], stage1_31[176], stage1_31[177], stage1_31[178], stage1_31[179]},
      {stage1_33[24], stage1_33[25], stage1_33[26], stage1_33[27], stage1_33[28], stage1_33[29]},
      {stage2_35[4],stage2_34[27],stage2_33[52],stage2_32[61],stage2_31[66]}
   );
   gpc615_5 gpc2804 (
      {stage1_31[180], stage1_31[181], stage1_31[182], stage1_31[183], stage1_31[184]},
      {stage1_32[138]},
      {stage1_33[30], stage1_33[31], stage1_33[32], stage1_33[33], stage1_33[34], stage1_33[35]},
      {stage2_35[5],stage2_34[28],stage2_33[53],stage2_32[62],stage2_31[67]}
   );
   gpc615_5 gpc2805 (
      {stage1_31[185], stage1_31[186], stage1_31[187], stage1_31[188], stage1_31[189]},
      {stage1_32[139]},
      {stage1_33[36], stage1_33[37], stage1_33[38], stage1_33[39], stage1_33[40], stage1_33[41]},
      {stage2_35[6],stage2_34[29],stage2_33[54],stage2_32[63],stage2_31[68]}
   );
   gpc615_5 gpc2806 (
      {stage1_31[190], stage1_31[191], stage1_31[192], stage1_31[193], stage1_31[194]},
      {stage1_32[140]},
      {stage1_33[42], stage1_33[43], stage1_33[44], stage1_33[45], stage1_33[46], stage1_33[47]},
      {stage2_35[7],stage2_34[30],stage2_33[55],stage2_32[64],stage2_31[69]}
   );
   gpc615_5 gpc2807 (
      {stage1_31[195], stage1_31[196], stage1_31[197], stage1_31[198], stage1_31[199]},
      {stage1_32[141]},
      {stage1_33[48], stage1_33[49], stage1_33[50], stage1_33[51], stage1_33[52], stage1_33[53]},
      {stage2_35[8],stage2_34[31],stage2_33[56],stage2_32[65],stage2_31[70]}
   );
   gpc615_5 gpc2808 (
      {stage1_31[200], stage1_31[201], stage1_31[202], stage1_31[203], stage1_31[204]},
      {stage1_32[142]},
      {stage1_33[54], stage1_33[55], stage1_33[56], stage1_33[57], stage1_33[58], stage1_33[59]},
      {stage2_35[9],stage2_34[32],stage2_33[57],stage2_32[66],stage2_31[71]}
   );
   gpc615_5 gpc2809 (
      {stage1_31[205], stage1_31[206], stage1_31[207], stage1_31[208], stage1_31[209]},
      {stage1_32[143]},
      {stage1_33[60], stage1_33[61], stage1_33[62], stage1_33[63], stage1_33[64], stage1_33[65]},
      {stage2_35[10],stage2_34[33],stage2_33[58],stage2_32[67],stage2_31[72]}
   );
   gpc615_5 gpc2810 (
      {stage1_31[210], stage1_31[211], stage1_31[212], stage1_31[213], stage1_31[214]},
      {stage1_32[144]},
      {stage1_33[66], stage1_33[67], stage1_33[68], stage1_33[69], stage1_33[70], 1'b0},
      {stage2_35[11],stage2_34[34],stage2_33[59],stage2_32[68],stage2_31[73]}
   );
   gpc1_1 gpc2811 (
      {stage1_0[60]},
      {stage2_0[12]}
   );
   gpc1_1 gpc2812 (
      {stage1_0[61]},
      {stage2_0[13]}
   );
   gpc1_1 gpc2813 (
      {stage1_0[62]},
      {stage2_0[14]}
   );
   gpc1_1 gpc2814 (
      {stage1_0[63]},
      {stage2_0[15]}
   );
   gpc1_1 gpc2815 (
      {stage1_0[64]},
      {stage2_0[16]}
   );
   gpc1_1 gpc2816 (
      {stage1_0[65]},
      {stage2_0[17]}
   );
   gpc1_1 gpc2817 (
      {stage1_0[66]},
      {stage2_0[18]}
   );
   gpc1_1 gpc2818 (
      {stage1_0[67]},
      {stage2_0[19]}
   );
   gpc1_1 gpc2819 (
      {stage1_0[68]},
      {stage2_0[20]}
   );
   gpc1_1 gpc2820 (
      {stage1_0[69]},
      {stage2_0[21]}
   );
   gpc1_1 gpc2821 (
      {stage1_0[70]},
      {stage2_0[22]}
   );
   gpc1_1 gpc2822 (
      {stage1_0[71]},
      {stage2_0[23]}
   );
   gpc1_1 gpc2823 (
      {stage1_0[72]},
      {stage2_0[24]}
   );
   gpc1_1 gpc2824 (
      {stage1_0[73]},
      {stage2_0[25]}
   );
   gpc1_1 gpc2825 (
      {stage1_0[74]},
      {stage2_0[26]}
   );
   gpc1_1 gpc2826 (
      {stage1_0[75]},
      {stage2_0[27]}
   );
   gpc1_1 gpc2827 (
      {stage1_0[76]},
      {stage2_0[28]}
   );
   gpc1_1 gpc2828 (
      {stage1_0[77]},
      {stage2_0[29]}
   );
   gpc1_1 gpc2829 (
      {stage1_0[78]},
      {stage2_0[30]}
   );
   gpc1_1 gpc2830 (
      {stage1_0[79]},
      {stage2_0[31]}
   );
   gpc1_1 gpc2831 (
      {stage1_0[80]},
      {stage2_0[32]}
   );
   gpc1_1 gpc2832 (
      {stage1_0[81]},
      {stage2_0[33]}
   );
   gpc1_1 gpc2833 (
      {stage1_0[82]},
      {stage2_0[34]}
   );
   gpc1_1 gpc2834 (
      {stage1_0[83]},
      {stage2_0[35]}
   );
   gpc1_1 gpc2835 (
      {stage1_0[84]},
      {stage2_0[36]}
   );
   gpc1_1 gpc2836 (
      {stage1_0[85]},
      {stage2_0[37]}
   );
   gpc1_1 gpc2837 (
      {stage1_0[86]},
      {stage2_0[38]}
   );
   gpc1_1 gpc2838 (
      {stage1_0[87]},
      {stage2_0[39]}
   );
   gpc1_1 gpc2839 (
      {stage1_0[88]},
      {stage2_0[40]}
   );
   gpc1_1 gpc2840 (
      {stage1_0[89]},
      {stage2_0[41]}
   );
   gpc1_1 gpc2841 (
      {stage1_0[90]},
      {stage2_0[42]}
   );
   gpc1_1 gpc2842 (
      {stage1_0[91]},
      {stage2_0[43]}
   );
   gpc1_1 gpc2843 (
      {stage1_0[92]},
      {stage2_0[44]}
   );
   gpc1_1 gpc2844 (
      {stage1_0[93]},
      {stage2_0[45]}
   );
   gpc1_1 gpc2845 (
      {stage1_0[94]},
      {stage2_0[46]}
   );
   gpc1_1 gpc2846 (
      {stage1_0[95]},
      {stage2_0[47]}
   );
   gpc1_1 gpc2847 (
      {stage1_0[96]},
      {stage2_0[48]}
   );
   gpc1_1 gpc2848 (
      {stage1_0[97]},
      {stage2_0[49]}
   );
   gpc1_1 gpc2849 (
      {stage1_0[98]},
      {stage2_0[50]}
   );
   gpc1_1 gpc2850 (
      {stage1_0[99]},
      {stage2_0[51]}
   );
   gpc1_1 gpc2851 (
      {stage1_0[100]},
      {stage2_0[52]}
   );
   gpc1_1 gpc2852 (
      {stage1_0[101]},
      {stage2_0[53]}
   );
   gpc1_1 gpc2853 (
      {stage1_0[102]},
      {stage2_0[54]}
   );
   gpc1_1 gpc2854 (
      {stage1_0[103]},
      {stage2_0[55]}
   );
   gpc1_1 gpc2855 (
      {stage1_0[104]},
      {stage2_0[56]}
   );
   gpc1_1 gpc2856 (
      {stage1_0[105]},
      {stage2_0[57]}
   );
   gpc1_1 gpc2857 (
      {stage1_0[106]},
      {stage2_0[58]}
   );
   gpc1_1 gpc2858 (
      {stage1_0[107]},
      {stage2_0[59]}
   );
   gpc1_1 gpc2859 (
      {stage1_0[108]},
      {stage2_0[60]}
   );
   gpc1_1 gpc2860 (
      {stage1_0[109]},
      {stage2_0[61]}
   );
   gpc1_1 gpc2861 (
      {stage1_0[110]},
      {stage2_0[62]}
   );
   gpc1_1 gpc2862 (
      {stage1_1[182]},
      {stage2_1[39]}
   );
   gpc1_1 gpc2863 (
      {stage1_1[183]},
      {stage2_1[40]}
   );
   gpc1_1 gpc2864 (
      {stage1_1[184]},
      {stage2_1[41]}
   );
   gpc1_1 gpc2865 (
      {stage1_1[185]},
      {stage2_1[42]}
   );
   gpc1_1 gpc2866 (
      {stage1_1[186]},
      {stage2_1[43]}
   );
   gpc1_1 gpc2867 (
      {stage1_1[187]},
      {stage2_1[44]}
   );
   gpc1_1 gpc2868 (
      {stage1_1[188]},
      {stage2_1[45]}
   );
   gpc1_1 gpc2869 (
      {stage1_1[189]},
      {stage2_1[46]}
   );
   gpc1_1 gpc2870 (
      {stage1_1[190]},
      {stage2_1[47]}
   );
   gpc1_1 gpc2871 (
      {stage1_1[191]},
      {stage2_1[48]}
   );
   gpc1_1 gpc2872 (
      {stage1_1[192]},
      {stage2_1[49]}
   );
   gpc1_1 gpc2873 (
      {stage1_1[193]},
      {stage2_1[50]}
   );
   gpc1_1 gpc2874 (
      {stage1_1[194]},
      {stage2_1[51]}
   );
   gpc1_1 gpc2875 (
      {stage1_1[195]},
      {stage2_1[52]}
   );
   gpc1_1 gpc2876 (
      {stage1_1[196]},
      {stage2_1[53]}
   );
   gpc1_1 gpc2877 (
      {stage1_1[197]},
      {stage2_1[54]}
   );
   gpc1_1 gpc2878 (
      {stage1_1[198]},
      {stage2_1[55]}
   );
   gpc1_1 gpc2879 (
      {stage1_2[152]},
      {stage2_2[59]}
   );
   gpc1_1 gpc2880 (
      {stage1_2[153]},
      {stage2_2[60]}
   );
   gpc1_1 gpc2881 (
      {stage1_2[154]},
      {stage2_2[61]}
   );
   gpc1_1 gpc2882 (
      {stage1_2[155]},
      {stage2_2[62]}
   );
   gpc1_1 gpc2883 (
      {stage1_2[156]},
      {stage2_2[63]}
   );
   gpc1_1 gpc2884 (
      {stage1_2[157]},
      {stage2_2[64]}
   );
   gpc1_1 gpc2885 (
      {stage1_2[158]},
      {stage2_2[65]}
   );
   gpc1_1 gpc2886 (
      {stage1_2[159]},
      {stage2_2[66]}
   );
   gpc1_1 gpc2887 (
      {stage1_2[160]},
      {stage2_2[67]}
   );
   gpc1_1 gpc2888 (
      {stage1_2[161]},
      {stage2_2[68]}
   );
   gpc1_1 gpc2889 (
      {stage1_2[162]},
      {stage2_2[69]}
   );
   gpc1_1 gpc2890 (
      {stage1_2[163]},
      {stage2_2[70]}
   );
   gpc1_1 gpc2891 (
      {stage1_2[164]},
      {stage2_2[71]}
   );
   gpc1_1 gpc2892 (
      {stage1_2[165]},
      {stage2_2[72]}
   );
   gpc1_1 gpc2893 (
      {stage1_2[166]},
      {stage2_2[73]}
   );
   gpc1_1 gpc2894 (
      {stage1_2[167]},
      {stage2_2[74]}
   );
   gpc1_1 gpc2895 (
      {stage1_2[168]},
      {stage2_2[75]}
   );
   gpc1_1 gpc2896 (
      {stage1_2[169]},
      {stage2_2[76]}
   );
   gpc1_1 gpc2897 (
      {stage1_2[170]},
      {stage2_2[77]}
   );
   gpc1_1 gpc2898 (
      {stage1_2[171]},
      {stage2_2[78]}
   );
   gpc1_1 gpc2899 (
      {stage1_2[172]},
      {stage2_2[79]}
   );
   gpc1_1 gpc2900 (
      {stage1_2[173]},
      {stage2_2[80]}
   );
   gpc1_1 gpc2901 (
      {stage1_2[174]},
      {stage2_2[81]}
   );
   gpc1_1 gpc2902 (
      {stage1_2[175]},
      {stage2_2[82]}
   );
   gpc1_1 gpc2903 (
      {stage1_2[176]},
      {stage2_2[83]}
   );
   gpc1_1 gpc2904 (
      {stage1_2[177]},
      {stage2_2[84]}
   );
   gpc1_1 gpc2905 (
      {stage1_2[178]},
      {stage2_2[85]}
   );
   gpc1_1 gpc2906 (
      {stage1_2[179]},
      {stage2_2[86]}
   );
   gpc1_1 gpc2907 (
      {stage1_2[180]},
      {stage2_2[87]}
   );
   gpc1_1 gpc2908 (
      {stage1_2[181]},
      {stage2_2[88]}
   );
   gpc1_1 gpc2909 (
      {stage1_2[182]},
      {stage2_2[89]}
   );
   gpc1_1 gpc2910 (
      {stage1_2[183]},
      {stage2_2[90]}
   );
   gpc1_1 gpc2911 (
      {stage1_2[184]},
      {stage2_2[91]}
   );
   gpc1_1 gpc2912 (
      {stage1_2[185]},
      {stage2_2[92]}
   );
   gpc1_1 gpc2913 (
      {stage1_2[186]},
      {stage2_2[93]}
   );
   gpc1_1 gpc2914 (
      {stage1_2[187]},
      {stage2_2[94]}
   );
   gpc1_1 gpc2915 (
      {stage1_4[217]},
      {stage2_4[91]}
   );
   gpc1_1 gpc2916 (
      {stage1_4[218]},
      {stage2_4[92]}
   );
   gpc1_1 gpc2917 (
      {stage1_4[219]},
      {stage2_4[93]}
   );
   gpc1_1 gpc2918 (
      {stage1_4[220]},
      {stage2_4[94]}
   );
   gpc1_1 gpc2919 (
      {stage1_4[221]},
      {stage2_4[95]}
   );
   gpc1_1 gpc2920 (
      {stage1_4[222]},
      {stage2_4[96]}
   );
   gpc1_1 gpc2921 (
      {stage1_4[223]},
      {stage2_4[97]}
   );
   gpc1_1 gpc2922 (
      {stage1_4[224]},
      {stage2_4[98]}
   );
   gpc1_1 gpc2923 (
      {stage1_4[225]},
      {stage2_4[99]}
   );
   gpc1_1 gpc2924 (
      {stage1_4[226]},
      {stage2_4[100]}
   );
   gpc1_1 gpc2925 (
      {stage1_4[227]},
      {stage2_4[101]}
   );
   gpc1_1 gpc2926 (
      {stage1_4[228]},
      {stage2_4[102]}
   );
   gpc1_1 gpc2927 (
      {stage1_4[229]},
      {stage2_4[103]}
   );
   gpc1_1 gpc2928 (
      {stage1_4[230]},
      {stage2_4[104]}
   );
   gpc1_1 gpc2929 (
      {stage1_4[231]},
      {stage2_4[105]}
   );
   gpc1_1 gpc2930 (
      {stage1_4[232]},
      {stage2_4[106]}
   );
   gpc1_1 gpc2931 (
      {stage1_4[233]},
      {stage2_4[107]}
   );
   gpc1_1 gpc2932 (
      {stage1_4[234]},
      {stage2_4[108]}
   );
   gpc1_1 gpc2933 (
      {stage1_4[235]},
      {stage2_4[109]}
   );
   gpc1_1 gpc2934 (
      {stage1_4[236]},
      {stage2_4[110]}
   );
   gpc1_1 gpc2935 (
      {stage1_4[237]},
      {stage2_4[111]}
   );
   gpc1_1 gpc2936 (
      {stage1_4[238]},
      {stage2_4[112]}
   );
   gpc1_1 gpc2937 (
      {stage1_4[239]},
      {stage2_4[113]}
   );
   gpc1_1 gpc2938 (
      {stage1_4[240]},
      {stage2_4[114]}
   );
   gpc1_1 gpc2939 (
      {stage1_4[241]},
      {stage2_4[115]}
   );
   gpc1_1 gpc2940 (
      {stage1_4[242]},
      {stage2_4[116]}
   );
   gpc1_1 gpc2941 (
      {stage1_4[243]},
      {stage2_4[117]}
   );
   gpc1_1 gpc2942 (
      {stage1_4[244]},
      {stage2_4[118]}
   );
   gpc1_1 gpc2943 (
      {stage1_7[166]},
      {stage2_7[89]}
   );
   gpc1_1 gpc2944 (
      {stage1_7[167]},
      {stage2_7[90]}
   );
   gpc1_1 gpc2945 (
      {stage1_7[168]},
      {stage2_7[91]}
   );
   gpc1_1 gpc2946 (
      {stage1_7[169]},
      {stage2_7[92]}
   );
   gpc1_1 gpc2947 (
      {stage1_7[170]},
      {stage2_7[93]}
   );
   gpc1_1 gpc2948 (
      {stage1_7[171]},
      {stage2_7[94]}
   );
   gpc1_1 gpc2949 (
      {stage1_7[172]},
      {stage2_7[95]}
   );
   gpc1_1 gpc2950 (
      {stage1_7[173]},
      {stage2_7[96]}
   );
   gpc1_1 gpc2951 (
      {stage1_7[174]},
      {stage2_7[97]}
   );
   gpc1_1 gpc2952 (
      {stage1_7[175]},
      {stage2_7[98]}
   );
   gpc1_1 gpc2953 (
      {stage1_7[176]},
      {stage2_7[99]}
   );
   gpc1_1 gpc2954 (
      {stage1_7[177]},
      {stage2_7[100]}
   );
   gpc1_1 gpc2955 (
      {stage1_7[178]},
      {stage2_7[101]}
   );
   gpc1_1 gpc2956 (
      {stage1_7[179]},
      {stage2_7[102]}
   );
   gpc1_1 gpc2957 (
      {stage1_7[180]},
      {stage2_7[103]}
   );
   gpc1_1 gpc2958 (
      {stage1_7[181]},
      {stage2_7[104]}
   );
   gpc1_1 gpc2959 (
      {stage1_7[182]},
      {stage2_7[105]}
   );
   gpc1_1 gpc2960 (
      {stage1_7[183]},
      {stage2_7[106]}
   );
   gpc1_1 gpc2961 (
      {stage1_7[184]},
      {stage2_7[107]}
   );
   gpc1_1 gpc2962 (
      {stage1_7[185]},
      {stage2_7[108]}
   );
   gpc1_1 gpc2963 (
      {stage1_9[210]},
      {stage2_9[106]}
   );
   gpc1_1 gpc2964 (
      {stage1_9[211]},
      {stage2_9[107]}
   );
   gpc1_1 gpc2965 (
      {stage1_11[161]},
      {stage2_11[71]}
   );
   gpc1_1 gpc2966 (
      {stage1_11[162]},
      {stage2_11[72]}
   );
   gpc1_1 gpc2967 (
      {stage1_11[163]},
      {stage2_11[73]}
   );
   gpc1_1 gpc2968 (
      {stage1_11[164]},
      {stage2_11[74]}
   );
   gpc1_1 gpc2969 (
      {stage1_11[165]},
      {stage2_11[75]}
   );
   gpc1_1 gpc2970 (
      {stage1_11[166]},
      {stage2_11[76]}
   );
   gpc1_1 gpc2971 (
      {stage1_11[167]},
      {stage2_11[77]}
   );
   gpc1_1 gpc2972 (
      {stage1_11[168]},
      {stage2_11[78]}
   );
   gpc1_1 gpc2973 (
      {stage1_11[169]},
      {stage2_11[79]}
   );
   gpc1_1 gpc2974 (
      {stage1_11[170]},
      {stage2_11[80]}
   );
   gpc1_1 gpc2975 (
      {stage1_11[171]},
      {stage2_11[81]}
   );
   gpc1_1 gpc2976 (
      {stage1_11[172]},
      {stage2_11[82]}
   );
   gpc1_1 gpc2977 (
      {stage1_11[173]},
      {stage2_11[83]}
   );
   gpc1_1 gpc2978 (
      {stage1_11[174]},
      {stage2_11[84]}
   );
   gpc1_1 gpc2979 (
      {stage1_11[175]},
      {stage2_11[85]}
   );
   gpc1_1 gpc2980 (
      {stage1_11[176]},
      {stage2_11[86]}
   );
   gpc1_1 gpc2981 (
      {stage1_11[177]},
      {stage2_11[87]}
   );
   gpc1_1 gpc2982 (
      {stage1_11[178]},
      {stage2_11[88]}
   );
   gpc1_1 gpc2983 (
      {stage1_11[179]},
      {stage2_11[89]}
   );
   gpc1_1 gpc2984 (
      {stage1_11[180]},
      {stage2_11[90]}
   );
   gpc1_1 gpc2985 (
      {stage1_11[181]},
      {stage2_11[91]}
   );
   gpc1_1 gpc2986 (
      {stage1_11[182]},
      {stage2_11[92]}
   );
   gpc1_1 gpc2987 (
      {stage1_11[183]},
      {stage2_11[93]}
   );
   gpc1_1 gpc2988 (
      {stage1_11[184]},
      {stage2_11[94]}
   );
   gpc1_1 gpc2989 (
      {stage1_11[185]},
      {stage2_11[95]}
   );
   gpc1_1 gpc2990 (
      {stage1_11[186]},
      {stage2_11[96]}
   );
   gpc1_1 gpc2991 (
      {stage1_11[187]},
      {stage2_11[97]}
   );
   gpc1_1 gpc2992 (
      {stage1_11[188]},
      {stage2_11[98]}
   );
   gpc1_1 gpc2993 (
      {stage1_11[189]},
      {stage2_11[99]}
   );
   gpc1_1 gpc2994 (
      {stage1_11[190]},
      {stage2_11[100]}
   );
   gpc1_1 gpc2995 (
      {stage1_11[191]},
      {stage2_11[101]}
   );
   gpc1_1 gpc2996 (
      {stage1_11[192]},
      {stage2_11[102]}
   );
   gpc1_1 gpc2997 (
      {stage1_11[193]},
      {stage2_11[103]}
   );
   gpc1_1 gpc2998 (
      {stage1_11[194]},
      {stage2_11[104]}
   );
   gpc1_1 gpc2999 (
      {stage1_11[195]},
      {stage2_11[105]}
   );
   gpc1_1 gpc3000 (
      {stage1_11[196]},
      {stage2_11[106]}
   );
   gpc1_1 gpc3001 (
      {stage1_11[197]},
      {stage2_11[107]}
   );
   gpc1_1 gpc3002 (
      {stage1_11[198]},
      {stage2_11[108]}
   );
   gpc1_1 gpc3003 (
      {stage1_11[199]},
      {stage2_11[109]}
   );
   gpc1_1 gpc3004 (
      {stage1_11[200]},
      {stage2_11[110]}
   );
   gpc1_1 gpc3005 (
      {stage1_11[201]},
      {stage2_11[111]}
   );
   gpc1_1 gpc3006 (
      {stage1_11[202]},
      {stage2_11[112]}
   );
   gpc1_1 gpc3007 (
      {stage1_11[203]},
      {stage2_11[113]}
   );
   gpc1_1 gpc3008 (
      {stage1_11[204]},
      {stage2_11[114]}
   );
   gpc1_1 gpc3009 (
      {stage1_11[205]},
      {stage2_11[115]}
   );
   gpc1_1 gpc3010 (
      {stage1_12[215]},
      {stage2_12[95]}
   );
   gpc1_1 gpc3011 (
      {stage1_12[216]},
      {stage2_12[96]}
   );
   gpc1_1 gpc3012 (
      {stage1_12[217]},
      {stage2_12[97]}
   );
   gpc1_1 gpc3013 (
      {stage1_12[218]},
      {stage2_12[98]}
   );
   gpc1_1 gpc3014 (
      {stage1_12[219]},
      {stage2_12[99]}
   );
   gpc1_1 gpc3015 (
      {stage1_12[220]},
      {stage2_12[100]}
   );
   gpc1_1 gpc3016 (
      {stage1_12[221]},
      {stage2_12[101]}
   );
   gpc1_1 gpc3017 (
      {stage1_13[198]},
      {stage2_13[90]}
   );
   gpc1_1 gpc3018 (
      {stage1_13[199]},
      {stage2_13[91]}
   );
   gpc1_1 gpc3019 (
      {stage1_13[200]},
      {stage2_13[92]}
   );
   gpc1_1 gpc3020 (
      {stage1_13[201]},
      {stage2_13[93]}
   );
   gpc1_1 gpc3021 (
      {stage1_13[202]},
      {stage2_13[94]}
   );
   gpc1_1 gpc3022 (
      {stage1_13[203]},
      {stage2_13[95]}
   );
   gpc1_1 gpc3023 (
      {stage1_13[204]},
      {stage2_13[96]}
   );
   gpc1_1 gpc3024 (
      {stage1_13[205]},
      {stage2_13[97]}
   );
   gpc1_1 gpc3025 (
      {stage1_13[206]},
      {stage2_13[98]}
   );
   gpc1_1 gpc3026 (
      {stage1_13[207]},
      {stage2_13[99]}
   );
   gpc1_1 gpc3027 (
      {stage1_13[208]},
      {stage2_13[100]}
   );
   gpc1_1 gpc3028 (
      {stage1_13[209]},
      {stage2_13[101]}
   );
   gpc1_1 gpc3029 (
      {stage1_13[210]},
      {stage2_13[102]}
   );
   gpc1_1 gpc3030 (
      {stage1_13[211]},
      {stage2_13[103]}
   );
   gpc1_1 gpc3031 (
      {stage1_13[212]},
      {stage2_13[104]}
   );
   gpc1_1 gpc3032 (
      {stage1_13[213]},
      {stage2_13[105]}
   );
   gpc1_1 gpc3033 (
      {stage1_13[214]},
      {stage2_13[106]}
   );
   gpc1_1 gpc3034 (
      {stage1_13[215]},
      {stage2_13[107]}
   );
   gpc1_1 gpc3035 (
      {stage1_13[216]},
      {stage2_13[108]}
   );
   gpc1_1 gpc3036 (
      {stage1_13[217]},
      {stage2_13[109]}
   );
   gpc1_1 gpc3037 (
      {stage1_13[218]},
      {stage2_13[110]}
   );
   gpc1_1 gpc3038 (
      {stage1_13[219]},
      {stage2_13[111]}
   );
   gpc1_1 gpc3039 (
      {stage1_13[220]},
      {stage2_13[112]}
   );
   gpc1_1 gpc3040 (
      {stage1_13[221]},
      {stage2_13[113]}
   );
   gpc1_1 gpc3041 (
      {stage1_13[222]},
      {stage2_13[114]}
   );
   gpc1_1 gpc3042 (
      {stage1_13[223]},
      {stage2_13[115]}
   );
   gpc1_1 gpc3043 (
      {stage1_13[224]},
      {stage2_13[116]}
   );
   gpc1_1 gpc3044 (
      {stage1_13[225]},
      {stage2_13[117]}
   );
   gpc1_1 gpc3045 (
      {stage1_13[226]},
      {stage2_13[118]}
   );
   gpc1_1 gpc3046 (
      {stage1_13[227]},
      {stage2_13[119]}
   );
   gpc1_1 gpc3047 (
      {stage1_13[228]},
      {stage2_13[120]}
   );
   gpc1_1 gpc3048 (
      {stage1_13[229]},
      {stage2_13[121]}
   );
   gpc1_1 gpc3049 (
      {stage1_13[230]},
      {stage2_13[122]}
   );
   gpc1_1 gpc3050 (
      {stage1_13[231]},
      {stage2_13[123]}
   );
   gpc1_1 gpc3051 (
      {stage1_15[222]},
      {stage2_15[83]}
   );
   gpc1_1 gpc3052 (
      {stage1_15[223]},
      {stage2_15[84]}
   );
   gpc1_1 gpc3053 (
      {stage1_15[224]},
      {stage2_15[85]}
   );
   gpc1_1 gpc3054 (
      {stage1_15[225]},
      {stage2_15[86]}
   );
   gpc1_1 gpc3055 (
      {stage1_15[226]},
      {stage2_15[87]}
   );
   gpc1_1 gpc3056 (
      {stage1_15[227]},
      {stage2_15[88]}
   );
   gpc1_1 gpc3057 (
      {stage1_15[228]},
      {stage2_15[89]}
   );
   gpc1_1 gpc3058 (
      {stage1_15[229]},
      {stage2_15[90]}
   );
   gpc1_1 gpc3059 (
      {stage1_15[230]},
      {stage2_15[91]}
   );
   gpc1_1 gpc3060 (
      {stage1_15[231]},
      {stage2_15[92]}
   );
   gpc1_1 gpc3061 (
      {stage1_15[232]},
      {stage2_15[93]}
   );
   gpc1_1 gpc3062 (
      {stage1_15[233]},
      {stage2_15[94]}
   );
   gpc1_1 gpc3063 (
      {stage1_15[234]},
      {stage2_15[95]}
   );
   gpc1_1 gpc3064 (
      {stage1_15[235]},
      {stage2_15[96]}
   );
   gpc1_1 gpc3065 (
      {stage1_15[236]},
      {stage2_15[97]}
   );
   gpc1_1 gpc3066 (
      {stage1_16[196]},
      {stage2_16[107]}
   );
   gpc1_1 gpc3067 (
      {stage1_16[197]},
      {stage2_16[108]}
   );
   gpc1_1 gpc3068 (
      {stage1_16[198]},
      {stage2_16[109]}
   );
   gpc1_1 gpc3069 (
      {stage1_16[199]},
      {stage2_16[110]}
   );
   gpc1_1 gpc3070 (
      {stage1_16[200]},
      {stage2_16[111]}
   );
   gpc1_1 gpc3071 (
      {stage1_16[201]},
      {stage2_16[112]}
   );
   gpc1_1 gpc3072 (
      {stage1_16[202]},
      {stage2_16[113]}
   );
   gpc1_1 gpc3073 (
      {stage1_16[203]},
      {stage2_16[114]}
   );
   gpc1_1 gpc3074 (
      {stage1_16[204]},
      {stage2_16[115]}
   );
   gpc1_1 gpc3075 (
      {stage1_16[205]},
      {stage2_16[116]}
   );
   gpc1_1 gpc3076 (
      {stage1_16[206]},
      {stage2_16[117]}
   );
   gpc1_1 gpc3077 (
      {stage1_16[207]},
      {stage2_16[118]}
   );
   gpc1_1 gpc3078 (
      {stage1_16[208]},
      {stage2_16[119]}
   );
   gpc1_1 gpc3079 (
      {stage1_16[209]},
      {stage2_16[120]}
   );
   gpc1_1 gpc3080 (
      {stage1_16[210]},
      {stage2_16[121]}
   );
   gpc1_1 gpc3081 (
      {stage1_16[211]},
      {stage2_16[122]}
   );
   gpc1_1 gpc3082 (
      {stage1_16[212]},
      {stage2_16[123]}
   );
   gpc1_1 gpc3083 (
      {stage1_16[213]},
      {stage2_16[124]}
   );
   gpc1_1 gpc3084 (
      {stage1_17[178]},
      {stage2_17[82]}
   );
   gpc1_1 gpc3085 (
      {stage1_17[179]},
      {stage2_17[83]}
   );
   gpc1_1 gpc3086 (
      {stage1_17[180]},
      {stage2_17[84]}
   );
   gpc1_1 gpc3087 (
      {stage1_17[181]},
      {stage2_17[85]}
   );
   gpc1_1 gpc3088 (
      {stage1_17[182]},
      {stage2_17[86]}
   );
   gpc1_1 gpc3089 (
      {stage1_17[183]},
      {stage2_17[87]}
   );
   gpc1_1 gpc3090 (
      {stage1_17[184]},
      {stage2_17[88]}
   );
   gpc1_1 gpc3091 (
      {stage1_17[185]},
      {stage2_17[89]}
   );
   gpc1_1 gpc3092 (
      {stage1_17[186]},
      {stage2_17[90]}
   );
   gpc1_1 gpc3093 (
      {stage1_17[187]},
      {stage2_17[91]}
   );
   gpc1_1 gpc3094 (
      {stage1_17[188]},
      {stage2_17[92]}
   );
   gpc1_1 gpc3095 (
      {stage1_17[189]},
      {stage2_17[93]}
   );
   gpc1_1 gpc3096 (
      {stage1_17[190]},
      {stage2_17[94]}
   );
   gpc1_1 gpc3097 (
      {stage1_17[191]},
      {stage2_17[95]}
   );
   gpc1_1 gpc3098 (
      {stage1_17[192]},
      {stage2_17[96]}
   );
   gpc1_1 gpc3099 (
      {stage1_17[193]},
      {stage2_17[97]}
   );
   gpc1_1 gpc3100 (
      {stage1_17[194]},
      {stage2_17[98]}
   );
   gpc1_1 gpc3101 (
      {stage1_17[195]},
      {stage2_17[99]}
   );
   gpc1_1 gpc3102 (
      {stage1_17[196]},
      {stage2_17[100]}
   );
   gpc1_1 gpc3103 (
      {stage1_17[197]},
      {stage2_17[101]}
   );
   gpc1_1 gpc3104 (
      {stage1_17[198]},
      {stage2_17[102]}
   );
   gpc1_1 gpc3105 (
      {stage1_17[199]},
      {stage2_17[103]}
   );
   gpc1_1 gpc3106 (
      {stage1_17[200]},
      {stage2_17[104]}
   );
   gpc1_1 gpc3107 (
      {stage1_17[201]},
      {stage2_17[105]}
   );
   gpc1_1 gpc3108 (
      {stage1_17[202]},
      {stage2_17[106]}
   );
   gpc1_1 gpc3109 (
      {stage1_17[203]},
      {stage2_17[107]}
   );
   gpc1_1 gpc3110 (
      {stage1_17[204]},
      {stage2_17[108]}
   );
   gpc1_1 gpc3111 (
      {stage1_17[205]},
      {stage2_17[109]}
   );
   gpc1_1 gpc3112 (
      {stage1_17[206]},
      {stage2_17[110]}
   );
   gpc1_1 gpc3113 (
      {stage1_17[207]},
      {stage2_17[111]}
   );
   gpc1_1 gpc3114 (
      {stage1_17[208]},
      {stage2_17[112]}
   );
   gpc1_1 gpc3115 (
      {stage1_17[209]},
      {stage2_17[113]}
   );
   gpc1_1 gpc3116 (
      {stage1_17[210]},
      {stage2_17[114]}
   );
   gpc1_1 gpc3117 (
      {stage1_17[211]},
      {stage2_17[115]}
   );
   gpc1_1 gpc3118 (
      {stage1_17[212]},
      {stage2_17[116]}
   );
   gpc1_1 gpc3119 (
      {stage1_17[213]},
      {stage2_17[117]}
   );
   gpc1_1 gpc3120 (
      {stage1_17[214]},
      {stage2_17[118]}
   );
   gpc1_1 gpc3121 (
      {stage1_17[215]},
      {stage2_17[119]}
   );
   gpc1_1 gpc3122 (
      {stage1_17[216]},
      {stage2_17[120]}
   );
   gpc1_1 gpc3123 (
      {stage1_17[217]},
      {stage2_17[121]}
   );
   gpc1_1 gpc3124 (
      {stage1_17[218]},
      {stage2_17[122]}
   );
   gpc1_1 gpc3125 (
      {stage1_17[219]},
      {stage2_17[123]}
   );
   gpc1_1 gpc3126 (
      {stage1_17[220]},
      {stage2_17[124]}
   );
   gpc1_1 gpc3127 (
      {stage1_17[221]},
      {stage2_17[125]}
   );
   gpc1_1 gpc3128 (
      {stage1_17[222]},
      {stage2_17[126]}
   );
   gpc1_1 gpc3129 (
      {stage1_17[223]},
      {stage2_17[127]}
   );
   gpc1_1 gpc3130 (
      {stage1_18[194]},
      {stage2_18[64]}
   );
   gpc1_1 gpc3131 (
      {stage1_18[195]},
      {stage2_18[65]}
   );
   gpc1_1 gpc3132 (
      {stage1_18[196]},
      {stage2_18[66]}
   );
   gpc1_1 gpc3133 (
      {stage1_18[197]},
      {stage2_18[67]}
   );
   gpc1_1 gpc3134 (
      {stage1_18[198]},
      {stage2_18[68]}
   );
   gpc1_1 gpc3135 (
      {stage1_18[199]},
      {stage2_18[69]}
   );
   gpc1_1 gpc3136 (
      {stage1_18[200]},
      {stage2_18[70]}
   );
   gpc1_1 gpc3137 (
      {stage1_18[201]},
      {stage2_18[71]}
   );
   gpc1_1 gpc3138 (
      {stage1_18[202]},
      {stage2_18[72]}
   );
   gpc1_1 gpc3139 (
      {stage1_19[261]},
      {stage2_19[96]}
   );
   gpc1_1 gpc3140 (
      {stage1_19[262]},
      {stage2_19[97]}
   );
   gpc1_1 gpc3141 (
      {stage1_20[211]},
      {stage2_20[107]}
   );
   gpc1_1 gpc3142 (
      {stage1_20[212]},
      {stage2_20[108]}
   );
   gpc1_1 gpc3143 (
      {stage1_20[213]},
      {stage2_20[109]}
   );
   gpc1_1 gpc3144 (
      {stage1_21[227]},
      {stage2_21[82]}
   );
   gpc1_1 gpc3145 (
      {stage1_21[228]},
      {stage2_21[83]}
   );
   gpc1_1 gpc3146 (
      {stage1_21[229]},
      {stage2_21[84]}
   );
   gpc1_1 gpc3147 (
      {stage1_21[230]},
      {stage2_21[85]}
   );
   gpc1_1 gpc3148 (
      {stage1_21[231]},
      {stage2_21[86]}
   );
   gpc1_1 gpc3149 (
      {stage1_21[232]},
      {stage2_21[87]}
   );
   gpc1_1 gpc3150 (
      {stage1_21[233]},
      {stage2_21[88]}
   );
   gpc1_1 gpc3151 (
      {stage1_21[234]},
      {stage2_21[89]}
   );
   gpc1_1 gpc3152 (
      {stage1_21[235]},
      {stage2_21[90]}
   );
   gpc1_1 gpc3153 (
      {stage1_21[236]},
      {stage2_21[91]}
   );
   gpc1_1 gpc3154 (
      {stage1_21[237]},
      {stage2_21[92]}
   );
   gpc1_1 gpc3155 (
      {stage1_21[238]},
      {stage2_21[93]}
   );
   gpc1_1 gpc3156 (
      {stage1_21[239]},
      {stage2_21[94]}
   );
   gpc1_1 gpc3157 (
      {stage1_21[240]},
      {stage2_21[95]}
   );
   gpc1_1 gpc3158 (
      {stage1_21[241]},
      {stage2_21[96]}
   );
   gpc1_1 gpc3159 (
      {stage1_21[242]},
      {stage2_21[97]}
   );
   gpc1_1 gpc3160 (
      {stage1_21[243]},
      {stage2_21[98]}
   );
   gpc1_1 gpc3161 (
      {stage1_21[244]},
      {stage2_21[99]}
   );
   gpc1_1 gpc3162 (
      {stage1_21[245]},
      {stage2_21[100]}
   );
   gpc1_1 gpc3163 (
      {stage1_21[246]},
      {stage2_21[101]}
   );
   gpc1_1 gpc3164 (
      {stage1_21[247]},
      {stage2_21[102]}
   );
   gpc1_1 gpc3165 (
      {stage1_21[248]},
      {stage2_21[103]}
   );
   gpc1_1 gpc3166 (
      {stage1_21[249]},
      {stage2_21[104]}
   );
   gpc1_1 gpc3167 (
      {stage1_21[250]},
      {stage2_21[105]}
   );
   gpc1_1 gpc3168 (
      {stage1_21[251]},
      {stage2_21[106]}
   );
   gpc1_1 gpc3169 (
      {stage1_21[252]},
      {stage2_21[107]}
   );
   gpc1_1 gpc3170 (
      {stage1_21[253]},
      {stage2_21[108]}
   );
   gpc1_1 gpc3171 (
      {stage1_21[254]},
      {stage2_21[109]}
   );
   gpc1_1 gpc3172 (
      {stage1_21[255]},
      {stage2_21[110]}
   );
   gpc1_1 gpc3173 (
      {stage1_21[256]},
      {stage2_21[111]}
   );
   gpc1_1 gpc3174 (
      {stage1_21[257]},
      {stage2_21[112]}
   );
   gpc1_1 gpc3175 (
      {stage1_21[258]},
      {stage2_21[113]}
   );
   gpc1_1 gpc3176 (
      {stage1_21[259]},
      {stage2_21[114]}
   );
   gpc1_1 gpc3177 (
      {stage1_21[260]},
      {stage2_21[115]}
   );
   gpc1_1 gpc3178 (
      {stage1_21[261]},
      {stage2_21[116]}
   );
   gpc1_1 gpc3179 (
      {stage1_21[262]},
      {stage2_21[117]}
   );
   gpc1_1 gpc3180 (
      {stage1_21[263]},
      {stage2_21[118]}
   );
   gpc1_1 gpc3181 (
      {stage1_21[264]},
      {stage2_21[119]}
   );
   gpc1_1 gpc3182 (
      {stage1_21[265]},
      {stage2_21[120]}
   );
   gpc1_1 gpc3183 (
      {stage1_21[266]},
      {stage2_21[121]}
   );
   gpc1_1 gpc3184 (
      {stage1_21[267]},
      {stage2_21[122]}
   );
   gpc1_1 gpc3185 (
      {stage1_21[268]},
      {stage2_21[123]}
   );
   gpc1_1 gpc3186 (
      {stage1_21[269]},
      {stage2_21[124]}
   );
   gpc1_1 gpc3187 (
      {stage1_22[268]},
      {stage2_22[89]}
   );
   gpc1_1 gpc3188 (
      {stage1_22[269]},
      {stage2_22[90]}
   );
   gpc1_1 gpc3189 (
      {stage1_22[270]},
      {stage2_22[91]}
   );
   gpc1_1 gpc3190 (
      {stage1_22[271]},
      {stage2_22[92]}
   );
   gpc1_1 gpc3191 (
      {stage1_22[272]},
      {stage2_22[93]}
   );
   gpc1_1 gpc3192 (
      {stage1_22[273]},
      {stage2_22[94]}
   );
   gpc1_1 gpc3193 (
      {stage1_23[146]},
      {stage2_23[103]}
   );
   gpc1_1 gpc3194 (
      {stage1_23[147]},
      {stage2_23[104]}
   );
   gpc1_1 gpc3195 (
      {stage1_23[148]},
      {stage2_23[105]}
   );
   gpc1_1 gpc3196 (
      {stage1_23[149]},
      {stage2_23[106]}
   );
   gpc1_1 gpc3197 (
      {stage1_23[150]},
      {stage2_23[107]}
   );
   gpc1_1 gpc3198 (
      {stage1_23[151]},
      {stage2_23[108]}
   );
   gpc1_1 gpc3199 (
      {stage1_23[152]},
      {stage2_23[109]}
   );
   gpc1_1 gpc3200 (
      {stage1_23[153]},
      {stage2_23[110]}
   );
   gpc1_1 gpc3201 (
      {stage1_23[154]},
      {stage2_23[111]}
   );
   gpc1_1 gpc3202 (
      {stage1_23[155]},
      {stage2_23[112]}
   );
   gpc1_1 gpc3203 (
      {stage1_23[156]},
      {stage2_23[113]}
   );
   gpc1_1 gpc3204 (
      {stage1_23[157]},
      {stage2_23[114]}
   );
   gpc1_1 gpc3205 (
      {stage1_23[158]},
      {stage2_23[115]}
   );
   gpc1_1 gpc3206 (
      {stage1_23[159]},
      {stage2_23[116]}
   );
   gpc1_1 gpc3207 (
      {stage1_23[160]},
      {stage2_23[117]}
   );
   gpc1_1 gpc3208 (
      {stage1_23[161]},
      {stage2_23[118]}
   );
   gpc1_1 gpc3209 (
      {stage1_23[162]},
      {stage2_23[119]}
   );
   gpc1_1 gpc3210 (
      {stage1_23[163]},
      {stage2_23[120]}
   );
   gpc1_1 gpc3211 (
      {stage1_23[164]},
      {stage2_23[121]}
   );
   gpc1_1 gpc3212 (
      {stage1_23[165]},
      {stage2_23[122]}
   );
   gpc1_1 gpc3213 (
      {stage1_24[217]},
      {stage2_24[86]}
   );
   gpc1_1 gpc3214 (
      {stage1_24[218]},
      {stage2_24[87]}
   );
   gpc1_1 gpc3215 (
      {stage1_24[219]},
      {stage2_24[88]}
   );
   gpc1_1 gpc3216 (
      {stage1_24[220]},
      {stage2_24[89]}
   );
   gpc1_1 gpc3217 (
      {stage1_25[255]},
      {stage2_25[84]}
   );
   gpc1_1 gpc3218 (
      {stage1_25[256]},
      {stage2_25[85]}
   );
   gpc1_1 gpc3219 (
      {stage1_25[257]},
      {stage2_25[86]}
   );
   gpc1_1 gpc3220 (
      {stage1_25[258]},
      {stage2_25[87]}
   );
   gpc1_1 gpc3221 (
      {stage1_25[259]},
      {stage2_25[88]}
   );
   gpc1_1 gpc3222 (
      {stage1_25[260]},
      {stage2_25[89]}
   );
   gpc1_1 gpc3223 (
      {stage1_25[261]},
      {stage2_25[90]}
   );
   gpc1_1 gpc3224 (
      {stage1_25[262]},
      {stage2_25[91]}
   );
   gpc1_1 gpc3225 (
      {stage1_25[263]},
      {stage2_25[92]}
   );
   gpc1_1 gpc3226 (
      {stage1_25[264]},
      {stage2_25[93]}
   );
   gpc1_1 gpc3227 (
      {stage1_25[265]},
      {stage2_25[94]}
   );
   gpc1_1 gpc3228 (
      {stage1_25[266]},
      {stage2_25[95]}
   );
   gpc1_1 gpc3229 (
      {stage1_25[267]},
      {stage2_25[96]}
   );
   gpc1_1 gpc3230 (
      {stage1_25[268]},
      {stage2_25[97]}
   );
   gpc1_1 gpc3231 (
      {stage1_25[269]},
      {stage2_25[98]}
   );
   gpc1_1 gpc3232 (
      {stage1_25[270]},
      {stage2_25[99]}
   );
   gpc1_1 gpc3233 (
      {stage1_25[271]},
      {stage2_25[100]}
   );
   gpc1_1 gpc3234 (
      {stage1_25[272]},
      {stage2_25[101]}
   );
   gpc1_1 gpc3235 (
      {stage1_25[273]},
      {stage2_25[102]}
   );
   gpc1_1 gpc3236 (
      {stage1_26[186]},
      {stage2_26[95]}
   );
   gpc1_1 gpc3237 (
      {stage1_26[187]},
      {stage2_26[96]}
   );
   gpc1_1 gpc3238 (
      {stage1_26[188]},
      {stage2_26[97]}
   );
   gpc1_1 gpc3239 (
      {stage1_26[189]},
      {stage2_26[98]}
   );
   gpc1_1 gpc3240 (
      {stage1_26[190]},
      {stage2_26[99]}
   );
   gpc1_1 gpc3241 (
      {stage1_27[196]},
      {stage2_27[81]}
   );
   gpc1_1 gpc3242 (
      {stage1_27[197]},
      {stage2_27[82]}
   );
   gpc1_1 gpc3243 (
      {stage1_27[198]},
      {stage2_27[83]}
   );
   gpc1_1 gpc3244 (
      {stage1_27[199]},
      {stage2_27[84]}
   );
   gpc1_1 gpc3245 (
      {stage1_28[149]},
      {stage2_28[72]}
   );
   gpc1_1 gpc3246 (
      {stage1_28[150]},
      {stage2_28[73]}
   );
   gpc1_1 gpc3247 (
      {stage1_28[151]},
      {stage2_28[74]}
   );
   gpc1_1 gpc3248 (
      {stage1_28[152]},
      {stage2_28[75]}
   );
   gpc1_1 gpc3249 (
      {stage1_28[153]},
      {stage2_28[76]}
   );
   gpc1_1 gpc3250 (
      {stage1_28[154]},
      {stage2_28[77]}
   );
   gpc1_1 gpc3251 (
      {stage1_28[155]},
      {stage2_28[78]}
   );
   gpc1_1 gpc3252 (
      {stage1_28[156]},
      {stage2_28[79]}
   );
   gpc1_1 gpc3253 (
      {stage1_28[157]},
      {stage2_28[80]}
   );
   gpc1_1 gpc3254 (
      {stage1_28[158]},
      {stage2_28[81]}
   );
   gpc1_1 gpc3255 (
      {stage1_28[159]},
      {stage2_28[82]}
   );
   gpc1_1 gpc3256 (
      {stage1_28[160]},
      {stage2_28[83]}
   );
   gpc1_1 gpc3257 (
      {stage1_28[161]},
      {stage2_28[84]}
   );
   gpc1_1 gpc3258 (
      {stage1_28[162]},
      {stage2_28[85]}
   );
   gpc1_1 gpc3259 (
      {stage1_28[163]},
      {stage2_28[86]}
   );
   gpc1_1 gpc3260 (
      {stage1_28[164]},
      {stage2_28[87]}
   );
   gpc1_1 gpc3261 (
      {stage1_28[165]},
      {stage2_28[88]}
   );
   gpc1_1 gpc3262 (
      {stage1_28[166]},
      {stage2_28[89]}
   );
   gpc1_1 gpc3263 (
      {stage1_28[167]},
      {stage2_28[90]}
   );
   gpc1_1 gpc3264 (
      {stage1_28[168]},
      {stage2_28[91]}
   );
   gpc1_1 gpc3265 (
      {stage1_28[169]},
      {stage2_28[92]}
   );
   gpc1_1 gpc3266 (
      {stage1_28[170]},
      {stage2_28[93]}
   );
   gpc1_1 gpc3267 (
      {stage1_28[171]},
      {stage2_28[94]}
   );
   gpc1_1 gpc3268 (
      {stage1_28[172]},
      {stage2_28[95]}
   );
   gpc1_1 gpc3269 (
      {stage1_28[173]},
      {stage2_28[96]}
   );
   gpc1_1 gpc3270 (
      {stage1_28[174]},
      {stage2_28[97]}
   );
   gpc1_1 gpc3271 (
      {stage1_28[175]},
      {stage2_28[98]}
   );
   gpc1_1 gpc3272 (
      {stage1_28[176]},
      {stage2_28[99]}
   );
   gpc1_1 gpc3273 (
      {stage1_28[177]},
      {stage2_28[100]}
   );
   gpc1_1 gpc3274 (
      {stage1_28[178]},
      {stage2_28[101]}
   );
   gpc1_1 gpc3275 (
      {stage1_28[179]},
      {stage2_28[102]}
   );
   gpc1_1 gpc3276 (
      {stage1_28[180]},
      {stage2_28[103]}
   );
   gpc1_1 gpc3277 (
      {stage1_28[181]},
      {stage2_28[104]}
   );
   gpc1_1 gpc3278 (
      {stage1_28[182]},
      {stage2_28[105]}
   );
   gpc1_1 gpc3279 (
      {stage1_28[183]},
      {stage2_28[106]}
   );
   gpc1_1 gpc3280 (
      {stage1_28[184]},
      {stage2_28[107]}
   );
   gpc1_1 gpc3281 (
      {stage1_28[185]},
      {stage2_28[108]}
   );
   gpc1_1 gpc3282 (
      {stage1_28[186]},
      {stage2_28[109]}
   );
   gpc1_1 gpc3283 (
      {stage1_28[187]},
      {stage2_28[110]}
   );
   gpc1_1 gpc3284 (
      {stage1_28[188]},
      {stage2_28[111]}
   );
   gpc1_1 gpc3285 (
      {stage1_28[189]},
      {stage2_28[112]}
   );
   gpc1_1 gpc3286 (
      {stage1_28[190]},
      {stage2_28[113]}
   );
   gpc1_1 gpc3287 (
      {stage1_28[191]},
      {stage2_28[114]}
   );
   gpc1_1 gpc3288 (
      {stage1_28[192]},
      {stage2_28[115]}
   );
   gpc1_1 gpc3289 (
      {stage1_28[193]},
      {stage2_28[116]}
   );
   gpc1_1 gpc3290 (
      {stage1_28[194]},
      {stage2_28[117]}
   );
   gpc1_1 gpc3291 (
      {stage1_28[195]},
      {stage2_28[118]}
   );
   gpc1_1 gpc3292 (
      {stage1_28[196]},
      {stage2_28[119]}
   );
   gpc1_1 gpc3293 (
      {stage1_28[197]},
      {stage2_28[120]}
   );
   gpc1_1 gpc3294 (
      {stage1_28[198]},
      {stage2_28[121]}
   );
   gpc1_1 gpc3295 (
      {stage1_28[199]},
      {stage2_28[122]}
   );
   gpc1_1 gpc3296 (
      {stage1_28[200]},
      {stage2_28[123]}
   );
   gpc1_1 gpc3297 (
      {stage1_28[201]},
      {stage2_28[124]}
   );
   gpc1_1 gpc3298 (
      {stage1_28[202]},
      {stage2_28[125]}
   );
   gpc1_1 gpc3299 (
      {stage1_28[203]},
      {stage2_28[126]}
   );
   gpc1_1 gpc3300 (
      {stage1_28[204]},
      {stage2_28[127]}
   );
   gpc1_1 gpc3301 (
      {stage1_28[205]},
      {stage2_28[128]}
   );
   gpc1_1 gpc3302 (
      {stage1_28[206]},
      {stage2_28[129]}
   );
   gpc1_1 gpc3303 (
      {stage1_28[207]},
      {stage2_28[130]}
   );
   gpc1_1 gpc3304 (
      {stage1_28[208]},
      {stage2_28[131]}
   );
   gpc1_1 gpc3305 (
      {stage1_28[209]},
      {stage2_28[132]}
   );
   gpc1_1 gpc3306 (
      {stage1_28[210]},
      {stage2_28[133]}
   );
   gpc1_1 gpc3307 (
      {stage1_28[211]},
      {stage2_28[134]}
   );
   gpc1_1 gpc3308 (
      {stage1_28[212]},
      {stage2_28[135]}
   );
   gpc1_1 gpc3309 (
      {stage1_28[213]},
      {stage2_28[136]}
   );
   gpc1_1 gpc3310 (
      {stage1_28[214]},
      {stage2_28[137]}
   );
   gpc1_1 gpc3311 (
      {stage1_28[215]},
      {stage2_28[138]}
   );
   gpc1_1 gpc3312 (
      {stage1_28[216]},
      {stage2_28[139]}
   );
   gpc1_1 gpc3313 (
      {stage1_28[217]},
      {stage2_28[140]}
   );
   gpc1_1 gpc3314 (
      {stage1_28[218]},
      {stage2_28[141]}
   );
   gpc1_1 gpc3315 (
      {stage1_28[219]},
      {stage2_28[142]}
   );
   gpc1_1 gpc3316 (
      {stage1_28[220]},
      {stage2_28[143]}
   );
   gpc1_1 gpc3317 (
      {stage1_28[221]},
      {stage2_28[144]}
   );
   gpc1_1 gpc3318 (
      {stage1_28[222]},
      {stage2_28[145]}
   );
   gpc1_1 gpc3319 (
      {stage1_28[223]},
      {stage2_28[146]}
   );
   gpc1_1 gpc3320 (
      {stage1_28[224]},
      {stage2_28[147]}
   );
   gpc1_1 gpc3321 (
      {stage1_28[225]},
      {stage2_28[148]}
   );
   gpc1_1 gpc3322 (
      {stage1_28[226]},
      {stage2_28[149]}
   );
   gpc1_1 gpc3323 (
      {stage1_28[227]},
      {stage2_28[150]}
   );
   gpc1_1 gpc3324 (
      {stage1_28[228]},
      {stage2_28[151]}
   );
   gpc1_1 gpc3325 (
      {stage1_28[229]},
      {stage2_28[152]}
   );
   gpc1_1 gpc3326 (
      {stage1_28[230]},
      {stage2_28[153]}
   );
   gpc1_1 gpc3327 (
      {stage1_28[231]},
      {stage2_28[154]}
   );
   gpc1_1 gpc3328 (
      {stage1_28[232]},
      {stage2_28[155]}
   );
   gpc1_1 gpc3329 (
      {stage1_28[233]},
      {stage2_28[156]}
   );
   gpc1_1 gpc3330 (
      {stage1_28[234]},
      {stage2_28[157]}
   );
   gpc1_1 gpc3331 (
      {stage1_28[235]},
      {stage2_28[158]}
   );
   gpc1_1 gpc3332 (
      {stage1_28[236]},
      {stage2_28[159]}
   );
   gpc1_1 gpc3333 (
      {stage1_28[237]},
      {stage2_28[160]}
   );
   gpc1_1 gpc3334 (
      {stage1_28[238]},
      {stage2_28[161]}
   );
   gpc1_1 gpc3335 (
      {stage1_28[239]},
      {stage2_28[162]}
   );
   gpc1_1 gpc3336 (
      {stage1_28[240]},
      {stage2_28[163]}
   );
   gpc1_1 gpc3337 (
      {stage1_28[241]},
      {stage2_28[164]}
   );
   gpc1_1 gpc3338 (
      {stage1_28[242]},
      {stage2_28[165]}
   );
   gpc1_1 gpc3339 (
      {stage1_28[243]},
      {stage2_28[166]}
   );
   gpc1_1 gpc3340 (
      {stage1_28[244]},
      {stage2_28[167]}
   );
   gpc1_1 gpc3341 (
      {stage1_28[245]},
      {stage2_28[168]}
   );
   gpc1_1 gpc3342 (
      {stage1_28[246]},
      {stage2_28[169]}
   );
   gpc1_1 gpc3343 (
      {stage1_28[247]},
      {stage2_28[170]}
   );
   gpc1_1 gpc3344 (
      {stage1_29[180]},
      {stage2_29[80]}
   );
   gpc1_1 gpc3345 (
      {stage1_29[181]},
      {stage2_29[81]}
   );
   gpc1_1 gpc3346 (
      {stage1_29[182]},
      {stage2_29[82]}
   );
   gpc1_1 gpc3347 (
      {stage1_29[183]},
      {stage2_29[83]}
   );
   gpc1_1 gpc3348 (
      {stage1_29[184]},
      {stage2_29[84]}
   );
   gpc1_1 gpc3349 (
      {stage1_29[185]},
      {stage2_29[85]}
   );
   gpc1_1 gpc3350 (
      {stage1_29[186]},
      {stage2_29[86]}
   );
   gpc1_1 gpc3351 (
      {stage1_29[187]},
      {stage2_29[87]}
   );
   gpc1_1 gpc3352 (
      {stage1_29[188]},
      {stage2_29[88]}
   );
   gpc1_1 gpc3353 (
      {stage1_29[189]},
      {stage2_29[89]}
   );
   gpc1_1 gpc3354 (
      {stage1_29[190]},
      {stage2_29[90]}
   );
   gpc1_1 gpc3355 (
      {stage1_29[191]},
      {stage2_29[91]}
   );
   gpc1_1 gpc3356 (
      {stage1_29[192]},
      {stage2_29[92]}
   );
   gpc1_1 gpc3357 (
      {stage1_29[193]},
      {stage2_29[93]}
   );
   gpc1_1 gpc3358 (
      {stage1_29[194]},
      {stage2_29[94]}
   );
   gpc1_1 gpc3359 (
      {stage1_29[195]},
      {stage2_29[95]}
   );
   gpc1_1 gpc3360 (
      {stage1_29[196]},
      {stage2_29[96]}
   );
   gpc1_1 gpc3361 (
      {stage1_29[197]},
      {stage2_29[97]}
   );
   gpc1_1 gpc3362 (
      {stage1_29[198]},
      {stage2_29[98]}
   );
   gpc1_1 gpc3363 (
      {stage1_29[199]},
      {stage2_29[99]}
   );
   gpc1_1 gpc3364 (
      {stage1_29[200]},
      {stage2_29[100]}
   );
   gpc1_1 gpc3365 (
      {stage1_29[201]},
      {stage2_29[101]}
   );
   gpc1_1 gpc3366 (
      {stage1_29[202]},
      {stage2_29[102]}
   );
   gpc1_1 gpc3367 (
      {stage1_29[203]},
      {stage2_29[103]}
   );
   gpc1_1 gpc3368 (
      {stage1_29[204]},
      {stage2_29[104]}
   );
   gpc1_1 gpc3369 (
      {stage1_29[205]},
      {stage2_29[105]}
   );
   gpc1_1 gpc3370 (
      {stage1_29[206]},
      {stage2_29[106]}
   );
   gpc1_1 gpc3371 (
      {stage1_29[207]},
      {stage2_29[107]}
   );
   gpc1_1 gpc3372 (
      {stage1_29[208]},
      {stage2_29[108]}
   );
   gpc1_1 gpc3373 (
      {stage1_29[209]},
      {stage2_29[109]}
   );
   gpc1_1 gpc3374 (
      {stage1_29[210]},
      {stage2_29[110]}
   );
   gpc1_1 gpc3375 (
      {stage1_29[211]},
      {stage2_29[111]}
   );
   gpc1_1 gpc3376 (
      {stage1_29[212]},
      {stage2_29[112]}
   );
   gpc1_1 gpc3377 (
      {stage1_29[213]},
      {stage2_29[113]}
   );
   gpc1_1 gpc3378 (
      {stage1_29[214]},
      {stage2_29[114]}
   );
   gpc1_1 gpc3379 (
      {stage1_29[215]},
      {stage2_29[115]}
   );
   gpc1_1 gpc3380 (
      {stage1_29[216]},
      {stage2_29[116]}
   );
   gpc1_1 gpc3381 (
      {stage1_29[217]},
      {stage2_29[117]}
   );
   gpc1_1 gpc3382 (
      {stage1_29[218]},
      {stage2_29[118]}
   );
   gpc1_1 gpc3383 (
      {stage1_29[219]},
      {stage2_29[119]}
   );
   gpc1_1 gpc3384 (
      {stage1_29[220]},
      {stage2_29[120]}
   );
   gpc1_1 gpc3385 (
      {stage1_29[221]},
      {stage2_29[121]}
   );
   gpc1_1 gpc3386 (
      {stage1_29[222]},
      {stage2_29[122]}
   );
   gpc1_1 gpc3387 (
      {stage1_29[223]},
      {stage2_29[123]}
   );
   gpc1_1 gpc3388 (
      {stage1_29[224]},
      {stage2_29[124]}
   );
   gpc1_1 gpc3389 (
      {stage1_29[225]},
      {stage2_29[125]}
   );
   gpc1_1 gpc3390 (
      {stage1_29[226]},
      {stage2_29[126]}
   );
   gpc1_1 gpc3391 (
      {stage1_29[227]},
      {stage2_29[127]}
   );
   gpc1_1 gpc3392 (
      {stage1_29[228]},
      {stage2_29[128]}
   );
   gpc1_1 gpc3393 (
      {stage1_29[229]},
      {stage2_29[129]}
   );
   gpc1_1 gpc3394 (
      {stage1_29[230]},
      {stage2_29[130]}
   );
   gpc1_1 gpc3395 (
      {stage1_29[231]},
      {stage2_29[131]}
   );
   gpc1_1 gpc3396 (
      {stage1_29[232]},
      {stage2_29[132]}
   );
   gpc1_1 gpc3397 (
      {stage1_29[233]},
      {stage2_29[133]}
   );
   gpc1_1 gpc3398 (
      {stage1_29[234]},
      {stage2_29[134]}
   );
   gpc1_1 gpc3399 (
      {stage1_29[235]},
      {stage2_29[135]}
   );
   gpc1_1 gpc3400 (
      {stage1_29[236]},
      {stage2_29[136]}
   );
   gpc1_1 gpc3401 (
      {stage1_29[237]},
      {stage2_29[137]}
   );
   gpc1_1 gpc3402 (
      {stage1_29[238]},
      {stage2_29[138]}
   );
   gpc1_1 gpc3403 (
      {stage1_29[239]},
      {stage2_29[139]}
   );
   gpc1_1 gpc3404 (
      {stage1_29[240]},
      {stage2_29[140]}
   );
   gpc1_1 gpc3405 (
      {stage1_29[241]},
      {stage2_29[141]}
   );
   gpc1_1 gpc3406 (
      {stage1_29[242]},
      {stage2_29[142]}
   );
   gpc1_1 gpc3407 (
      {stage1_30[192]},
      {stage2_30[77]}
   );
   gpc1_1 gpc3408 (
      {stage1_30[193]},
      {stage2_30[78]}
   );
   gpc1_1 gpc3409 (
      {stage1_30[194]},
      {stage2_30[79]}
   );
   gpc1_1 gpc3410 (
      {stage1_30[195]},
      {stage2_30[80]}
   );
   gpc1_1 gpc3411 (
      {stage1_30[196]},
      {stage2_30[81]}
   );
   gpc1_1 gpc3412 (
      {stage1_30[197]},
      {stage2_30[82]}
   );
   gpc1_1 gpc3413 (
      {stage1_30[198]},
      {stage2_30[83]}
   );
   gpc1_1 gpc3414 (
      {stage1_30[199]},
      {stage2_30[84]}
   );
   gpc1_1 gpc3415 (
      {stage1_30[200]},
      {stage2_30[85]}
   );
   gpc1_1 gpc3416 (
      {stage1_30[201]},
      {stage2_30[86]}
   );
   gpc1_1 gpc3417 (
      {stage1_30[202]},
      {stage2_30[87]}
   );
   gpc1_1 gpc3418 (
      {stage1_30[203]},
      {stage2_30[88]}
   );
   gpc1_1 gpc3419 (
      {stage1_30[204]},
      {stage2_30[89]}
   );
   gpc1_1 gpc3420 (
      {stage1_30[205]},
      {stage2_30[90]}
   );
   gpc1_1 gpc3421 (
      {stage1_30[206]},
      {stage2_30[91]}
   );
   gpc1_1 gpc3422 (
      {stage1_31[215]},
      {stage2_31[74]}
   );
   gpc1_1 gpc3423 (
      {stage1_31[216]},
      {stage2_31[75]}
   );
   gpc1_1 gpc3424 (
      {stage1_31[217]},
      {stage2_31[76]}
   );
   gpc1_1 gpc3425 (
      {stage1_31[218]},
      {stage2_31[77]}
   );
   gpc1_1 gpc3426 (
      {stage1_31[219]},
      {stage2_31[78]}
   );
   gpc1_1 gpc3427 (
      {stage1_31[220]},
      {stage2_31[79]}
   );
   gpc1_1 gpc3428 (
      {stage1_31[221]},
      {stage2_31[80]}
   );
   gpc1_1 gpc3429 (
      {stage1_31[222]},
      {stage2_31[81]}
   );
   gpc1_1 gpc3430 (
      {stage1_31[223]},
      {stage2_31[82]}
   );
   gpc1_1 gpc3431 (
      {stage1_31[224]},
      {stage2_31[83]}
   );
   gpc1_1 gpc3432 (
      {stage1_31[225]},
      {stage2_31[84]}
   );
   gpc1_1 gpc3433 (
      {stage1_31[226]},
      {stage2_31[85]}
   );
   gpc1_1 gpc3434 (
      {stage1_31[227]},
      {stage2_31[86]}
   );
   gpc1_1 gpc3435 (
      {stage1_31[228]},
      {stage2_31[87]}
   );
   gpc1_1 gpc3436 (
      {stage1_31[229]},
      {stage2_31[88]}
   );
   gpc1_1 gpc3437 (
      {stage1_31[230]},
      {stage2_31[89]}
   );
   gpc1_1 gpc3438 (
      {stage1_31[231]},
      {stage2_31[90]}
   );
   gpc1_1 gpc3439 (
      {stage1_31[232]},
      {stage2_31[91]}
   );
   gpc1_1 gpc3440 (
      {stage1_31[233]},
      {stage2_31[92]}
   );
   gpc1_1 gpc3441 (
      {stage1_31[234]},
      {stage2_31[93]}
   );
   gpc1_1 gpc3442 (
      {stage1_31[235]},
      {stage2_31[94]}
   );
   gpc1_1 gpc3443 (
      {stage1_31[236]},
      {stage2_31[95]}
   );
   gpc1_1 gpc3444 (
      {stage1_31[237]},
      {stage2_31[96]}
   );
   gpc1_1 gpc3445 (
      {stage1_31[238]},
      {stage2_31[97]}
   );
   gpc1_1 gpc3446 (
      {stage1_31[239]},
      {stage2_31[98]}
   );
   gpc1_1 gpc3447 (
      {stage1_31[240]},
      {stage2_31[99]}
   );
   gpc1_1 gpc3448 (
      {stage1_31[241]},
      {stage2_31[100]}
   );
   gpc1_1 gpc3449 (
      {stage1_31[242]},
      {stage2_31[101]}
   );
   gpc1_1 gpc3450 (
      {stage1_32[145]},
      {stage2_32[69]}
   );
   gpc1_1 gpc3451 (
      {stage1_32[146]},
      {stage2_32[70]}
   );
   gpc1_1 gpc3452 (
      {stage1_32[147]},
      {stage2_32[71]}
   );
   gpc1_1 gpc3453 (
      {stage1_32[148]},
      {stage2_32[72]}
   );
   gpc1_1 gpc3454 (
      {stage1_32[149]},
      {stage2_32[73]}
   );
   gpc1163_5 gpc3455 (
      {stage2_0[0], stage2_0[1], stage2_0[2]},
      {stage2_1[0], stage2_1[1], stage2_1[2], stage2_1[3], stage2_1[4], stage2_1[5]},
      {stage2_2[0]},
      {stage2_3[0]},
      {stage3_4[0],stage3_3[0],stage3_2[0],stage3_1[0],stage3_0[0]}
   );
   gpc606_5 gpc3456 (
      {stage2_0[3], stage2_0[4], stage2_0[5], stage2_0[6], stage2_0[7], stage2_0[8]},
      {stage2_2[1], stage2_2[2], stage2_2[3], stage2_2[4], stage2_2[5], stage2_2[6]},
      {stage3_4[1],stage3_3[1],stage3_2[1],stage3_1[1],stage3_0[1]}
   );
   gpc606_5 gpc3457 (
      {stage2_0[9], stage2_0[10], stage2_0[11], stage2_0[12], stage2_0[13], stage2_0[14]},
      {stage2_2[7], stage2_2[8], stage2_2[9], stage2_2[10], stage2_2[11], stage2_2[12]},
      {stage3_4[2],stage3_3[2],stage3_2[2],stage3_1[2],stage3_0[2]}
   );
   gpc606_5 gpc3458 (
      {stage2_0[15], stage2_0[16], stage2_0[17], stage2_0[18], stage2_0[19], stage2_0[20]},
      {stage2_2[13], stage2_2[14], stage2_2[15], stage2_2[16], stage2_2[17], stage2_2[18]},
      {stage3_4[3],stage3_3[3],stage3_2[3],stage3_1[3],stage3_0[3]}
   );
   gpc606_5 gpc3459 (
      {stage2_0[21], stage2_0[22], stage2_0[23], stage2_0[24], stage2_0[25], stage2_0[26]},
      {stage2_2[19], stage2_2[20], stage2_2[21], stage2_2[22], stage2_2[23], stage2_2[24]},
      {stage3_4[4],stage3_3[4],stage3_2[4],stage3_1[4],stage3_0[4]}
   );
   gpc606_5 gpc3460 (
      {stage2_0[27], stage2_0[28], stage2_0[29], stage2_0[30], stage2_0[31], stage2_0[32]},
      {stage2_2[25], stage2_2[26], stage2_2[27], stage2_2[28], stage2_2[29], stage2_2[30]},
      {stage3_4[5],stage3_3[5],stage3_2[5],stage3_1[5],stage3_0[5]}
   );
   gpc606_5 gpc3461 (
      {stage2_0[33], stage2_0[34], stage2_0[35], stage2_0[36], stage2_0[37], stage2_0[38]},
      {stage2_2[31], stage2_2[32], stage2_2[33], stage2_2[34], stage2_2[35], stage2_2[36]},
      {stage3_4[6],stage3_3[6],stage3_2[6],stage3_1[6],stage3_0[6]}
   );
   gpc606_5 gpc3462 (
      {stage2_0[39], stage2_0[40], stage2_0[41], stage2_0[42], stage2_0[43], stage2_0[44]},
      {stage2_2[37], stage2_2[38], stage2_2[39], stage2_2[40], stage2_2[41], stage2_2[42]},
      {stage3_4[7],stage3_3[7],stage3_2[7],stage3_1[7],stage3_0[7]}
   );
   gpc606_5 gpc3463 (
      {stage2_0[45], stage2_0[46], stage2_0[47], stage2_0[48], stage2_0[49], stage2_0[50]},
      {stage2_2[43], stage2_2[44], stage2_2[45], stage2_2[46], stage2_2[47], stage2_2[48]},
      {stage3_4[8],stage3_3[8],stage3_2[8],stage3_1[8],stage3_0[8]}
   );
   gpc606_5 gpc3464 (
      {stage2_0[51], stage2_0[52], stage2_0[53], stage2_0[54], stage2_0[55], stage2_0[56]},
      {stage2_2[49], stage2_2[50], stage2_2[51], stage2_2[52], stage2_2[53], stage2_2[54]},
      {stage3_4[9],stage3_3[9],stage3_2[9],stage3_1[9],stage3_0[9]}
   );
   gpc606_5 gpc3465 (
      {stage2_0[57], stage2_0[58], stage2_0[59], stage2_0[60], stage2_0[61], stage2_0[62]},
      {stage2_2[55], stage2_2[56], stage2_2[57], stage2_2[58], stage2_2[59], stage2_2[60]},
      {stage3_4[10],stage3_3[10],stage3_2[10],stage3_1[10],stage3_0[10]}
   );
   gpc606_5 gpc3466 (
      {stage2_1[6], stage2_1[7], stage2_1[8], stage2_1[9], stage2_1[10], stage2_1[11]},
      {stage2_3[1], stage2_3[2], stage2_3[3], stage2_3[4], stage2_3[5], stage2_3[6]},
      {stage3_5[0],stage3_4[11],stage3_3[11],stage3_2[11],stage3_1[11]}
   );
   gpc606_5 gpc3467 (
      {stage2_1[12], stage2_1[13], stage2_1[14], stage2_1[15], stage2_1[16], stage2_1[17]},
      {stage2_3[7], stage2_3[8], stage2_3[9], stage2_3[10], stage2_3[11], stage2_3[12]},
      {stage3_5[1],stage3_4[12],stage3_3[12],stage3_2[12],stage3_1[12]}
   );
   gpc606_5 gpc3468 (
      {stage2_1[18], stage2_1[19], stage2_1[20], stage2_1[21], stage2_1[22], stage2_1[23]},
      {stage2_3[13], stage2_3[14], stage2_3[15], stage2_3[16], stage2_3[17], stage2_3[18]},
      {stage3_5[2],stage3_4[13],stage3_3[13],stage3_2[13],stage3_1[13]}
   );
   gpc606_5 gpc3469 (
      {stage2_1[24], stage2_1[25], stage2_1[26], stage2_1[27], stage2_1[28], stage2_1[29]},
      {stage2_3[19], stage2_3[20], stage2_3[21], stage2_3[22], stage2_3[23], stage2_3[24]},
      {stage3_5[3],stage3_4[14],stage3_3[14],stage3_2[14],stage3_1[14]}
   );
   gpc606_5 gpc3470 (
      {stage2_1[30], stage2_1[31], stage2_1[32], stage2_1[33], stage2_1[34], stage2_1[35]},
      {stage2_3[25], stage2_3[26], stage2_3[27], stage2_3[28], stage2_3[29], stage2_3[30]},
      {stage3_5[4],stage3_4[15],stage3_3[15],stage3_2[15],stage3_1[15]}
   );
   gpc606_5 gpc3471 (
      {stage2_1[36], stage2_1[37], stage2_1[38], stage2_1[39], stage2_1[40], stage2_1[41]},
      {stage2_3[31], stage2_3[32], stage2_3[33], stage2_3[34], stage2_3[35], stage2_3[36]},
      {stage3_5[5],stage3_4[16],stage3_3[16],stage3_2[16],stage3_1[16]}
   );
   gpc606_5 gpc3472 (
      {stage2_1[42], stage2_1[43], stage2_1[44], stage2_1[45], stage2_1[46], stage2_1[47]},
      {stage2_3[37], stage2_3[38], stage2_3[39], stage2_3[40], stage2_3[41], stage2_3[42]},
      {stage3_5[6],stage3_4[17],stage3_3[17],stage3_2[17],stage3_1[17]}
   );
   gpc615_5 gpc3473 (
      {stage2_2[61], stage2_2[62], stage2_2[63], stage2_2[64], stage2_2[65]},
      {stage2_3[43]},
      {stage2_4[0], stage2_4[1], stage2_4[2], stage2_4[3], stage2_4[4], stage2_4[5]},
      {stage3_6[0],stage3_5[7],stage3_4[18],stage3_3[18],stage3_2[18]}
   );
   gpc615_5 gpc3474 (
      {stage2_2[66], stage2_2[67], stage2_2[68], stage2_2[69], stage2_2[70]},
      {stage2_3[44]},
      {stage2_4[6], stage2_4[7], stage2_4[8], stage2_4[9], stage2_4[10], stage2_4[11]},
      {stage3_6[1],stage3_5[8],stage3_4[19],stage3_3[19],stage3_2[19]}
   );
   gpc615_5 gpc3475 (
      {stage2_2[71], stage2_2[72], stage2_2[73], stage2_2[74], stage2_2[75]},
      {stage2_3[45]},
      {stage2_4[12], stage2_4[13], stage2_4[14], stage2_4[15], stage2_4[16], stage2_4[17]},
      {stage3_6[2],stage3_5[9],stage3_4[20],stage3_3[20],stage3_2[20]}
   );
   gpc615_5 gpc3476 (
      {stage2_2[76], stage2_2[77], stage2_2[78], stage2_2[79], stage2_2[80]},
      {stage2_3[46]},
      {stage2_4[18], stage2_4[19], stage2_4[20], stage2_4[21], stage2_4[22], stage2_4[23]},
      {stage3_6[3],stage3_5[10],stage3_4[21],stage3_3[21],stage3_2[21]}
   );
   gpc615_5 gpc3477 (
      {stage2_3[47], stage2_3[48], stage2_3[49], stage2_3[50], stage2_3[51]},
      {stage2_4[24]},
      {stage2_5[0], stage2_5[1], stage2_5[2], stage2_5[3], stage2_5[4], stage2_5[5]},
      {stage3_7[0],stage3_6[4],stage3_5[11],stage3_4[22],stage3_3[22]}
   );
   gpc615_5 gpc3478 (
      {stage2_3[52], stage2_3[53], stage2_3[54], stage2_3[55], stage2_3[56]},
      {stage2_4[25]},
      {stage2_5[6], stage2_5[7], stage2_5[8], stage2_5[9], stage2_5[10], stage2_5[11]},
      {stage3_7[1],stage3_6[5],stage3_5[12],stage3_4[23],stage3_3[23]}
   );
   gpc615_5 gpc3479 (
      {stage2_3[57], stage2_3[58], stage2_3[59], stage2_3[60], stage2_3[61]},
      {stage2_4[26]},
      {stage2_5[12], stage2_5[13], stage2_5[14], stage2_5[15], stage2_5[16], stage2_5[17]},
      {stage3_7[2],stage3_6[6],stage3_5[13],stage3_4[24],stage3_3[24]}
   );
   gpc615_5 gpc3480 (
      {stage2_3[62], stage2_3[63], stage2_3[64], stage2_3[65], stage2_3[66]},
      {stage2_4[27]},
      {stage2_5[18], stage2_5[19], stage2_5[20], stage2_5[21], stage2_5[22], stage2_5[23]},
      {stage3_7[3],stage3_6[7],stage3_5[14],stage3_4[25],stage3_3[25]}
   );
   gpc615_5 gpc3481 (
      {stage2_3[67], stage2_3[68], stage2_3[69], stage2_3[70], stage2_3[71]},
      {stage2_4[28]},
      {stage2_5[24], stage2_5[25], stage2_5[26], stage2_5[27], stage2_5[28], stage2_5[29]},
      {stage3_7[4],stage3_6[8],stage3_5[15],stage3_4[26],stage3_3[26]}
   );
   gpc615_5 gpc3482 (
      {stage2_3[72], stage2_3[73], stage2_3[74], stage2_3[75], stage2_3[76]},
      {stage2_4[29]},
      {stage2_5[30], stage2_5[31], stage2_5[32], stage2_5[33], stage2_5[34], stage2_5[35]},
      {stage3_7[5],stage3_6[9],stage3_5[16],stage3_4[27],stage3_3[27]}
   );
   gpc606_5 gpc3483 (
      {stage2_4[30], stage2_4[31], stage2_4[32], stage2_4[33], stage2_4[34], stage2_4[35]},
      {stage2_6[0], stage2_6[1], stage2_6[2], stage2_6[3], stage2_6[4], stage2_6[5]},
      {stage3_8[0],stage3_7[6],stage3_6[10],stage3_5[17],stage3_4[28]}
   );
   gpc606_5 gpc3484 (
      {stage2_4[36], stage2_4[37], stage2_4[38], stage2_4[39], stage2_4[40], stage2_4[41]},
      {stage2_6[6], stage2_6[7], stage2_6[8], stage2_6[9], stage2_6[10], stage2_6[11]},
      {stage3_8[1],stage3_7[7],stage3_6[11],stage3_5[18],stage3_4[29]}
   );
   gpc606_5 gpc3485 (
      {stage2_4[42], stage2_4[43], stage2_4[44], stage2_4[45], stage2_4[46], stage2_4[47]},
      {stage2_6[12], stage2_6[13], stage2_6[14], stage2_6[15], stage2_6[16], stage2_6[17]},
      {stage3_8[2],stage3_7[8],stage3_6[12],stage3_5[19],stage3_4[30]}
   );
   gpc606_5 gpc3486 (
      {stage2_4[48], stage2_4[49], stage2_4[50], stage2_4[51], stage2_4[52], stage2_4[53]},
      {stage2_6[18], stage2_6[19], stage2_6[20], stage2_6[21], stage2_6[22], stage2_6[23]},
      {stage3_8[3],stage3_7[9],stage3_6[13],stage3_5[20],stage3_4[31]}
   );
   gpc606_5 gpc3487 (
      {stage2_4[54], stage2_4[55], stage2_4[56], stage2_4[57], stage2_4[58], stage2_4[59]},
      {stage2_6[24], stage2_6[25], stage2_6[26], stage2_6[27], stage2_6[28], stage2_6[29]},
      {stage3_8[4],stage3_7[10],stage3_6[14],stage3_5[21],stage3_4[32]}
   );
   gpc606_5 gpc3488 (
      {stage2_4[60], stage2_4[61], stage2_4[62], stage2_4[63], stage2_4[64], stage2_4[65]},
      {stage2_6[30], stage2_6[31], stage2_6[32], stage2_6[33], stage2_6[34], stage2_6[35]},
      {stage3_8[5],stage3_7[11],stage3_6[15],stage3_5[22],stage3_4[33]}
   );
   gpc606_5 gpc3489 (
      {stage2_4[66], stage2_4[67], stage2_4[68], stage2_4[69], stage2_4[70], stage2_4[71]},
      {stage2_6[36], stage2_6[37], stage2_6[38], stage2_6[39], stage2_6[40], stage2_6[41]},
      {stage3_8[6],stage3_7[12],stage3_6[16],stage3_5[23],stage3_4[34]}
   );
   gpc606_5 gpc3490 (
      {stage2_4[72], stage2_4[73], stage2_4[74], stage2_4[75], stage2_4[76], stage2_4[77]},
      {stage2_6[42], stage2_6[43], stage2_6[44], stage2_6[45], stage2_6[46], stage2_6[47]},
      {stage3_8[7],stage3_7[13],stage3_6[17],stage3_5[24],stage3_4[35]}
   );
   gpc606_5 gpc3491 (
      {stage2_4[78], stage2_4[79], stage2_4[80], stage2_4[81], stage2_4[82], stage2_4[83]},
      {stage2_6[48], stage2_6[49], stage2_6[50], stage2_6[51], stage2_6[52], stage2_6[53]},
      {stage3_8[8],stage3_7[14],stage3_6[18],stage3_5[25],stage3_4[36]}
   );
   gpc606_5 gpc3492 (
      {stage2_4[84], stage2_4[85], stage2_4[86], stage2_4[87], stage2_4[88], stage2_4[89]},
      {stage2_6[54], stage2_6[55], stage2_6[56], stage2_6[57], stage2_6[58], stage2_6[59]},
      {stage3_8[9],stage3_7[15],stage3_6[19],stage3_5[26],stage3_4[37]}
   );
   gpc606_5 gpc3493 (
      {stage2_4[90], stage2_4[91], stage2_4[92], stage2_4[93], stage2_4[94], stage2_4[95]},
      {stage2_6[60], stage2_6[61], stage2_6[62], stage2_6[63], stage2_6[64], stage2_6[65]},
      {stage3_8[10],stage3_7[16],stage3_6[20],stage3_5[27],stage3_4[38]}
   );
   gpc606_5 gpc3494 (
      {stage2_4[96], stage2_4[97], stage2_4[98], stage2_4[99], stage2_4[100], stage2_4[101]},
      {stage2_6[66], stage2_6[67], stage2_6[68], stage2_6[69], stage2_6[70], stage2_6[71]},
      {stage3_8[11],stage3_7[17],stage3_6[21],stage3_5[28],stage3_4[39]}
   );
   gpc606_5 gpc3495 (
      {stage2_4[102], stage2_4[103], stage2_4[104], stage2_4[105], stage2_4[106], stage2_4[107]},
      {stage2_6[72], stage2_6[73], stage2_6[74], stage2_6[75], stage2_6[76], stage2_6[77]},
      {stage3_8[12],stage3_7[18],stage3_6[22],stage3_5[29],stage3_4[40]}
   );
   gpc606_5 gpc3496 (
      {stage2_4[108], stage2_4[109], stage2_4[110], stage2_4[111], stage2_4[112], stage2_4[113]},
      {stage2_6[78], stage2_6[79], stage2_6[80], stage2_6[81], stage2_6[82], stage2_6[83]},
      {stage3_8[13],stage3_7[19],stage3_6[23],stage3_5[30],stage3_4[41]}
   );
   gpc606_5 gpc3497 (
      {stage2_5[36], stage2_5[37], stage2_5[38], stage2_5[39], stage2_5[40], stage2_5[41]},
      {stage2_7[0], stage2_7[1], stage2_7[2], stage2_7[3], stage2_7[4], stage2_7[5]},
      {stage3_9[0],stage3_8[14],stage3_7[20],stage3_6[24],stage3_5[31]}
   );
   gpc606_5 gpc3498 (
      {stage2_5[42], stage2_5[43], stage2_5[44], stage2_5[45], stage2_5[46], stage2_5[47]},
      {stage2_7[6], stage2_7[7], stage2_7[8], stage2_7[9], stage2_7[10], stage2_7[11]},
      {stage3_9[1],stage3_8[15],stage3_7[21],stage3_6[25],stage3_5[32]}
   );
   gpc606_5 gpc3499 (
      {stage2_5[48], stage2_5[49], stage2_5[50], stage2_5[51], stage2_5[52], stage2_5[53]},
      {stage2_7[12], stage2_7[13], stage2_7[14], stage2_7[15], stage2_7[16], stage2_7[17]},
      {stage3_9[2],stage3_8[16],stage3_7[22],stage3_6[26],stage3_5[33]}
   );
   gpc606_5 gpc3500 (
      {stage2_5[54], stage2_5[55], stage2_5[56], stage2_5[57], stage2_5[58], stage2_5[59]},
      {stage2_7[18], stage2_7[19], stage2_7[20], stage2_7[21], stage2_7[22], stage2_7[23]},
      {stage3_9[3],stage3_8[17],stage3_7[23],stage3_6[27],stage3_5[34]}
   );
   gpc606_5 gpc3501 (
      {stage2_5[60], stage2_5[61], stage2_5[62], stage2_5[63], stage2_5[64], stage2_5[65]},
      {stage2_7[24], stage2_7[25], stage2_7[26], stage2_7[27], stage2_7[28], stage2_7[29]},
      {stage3_9[4],stage3_8[18],stage3_7[24],stage3_6[28],stage3_5[35]}
   );
   gpc606_5 gpc3502 (
      {stage2_5[66], stage2_5[67], stage2_5[68], stage2_5[69], stage2_5[70], stage2_5[71]},
      {stage2_7[30], stage2_7[31], stage2_7[32], stage2_7[33], stage2_7[34], stage2_7[35]},
      {stage3_9[5],stage3_8[19],stage3_7[25],stage3_6[29],stage3_5[36]}
   );
   gpc615_5 gpc3503 (
      {stage2_6[84], stage2_6[85], stage2_6[86], stage2_6[87], stage2_6[88]},
      {stage2_7[36]},
      {stage2_8[0], stage2_8[1], stage2_8[2], stage2_8[3], stage2_8[4], stage2_8[5]},
      {stage3_10[0],stage3_9[6],stage3_8[20],stage3_7[26],stage3_6[30]}
   );
   gpc615_5 gpc3504 (
      {stage2_7[37], stage2_7[38], stage2_7[39], stage2_7[40], stage2_7[41]},
      {stage2_8[6]},
      {stage2_9[0], stage2_9[1], stage2_9[2], stage2_9[3], stage2_9[4], stage2_9[5]},
      {stage3_11[0],stage3_10[1],stage3_9[7],stage3_8[21],stage3_7[27]}
   );
   gpc615_5 gpc3505 (
      {stage2_7[42], stage2_7[43], stage2_7[44], stage2_7[45], stage2_7[46]},
      {stage2_8[7]},
      {stage2_9[6], stage2_9[7], stage2_9[8], stage2_9[9], stage2_9[10], stage2_9[11]},
      {stage3_11[1],stage3_10[2],stage3_9[8],stage3_8[22],stage3_7[28]}
   );
   gpc615_5 gpc3506 (
      {stage2_7[47], stage2_7[48], stage2_7[49], stage2_7[50], stage2_7[51]},
      {stage2_8[8]},
      {stage2_9[12], stage2_9[13], stage2_9[14], stage2_9[15], stage2_9[16], stage2_9[17]},
      {stage3_11[2],stage3_10[3],stage3_9[9],stage3_8[23],stage3_7[29]}
   );
   gpc615_5 gpc3507 (
      {stage2_7[52], stage2_7[53], stage2_7[54], stage2_7[55], stage2_7[56]},
      {stage2_8[9]},
      {stage2_9[18], stage2_9[19], stage2_9[20], stage2_9[21], stage2_9[22], stage2_9[23]},
      {stage3_11[3],stage3_10[4],stage3_9[10],stage3_8[24],stage3_7[30]}
   );
   gpc615_5 gpc3508 (
      {stage2_7[57], stage2_7[58], stage2_7[59], stage2_7[60], stage2_7[61]},
      {stage2_8[10]},
      {stage2_9[24], stage2_9[25], stage2_9[26], stage2_9[27], stage2_9[28], stage2_9[29]},
      {stage3_11[4],stage3_10[5],stage3_9[11],stage3_8[25],stage3_7[31]}
   );
   gpc615_5 gpc3509 (
      {stage2_7[62], stage2_7[63], stage2_7[64], stage2_7[65], stage2_7[66]},
      {stage2_8[11]},
      {stage2_9[30], stage2_9[31], stage2_9[32], stage2_9[33], stage2_9[34], stage2_9[35]},
      {stage3_11[5],stage3_10[6],stage3_9[12],stage3_8[26],stage3_7[32]}
   );
   gpc615_5 gpc3510 (
      {stage2_7[67], stage2_7[68], stage2_7[69], stage2_7[70], stage2_7[71]},
      {stage2_8[12]},
      {stage2_9[36], stage2_9[37], stage2_9[38], stage2_9[39], stage2_9[40], stage2_9[41]},
      {stage3_11[6],stage3_10[7],stage3_9[13],stage3_8[27],stage3_7[33]}
   );
   gpc615_5 gpc3511 (
      {stage2_7[72], stage2_7[73], stage2_7[74], stage2_7[75], stage2_7[76]},
      {stage2_8[13]},
      {stage2_9[42], stage2_9[43], stage2_9[44], stage2_9[45], stage2_9[46], stage2_9[47]},
      {stage3_11[7],stage3_10[8],stage3_9[14],stage3_8[28],stage3_7[34]}
   );
   gpc615_5 gpc3512 (
      {stage2_7[77], stage2_7[78], stage2_7[79], stage2_7[80], stage2_7[81]},
      {stage2_8[14]},
      {stage2_9[48], stage2_9[49], stage2_9[50], stage2_9[51], stage2_9[52], stage2_9[53]},
      {stage3_11[8],stage3_10[9],stage3_9[15],stage3_8[29],stage3_7[35]}
   );
   gpc615_5 gpc3513 (
      {stage2_7[82], stage2_7[83], stage2_7[84], stage2_7[85], stage2_7[86]},
      {stage2_8[15]},
      {stage2_9[54], stage2_9[55], stage2_9[56], stage2_9[57], stage2_9[58], stage2_9[59]},
      {stage3_11[9],stage3_10[10],stage3_9[16],stage3_8[30],stage3_7[36]}
   );
   gpc615_5 gpc3514 (
      {stage2_7[87], stage2_7[88], stage2_7[89], stage2_7[90], stage2_7[91]},
      {stage2_8[16]},
      {stage2_9[60], stage2_9[61], stage2_9[62], stage2_9[63], stage2_9[64], stage2_9[65]},
      {stage3_11[10],stage3_10[11],stage3_9[17],stage3_8[31],stage3_7[37]}
   );
   gpc615_5 gpc3515 (
      {stage2_7[92], stage2_7[93], stage2_7[94], stage2_7[95], stage2_7[96]},
      {stage2_8[17]},
      {stage2_9[66], stage2_9[67], stage2_9[68], stage2_9[69], stage2_9[70], stage2_9[71]},
      {stage3_11[11],stage3_10[12],stage3_9[18],stage3_8[32],stage3_7[38]}
   );
   gpc615_5 gpc3516 (
      {stage2_7[97], stage2_7[98], stage2_7[99], stage2_7[100], stage2_7[101]},
      {stage2_8[18]},
      {stage2_9[72], stage2_9[73], stage2_9[74], stage2_9[75], stage2_9[76], stage2_9[77]},
      {stage3_11[12],stage3_10[13],stage3_9[19],stage3_8[33],stage3_7[39]}
   );
   gpc606_5 gpc3517 (
      {stage2_8[19], stage2_8[20], stage2_8[21], stage2_8[22], stage2_8[23], stage2_8[24]},
      {stage2_10[0], stage2_10[1], stage2_10[2], stage2_10[3], stage2_10[4], stage2_10[5]},
      {stage3_12[0],stage3_11[13],stage3_10[14],stage3_9[20],stage3_8[34]}
   );
   gpc606_5 gpc3518 (
      {stage2_8[25], stage2_8[26], stage2_8[27], stage2_8[28], stage2_8[29], stage2_8[30]},
      {stage2_10[6], stage2_10[7], stage2_10[8], stage2_10[9], stage2_10[10], stage2_10[11]},
      {stage3_12[1],stage3_11[14],stage3_10[15],stage3_9[21],stage3_8[35]}
   );
   gpc606_5 gpc3519 (
      {stage2_8[31], stage2_8[32], stage2_8[33], stage2_8[34], stage2_8[35], stage2_8[36]},
      {stage2_10[12], stage2_10[13], stage2_10[14], stage2_10[15], stage2_10[16], stage2_10[17]},
      {stage3_12[2],stage3_11[15],stage3_10[16],stage3_9[22],stage3_8[36]}
   );
   gpc606_5 gpc3520 (
      {stage2_8[37], stage2_8[38], stage2_8[39], stage2_8[40], stage2_8[41], stage2_8[42]},
      {stage2_10[18], stage2_10[19], stage2_10[20], stage2_10[21], stage2_10[22], stage2_10[23]},
      {stage3_12[3],stage3_11[16],stage3_10[17],stage3_9[23],stage3_8[37]}
   );
   gpc615_5 gpc3521 (
      {stage2_9[78], stage2_9[79], stage2_9[80], stage2_9[81], stage2_9[82]},
      {stage2_10[24]},
      {stage2_11[0], stage2_11[1], stage2_11[2], stage2_11[3], stage2_11[4], stage2_11[5]},
      {stage3_13[0],stage3_12[4],stage3_11[17],stage3_10[18],stage3_9[24]}
   );
   gpc606_5 gpc3522 (
      {stage2_10[25], stage2_10[26], stage2_10[27], stage2_10[28], stage2_10[29], stage2_10[30]},
      {stage2_12[0], stage2_12[1], stage2_12[2], stage2_12[3], stage2_12[4], stage2_12[5]},
      {stage3_14[0],stage3_13[1],stage3_12[5],stage3_11[18],stage3_10[19]}
   );
   gpc606_5 gpc3523 (
      {stage2_10[31], stage2_10[32], stage2_10[33], stage2_10[34], stage2_10[35], stage2_10[36]},
      {stage2_12[6], stage2_12[7], stage2_12[8], stage2_12[9], stage2_12[10], stage2_12[11]},
      {stage3_14[1],stage3_13[2],stage3_12[6],stage3_11[19],stage3_10[20]}
   );
   gpc606_5 gpc3524 (
      {stage2_10[37], stage2_10[38], stage2_10[39], stage2_10[40], stage2_10[41], stage2_10[42]},
      {stage2_12[12], stage2_12[13], stage2_12[14], stage2_12[15], stage2_12[16], stage2_12[17]},
      {stage3_14[2],stage3_13[3],stage3_12[7],stage3_11[20],stage3_10[21]}
   );
   gpc606_5 gpc3525 (
      {stage2_10[43], stage2_10[44], stage2_10[45], stage2_10[46], stage2_10[47], stage2_10[48]},
      {stage2_12[18], stage2_12[19], stage2_12[20], stage2_12[21], stage2_12[22], stage2_12[23]},
      {stage3_14[3],stage3_13[4],stage3_12[8],stage3_11[21],stage3_10[22]}
   );
   gpc606_5 gpc3526 (
      {stage2_10[49], stage2_10[50], stage2_10[51], stage2_10[52], stage2_10[53], stage2_10[54]},
      {stage2_12[24], stage2_12[25], stage2_12[26], stage2_12[27], stage2_12[28], stage2_12[29]},
      {stage3_14[4],stage3_13[5],stage3_12[9],stage3_11[22],stage3_10[23]}
   );
   gpc606_5 gpc3527 (
      {stage2_10[55], stage2_10[56], stage2_10[57], stage2_10[58], stage2_10[59], stage2_10[60]},
      {stage2_12[30], stage2_12[31], stage2_12[32], stage2_12[33], stage2_12[34], stage2_12[35]},
      {stage3_14[5],stage3_13[6],stage3_12[10],stage3_11[23],stage3_10[24]}
   );
   gpc606_5 gpc3528 (
      {stage2_10[61], stage2_10[62], stage2_10[63], stage2_10[64], stage2_10[65], stage2_10[66]},
      {stage2_12[36], stage2_12[37], stage2_12[38], stage2_12[39], stage2_12[40], stage2_12[41]},
      {stage3_14[6],stage3_13[7],stage3_12[11],stage3_11[24],stage3_10[25]}
   );
   gpc615_5 gpc3529 (
      {stage2_10[67], stage2_10[68], stage2_10[69], stage2_10[70], stage2_10[71]},
      {stage2_11[6]},
      {stage2_12[42], stage2_12[43], stage2_12[44], stage2_12[45], stage2_12[46], stage2_12[47]},
      {stage3_14[7],stage3_13[8],stage3_12[12],stage3_11[25],stage3_10[26]}
   );
   gpc615_5 gpc3530 (
      {stage2_10[72], stage2_10[73], stage2_10[74], stage2_10[75], stage2_10[76]},
      {stage2_11[7]},
      {stage2_12[48], stage2_12[49], stage2_12[50], stage2_12[51], stage2_12[52], stage2_12[53]},
      {stage3_14[8],stage3_13[9],stage3_12[13],stage3_11[26],stage3_10[27]}
   );
   gpc615_5 gpc3531 (
      {stage2_10[77], stage2_10[78], stage2_10[79], stage2_10[80], stage2_10[81]},
      {stage2_11[8]},
      {stage2_12[54], stage2_12[55], stage2_12[56], stage2_12[57], stage2_12[58], stage2_12[59]},
      {stage3_14[9],stage3_13[10],stage3_12[14],stage3_11[27],stage3_10[28]}
   );
   gpc615_5 gpc3532 (
      {stage2_10[82], stage2_10[83], stage2_10[84], stage2_10[85], stage2_10[86]},
      {stage2_11[9]},
      {stage2_12[60], stage2_12[61], stage2_12[62], stage2_12[63], stage2_12[64], stage2_12[65]},
      {stage3_14[10],stage3_13[11],stage3_12[15],stage3_11[28],stage3_10[29]}
   );
   gpc615_5 gpc3533 (
      {stage2_11[10], stage2_11[11], stage2_11[12], stage2_11[13], stage2_11[14]},
      {stage2_12[66]},
      {stage2_13[0], stage2_13[1], stage2_13[2], stage2_13[3], stage2_13[4], stage2_13[5]},
      {stage3_15[0],stage3_14[11],stage3_13[12],stage3_12[16],stage3_11[29]}
   );
   gpc615_5 gpc3534 (
      {stage2_11[15], stage2_11[16], stage2_11[17], stage2_11[18], stage2_11[19]},
      {stage2_12[67]},
      {stage2_13[6], stage2_13[7], stage2_13[8], stage2_13[9], stage2_13[10], stage2_13[11]},
      {stage3_15[1],stage3_14[12],stage3_13[13],stage3_12[17],stage3_11[30]}
   );
   gpc615_5 gpc3535 (
      {stage2_11[20], stage2_11[21], stage2_11[22], stage2_11[23], stage2_11[24]},
      {stage2_12[68]},
      {stage2_13[12], stage2_13[13], stage2_13[14], stage2_13[15], stage2_13[16], stage2_13[17]},
      {stage3_15[2],stage3_14[13],stage3_13[14],stage3_12[18],stage3_11[31]}
   );
   gpc615_5 gpc3536 (
      {stage2_11[25], stage2_11[26], stage2_11[27], stage2_11[28], stage2_11[29]},
      {stage2_12[69]},
      {stage2_13[18], stage2_13[19], stage2_13[20], stage2_13[21], stage2_13[22], stage2_13[23]},
      {stage3_15[3],stage3_14[14],stage3_13[15],stage3_12[19],stage3_11[32]}
   );
   gpc615_5 gpc3537 (
      {stage2_11[30], stage2_11[31], stage2_11[32], stage2_11[33], stage2_11[34]},
      {stage2_12[70]},
      {stage2_13[24], stage2_13[25], stage2_13[26], stage2_13[27], stage2_13[28], stage2_13[29]},
      {stage3_15[4],stage3_14[15],stage3_13[16],stage3_12[20],stage3_11[33]}
   );
   gpc615_5 gpc3538 (
      {stage2_11[35], stage2_11[36], stage2_11[37], stage2_11[38], stage2_11[39]},
      {stage2_12[71]},
      {stage2_13[30], stage2_13[31], stage2_13[32], stage2_13[33], stage2_13[34], stage2_13[35]},
      {stage3_15[5],stage3_14[16],stage3_13[17],stage3_12[21],stage3_11[34]}
   );
   gpc615_5 gpc3539 (
      {stage2_11[40], stage2_11[41], stage2_11[42], stage2_11[43], stage2_11[44]},
      {stage2_12[72]},
      {stage2_13[36], stage2_13[37], stage2_13[38], stage2_13[39], stage2_13[40], stage2_13[41]},
      {stage3_15[6],stage3_14[17],stage3_13[18],stage3_12[22],stage3_11[35]}
   );
   gpc615_5 gpc3540 (
      {stage2_11[45], stage2_11[46], stage2_11[47], stage2_11[48], stage2_11[49]},
      {stage2_12[73]},
      {stage2_13[42], stage2_13[43], stage2_13[44], stage2_13[45], stage2_13[46], stage2_13[47]},
      {stage3_15[7],stage3_14[18],stage3_13[19],stage3_12[23],stage3_11[36]}
   );
   gpc615_5 gpc3541 (
      {stage2_11[50], stage2_11[51], stage2_11[52], stage2_11[53], stage2_11[54]},
      {stage2_12[74]},
      {stage2_13[48], stage2_13[49], stage2_13[50], stage2_13[51], stage2_13[52], stage2_13[53]},
      {stage3_15[8],stage3_14[19],stage3_13[20],stage3_12[24],stage3_11[37]}
   );
   gpc615_5 gpc3542 (
      {stage2_11[55], stage2_11[56], stage2_11[57], stage2_11[58], stage2_11[59]},
      {stage2_12[75]},
      {stage2_13[54], stage2_13[55], stage2_13[56], stage2_13[57], stage2_13[58], stage2_13[59]},
      {stage3_15[9],stage3_14[20],stage3_13[21],stage3_12[25],stage3_11[38]}
   );
   gpc615_5 gpc3543 (
      {stage2_11[60], stage2_11[61], stage2_11[62], stage2_11[63], stage2_11[64]},
      {stage2_12[76]},
      {stage2_13[60], stage2_13[61], stage2_13[62], stage2_13[63], stage2_13[64], stage2_13[65]},
      {stage3_15[10],stage3_14[21],stage3_13[22],stage3_12[26],stage3_11[39]}
   );
   gpc615_5 gpc3544 (
      {stage2_11[65], stage2_11[66], stage2_11[67], stage2_11[68], stage2_11[69]},
      {stage2_12[77]},
      {stage2_13[66], stage2_13[67], stage2_13[68], stage2_13[69], stage2_13[70], stage2_13[71]},
      {stage3_15[11],stage3_14[22],stage3_13[23],stage3_12[27],stage3_11[40]}
   );
   gpc615_5 gpc3545 (
      {stage2_11[70], stage2_11[71], stage2_11[72], stage2_11[73], stage2_11[74]},
      {stage2_12[78]},
      {stage2_13[72], stage2_13[73], stage2_13[74], stage2_13[75], stage2_13[76], stage2_13[77]},
      {stage3_15[12],stage3_14[23],stage3_13[24],stage3_12[28],stage3_11[41]}
   );
   gpc615_5 gpc3546 (
      {stage2_11[75], stage2_11[76], stage2_11[77], stage2_11[78], stage2_11[79]},
      {stage2_12[79]},
      {stage2_13[78], stage2_13[79], stage2_13[80], stage2_13[81], stage2_13[82], stage2_13[83]},
      {stage3_15[13],stage3_14[24],stage3_13[25],stage3_12[29],stage3_11[42]}
   );
   gpc615_5 gpc3547 (
      {stage2_11[80], stage2_11[81], stage2_11[82], stage2_11[83], stage2_11[84]},
      {stage2_12[80]},
      {stage2_13[84], stage2_13[85], stage2_13[86], stage2_13[87], stage2_13[88], stage2_13[89]},
      {stage3_15[14],stage3_14[25],stage3_13[26],stage3_12[30],stage3_11[43]}
   );
   gpc615_5 gpc3548 (
      {stage2_11[85], stage2_11[86], stage2_11[87], stage2_11[88], stage2_11[89]},
      {stage2_12[81]},
      {stage2_13[90], stage2_13[91], stage2_13[92], stage2_13[93], stage2_13[94], stage2_13[95]},
      {stage3_15[15],stage3_14[26],stage3_13[27],stage3_12[31],stage3_11[44]}
   );
   gpc615_5 gpc3549 (
      {stage2_11[90], stage2_11[91], stage2_11[92], stage2_11[93], stage2_11[94]},
      {stage2_12[82]},
      {stage2_13[96], stage2_13[97], stage2_13[98], stage2_13[99], stage2_13[100], stage2_13[101]},
      {stage3_15[16],stage3_14[27],stage3_13[28],stage3_12[32],stage3_11[45]}
   );
   gpc615_5 gpc3550 (
      {stage2_11[95], stage2_11[96], stage2_11[97], stage2_11[98], stage2_11[99]},
      {stage2_12[83]},
      {stage2_13[102], stage2_13[103], stage2_13[104], stage2_13[105], stage2_13[106], stage2_13[107]},
      {stage3_15[17],stage3_14[28],stage3_13[29],stage3_12[33],stage3_11[46]}
   );
   gpc615_5 gpc3551 (
      {stage2_11[100], stage2_11[101], stage2_11[102], stage2_11[103], stage2_11[104]},
      {stage2_12[84]},
      {stage2_13[108], stage2_13[109], stage2_13[110], stage2_13[111], stage2_13[112], stage2_13[113]},
      {stage3_15[18],stage3_14[29],stage3_13[30],stage3_12[34],stage3_11[47]}
   );
   gpc615_5 gpc3552 (
      {stage2_11[105], stage2_11[106], stage2_11[107], stage2_11[108], stage2_11[109]},
      {stage2_12[85]},
      {stage2_13[114], stage2_13[115], stage2_13[116], stage2_13[117], stage2_13[118], stage2_13[119]},
      {stage3_15[19],stage3_14[30],stage3_13[31],stage3_12[35],stage3_11[48]}
   );
   gpc606_5 gpc3553 (
      {stage2_12[86], stage2_12[87], stage2_12[88], stage2_12[89], stage2_12[90], stage2_12[91]},
      {stage2_14[0], stage2_14[1], stage2_14[2], stage2_14[3], stage2_14[4], stage2_14[5]},
      {stage3_16[0],stage3_15[20],stage3_14[31],stage3_13[32],stage3_12[36]}
   );
   gpc615_5 gpc3554 (
      {stage2_14[6], stage2_14[7], stage2_14[8], stage2_14[9], stage2_14[10]},
      {stage2_15[0]},
      {stage2_16[0], stage2_16[1], stage2_16[2], stage2_16[3], stage2_16[4], stage2_16[5]},
      {stage3_18[0],stage3_17[0],stage3_16[1],stage3_15[21],stage3_14[32]}
   );
   gpc615_5 gpc3555 (
      {stage2_14[11], stage2_14[12], stage2_14[13], stage2_14[14], stage2_14[15]},
      {stage2_15[1]},
      {stage2_16[6], stage2_16[7], stage2_16[8], stage2_16[9], stage2_16[10], stage2_16[11]},
      {stage3_18[1],stage3_17[1],stage3_16[2],stage3_15[22],stage3_14[33]}
   );
   gpc615_5 gpc3556 (
      {stage2_14[16], stage2_14[17], stage2_14[18], stage2_14[19], stage2_14[20]},
      {stage2_15[2]},
      {stage2_16[12], stage2_16[13], stage2_16[14], stage2_16[15], stage2_16[16], stage2_16[17]},
      {stage3_18[2],stage3_17[2],stage3_16[3],stage3_15[23],stage3_14[34]}
   );
   gpc615_5 gpc3557 (
      {stage2_14[21], stage2_14[22], stage2_14[23], stage2_14[24], stage2_14[25]},
      {stage2_15[3]},
      {stage2_16[18], stage2_16[19], stage2_16[20], stage2_16[21], stage2_16[22], stage2_16[23]},
      {stage3_18[3],stage3_17[3],stage3_16[4],stage3_15[24],stage3_14[35]}
   );
   gpc615_5 gpc3558 (
      {stage2_14[26], stage2_14[27], stage2_14[28], stage2_14[29], stage2_14[30]},
      {stage2_15[4]},
      {stage2_16[24], stage2_16[25], stage2_16[26], stage2_16[27], stage2_16[28], stage2_16[29]},
      {stage3_18[4],stage3_17[4],stage3_16[5],stage3_15[25],stage3_14[36]}
   );
   gpc615_5 gpc3559 (
      {stage2_14[31], stage2_14[32], stage2_14[33], stage2_14[34], stage2_14[35]},
      {stage2_15[5]},
      {stage2_16[30], stage2_16[31], stage2_16[32], stage2_16[33], stage2_16[34], stage2_16[35]},
      {stage3_18[5],stage3_17[5],stage3_16[6],stage3_15[26],stage3_14[37]}
   );
   gpc615_5 gpc3560 (
      {stage2_14[36], stage2_14[37], stage2_14[38], stage2_14[39], stage2_14[40]},
      {stage2_15[6]},
      {stage2_16[36], stage2_16[37], stage2_16[38], stage2_16[39], stage2_16[40], stage2_16[41]},
      {stage3_18[6],stage3_17[6],stage3_16[7],stage3_15[27],stage3_14[38]}
   );
   gpc615_5 gpc3561 (
      {stage2_14[41], stage2_14[42], stage2_14[43], stage2_14[44], stage2_14[45]},
      {stage2_15[7]},
      {stage2_16[42], stage2_16[43], stage2_16[44], stage2_16[45], stage2_16[46], stage2_16[47]},
      {stage3_18[7],stage3_17[7],stage3_16[8],stage3_15[28],stage3_14[39]}
   );
   gpc615_5 gpc3562 (
      {stage2_14[46], stage2_14[47], stage2_14[48], stage2_14[49], stage2_14[50]},
      {stage2_15[8]},
      {stage2_16[48], stage2_16[49], stage2_16[50], stage2_16[51], stage2_16[52], stage2_16[53]},
      {stage3_18[8],stage3_17[8],stage3_16[9],stage3_15[29],stage3_14[40]}
   );
   gpc615_5 gpc3563 (
      {stage2_14[51], stage2_14[52], stage2_14[53], stage2_14[54], stage2_14[55]},
      {stage2_15[9]},
      {stage2_16[54], stage2_16[55], stage2_16[56], stage2_16[57], stage2_16[58], stage2_16[59]},
      {stage3_18[9],stage3_17[9],stage3_16[10],stage3_15[30],stage3_14[41]}
   );
   gpc615_5 gpc3564 (
      {stage2_15[10], stage2_15[11], stage2_15[12], stage2_15[13], stage2_15[14]},
      {stage2_16[60]},
      {stage2_17[0], stage2_17[1], stage2_17[2], stage2_17[3], stage2_17[4], stage2_17[5]},
      {stage3_19[0],stage3_18[10],stage3_17[10],stage3_16[11],stage3_15[31]}
   );
   gpc615_5 gpc3565 (
      {stage2_15[15], stage2_15[16], stage2_15[17], stage2_15[18], stage2_15[19]},
      {stage2_16[61]},
      {stage2_17[6], stage2_17[7], stage2_17[8], stage2_17[9], stage2_17[10], stage2_17[11]},
      {stage3_19[1],stage3_18[11],stage3_17[11],stage3_16[12],stage3_15[32]}
   );
   gpc615_5 gpc3566 (
      {stage2_15[20], stage2_15[21], stage2_15[22], stage2_15[23], stage2_15[24]},
      {stage2_16[62]},
      {stage2_17[12], stage2_17[13], stage2_17[14], stage2_17[15], stage2_17[16], stage2_17[17]},
      {stage3_19[2],stage3_18[12],stage3_17[12],stage3_16[13],stage3_15[33]}
   );
   gpc615_5 gpc3567 (
      {stage2_15[25], stage2_15[26], stage2_15[27], stage2_15[28], stage2_15[29]},
      {stage2_16[63]},
      {stage2_17[18], stage2_17[19], stage2_17[20], stage2_17[21], stage2_17[22], stage2_17[23]},
      {stage3_19[3],stage3_18[13],stage3_17[13],stage3_16[14],stage3_15[34]}
   );
   gpc615_5 gpc3568 (
      {stage2_15[30], stage2_15[31], stage2_15[32], stage2_15[33], stage2_15[34]},
      {stage2_16[64]},
      {stage2_17[24], stage2_17[25], stage2_17[26], stage2_17[27], stage2_17[28], stage2_17[29]},
      {stage3_19[4],stage3_18[14],stage3_17[14],stage3_16[15],stage3_15[35]}
   );
   gpc615_5 gpc3569 (
      {stage2_15[35], stage2_15[36], stage2_15[37], stage2_15[38], stage2_15[39]},
      {stage2_16[65]},
      {stage2_17[30], stage2_17[31], stage2_17[32], stage2_17[33], stage2_17[34], stage2_17[35]},
      {stage3_19[5],stage3_18[15],stage3_17[15],stage3_16[16],stage3_15[36]}
   );
   gpc615_5 gpc3570 (
      {stage2_15[40], stage2_15[41], stage2_15[42], stage2_15[43], stage2_15[44]},
      {stage2_16[66]},
      {stage2_17[36], stage2_17[37], stage2_17[38], stage2_17[39], stage2_17[40], stage2_17[41]},
      {stage3_19[6],stage3_18[16],stage3_17[16],stage3_16[17],stage3_15[37]}
   );
   gpc615_5 gpc3571 (
      {stage2_15[45], stage2_15[46], stage2_15[47], stage2_15[48], stage2_15[49]},
      {stage2_16[67]},
      {stage2_17[42], stage2_17[43], stage2_17[44], stage2_17[45], stage2_17[46], stage2_17[47]},
      {stage3_19[7],stage3_18[17],stage3_17[17],stage3_16[18],stage3_15[38]}
   );
   gpc615_5 gpc3572 (
      {stage2_15[50], stage2_15[51], stage2_15[52], stage2_15[53], stage2_15[54]},
      {stage2_16[68]},
      {stage2_17[48], stage2_17[49], stage2_17[50], stage2_17[51], stage2_17[52], stage2_17[53]},
      {stage3_19[8],stage3_18[18],stage3_17[18],stage3_16[19],stage3_15[39]}
   );
   gpc615_5 gpc3573 (
      {stage2_15[55], stage2_15[56], stage2_15[57], stage2_15[58], stage2_15[59]},
      {stage2_16[69]},
      {stage2_17[54], stage2_17[55], stage2_17[56], stage2_17[57], stage2_17[58], stage2_17[59]},
      {stage3_19[9],stage3_18[19],stage3_17[19],stage3_16[20],stage3_15[40]}
   );
   gpc615_5 gpc3574 (
      {stage2_15[60], stage2_15[61], stage2_15[62], stage2_15[63], stage2_15[64]},
      {stage2_16[70]},
      {stage2_17[60], stage2_17[61], stage2_17[62], stage2_17[63], stage2_17[64], stage2_17[65]},
      {stage3_19[10],stage3_18[20],stage3_17[20],stage3_16[21],stage3_15[41]}
   );
   gpc615_5 gpc3575 (
      {stage2_15[65], stage2_15[66], stage2_15[67], stage2_15[68], stage2_15[69]},
      {stage2_16[71]},
      {stage2_17[66], stage2_17[67], stage2_17[68], stage2_17[69], stage2_17[70], stage2_17[71]},
      {stage3_19[11],stage3_18[21],stage3_17[21],stage3_16[22],stage3_15[42]}
   );
   gpc135_4 gpc3576 (
      {stage2_16[72], stage2_16[73], stage2_16[74], stage2_16[75], stage2_16[76]},
      {stage2_17[72], stage2_17[73], stage2_17[74]},
      {stage2_18[0]},
      {stage3_19[12],stage3_18[22],stage3_17[22],stage3_16[23]}
   );
   gpc606_5 gpc3577 (
      {stage2_16[77], stage2_16[78], stage2_16[79], stage2_16[80], stage2_16[81], stage2_16[82]},
      {stage2_18[1], stage2_18[2], stage2_18[3], stage2_18[4], stage2_18[5], stage2_18[6]},
      {stage3_20[0],stage3_19[13],stage3_18[23],stage3_17[23],stage3_16[24]}
   );
   gpc606_5 gpc3578 (
      {stage2_18[7], stage2_18[8], stage2_18[9], stage2_18[10], stage2_18[11], stage2_18[12]},
      {stage2_20[0], stage2_20[1], stage2_20[2], stage2_20[3], stage2_20[4], stage2_20[5]},
      {stage3_22[0],stage3_21[0],stage3_20[1],stage3_19[14],stage3_18[24]}
   );
   gpc606_5 gpc3579 (
      {stage2_18[13], stage2_18[14], stage2_18[15], stage2_18[16], stage2_18[17], stage2_18[18]},
      {stage2_20[6], stage2_20[7], stage2_20[8], stage2_20[9], stage2_20[10], stage2_20[11]},
      {stage3_22[1],stage3_21[1],stage3_20[2],stage3_19[15],stage3_18[25]}
   );
   gpc606_5 gpc3580 (
      {stage2_18[19], stage2_18[20], stage2_18[21], stage2_18[22], stage2_18[23], stage2_18[24]},
      {stage2_20[12], stage2_20[13], stage2_20[14], stage2_20[15], stage2_20[16], stage2_20[17]},
      {stage3_22[2],stage3_21[2],stage3_20[3],stage3_19[16],stage3_18[26]}
   );
   gpc606_5 gpc3581 (
      {stage2_18[25], stage2_18[26], stage2_18[27], stage2_18[28], stage2_18[29], stage2_18[30]},
      {stage2_20[18], stage2_20[19], stage2_20[20], stage2_20[21], stage2_20[22], stage2_20[23]},
      {stage3_22[3],stage3_21[3],stage3_20[4],stage3_19[17],stage3_18[27]}
   );
   gpc606_5 gpc3582 (
      {stage2_18[31], stage2_18[32], stage2_18[33], stage2_18[34], stage2_18[35], stage2_18[36]},
      {stage2_20[24], stage2_20[25], stage2_20[26], stage2_20[27], stage2_20[28], stage2_20[29]},
      {stage3_22[4],stage3_21[4],stage3_20[5],stage3_19[18],stage3_18[28]}
   );
   gpc606_5 gpc3583 (
      {stage2_18[37], stage2_18[38], stage2_18[39], stage2_18[40], stage2_18[41], stage2_18[42]},
      {stage2_20[30], stage2_20[31], stage2_20[32], stage2_20[33], stage2_20[34], stage2_20[35]},
      {stage3_22[5],stage3_21[5],stage3_20[6],stage3_19[19],stage3_18[29]}
   );
   gpc606_5 gpc3584 (
      {stage2_18[43], stage2_18[44], stage2_18[45], stage2_18[46], stage2_18[47], stage2_18[48]},
      {stage2_20[36], stage2_20[37], stage2_20[38], stage2_20[39], stage2_20[40], stage2_20[41]},
      {stage3_22[6],stage3_21[6],stage3_20[7],stage3_19[20],stage3_18[30]}
   );
   gpc606_5 gpc3585 (
      {stage2_18[49], stage2_18[50], stage2_18[51], stage2_18[52], stage2_18[53], stage2_18[54]},
      {stage2_20[42], stage2_20[43], stage2_20[44], stage2_20[45], stage2_20[46], stage2_20[47]},
      {stage3_22[7],stage3_21[7],stage3_20[8],stage3_19[21],stage3_18[31]}
   );
   gpc606_5 gpc3586 (
      {stage2_18[55], stage2_18[56], stage2_18[57], stage2_18[58], stage2_18[59], stage2_18[60]},
      {stage2_20[48], stage2_20[49], stage2_20[50], stage2_20[51], stage2_20[52], stage2_20[53]},
      {stage3_22[8],stage3_21[8],stage3_20[9],stage3_19[22],stage3_18[32]}
   );
   gpc606_5 gpc3587 (
      {stage2_18[61], stage2_18[62], stage2_18[63], stage2_18[64], stage2_18[65], stage2_18[66]},
      {stage2_20[54], stage2_20[55], stage2_20[56], stage2_20[57], stage2_20[58], stage2_20[59]},
      {stage3_22[9],stage3_21[9],stage3_20[10],stage3_19[23],stage3_18[33]}
   );
   gpc606_5 gpc3588 (
      {stage2_18[67], stage2_18[68], stage2_18[69], stage2_18[70], stage2_18[71], stage2_18[72]},
      {stage2_20[60], stage2_20[61], stage2_20[62], stage2_20[63], stage2_20[64], stage2_20[65]},
      {stage3_22[10],stage3_21[10],stage3_20[11],stage3_19[24],stage3_18[34]}
   );
   gpc606_5 gpc3589 (
      {stage2_19[0], stage2_19[1], stage2_19[2], stage2_19[3], stage2_19[4], stage2_19[5]},
      {stage2_21[0], stage2_21[1], stage2_21[2], stage2_21[3], stage2_21[4], stage2_21[5]},
      {stage3_23[0],stage3_22[11],stage3_21[11],stage3_20[12],stage3_19[25]}
   );
   gpc606_5 gpc3590 (
      {stage2_19[6], stage2_19[7], stage2_19[8], stage2_19[9], stage2_19[10], stage2_19[11]},
      {stage2_21[6], stage2_21[7], stage2_21[8], stage2_21[9], stage2_21[10], stage2_21[11]},
      {stage3_23[1],stage3_22[12],stage3_21[12],stage3_20[13],stage3_19[26]}
   );
   gpc606_5 gpc3591 (
      {stage2_19[12], stage2_19[13], stage2_19[14], stage2_19[15], stage2_19[16], stage2_19[17]},
      {stage2_21[12], stage2_21[13], stage2_21[14], stage2_21[15], stage2_21[16], stage2_21[17]},
      {stage3_23[2],stage3_22[13],stage3_21[13],stage3_20[14],stage3_19[27]}
   );
   gpc606_5 gpc3592 (
      {stage2_19[18], stage2_19[19], stage2_19[20], stage2_19[21], stage2_19[22], stage2_19[23]},
      {stage2_21[18], stage2_21[19], stage2_21[20], stage2_21[21], stage2_21[22], stage2_21[23]},
      {stage3_23[3],stage3_22[14],stage3_21[14],stage3_20[15],stage3_19[28]}
   );
   gpc606_5 gpc3593 (
      {stage2_19[24], stage2_19[25], stage2_19[26], stage2_19[27], stage2_19[28], stage2_19[29]},
      {stage2_21[24], stage2_21[25], stage2_21[26], stage2_21[27], stage2_21[28], stage2_21[29]},
      {stage3_23[4],stage3_22[15],stage3_21[15],stage3_20[16],stage3_19[29]}
   );
   gpc606_5 gpc3594 (
      {stage2_19[30], stage2_19[31], stage2_19[32], stage2_19[33], stage2_19[34], stage2_19[35]},
      {stage2_21[30], stage2_21[31], stage2_21[32], stage2_21[33], stage2_21[34], stage2_21[35]},
      {stage3_23[5],stage3_22[16],stage3_21[16],stage3_20[17],stage3_19[30]}
   );
   gpc606_5 gpc3595 (
      {stage2_19[36], stage2_19[37], stage2_19[38], stage2_19[39], stage2_19[40], stage2_19[41]},
      {stage2_21[36], stage2_21[37], stage2_21[38], stage2_21[39], stage2_21[40], stage2_21[41]},
      {stage3_23[6],stage3_22[17],stage3_21[17],stage3_20[18],stage3_19[31]}
   );
   gpc606_5 gpc3596 (
      {stage2_19[42], stage2_19[43], stage2_19[44], stage2_19[45], stage2_19[46], stage2_19[47]},
      {stage2_21[42], stage2_21[43], stage2_21[44], stage2_21[45], stage2_21[46], stage2_21[47]},
      {stage3_23[7],stage3_22[18],stage3_21[18],stage3_20[19],stage3_19[32]}
   );
   gpc606_5 gpc3597 (
      {stage2_19[48], stage2_19[49], stage2_19[50], stage2_19[51], stage2_19[52], stage2_19[53]},
      {stage2_21[48], stage2_21[49], stage2_21[50], stage2_21[51], stage2_21[52], stage2_21[53]},
      {stage3_23[8],stage3_22[19],stage3_21[19],stage3_20[20],stage3_19[33]}
   );
   gpc615_5 gpc3598 (
      {stage2_19[54], stage2_19[55], stage2_19[56], stage2_19[57], stage2_19[58]},
      {stage2_20[66]},
      {stage2_21[54], stage2_21[55], stage2_21[56], stage2_21[57], stage2_21[58], stage2_21[59]},
      {stage3_23[9],stage3_22[20],stage3_21[20],stage3_20[21],stage3_19[34]}
   );
   gpc615_5 gpc3599 (
      {stage2_19[59], stage2_19[60], stage2_19[61], stage2_19[62], stage2_19[63]},
      {stage2_20[67]},
      {stage2_21[60], stage2_21[61], stage2_21[62], stage2_21[63], stage2_21[64], stage2_21[65]},
      {stage3_23[10],stage3_22[21],stage3_21[21],stage3_20[22],stage3_19[35]}
   );
   gpc606_5 gpc3600 (
      {stage2_20[68], stage2_20[69], stage2_20[70], stage2_20[71], stage2_20[72], stage2_20[73]},
      {stage2_22[0], stage2_22[1], stage2_22[2], stage2_22[3], stage2_22[4], stage2_22[5]},
      {stage3_24[0],stage3_23[11],stage3_22[22],stage3_21[22],stage3_20[23]}
   );
   gpc606_5 gpc3601 (
      {stage2_20[74], stage2_20[75], stage2_20[76], stage2_20[77], stage2_20[78], stage2_20[79]},
      {stage2_22[6], stage2_22[7], stage2_22[8], stage2_22[9], stage2_22[10], stage2_22[11]},
      {stage3_24[1],stage3_23[12],stage3_22[23],stage3_21[23],stage3_20[24]}
   );
   gpc606_5 gpc3602 (
      {stage2_20[80], stage2_20[81], stage2_20[82], stage2_20[83], stage2_20[84], stage2_20[85]},
      {stage2_22[12], stage2_22[13], stage2_22[14], stage2_22[15], stage2_22[16], stage2_22[17]},
      {stage3_24[2],stage3_23[13],stage3_22[24],stage3_21[24],stage3_20[25]}
   );
   gpc606_5 gpc3603 (
      {stage2_20[86], stage2_20[87], stage2_20[88], stage2_20[89], stage2_20[90], stage2_20[91]},
      {stage2_22[18], stage2_22[19], stage2_22[20], stage2_22[21], stage2_22[22], stage2_22[23]},
      {stage3_24[3],stage3_23[14],stage3_22[25],stage3_21[25],stage3_20[26]}
   );
   gpc606_5 gpc3604 (
      {stage2_20[92], stage2_20[93], stage2_20[94], stage2_20[95], stage2_20[96], stage2_20[97]},
      {stage2_22[24], stage2_22[25], stage2_22[26], stage2_22[27], stage2_22[28], stage2_22[29]},
      {stage3_24[4],stage3_23[15],stage3_22[26],stage3_21[26],stage3_20[27]}
   );
   gpc606_5 gpc3605 (
      {stage2_20[98], stage2_20[99], stage2_20[100], stage2_20[101], stage2_20[102], stage2_20[103]},
      {stage2_22[30], stage2_22[31], stage2_22[32], stage2_22[33], stage2_22[34], stage2_22[35]},
      {stage3_24[5],stage3_23[16],stage3_22[27],stage3_21[27],stage3_20[28]}
   );
   gpc606_5 gpc3606 (
      {stage2_20[104], stage2_20[105], stage2_20[106], stage2_20[107], stage2_20[108], stage2_20[109]},
      {stage2_22[36], stage2_22[37], stage2_22[38], stage2_22[39], stage2_22[40], stage2_22[41]},
      {stage3_24[6],stage3_23[17],stage3_22[28],stage3_21[28],stage3_20[29]}
   );
   gpc606_5 gpc3607 (
      {stage2_21[66], stage2_21[67], stage2_21[68], stage2_21[69], stage2_21[70], stage2_21[71]},
      {stage2_23[0], stage2_23[1], stage2_23[2], stage2_23[3], stage2_23[4], stage2_23[5]},
      {stage3_25[0],stage3_24[7],stage3_23[18],stage3_22[29],stage3_21[29]}
   );
   gpc606_5 gpc3608 (
      {stage2_21[72], stage2_21[73], stage2_21[74], stage2_21[75], stage2_21[76], stage2_21[77]},
      {stage2_23[6], stage2_23[7], stage2_23[8], stage2_23[9], stage2_23[10], stage2_23[11]},
      {stage3_25[1],stage3_24[8],stage3_23[19],stage3_22[30],stage3_21[30]}
   );
   gpc606_5 gpc3609 (
      {stage2_21[78], stage2_21[79], stage2_21[80], stage2_21[81], stage2_21[82], stage2_21[83]},
      {stage2_23[12], stage2_23[13], stage2_23[14], stage2_23[15], stage2_23[16], stage2_23[17]},
      {stage3_25[2],stage3_24[9],stage3_23[20],stage3_22[31],stage3_21[31]}
   );
   gpc606_5 gpc3610 (
      {stage2_21[84], stage2_21[85], stage2_21[86], stage2_21[87], stage2_21[88], stage2_21[89]},
      {stage2_23[18], stage2_23[19], stage2_23[20], stage2_23[21], stage2_23[22], stage2_23[23]},
      {stage3_25[3],stage3_24[10],stage3_23[21],stage3_22[32],stage3_21[32]}
   );
   gpc606_5 gpc3611 (
      {stage2_21[90], stage2_21[91], stage2_21[92], stage2_21[93], stage2_21[94], stage2_21[95]},
      {stage2_23[24], stage2_23[25], stage2_23[26], stage2_23[27], stage2_23[28], stage2_23[29]},
      {stage3_25[4],stage3_24[11],stage3_23[22],stage3_22[33],stage3_21[33]}
   );
   gpc615_5 gpc3612 (
      {stage2_22[42], stage2_22[43], stage2_22[44], stage2_22[45], stage2_22[46]},
      {stage2_23[30]},
      {stage2_24[0], stage2_24[1], stage2_24[2], stage2_24[3], stage2_24[4], stage2_24[5]},
      {stage3_26[0],stage3_25[5],stage3_24[12],stage3_23[23],stage3_22[34]}
   );
   gpc615_5 gpc3613 (
      {stage2_22[47], stage2_22[48], stage2_22[49], stage2_22[50], stage2_22[51]},
      {stage2_23[31]},
      {stage2_24[6], stage2_24[7], stage2_24[8], stage2_24[9], stage2_24[10], stage2_24[11]},
      {stage3_26[1],stage3_25[6],stage3_24[13],stage3_23[24],stage3_22[35]}
   );
   gpc615_5 gpc3614 (
      {stage2_22[52], stage2_22[53], stage2_22[54], stage2_22[55], stage2_22[56]},
      {stage2_23[32]},
      {stage2_24[12], stage2_24[13], stage2_24[14], stage2_24[15], stage2_24[16], stage2_24[17]},
      {stage3_26[2],stage3_25[7],stage3_24[14],stage3_23[25],stage3_22[36]}
   );
   gpc615_5 gpc3615 (
      {stage2_22[57], stage2_22[58], stage2_22[59], stage2_22[60], stage2_22[61]},
      {stage2_23[33]},
      {stage2_24[18], stage2_24[19], stage2_24[20], stage2_24[21], stage2_24[22], stage2_24[23]},
      {stage3_26[3],stage3_25[8],stage3_24[15],stage3_23[26],stage3_22[37]}
   );
   gpc615_5 gpc3616 (
      {stage2_22[62], stage2_22[63], stage2_22[64], stage2_22[65], stage2_22[66]},
      {stage2_23[34]},
      {stage2_24[24], stage2_24[25], stage2_24[26], stage2_24[27], stage2_24[28], stage2_24[29]},
      {stage3_26[4],stage3_25[9],stage3_24[16],stage3_23[27],stage3_22[38]}
   );
   gpc615_5 gpc3617 (
      {stage2_22[67], stage2_22[68], stage2_22[69], stage2_22[70], stage2_22[71]},
      {stage2_23[35]},
      {stage2_24[30], stage2_24[31], stage2_24[32], stage2_24[33], stage2_24[34], stage2_24[35]},
      {stage3_26[5],stage3_25[10],stage3_24[17],stage3_23[28],stage3_22[39]}
   );
   gpc615_5 gpc3618 (
      {stage2_22[72], stage2_22[73], stage2_22[74], stage2_22[75], stage2_22[76]},
      {stage2_23[36]},
      {stage2_24[36], stage2_24[37], stage2_24[38], stage2_24[39], stage2_24[40], stage2_24[41]},
      {stage3_26[6],stage3_25[11],stage3_24[18],stage3_23[29],stage3_22[40]}
   );
   gpc615_5 gpc3619 (
      {stage2_22[77], stage2_22[78], stage2_22[79], stage2_22[80], stage2_22[81]},
      {stage2_23[37]},
      {stage2_24[42], stage2_24[43], stage2_24[44], stage2_24[45], stage2_24[46], stage2_24[47]},
      {stage3_26[7],stage3_25[12],stage3_24[19],stage3_23[30],stage3_22[41]}
   );
   gpc615_5 gpc3620 (
      {stage2_22[82], stage2_22[83], stage2_22[84], stage2_22[85], stage2_22[86]},
      {stage2_23[38]},
      {stage2_24[48], stage2_24[49], stage2_24[50], stage2_24[51], stage2_24[52], stage2_24[53]},
      {stage3_26[8],stage3_25[13],stage3_24[20],stage3_23[31],stage3_22[42]}
   );
   gpc606_5 gpc3621 (
      {stage2_23[39], stage2_23[40], stage2_23[41], stage2_23[42], stage2_23[43], stage2_23[44]},
      {stage2_25[0], stage2_25[1], stage2_25[2], stage2_25[3], stage2_25[4], stage2_25[5]},
      {stage3_27[0],stage3_26[9],stage3_25[14],stage3_24[21],stage3_23[32]}
   );
   gpc606_5 gpc3622 (
      {stage2_23[45], stage2_23[46], stage2_23[47], stage2_23[48], stage2_23[49], stage2_23[50]},
      {stage2_25[6], stage2_25[7], stage2_25[8], stage2_25[9], stage2_25[10], stage2_25[11]},
      {stage3_27[1],stage3_26[10],stage3_25[15],stage3_24[22],stage3_23[33]}
   );
   gpc606_5 gpc3623 (
      {stage2_23[51], stage2_23[52], stage2_23[53], stage2_23[54], stage2_23[55], stage2_23[56]},
      {stage2_25[12], stage2_25[13], stage2_25[14], stage2_25[15], stage2_25[16], stage2_25[17]},
      {stage3_27[2],stage3_26[11],stage3_25[16],stage3_24[23],stage3_23[34]}
   );
   gpc606_5 gpc3624 (
      {stage2_23[57], stage2_23[58], stage2_23[59], stage2_23[60], stage2_23[61], stage2_23[62]},
      {stage2_25[18], stage2_25[19], stage2_25[20], stage2_25[21], stage2_25[22], stage2_25[23]},
      {stage3_27[3],stage3_26[12],stage3_25[17],stage3_24[24],stage3_23[35]}
   );
   gpc606_5 gpc3625 (
      {stage2_23[63], stage2_23[64], stage2_23[65], stage2_23[66], stage2_23[67], stage2_23[68]},
      {stage2_25[24], stage2_25[25], stage2_25[26], stage2_25[27], stage2_25[28], stage2_25[29]},
      {stage3_27[4],stage3_26[13],stage3_25[18],stage3_24[25],stage3_23[36]}
   );
   gpc606_5 gpc3626 (
      {stage2_23[69], stage2_23[70], stage2_23[71], stage2_23[72], stage2_23[73], stage2_23[74]},
      {stage2_25[30], stage2_25[31], stage2_25[32], stage2_25[33], stage2_25[34], stage2_25[35]},
      {stage3_27[5],stage3_26[14],stage3_25[19],stage3_24[26],stage3_23[37]}
   );
   gpc606_5 gpc3627 (
      {stage2_23[75], stage2_23[76], stage2_23[77], stage2_23[78], stage2_23[79], stage2_23[80]},
      {stage2_25[36], stage2_25[37], stage2_25[38], stage2_25[39], stage2_25[40], stage2_25[41]},
      {stage3_27[6],stage3_26[15],stage3_25[20],stage3_24[27],stage3_23[38]}
   );
   gpc606_5 gpc3628 (
      {stage2_23[81], stage2_23[82], stage2_23[83], stage2_23[84], stage2_23[85], stage2_23[86]},
      {stage2_25[42], stage2_25[43], stage2_25[44], stage2_25[45], stage2_25[46], stage2_25[47]},
      {stage3_27[7],stage3_26[16],stage3_25[21],stage3_24[28],stage3_23[39]}
   );
   gpc606_5 gpc3629 (
      {stage2_23[87], stage2_23[88], stage2_23[89], stage2_23[90], stage2_23[91], stage2_23[92]},
      {stage2_25[48], stage2_25[49], stage2_25[50], stage2_25[51], stage2_25[52], stage2_25[53]},
      {stage3_27[8],stage3_26[17],stage3_25[22],stage3_24[29],stage3_23[40]}
   );
   gpc606_5 gpc3630 (
      {stage2_23[93], stage2_23[94], stage2_23[95], stage2_23[96], stage2_23[97], stage2_23[98]},
      {stage2_25[54], stage2_25[55], stage2_25[56], stage2_25[57], stage2_25[58], stage2_25[59]},
      {stage3_27[9],stage3_26[18],stage3_25[23],stage3_24[30],stage3_23[41]}
   );
   gpc606_5 gpc3631 (
      {stage2_23[99], stage2_23[100], stage2_23[101], stage2_23[102], stage2_23[103], stage2_23[104]},
      {stage2_25[60], stage2_25[61], stage2_25[62], stage2_25[63], stage2_25[64], stage2_25[65]},
      {stage3_27[10],stage3_26[19],stage3_25[24],stage3_24[31],stage3_23[42]}
   );
   gpc606_5 gpc3632 (
      {stage2_23[105], stage2_23[106], stage2_23[107], stage2_23[108], stage2_23[109], stage2_23[110]},
      {stage2_25[66], stage2_25[67], stage2_25[68], stage2_25[69], stage2_25[70], stage2_25[71]},
      {stage3_27[11],stage3_26[20],stage3_25[25],stage3_24[32],stage3_23[43]}
   );
   gpc606_5 gpc3633 (
      {stage2_23[111], stage2_23[112], stage2_23[113], stage2_23[114], stage2_23[115], stage2_23[116]},
      {stage2_25[72], stage2_25[73], stage2_25[74], stage2_25[75], stage2_25[76], stage2_25[77]},
      {stage3_27[12],stage3_26[21],stage3_25[26],stage3_24[33],stage3_23[44]}
   );
   gpc606_5 gpc3634 (
      {stage2_23[117], stage2_23[118], stage2_23[119], stage2_23[120], stage2_23[121], stage2_23[122]},
      {stage2_25[78], stage2_25[79], stage2_25[80], stage2_25[81], stage2_25[82], stage2_25[83]},
      {stage3_27[13],stage3_26[22],stage3_25[27],stage3_24[34],stage3_23[45]}
   );
   gpc606_5 gpc3635 (
      {stage2_24[54], stage2_24[55], stage2_24[56], stage2_24[57], stage2_24[58], stage2_24[59]},
      {stage2_26[0], stage2_26[1], stage2_26[2], stage2_26[3], stage2_26[4], stage2_26[5]},
      {stage3_28[0],stage3_27[14],stage3_26[23],stage3_25[28],stage3_24[35]}
   );
   gpc606_5 gpc3636 (
      {stage2_24[60], stage2_24[61], stage2_24[62], stage2_24[63], stage2_24[64], stage2_24[65]},
      {stage2_26[6], stage2_26[7], stage2_26[8], stage2_26[9], stage2_26[10], stage2_26[11]},
      {stage3_28[1],stage3_27[15],stage3_26[24],stage3_25[29],stage3_24[36]}
   );
   gpc1163_5 gpc3637 (
      {stage2_26[12], stage2_26[13], stage2_26[14]},
      {stage2_27[0], stage2_27[1], stage2_27[2], stage2_27[3], stage2_27[4], stage2_27[5]},
      {stage2_28[0]},
      {stage2_29[0]},
      {stage3_30[0],stage3_29[0],stage3_28[2],stage3_27[16],stage3_26[25]}
   );
   gpc606_5 gpc3638 (
      {stage2_26[15], stage2_26[16], stage2_26[17], stage2_26[18], stage2_26[19], stage2_26[20]},
      {stage2_28[1], stage2_28[2], stage2_28[3], stage2_28[4], stage2_28[5], stage2_28[6]},
      {stage3_30[1],stage3_29[1],stage3_28[3],stage3_27[17],stage3_26[26]}
   );
   gpc606_5 gpc3639 (
      {stage2_26[21], stage2_26[22], stage2_26[23], stage2_26[24], stage2_26[25], stage2_26[26]},
      {stage2_28[7], stage2_28[8], stage2_28[9], stage2_28[10], stage2_28[11], stage2_28[12]},
      {stage3_30[2],stage3_29[2],stage3_28[4],stage3_27[18],stage3_26[27]}
   );
   gpc606_5 gpc3640 (
      {stage2_26[27], stage2_26[28], stage2_26[29], stage2_26[30], stage2_26[31], stage2_26[32]},
      {stage2_28[13], stage2_28[14], stage2_28[15], stage2_28[16], stage2_28[17], stage2_28[18]},
      {stage3_30[3],stage3_29[3],stage3_28[5],stage3_27[19],stage3_26[28]}
   );
   gpc606_5 gpc3641 (
      {stage2_26[33], stage2_26[34], stage2_26[35], stage2_26[36], stage2_26[37], stage2_26[38]},
      {stage2_28[19], stage2_28[20], stage2_28[21], stage2_28[22], stage2_28[23], stage2_28[24]},
      {stage3_30[4],stage3_29[4],stage3_28[6],stage3_27[20],stage3_26[29]}
   );
   gpc606_5 gpc3642 (
      {stage2_26[39], stage2_26[40], stage2_26[41], stage2_26[42], stage2_26[43], stage2_26[44]},
      {stage2_28[25], stage2_28[26], stage2_28[27], stage2_28[28], stage2_28[29], stage2_28[30]},
      {stage3_30[5],stage3_29[5],stage3_28[7],stage3_27[21],stage3_26[30]}
   );
   gpc606_5 gpc3643 (
      {stage2_26[45], stage2_26[46], stage2_26[47], stage2_26[48], stage2_26[49], stage2_26[50]},
      {stage2_28[31], stage2_28[32], stage2_28[33], stage2_28[34], stage2_28[35], stage2_28[36]},
      {stage3_30[6],stage3_29[6],stage3_28[8],stage3_27[22],stage3_26[31]}
   );
   gpc606_5 gpc3644 (
      {stage2_26[51], stage2_26[52], stage2_26[53], stage2_26[54], stage2_26[55], stage2_26[56]},
      {stage2_28[37], stage2_28[38], stage2_28[39], stage2_28[40], stage2_28[41], stage2_28[42]},
      {stage3_30[7],stage3_29[7],stage3_28[9],stage3_27[23],stage3_26[32]}
   );
   gpc606_5 gpc3645 (
      {stage2_26[57], stage2_26[58], stage2_26[59], stage2_26[60], stage2_26[61], stage2_26[62]},
      {stage2_28[43], stage2_28[44], stage2_28[45], stage2_28[46], stage2_28[47], stage2_28[48]},
      {stage3_30[8],stage3_29[8],stage3_28[10],stage3_27[24],stage3_26[33]}
   );
   gpc606_5 gpc3646 (
      {stage2_26[63], stage2_26[64], stage2_26[65], stage2_26[66], stage2_26[67], stage2_26[68]},
      {stage2_28[49], stage2_28[50], stage2_28[51], stage2_28[52], stage2_28[53], stage2_28[54]},
      {stage3_30[9],stage3_29[9],stage3_28[11],stage3_27[25],stage3_26[34]}
   );
   gpc606_5 gpc3647 (
      {stage2_26[69], stage2_26[70], stage2_26[71], stage2_26[72], stage2_26[73], stage2_26[74]},
      {stage2_28[55], stage2_28[56], stage2_28[57], stage2_28[58], stage2_28[59], stage2_28[60]},
      {stage3_30[10],stage3_29[10],stage3_28[12],stage3_27[26],stage3_26[35]}
   );
   gpc606_5 gpc3648 (
      {stage2_26[75], stage2_26[76], stage2_26[77], stage2_26[78], stage2_26[79], stage2_26[80]},
      {stage2_28[61], stage2_28[62], stage2_28[63], stage2_28[64], stage2_28[65], stage2_28[66]},
      {stage3_30[11],stage3_29[11],stage3_28[13],stage3_27[27],stage3_26[36]}
   );
   gpc606_5 gpc3649 (
      {stage2_26[81], stage2_26[82], stage2_26[83], stage2_26[84], stage2_26[85], stage2_26[86]},
      {stage2_28[67], stage2_28[68], stage2_28[69], stage2_28[70], stage2_28[71], stage2_28[72]},
      {stage3_30[12],stage3_29[12],stage3_28[14],stage3_27[28],stage3_26[37]}
   );
   gpc606_5 gpc3650 (
      {stage2_27[6], stage2_27[7], stage2_27[8], stage2_27[9], stage2_27[10], stage2_27[11]},
      {stage2_29[1], stage2_29[2], stage2_29[3], stage2_29[4], stage2_29[5], stage2_29[6]},
      {stage3_31[0],stage3_30[13],stage3_29[13],stage3_28[15],stage3_27[29]}
   );
   gpc615_5 gpc3651 (
      {stage2_27[12], stage2_27[13], stage2_27[14], stage2_27[15], stage2_27[16]},
      {stage2_28[73]},
      {stage2_29[7], stage2_29[8], stage2_29[9], stage2_29[10], stage2_29[11], stage2_29[12]},
      {stage3_31[1],stage3_30[14],stage3_29[14],stage3_28[16],stage3_27[30]}
   );
   gpc615_5 gpc3652 (
      {stage2_27[17], stage2_27[18], stage2_27[19], stage2_27[20], stage2_27[21]},
      {stage2_28[74]},
      {stage2_29[13], stage2_29[14], stage2_29[15], stage2_29[16], stage2_29[17], stage2_29[18]},
      {stage3_31[2],stage3_30[15],stage3_29[15],stage3_28[17],stage3_27[31]}
   );
   gpc615_5 gpc3653 (
      {stage2_27[22], stage2_27[23], stage2_27[24], stage2_27[25], stage2_27[26]},
      {stage2_28[75]},
      {stage2_29[19], stage2_29[20], stage2_29[21], stage2_29[22], stage2_29[23], stage2_29[24]},
      {stage3_31[3],stage3_30[16],stage3_29[16],stage3_28[18],stage3_27[32]}
   );
   gpc615_5 gpc3654 (
      {stage2_27[27], stage2_27[28], stage2_27[29], stage2_27[30], stage2_27[31]},
      {stage2_28[76]},
      {stage2_29[25], stage2_29[26], stage2_29[27], stage2_29[28], stage2_29[29], stage2_29[30]},
      {stage3_31[4],stage3_30[17],stage3_29[17],stage3_28[19],stage3_27[33]}
   );
   gpc615_5 gpc3655 (
      {stage2_27[32], stage2_27[33], stage2_27[34], stage2_27[35], stage2_27[36]},
      {stage2_28[77]},
      {stage2_29[31], stage2_29[32], stage2_29[33], stage2_29[34], stage2_29[35], stage2_29[36]},
      {stage3_31[5],stage3_30[18],stage3_29[18],stage3_28[20],stage3_27[34]}
   );
   gpc615_5 gpc3656 (
      {stage2_27[37], stage2_27[38], stage2_27[39], stage2_27[40], stage2_27[41]},
      {stage2_28[78]},
      {stage2_29[37], stage2_29[38], stage2_29[39], stage2_29[40], stage2_29[41], stage2_29[42]},
      {stage3_31[6],stage3_30[19],stage3_29[19],stage3_28[21],stage3_27[35]}
   );
   gpc615_5 gpc3657 (
      {stage2_27[42], stage2_27[43], stage2_27[44], stage2_27[45], stage2_27[46]},
      {stage2_28[79]},
      {stage2_29[43], stage2_29[44], stage2_29[45], stage2_29[46], stage2_29[47], stage2_29[48]},
      {stage3_31[7],stage3_30[20],stage3_29[20],stage3_28[22],stage3_27[36]}
   );
   gpc615_5 gpc3658 (
      {stage2_27[47], stage2_27[48], stage2_27[49], stage2_27[50], stage2_27[51]},
      {stage2_28[80]},
      {stage2_29[49], stage2_29[50], stage2_29[51], stage2_29[52], stage2_29[53], stage2_29[54]},
      {stage3_31[8],stage3_30[21],stage3_29[21],stage3_28[23],stage3_27[37]}
   );
   gpc615_5 gpc3659 (
      {stage2_27[52], stage2_27[53], stage2_27[54], stage2_27[55], stage2_27[56]},
      {stage2_28[81]},
      {stage2_29[55], stage2_29[56], stage2_29[57], stage2_29[58], stage2_29[59], stage2_29[60]},
      {stage3_31[9],stage3_30[22],stage3_29[22],stage3_28[24],stage3_27[38]}
   );
   gpc615_5 gpc3660 (
      {stage2_27[57], stage2_27[58], stage2_27[59], stage2_27[60], stage2_27[61]},
      {stage2_28[82]},
      {stage2_29[61], stage2_29[62], stage2_29[63], stage2_29[64], stage2_29[65], stage2_29[66]},
      {stage3_31[10],stage3_30[23],stage3_29[23],stage3_28[25],stage3_27[39]}
   );
   gpc615_5 gpc3661 (
      {stage2_27[62], stage2_27[63], stage2_27[64], stage2_27[65], stage2_27[66]},
      {stage2_28[83]},
      {stage2_29[67], stage2_29[68], stage2_29[69], stage2_29[70], stage2_29[71], stage2_29[72]},
      {stage3_31[11],stage3_30[24],stage3_29[24],stage3_28[26],stage3_27[40]}
   );
   gpc615_5 gpc3662 (
      {stage2_27[67], stage2_27[68], stage2_27[69], stage2_27[70], stage2_27[71]},
      {stage2_28[84]},
      {stage2_29[73], stage2_29[74], stage2_29[75], stage2_29[76], stage2_29[77], stage2_29[78]},
      {stage3_31[12],stage3_30[25],stage3_29[25],stage3_28[27],stage3_27[41]}
   );
   gpc606_5 gpc3663 (
      {stage2_28[85], stage2_28[86], stage2_28[87], stage2_28[88], stage2_28[89], stage2_28[90]},
      {stage2_30[0], stage2_30[1], stage2_30[2], stage2_30[3], stage2_30[4], stage2_30[5]},
      {stage3_32[0],stage3_31[13],stage3_30[26],stage3_29[26],stage3_28[28]}
   );
   gpc606_5 gpc3664 (
      {stage2_28[91], stage2_28[92], stage2_28[93], stage2_28[94], stage2_28[95], stage2_28[96]},
      {stage2_30[6], stage2_30[7], stage2_30[8], stage2_30[9], stage2_30[10], stage2_30[11]},
      {stage3_32[1],stage3_31[14],stage3_30[27],stage3_29[27],stage3_28[29]}
   );
   gpc606_5 gpc3665 (
      {stage2_28[97], stage2_28[98], stage2_28[99], stage2_28[100], stage2_28[101], stage2_28[102]},
      {stage2_30[12], stage2_30[13], stage2_30[14], stage2_30[15], stage2_30[16], stage2_30[17]},
      {stage3_32[2],stage3_31[15],stage3_30[28],stage3_29[28],stage3_28[30]}
   );
   gpc606_5 gpc3666 (
      {stage2_28[103], stage2_28[104], stage2_28[105], stage2_28[106], stage2_28[107], stage2_28[108]},
      {stage2_30[18], stage2_30[19], stage2_30[20], stage2_30[21], stage2_30[22], stage2_30[23]},
      {stage3_32[3],stage3_31[16],stage3_30[29],stage3_29[29],stage3_28[31]}
   );
   gpc606_5 gpc3667 (
      {stage2_28[109], stage2_28[110], stage2_28[111], stage2_28[112], stage2_28[113], stage2_28[114]},
      {stage2_30[24], stage2_30[25], stage2_30[26], stage2_30[27], stage2_30[28], stage2_30[29]},
      {stage3_32[4],stage3_31[17],stage3_30[30],stage3_29[30],stage3_28[32]}
   );
   gpc606_5 gpc3668 (
      {stage2_28[115], stage2_28[116], stage2_28[117], stage2_28[118], stage2_28[119], stage2_28[120]},
      {stage2_30[30], stage2_30[31], stage2_30[32], stage2_30[33], stage2_30[34], stage2_30[35]},
      {stage3_32[5],stage3_31[18],stage3_30[31],stage3_29[31],stage3_28[33]}
   );
   gpc606_5 gpc3669 (
      {stage2_28[121], stage2_28[122], stage2_28[123], stage2_28[124], stage2_28[125], stage2_28[126]},
      {stage2_30[36], stage2_30[37], stage2_30[38], stage2_30[39], stage2_30[40], stage2_30[41]},
      {stage3_32[6],stage3_31[19],stage3_30[32],stage3_29[32],stage3_28[34]}
   );
   gpc606_5 gpc3670 (
      {stage2_28[127], stage2_28[128], stage2_28[129], stage2_28[130], stage2_28[131], stage2_28[132]},
      {stage2_30[42], stage2_30[43], stage2_30[44], stage2_30[45], stage2_30[46], stage2_30[47]},
      {stage3_32[7],stage3_31[20],stage3_30[33],stage3_29[33],stage3_28[35]}
   );
   gpc606_5 gpc3671 (
      {stage2_29[79], stage2_29[80], stage2_29[81], stage2_29[82], stage2_29[83], stage2_29[84]},
      {stage2_31[0], stage2_31[1], stage2_31[2], stage2_31[3], stage2_31[4], stage2_31[5]},
      {stage3_33[0],stage3_32[8],stage3_31[21],stage3_30[34],stage3_29[34]}
   );
   gpc606_5 gpc3672 (
      {stage2_29[85], stage2_29[86], stage2_29[87], stage2_29[88], stage2_29[89], stage2_29[90]},
      {stage2_31[6], stage2_31[7], stage2_31[8], stage2_31[9], stage2_31[10], stage2_31[11]},
      {stage3_33[1],stage3_32[9],stage3_31[22],stage3_30[35],stage3_29[35]}
   );
   gpc606_5 gpc3673 (
      {stage2_29[91], stage2_29[92], stage2_29[93], stage2_29[94], stage2_29[95], stage2_29[96]},
      {stage2_31[12], stage2_31[13], stage2_31[14], stage2_31[15], stage2_31[16], stage2_31[17]},
      {stage3_33[2],stage3_32[10],stage3_31[23],stage3_30[36],stage3_29[36]}
   );
   gpc606_5 gpc3674 (
      {stage2_29[97], stage2_29[98], stage2_29[99], stage2_29[100], stage2_29[101], stage2_29[102]},
      {stage2_31[18], stage2_31[19], stage2_31[20], stage2_31[21], stage2_31[22], stage2_31[23]},
      {stage3_33[3],stage3_32[11],stage3_31[24],stage3_30[37],stage3_29[37]}
   );
   gpc606_5 gpc3675 (
      {stage2_29[103], stage2_29[104], stage2_29[105], stage2_29[106], stage2_29[107], stage2_29[108]},
      {stage2_31[24], stage2_31[25], stage2_31[26], stage2_31[27], stage2_31[28], stage2_31[29]},
      {stage3_33[4],stage3_32[12],stage3_31[25],stage3_30[38],stage3_29[38]}
   );
   gpc606_5 gpc3676 (
      {stage2_29[109], stage2_29[110], stage2_29[111], stage2_29[112], stage2_29[113], stage2_29[114]},
      {stage2_31[30], stage2_31[31], stage2_31[32], stage2_31[33], stage2_31[34], stage2_31[35]},
      {stage3_33[5],stage3_32[13],stage3_31[26],stage3_30[39],stage3_29[39]}
   );
   gpc606_5 gpc3677 (
      {stage2_29[115], stage2_29[116], stage2_29[117], stage2_29[118], stage2_29[119], stage2_29[120]},
      {stage2_31[36], stage2_31[37], stage2_31[38], stage2_31[39], stage2_31[40], stage2_31[41]},
      {stage3_33[6],stage3_32[14],stage3_31[27],stage3_30[40],stage3_29[40]}
   );
   gpc606_5 gpc3678 (
      {stage2_29[121], stage2_29[122], stage2_29[123], stage2_29[124], stage2_29[125], stage2_29[126]},
      {stage2_31[42], stage2_31[43], stage2_31[44], stage2_31[45], stage2_31[46], stage2_31[47]},
      {stage3_33[7],stage3_32[15],stage3_31[28],stage3_30[41],stage3_29[41]}
   );
   gpc606_5 gpc3679 (
      {stage2_30[48], stage2_30[49], stage2_30[50], stage2_30[51], stage2_30[52], stage2_30[53]},
      {stage2_32[0], stage2_32[1], stage2_32[2], stage2_32[3], stage2_32[4], stage2_32[5]},
      {stage3_34[0],stage3_33[8],stage3_32[16],stage3_31[29],stage3_30[42]}
   );
   gpc606_5 gpc3680 (
      {stage2_30[54], stage2_30[55], stage2_30[56], stage2_30[57], stage2_30[58], stage2_30[59]},
      {stage2_32[6], stage2_32[7], stage2_32[8], stage2_32[9], stage2_32[10], stage2_32[11]},
      {stage3_34[1],stage3_33[9],stage3_32[17],stage3_31[30],stage3_30[43]}
   );
   gpc606_5 gpc3681 (
      {stage2_30[60], stage2_30[61], stage2_30[62], stage2_30[63], stage2_30[64], stage2_30[65]},
      {stage2_32[12], stage2_32[13], stage2_32[14], stage2_32[15], stage2_32[16], stage2_32[17]},
      {stage3_34[2],stage3_33[10],stage3_32[18],stage3_31[31],stage3_30[44]}
   );
   gpc615_5 gpc3682 (
      {stage2_31[48], stage2_31[49], stage2_31[50], stage2_31[51], stage2_31[52]},
      {stage2_32[18]},
      {stage2_33[0], stage2_33[1], stage2_33[2], stage2_33[3], stage2_33[4], stage2_33[5]},
      {stage3_35[0],stage3_34[3],stage3_33[11],stage3_32[19],stage3_31[32]}
   );
   gpc615_5 gpc3683 (
      {stage2_31[53], stage2_31[54], stage2_31[55], stage2_31[56], stage2_31[57]},
      {stage2_32[19]},
      {stage2_33[6], stage2_33[7], stage2_33[8], stage2_33[9], stage2_33[10], stage2_33[11]},
      {stage3_35[1],stage3_34[4],stage3_33[12],stage3_32[20],stage3_31[33]}
   );
   gpc615_5 gpc3684 (
      {stage2_31[58], stage2_31[59], stage2_31[60], stage2_31[61], stage2_31[62]},
      {stage2_32[20]},
      {stage2_33[12], stage2_33[13], stage2_33[14], stage2_33[15], stage2_33[16], stage2_33[17]},
      {stage3_35[2],stage3_34[5],stage3_33[13],stage3_32[21],stage3_31[34]}
   );
   gpc615_5 gpc3685 (
      {stage2_31[63], stage2_31[64], stage2_31[65], stage2_31[66], stage2_31[67]},
      {stage2_32[21]},
      {stage2_33[18], stage2_33[19], stage2_33[20], stage2_33[21], stage2_33[22], stage2_33[23]},
      {stage3_35[3],stage3_34[6],stage3_33[14],stage3_32[22],stage3_31[35]}
   );
   gpc615_5 gpc3686 (
      {stage2_31[68], stage2_31[69], stage2_31[70], stage2_31[71], stage2_31[72]},
      {stage2_32[22]},
      {stage2_33[24], stage2_33[25], stage2_33[26], stage2_33[27], stage2_33[28], stage2_33[29]},
      {stage3_35[4],stage3_34[7],stage3_33[15],stage3_32[23],stage3_31[36]}
   );
   gpc615_5 gpc3687 (
      {stage2_31[73], stage2_31[74], stage2_31[75], stage2_31[76], stage2_31[77]},
      {stage2_32[23]},
      {stage2_33[30], stage2_33[31], stage2_33[32], stage2_33[33], stage2_33[34], stage2_33[35]},
      {stage3_35[5],stage3_34[8],stage3_33[16],stage3_32[24],stage3_31[37]}
   );
   gpc615_5 gpc3688 (
      {stage2_31[78], stage2_31[79], stage2_31[80], stage2_31[81], stage2_31[82]},
      {stage2_32[24]},
      {stage2_33[36], stage2_33[37], stage2_33[38], stage2_33[39], stage2_33[40], stage2_33[41]},
      {stage3_35[6],stage3_34[9],stage3_33[17],stage3_32[25],stage3_31[38]}
   );
   gpc606_5 gpc3689 (
      {stage2_32[25], stage2_32[26], stage2_32[27], stage2_32[28], stage2_32[29], stage2_32[30]},
      {stage2_34[0], stage2_34[1], stage2_34[2], stage2_34[3], stage2_34[4], stage2_34[5]},
      {stage3_36[0],stage3_35[7],stage3_34[10],stage3_33[18],stage3_32[26]}
   );
   gpc615_5 gpc3690 (
      {stage2_32[31], stage2_32[32], stage2_32[33], stage2_32[34], stage2_32[35]},
      {stage2_33[42]},
      {stage2_34[6], stage2_34[7], stage2_34[8], stage2_34[9], stage2_34[10], stage2_34[11]},
      {stage3_36[1],stage3_35[8],stage3_34[11],stage3_33[19],stage3_32[27]}
   );
   gpc615_5 gpc3691 (
      {stage2_32[36], stage2_32[37], stage2_32[38], stage2_32[39], stage2_32[40]},
      {stage2_33[43]},
      {stage2_34[12], stage2_34[13], stage2_34[14], stage2_34[15], stage2_34[16], stage2_34[17]},
      {stage3_36[2],stage3_35[9],stage3_34[12],stage3_33[20],stage3_32[28]}
   );
   gpc615_5 gpc3692 (
      {stage2_32[41], stage2_32[42], stage2_32[43], stage2_32[44], stage2_32[45]},
      {stage2_33[44]},
      {stage2_34[18], stage2_34[19], stage2_34[20], stage2_34[21], stage2_34[22], stage2_34[23]},
      {stage3_36[3],stage3_35[10],stage3_34[13],stage3_33[21],stage3_32[29]}
   );
   gpc606_5 gpc3693 (
      {stage2_33[45], stage2_33[46], stage2_33[47], stage2_33[48], stage2_33[49], stage2_33[50]},
      {stage2_35[0], stage2_35[1], stage2_35[2], stage2_35[3], stage2_35[4], stage2_35[5]},
      {stage3_37[0],stage3_36[4],stage3_35[11],stage3_34[14],stage3_33[22]}
   );
   gpc606_5 gpc3694 (
      {stage2_33[51], stage2_33[52], stage2_33[53], stage2_33[54], stage2_33[55], stage2_33[56]},
      {stage2_35[6], stage2_35[7], stage2_35[8], stage2_35[9], stage2_35[10], stage2_35[11]},
      {stage3_37[1],stage3_36[5],stage3_35[12],stage3_34[15],stage3_33[23]}
   );
   gpc1_1 gpc3695 (
      {stage2_1[48]},
      {stage3_1[18]}
   );
   gpc1_1 gpc3696 (
      {stage2_1[49]},
      {stage3_1[19]}
   );
   gpc1_1 gpc3697 (
      {stage2_1[50]},
      {stage3_1[20]}
   );
   gpc1_1 gpc3698 (
      {stage2_1[51]},
      {stage3_1[21]}
   );
   gpc1_1 gpc3699 (
      {stage2_1[52]},
      {stage3_1[22]}
   );
   gpc1_1 gpc3700 (
      {stage2_1[53]},
      {stage3_1[23]}
   );
   gpc1_1 gpc3701 (
      {stage2_1[54]},
      {stage3_1[24]}
   );
   gpc1_1 gpc3702 (
      {stage2_1[55]},
      {stage3_1[25]}
   );
   gpc1_1 gpc3703 (
      {stage2_2[81]},
      {stage3_2[22]}
   );
   gpc1_1 gpc3704 (
      {stage2_2[82]},
      {stage3_2[23]}
   );
   gpc1_1 gpc3705 (
      {stage2_2[83]},
      {stage3_2[24]}
   );
   gpc1_1 gpc3706 (
      {stage2_2[84]},
      {stage3_2[25]}
   );
   gpc1_1 gpc3707 (
      {stage2_2[85]},
      {stage3_2[26]}
   );
   gpc1_1 gpc3708 (
      {stage2_2[86]},
      {stage3_2[27]}
   );
   gpc1_1 gpc3709 (
      {stage2_2[87]},
      {stage3_2[28]}
   );
   gpc1_1 gpc3710 (
      {stage2_2[88]},
      {stage3_2[29]}
   );
   gpc1_1 gpc3711 (
      {stage2_2[89]},
      {stage3_2[30]}
   );
   gpc1_1 gpc3712 (
      {stage2_2[90]},
      {stage3_2[31]}
   );
   gpc1_1 gpc3713 (
      {stage2_2[91]},
      {stage3_2[32]}
   );
   gpc1_1 gpc3714 (
      {stage2_2[92]},
      {stage3_2[33]}
   );
   gpc1_1 gpc3715 (
      {stage2_2[93]},
      {stage3_2[34]}
   );
   gpc1_1 gpc3716 (
      {stage2_2[94]},
      {stage3_2[35]}
   );
   gpc1_1 gpc3717 (
      {stage2_4[114]},
      {stage3_4[42]}
   );
   gpc1_1 gpc3718 (
      {stage2_4[115]},
      {stage3_4[43]}
   );
   gpc1_1 gpc3719 (
      {stage2_4[116]},
      {stage3_4[44]}
   );
   gpc1_1 gpc3720 (
      {stage2_4[117]},
      {stage3_4[45]}
   );
   gpc1_1 gpc3721 (
      {stage2_4[118]},
      {stage3_4[46]}
   );
   gpc1_1 gpc3722 (
      {stage2_5[72]},
      {stage3_5[37]}
   );
   gpc1_1 gpc3723 (
      {stage2_5[73]},
      {stage3_5[38]}
   );
   gpc1_1 gpc3724 (
      {stage2_5[74]},
      {stage3_5[39]}
   );
   gpc1_1 gpc3725 (
      {stage2_5[75]},
      {stage3_5[40]}
   );
   gpc1_1 gpc3726 (
      {stage2_5[76]},
      {stage3_5[41]}
   );
   gpc1_1 gpc3727 (
      {stage2_5[77]},
      {stage3_5[42]}
   );
   gpc1_1 gpc3728 (
      {stage2_5[78]},
      {stage3_5[43]}
   );
   gpc1_1 gpc3729 (
      {stage2_5[79]},
      {stage3_5[44]}
   );
   gpc1_1 gpc3730 (
      {stage2_5[80]},
      {stage3_5[45]}
   );
   gpc1_1 gpc3731 (
      {stage2_5[81]},
      {stage3_5[46]}
   );
   gpc1_1 gpc3732 (
      {stage2_5[82]},
      {stage3_5[47]}
   );
   gpc1_1 gpc3733 (
      {stage2_5[83]},
      {stage3_5[48]}
   );
   gpc1_1 gpc3734 (
      {stage2_5[84]},
      {stage3_5[49]}
   );
   gpc1_1 gpc3735 (
      {stage2_5[85]},
      {stage3_5[50]}
   );
   gpc1_1 gpc3736 (
      {stage2_5[86]},
      {stage3_5[51]}
   );
   gpc1_1 gpc3737 (
      {stage2_5[87]},
      {stage3_5[52]}
   );
   gpc1_1 gpc3738 (
      {stage2_5[88]},
      {stage3_5[53]}
   );
   gpc1_1 gpc3739 (
      {stage2_5[89]},
      {stage3_5[54]}
   );
   gpc1_1 gpc3740 (
      {stage2_5[90]},
      {stage3_5[55]}
   );
   gpc1_1 gpc3741 (
      {stage2_5[91]},
      {stage3_5[56]}
   );
   gpc1_1 gpc3742 (
      {stage2_5[92]},
      {stage3_5[57]}
   );
   gpc1_1 gpc3743 (
      {stage2_5[93]},
      {stage3_5[58]}
   );
   gpc1_1 gpc3744 (
      {stage2_6[89]},
      {stage3_6[31]}
   );
   gpc1_1 gpc3745 (
      {stage2_6[90]},
      {stage3_6[32]}
   );
   gpc1_1 gpc3746 (
      {stage2_6[91]},
      {stage3_6[33]}
   );
   gpc1_1 gpc3747 (
      {stage2_6[92]},
      {stage3_6[34]}
   );
   gpc1_1 gpc3748 (
      {stage2_6[93]},
      {stage3_6[35]}
   );
   gpc1_1 gpc3749 (
      {stage2_6[94]},
      {stage3_6[36]}
   );
   gpc1_1 gpc3750 (
      {stage2_6[95]},
      {stage3_6[37]}
   );
   gpc1_1 gpc3751 (
      {stage2_7[102]},
      {stage3_7[40]}
   );
   gpc1_1 gpc3752 (
      {stage2_7[103]},
      {stage3_7[41]}
   );
   gpc1_1 gpc3753 (
      {stage2_7[104]},
      {stage3_7[42]}
   );
   gpc1_1 gpc3754 (
      {stage2_7[105]},
      {stage3_7[43]}
   );
   gpc1_1 gpc3755 (
      {stage2_7[106]},
      {stage3_7[44]}
   );
   gpc1_1 gpc3756 (
      {stage2_7[107]},
      {stage3_7[45]}
   );
   gpc1_1 gpc3757 (
      {stage2_7[108]},
      {stage3_7[46]}
   );
   gpc1_1 gpc3758 (
      {stage2_8[43]},
      {stage3_8[38]}
   );
   gpc1_1 gpc3759 (
      {stage2_8[44]},
      {stage3_8[39]}
   );
   gpc1_1 gpc3760 (
      {stage2_8[45]},
      {stage3_8[40]}
   );
   gpc1_1 gpc3761 (
      {stage2_8[46]},
      {stage3_8[41]}
   );
   gpc1_1 gpc3762 (
      {stage2_8[47]},
      {stage3_8[42]}
   );
   gpc1_1 gpc3763 (
      {stage2_8[48]},
      {stage3_8[43]}
   );
   gpc1_1 gpc3764 (
      {stage2_8[49]},
      {stage3_8[44]}
   );
   gpc1_1 gpc3765 (
      {stage2_8[50]},
      {stage3_8[45]}
   );
   gpc1_1 gpc3766 (
      {stage2_8[51]},
      {stage3_8[46]}
   );
   gpc1_1 gpc3767 (
      {stage2_8[52]},
      {stage3_8[47]}
   );
   gpc1_1 gpc3768 (
      {stage2_8[53]},
      {stage3_8[48]}
   );
   gpc1_1 gpc3769 (
      {stage2_8[54]},
      {stage3_8[49]}
   );
   gpc1_1 gpc3770 (
      {stage2_8[55]},
      {stage3_8[50]}
   );
   gpc1_1 gpc3771 (
      {stage2_8[56]},
      {stage3_8[51]}
   );
   gpc1_1 gpc3772 (
      {stage2_8[57]},
      {stage3_8[52]}
   );
   gpc1_1 gpc3773 (
      {stage2_8[58]},
      {stage3_8[53]}
   );
   gpc1_1 gpc3774 (
      {stage2_8[59]},
      {stage3_8[54]}
   );
   gpc1_1 gpc3775 (
      {stage2_8[60]},
      {stage3_8[55]}
   );
   gpc1_1 gpc3776 (
      {stage2_8[61]},
      {stage3_8[56]}
   );
   gpc1_1 gpc3777 (
      {stage2_8[62]},
      {stage3_8[57]}
   );
   gpc1_1 gpc3778 (
      {stage2_8[63]},
      {stage3_8[58]}
   );
   gpc1_1 gpc3779 (
      {stage2_8[64]},
      {stage3_8[59]}
   );
   gpc1_1 gpc3780 (
      {stage2_8[65]},
      {stage3_8[60]}
   );
   gpc1_1 gpc3781 (
      {stage2_8[66]},
      {stage3_8[61]}
   );
   gpc1_1 gpc3782 (
      {stage2_8[67]},
      {stage3_8[62]}
   );
   gpc1_1 gpc3783 (
      {stage2_8[68]},
      {stage3_8[63]}
   );
   gpc1_1 gpc3784 (
      {stage2_8[69]},
      {stage3_8[64]}
   );
   gpc1_1 gpc3785 (
      {stage2_8[70]},
      {stage3_8[65]}
   );
   gpc1_1 gpc3786 (
      {stage2_8[71]},
      {stage3_8[66]}
   );
   gpc1_1 gpc3787 (
      {stage2_8[72]},
      {stage3_8[67]}
   );
   gpc1_1 gpc3788 (
      {stage2_8[73]},
      {stage3_8[68]}
   );
   gpc1_1 gpc3789 (
      {stage2_8[74]},
      {stage3_8[69]}
   );
   gpc1_1 gpc3790 (
      {stage2_8[75]},
      {stage3_8[70]}
   );
   gpc1_1 gpc3791 (
      {stage2_8[76]},
      {stage3_8[71]}
   );
   gpc1_1 gpc3792 (
      {stage2_8[77]},
      {stage3_8[72]}
   );
   gpc1_1 gpc3793 (
      {stage2_8[78]},
      {stage3_8[73]}
   );
   gpc1_1 gpc3794 (
      {stage2_8[79]},
      {stage3_8[74]}
   );
   gpc1_1 gpc3795 (
      {stage2_8[80]},
      {stage3_8[75]}
   );
   gpc1_1 gpc3796 (
      {stage2_8[81]},
      {stage3_8[76]}
   );
   gpc1_1 gpc3797 (
      {stage2_8[82]},
      {stage3_8[77]}
   );
   gpc1_1 gpc3798 (
      {stage2_8[83]},
      {stage3_8[78]}
   );
   gpc1_1 gpc3799 (
      {stage2_8[84]},
      {stage3_8[79]}
   );
   gpc1_1 gpc3800 (
      {stage2_8[85]},
      {stage3_8[80]}
   );
   gpc1_1 gpc3801 (
      {stage2_8[86]},
      {stage3_8[81]}
   );
   gpc1_1 gpc3802 (
      {stage2_8[87]},
      {stage3_8[82]}
   );
   gpc1_1 gpc3803 (
      {stage2_8[88]},
      {stage3_8[83]}
   );
   gpc1_1 gpc3804 (
      {stage2_8[89]},
      {stage3_8[84]}
   );
   gpc1_1 gpc3805 (
      {stage2_8[90]},
      {stage3_8[85]}
   );
   gpc1_1 gpc3806 (
      {stage2_8[91]},
      {stage3_8[86]}
   );
   gpc1_1 gpc3807 (
      {stage2_8[92]},
      {stage3_8[87]}
   );
   gpc1_1 gpc3808 (
      {stage2_8[93]},
      {stage3_8[88]}
   );
   gpc1_1 gpc3809 (
      {stage2_8[94]},
      {stage3_8[89]}
   );
   gpc1_1 gpc3810 (
      {stage2_8[95]},
      {stage3_8[90]}
   );
   gpc1_1 gpc3811 (
      {stage2_8[96]},
      {stage3_8[91]}
   );
   gpc1_1 gpc3812 (
      {stage2_8[97]},
      {stage3_8[92]}
   );
   gpc1_1 gpc3813 (
      {stage2_9[83]},
      {stage3_9[25]}
   );
   gpc1_1 gpc3814 (
      {stage2_9[84]},
      {stage3_9[26]}
   );
   gpc1_1 gpc3815 (
      {stage2_9[85]},
      {stage3_9[27]}
   );
   gpc1_1 gpc3816 (
      {stage2_9[86]},
      {stage3_9[28]}
   );
   gpc1_1 gpc3817 (
      {stage2_9[87]},
      {stage3_9[29]}
   );
   gpc1_1 gpc3818 (
      {stage2_9[88]},
      {stage3_9[30]}
   );
   gpc1_1 gpc3819 (
      {stage2_9[89]},
      {stage3_9[31]}
   );
   gpc1_1 gpc3820 (
      {stage2_9[90]},
      {stage3_9[32]}
   );
   gpc1_1 gpc3821 (
      {stage2_9[91]},
      {stage3_9[33]}
   );
   gpc1_1 gpc3822 (
      {stage2_9[92]},
      {stage3_9[34]}
   );
   gpc1_1 gpc3823 (
      {stage2_9[93]},
      {stage3_9[35]}
   );
   gpc1_1 gpc3824 (
      {stage2_9[94]},
      {stage3_9[36]}
   );
   gpc1_1 gpc3825 (
      {stage2_9[95]},
      {stage3_9[37]}
   );
   gpc1_1 gpc3826 (
      {stage2_9[96]},
      {stage3_9[38]}
   );
   gpc1_1 gpc3827 (
      {stage2_9[97]},
      {stage3_9[39]}
   );
   gpc1_1 gpc3828 (
      {stage2_9[98]},
      {stage3_9[40]}
   );
   gpc1_1 gpc3829 (
      {stage2_9[99]},
      {stage3_9[41]}
   );
   gpc1_1 gpc3830 (
      {stage2_9[100]},
      {stage3_9[42]}
   );
   gpc1_1 gpc3831 (
      {stage2_9[101]},
      {stage3_9[43]}
   );
   gpc1_1 gpc3832 (
      {stage2_9[102]},
      {stage3_9[44]}
   );
   gpc1_1 gpc3833 (
      {stage2_9[103]},
      {stage3_9[45]}
   );
   gpc1_1 gpc3834 (
      {stage2_9[104]},
      {stage3_9[46]}
   );
   gpc1_1 gpc3835 (
      {stage2_9[105]},
      {stage3_9[47]}
   );
   gpc1_1 gpc3836 (
      {stage2_9[106]},
      {stage3_9[48]}
   );
   gpc1_1 gpc3837 (
      {stage2_9[107]},
      {stage3_9[49]}
   );
   gpc1_1 gpc3838 (
      {stage2_10[87]},
      {stage3_10[30]}
   );
   gpc1_1 gpc3839 (
      {stage2_10[88]},
      {stage3_10[31]}
   );
   gpc1_1 gpc3840 (
      {stage2_10[89]},
      {stage3_10[32]}
   );
   gpc1_1 gpc3841 (
      {stage2_10[90]},
      {stage3_10[33]}
   );
   gpc1_1 gpc3842 (
      {stage2_10[91]},
      {stage3_10[34]}
   );
   gpc1_1 gpc3843 (
      {stage2_10[92]},
      {stage3_10[35]}
   );
   gpc1_1 gpc3844 (
      {stage2_10[93]},
      {stage3_10[36]}
   );
   gpc1_1 gpc3845 (
      {stage2_10[94]},
      {stage3_10[37]}
   );
   gpc1_1 gpc3846 (
      {stage2_11[110]},
      {stage3_11[49]}
   );
   gpc1_1 gpc3847 (
      {stage2_11[111]},
      {stage3_11[50]}
   );
   gpc1_1 gpc3848 (
      {stage2_11[112]},
      {stage3_11[51]}
   );
   gpc1_1 gpc3849 (
      {stage2_11[113]},
      {stage3_11[52]}
   );
   gpc1_1 gpc3850 (
      {stage2_11[114]},
      {stage3_11[53]}
   );
   gpc1_1 gpc3851 (
      {stage2_11[115]},
      {stage3_11[54]}
   );
   gpc1_1 gpc3852 (
      {stage2_12[92]},
      {stage3_12[37]}
   );
   gpc1_1 gpc3853 (
      {stage2_12[93]},
      {stage3_12[38]}
   );
   gpc1_1 gpc3854 (
      {stage2_12[94]},
      {stage3_12[39]}
   );
   gpc1_1 gpc3855 (
      {stage2_12[95]},
      {stage3_12[40]}
   );
   gpc1_1 gpc3856 (
      {stage2_12[96]},
      {stage3_12[41]}
   );
   gpc1_1 gpc3857 (
      {stage2_12[97]},
      {stage3_12[42]}
   );
   gpc1_1 gpc3858 (
      {stage2_12[98]},
      {stage3_12[43]}
   );
   gpc1_1 gpc3859 (
      {stage2_12[99]},
      {stage3_12[44]}
   );
   gpc1_1 gpc3860 (
      {stage2_12[100]},
      {stage3_12[45]}
   );
   gpc1_1 gpc3861 (
      {stage2_12[101]},
      {stage3_12[46]}
   );
   gpc1_1 gpc3862 (
      {stage2_13[120]},
      {stage3_13[33]}
   );
   gpc1_1 gpc3863 (
      {stage2_13[121]},
      {stage3_13[34]}
   );
   gpc1_1 gpc3864 (
      {stage2_13[122]},
      {stage3_13[35]}
   );
   gpc1_1 gpc3865 (
      {stage2_13[123]},
      {stage3_13[36]}
   );
   gpc1_1 gpc3866 (
      {stage2_14[56]},
      {stage3_14[42]}
   );
   gpc1_1 gpc3867 (
      {stage2_14[57]},
      {stage3_14[43]}
   );
   gpc1_1 gpc3868 (
      {stage2_14[58]},
      {stage3_14[44]}
   );
   gpc1_1 gpc3869 (
      {stage2_14[59]},
      {stage3_14[45]}
   );
   gpc1_1 gpc3870 (
      {stage2_14[60]},
      {stage3_14[46]}
   );
   gpc1_1 gpc3871 (
      {stage2_14[61]},
      {stage3_14[47]}
   );
   gpc1_1 gpc3872 (
      {stage2_14[62]},
      {stage3_14[48]}
   );
   gpc1_1 gpc3873 (
      {stage2_14[63]},
      {stage3_14[49]}
   );
   gpc1_1 gpc3874 (
      {stage2_14[64]},
      {stage3_14[50]}
   );
   gpc1_1 gpc3875 (
      {stage2_14[65]},
      {stage3_14[51]}
   );
   gpc1_1 gpc3876 (
      {stage2_14[66]},
      {stage3_14[52]}
   );
   gpc1_1 gpc3877 (
      {stage2_14[67]},
      {stage3_14[53]}
   );
   gpc1_1 gpc3878 (
      {stage2_14[68]},
      {stage3_14[54]}
   );
   gpc1_1 gpc3879 (
      {stage2_14[69]},
      {stage3_14[55]}
   );
   gpc1_1 gpc3880 (
      {stage2_15[70]},
      {stage3_15[43]}
   );
   gpc1_1 gpc3881 (
      {stage2_15[71]},
      {stage3_15[44]}
   );
   gpc1_1 gpc3882 (
      {stage2_15[72]},
      {stage3_15[45]}
   );
   gpc1_1 gpc3883 (
      {stage2_15[73]},
      {stage3_15[46]}
   );
   gpc1_1 gpc3884 (
      {stage2_15[74]},
      {stage3_15[47]}
   );
   gpc1_1 gpc3885 (
      {stage2_15[75]},
      {stage3_15[48]}
   );
   gpc1_1 gpc3886 (
      {stage2_15[76]},
      {stage3_15[49]}
   );
   gpc1_1 gpc3887 (
      {stage2_15[77]},
      {stage3_15[50]}
   );
   gpc1_1 gpc3888 (
      {stage2_15[78]},
      {stage3_15[51]}
   );
   gpc1_1 gpc3889 (
      {stage2_15[79]},
      {stage3_15[52]}
   );
   gpc1_1 gpc3890 (
      {stage2_15[80]},
      {stage3_15[53]}
   );
   gpc1_1 gpc3891 (
      {stage2_15[81]},
      {stage3_15[54]}
   );
   gpc1_1 gpc3892 (
      {stage2_15[82]},
      {stage3_15[55]}
   );
   gpc1_1 gpc3893 (
      {stage2_15[83]},
      {stage3_15[56]}
   );
   gpc1_1 gpc3894 (
      {stage2_15[84]},
      {stage3_15[57]}
   );
   gpc1_1 gpc3895 (
      {stage2_15[85]},
      {stage3_15[58]}
   );
   gpc1_1 gpc3896 (
      {stage2_15[86]},
      {stage3_15[59]}
   );
   gpc1_1 gpc3897 (
      {stage2_15[87]},
      {stage3_15[60]}
   );
   gpc1_1 gpc3898 (
      {stage2_15[88]},
      {stage3_15[61]}
   );
   gpc1_1 gpc3899 (
      {stage2_15[89]},
      {stage3_15[62]}
   );
   gpc1_1 gpc3900 (
      {stage2_15[90]},
      {stage3_15[63]}
   );
   gpc1_1 gpc3901 (
      {stage2_15[91]},
      {stage3_15[64]}
   );
   gpc1_1 gpc3902 (
      {stage2_15[92]},
      {stage3_15[65]}
   );
   gpc1_1 gpc3903 (
      {stage2_15[93]},
      {stage3_15[66]}
   );
   gpc1_1 gpc3904 (
      {stage2_15[94]},
      {stage3_15[67]}
   );
   gpc1_1 gpc3905 (
      {stage2_15[95]},
      {stage3_15[68]}
   );
   gpc1_1 gpc3906 (
      {stage2_15[96]},
      {stage3_15[69]}
   );
   gpc1_1 gpc3907 (
      {stage2_15[97]},
      {stage3_15[70]}
   );
   gpc1_1 gpc3908 (
      {stage2_16[83]},
      {stage3_16[25]}
   );
   gpc1_1 gpc3909 (
      {stage2_16[84]},
      {stage3_16[26]}
   );
   gpc1_1 gpc3910 (
      {stage2_16[85]},
      {stage3_16[27]}
   );
   gpc1_1 gpc3911 (
      {stage2_16[86]},
      {stage3_16[28]}
   );
   gpc1_1 gpc3912 (
      {stage2_16[87]},
      {stage3_16[29]}
   );
   gpc1_1 gpc3913 (
      {stage2_16[88]},
      {stage3_16[30]}
   );
   gpc1_1 gpc3914 (
      {stage2_16[89]},
      {stage3_16[31]}
   );
   gpc1_1 gpc3915 (
      {stage2_16[90]},
      {stage3_16[32]}
   );
   gpc1_1 gpc3916 (
      {stage2_16[91]},
      {stage3_16[33]}
   );
   gpc1_1 gpc3917 (
      {stage2_16[92]},
      {stage3_16[34]}
   );
   gpc1_1 gpc3918 (
      {stage2_16[93]},
      {stage3_16[35]}
   );
   gpc1_1 gpc3919 (
      {stage2_16[94]},
      {stage3_16[36]}
   );
   gpc1_1 gpc3920 (
      {stage2_16[95]},
      {stage3_16[37]}
   );
   gpc1_1 gpc3921 (
      {stage2_16[96]},
      {stage3_16[38]}
   );
   gpc1_1 gpc3922 (
      {stage2_16[97]},
      {stage3_16[39]}
   );
   gpc1_1 gpc3923 (
      {stage2_16[98]},
      {stage3_16[40]}
   );
   gpc1_1 gpc3924 (
      {stage2_16[99]},
      {stage3_16[41]}
   );
   gpc1_1 gpc3925 (
      {stage2_16[100]},
      {stage3_16[42]}
   );
   gpc1_1 gpc3926 (
      {stage2_16[101]},
      {stage3_16[43]}
   );
   gpc1_1 gpc3927 (
      {stage2_16[102]},
      {stage3_16[44]}
   );
   gpc1_1 gpc3928 (
      {stage2_16[103]},
      {stage3_16[45]}
   );
   gpc1_1 gpc3929 (
      {stage2_16[104]},
      {stage3_16[46]}
   );
   gpc1_1 gpc3930 (
      {stage2_16[105]},
      {stage3_16[47]}
   );
   gpc1_1 gpc3931 (
      {stage2_16[106]},
      {stage3_16[48]}
   );
   gpc1_1 gpc3932 (
      {stage2_16[107]},
      {stage3_16[49]}
   );
   gpc1_1 gpc3933 (
      {stage2_16[108]},
      {stage3_16[50]}
   );
   gpc1_1 gpc3934 (
      {stage2_16[109]},
      {stage3_16[51]}
   );
   gpc1_1 gpc3935 (
      {stage2_16[110]},
      {stage3_16[52]}
   );
   gpc1_1 gpc3936 (
      {stage2_16[111]},
      {stage3_16[53]}
   );
   gpc1_1 gpc3937 (
      {stage2_16[112]},
      {stage3_16[54]}
   );
   gpc1_1 gpc3938 (
      {stage2_16[113]},
      {stage3_16[55]}
   );
   gpc1_1 gpc3939 (
      {stage2_16[114]},
      {stage3_16[56]}
   );
   gpc1_1 gpc3940 (
      {stage2_16[115]},
      {stage3_16[57]}
   );
   gpc1_1 gpc3941 (
      {stage2_16[116]},
      {stage3_16[58]}
   );
   gpc1_1 gpc3942 (
      {stage2_16[117]},
      {stage3_16[59]}
   );
   gpc1_1 gpc3943 (
      {stage2_16[118]},
      {stage3_16[60]}
   );
   gpc1_1 gpc3944 (
      {stage2_16[119]},
      {stage3_16[61]}
   );
   gpc1_1 gpc3945 (
      {stage2_16[120]},
      {stage3_16[62]}
   );
   gpc1_1 gpc3946 (
      {stage2_16[121]},
      {stage3_16[63]}
   );
   gpc1_1 gpc3947 (
      {stage2_16[122]},
      {stage3_16[64]}
   );
   gpc1_1 gpc3948 (
      {stage2_16[123]},
      {stage3_16[65]}
   );
   gpc1_1 gpc3949 (
      {stage2_16[124]},
      {stage3_16[66]}
   );
   gpc1_1 gpc3950 (
      {stage2_17[75]},
      {stage3_17[24]}
   );
   gpc1_1 gpc3951 (
      {stage2_17[76]},
      {stage3_17[25]}
   );
   gpc1_1 gpc3952 (
      {stage2_17[77]},
      {stage3_17[26]}
   );
   gpc1_1 gpc3953 (
      {stage2_17[78]},
      {stage3_17[27]}
   );
   gpc1_1 gpc3954 (
      {stage2_17[79]},
      {stage3_17[28]}
   );
   gpc1_1 gpc3955 (
      {stage2_17[80]},
      {stage3_17[29]}
   );
   gpc1_1 gpc3956 (
      {stage2_17[81]},
      {stage3_17[30]}
   );
   gpc1_1 gpc3957 (
      {stage2_17[82]},
      {stage3_17[31]}
   );
   gpc1_1 gpc3958 (
      {stage2_17[83]},
      {stage3_17[32]}
   );
   gpc1_1 gpc3959 (
      {stage2_17[84]},
      {stage3_17[33]}
   );
   gpc1_1 gpc3960 (
      {stage2_17[85]},
      {stage3_17[34]}
   );
   gpc1_1 gpc3961 (
      {stage2_17[86]},
      {stage3_17[35]}
   );
   gpc1_1 gpc3962 (
      {stage2_17[87]},
      {stage3_17[36]}
   );
   gpc1_1 gpc3963 (
      {stage2_17[88]},
      {stage3_17[37]}
   );
   gpc1_1 gpc3964 (
      {stage2_17[89]},
      {stage3_17[38]}
   );
   gpc1_1 gpc3965 (
      {stage2_17[90]},
      {stage3_17[39]}
   );
   gpc1_1 gpc3966 (
      {stage2_17[91]},
      {stage3_17[40]}
   );
   gpc1_1 gpc3967 (
      {stage2_17[92]},
      {stage3_17[41]}
   );
   gpc1_1 gpc3968 (
      {stage2_17[93]},
      {stage3_17[42]}
   );
   gpc1_1 gpc3969 (
      {stage2_17[94]},
      {stage3_17[43]}
   );
   gpc1_1 gpc3970 (
      {stage2_17[95]},
      {stage3_17[44]}
   );
   gpc1_1 gpc3971 (
      {stage2_17[96]},
      {stage3_17[45]}
   );
   gpc1_1 gpc3972 (
      {stage2_17[97]},
      {stage3_17[46]}
   );
   gpc1_1 gpc3973 (
      {stage2_17[98]},
      {stage3_17[47]}
   );
   gpc1_1 gpc3974 (
      {stage2_17[99]},
      {stage3_17[48]}
   );
   gpc1_1 gpc3975 (
      {stage2_17[100]},
      {stage3_17[49]}
   );
   gpc1_1 gpc3976 (
      {stage2_17[101]},
      {stage3_17[50]}
   );
   gpc1_1 gpc3977 (
      {stage2_17[102]},
      {stage3_17[51]}
   );
   gpc1_1 gpc3978 (
      {stage2_17[103]},
      {stage3_17[52]}
   );
   gpc1_1 gpc3979 (
      {stage2_17[104]},
      {stage3_17[53]}
   );
   gpc1_1 gpc3980 (
      {stage2_17[105]},
      {stage3_17[54]}
   );
   gpc1_1 gpc3981 (
      {stage2_17[106]},
      {stage3_17[55]}
   );
   gpc1_1 gpc3982 (
      {stage2_17[107]},
      {stage3_17[56]}
   );
   gpc1_1 gpc3983 (
      {stage2_17[108]},
      {stage3_17[57]}
   );
   gpc1_1 gpc3984 (
      {stage2_17[109]},
      {stage3_17[58]}
   );
   gpc1_1 gpc3985 (
      {stage2_17[110]},
      {stage3_17[59]}
   );
   gpc1_1 gpc3986 (
      {stage2_17[111]},
      {stage3_17[60]}
   );
   gpc1_1 gpc3987 (
      {stage2_17[112]},
      {stage3_17[61]}
   );
   gpc1_1 gpc3988 (
      {stage2_17[113]},
      {stage3_17[62]}
   );
   gpc1_1 gpc3989 (
      {stage2_17[114]},
      {stage3_17[63]}
   );
   gpc1_1 gpc3990 (
      {stage2_17[115]},
      {stage3_17[64]}
   );
   gpc1_1 gpc3991 (
      {stage2_17[116]},
      {stage3_17[65]}
   );
   gpc1_1 gpc3992 (
      {stage2_17[117]},
      {stage3_17[66]}
   );
   gpc1_1 gpc3993 (
      {stage2_17[118]},
      {stage3_17[67]}
   );
   gpc1_1 gpc3994 (
      {stage2_17[119]},
      {stage3_17[68]}
   );
   gpc1_1 gpc3995 (
      {stage2_17[120]},
      {stage3_17[69]}
   );
   gpc1_1 gpc3996 (
      {stage2_17[121]},
      {stage3_17[70]}
   );
   gpc1_1 gpc3997 (
      {stage2_17[122]},
      {stage3_17[71]}
   );
   gpc1_1 gpc3998 (
      {stage2_17[123]},
      {stage3_17[72]}
   );
   gpc1_1 gpc3999 (
      {stage2_17[124]},
      {stage3_17[73]}
   );
   gpc1_1 gpc4000 (
      {stage2_17[125]},
      {stage3_17[74]}
   );
   gpc1_1 gpc4001 (
      {stage2_17[126]},
      {stage3_17[75]}
   );
   gpc1_1 gpc4002 (
      {stage2_17[127]},
      {stage3_17[76]}
   );
   gpc1_1 gpc4003 (
      {stage2_19[64]},
      {stage3_19[36]}
   );
   gpc1_1 gpc4004 (
      {stage2_19[65]},
      {stage3_19[37]}
   );
   gpc1_1 gpc4005 (
      {stage2_19[66]},
      {stage3_19[38]}
   );
   gpc1_1 gpc4006 (
      {stage2_19[67]},
      {stage3_19[39]}
   );
   gpc1_1 gpc4007 (
      {stage2_19[68]},
      {stage3_19[40]}
   );
   gpc1_1 gpc4008 (
      {stage2_19[69]},
      {stage3_19[41]}
   );
   gpc1_1 gpc4009 (
      {stage2_19[70]},
      {stage3_19[42]}
   );
   gpc1_1 gpc4010 (
      {stage2_19[71]},
      {stage3_19[43]}
   );
   gpc1_1 gpc4011 (
      {stage2_19[72]},
      {stage3_19[44]}
   );
   gpc1_1 gpc4012 (
      {stage2_19[73]},
      {stage3_19[45]}
   );
   gpc1_1 gpc4013 (
      {stage2_19[74]},
      {stage3_19[46]}
   );
   gpc1_1 gpc4014 (
      {stage2_19[75]},
      {stage3_19[47]}
   );
   gpc1_1 gpc4015 (
      {stage2_19[76]},
      {stage3_19[48]}
   );
   gpc1_1 gpc4016 (
      {stage2_19[77]},
      {stage3_19[49]}
   );
   gpc1_1 gpc4017 (
      {stage2_19[78]},
      {stage3_19[50]}
   );
   gpc1_1 gpc4018 (
      {stage2_19[79]},
      {stage3_19[51]}
   );
   gpc1_1 gpc4019 (
      {stage2_19[80]},
      {stage3_19[52]}
   );
   gpc1_1 gpc4020 (
      {stage2_19[81]},
      {stage3_19[53]}
   );
   gpc1_1 gpc4021 (
      {stage2_19[82]},
      {stage3_19[54]}
   );
   gpc1_1 gpc4022 (
      {stage2_19[83]},
      {stage3_19[55]}
   );
   gpc1_1 gpc4023 (
      {stage2_19[84]},
      {stage3_19[56]}
   );
   gpc1_1 gpc4024 (
      {stage2_19[85]},
      {stage3_19[57]}
   );
   gpc1_1 gpc4025 (
      {stage2_19[86]},
      {stage3_19[58]}
   );
   gpc1_1 gpc4026 (
      {stage2_19[87]},
      {stage3_19[59]}
   );
   gpc1_1 gpc4027 (
      {stage2_19[88]},
      {stage3_19[60]}
   );
   gpc1_1 gpc4028 (
      {stage2_19[89]},
      {stage3_19[61]}
   );
   gpc1_1 gpc4029 (
      {stage2_19[90]},
      {stage3_19[62]}
   );
   gpc1_1 gpc4030 (
      {stage2_19[91]},
      {stage3_19[63]}
   );
   gpc1_1 gpc4031 (
      {stage2_19[92]},
      {stage3_19[64]}
   );
   gpc1_1 gpc4032 (
      {stage2_19[93]},
      {stage3_19[65]}
   );
   gpc1_1 gpc4033 (
      {stage2_19[94]},
      {stage3_19[66]}
   );
   gpc1_1 gpc4034 (
      {stage2_19[95]},
      {stage3_19[67]}
   );
   gpc1_1 gpc4035 (
      {stage2_19[96]},
      {stage3_19[68]}
   );
   gpc1_1 gpc4036 (
      {stage2_19[97]},
      {stage3_19[69]}
   );
   gpc1_1 gpc4037 (
      {stage2_21[96]},
      {stage3_21[34]}
   );
   gpc1_1 gpc4038 (
      {stage2_21[97]},
      {stage3_21[35]}
   );
   gpc1_1 gpc4039 (
      {stage2_21[98]},
      {stage3_21[36]}
   );
   gpc1_1 gpc4040 (
      {stage2_21[99]},
      {stage3_21[37]}
   );
   gpc1_1 gpc4041 (
      {stage2_21[100]},
      {stage3_21[38]}
   );
   gpc1_1 gpc4042 (
      {stage2_21[101]},
      {stage3_21[39]}
   );
   gpc1_1 gpc4043 (
      {stage2_21[102]},
      {stage3_21[40]}
   );
   gpc1_1 gpc4044 (
      {stage2_21[103]},
      {stage3_21[41]}
   );
   gpc1_1 gpc4045 (
      {stage2_21[104]},
      {stage3_21[42]}
   );
   gpc1_1 gpc4046 (
      {stage2_21[105]},
      {stage3_21[43]}
   );
   gpc1_1 gpc4047 (
      {stage2_21[106]},
      {stage3_21[44]}
   );
   gpc1_1 gpc4048 (
      {stage2_21[107]},
      {stage3_21[45]}
   );
   gpc1_1 gpc4049 (
      {stage2_21[108]},
      {stage3_21[46]}
   );
   gpc1_1 gpc4050 (
      {stage2_21[109]},
      {stage3_21[47]}
   );
   gpc1_1 gpc4051 (
      {stage2_21[110]},
      {stage3_21[48]}
   );
   gpc1_1 gpc4052 (
      {stage2_21[111]},
      {stage3_21[49]}
   );
   gpc1_1 gpc4053 (
      {stage2_21[112]},
      {stage3_21[50]}
   );
   gpc1_1 gpc4054 (
      {stage2_21[113]},
      {stage3_21[51]}
   );
   gpc1_1 gpc4055 (
      {stage2_21[114]},
      {stage3_21[52]}
   );
   gpc1_1 gpc4056 (
      {stage2_21[115]},
      {stage3_21[53]}
   );
   gpc1_1 gpc4057 (
      {stage2_21[116]},
      {stage3_21[54]}
   );
   gpc1_1 gpc4058 (
      {stage2_21[117]},
      {stage3_21[55]}
   );
   gpc1_1 gpc4059 (
      {stage2_21[118]},
      {stage3_21[56]}
   );
   gpc1_1 gpc4060 (
      {stage2_21[119]},
      {stage3_21[57]}
   );
   gpc1_1 gpc4061 (
      {stage2_21[120]},
      {stage3_21[58]}
   );
   gpc1_1 gpc4062 (
      {stage2_21[121]},
      {stage3_21[59]}
   );
   gpc1_1 gpc4063 (
      {stage2_21[122]},
      {stage3_21[60]}
   );
   gpc1_1 gpc4064 (
      {stage2_21[123]},
      {stage3_21[61]}
   );
   gpc1_1 gpc4065 (
      {stage2_21[124]},
      {stage3_21[62]}
   );
   gpc1_1 gpc4066 (
      {stage2_22[87]},
      {stage3_22[43]}
   );
   gpc1_1 gpc4067 (
      {stage2_22[88]},
      {stage3_22[44]}
   );
   gpc1_1 gpc4068 (
      {stage2_22[89]},
      {stage3_22[45]}
   );
   gpc1_1 gpc4069 (
      {stage2_22[90]},
      {stage3_22[46]}
   );
   gpc1_1 gpc4070 (
      {stage2_22[91]},
      {stage3_22[47]}
   );
   gpc1_1 gpc4071 (
      {stage2_22[92]},
      {stage3_22[48]}
   );
   gpc1_1 gpc4072 (
      {stage2_22[93]},
      {stage3_22[49]}
   );
   gpc1_1 gpc4073 (
      {stage2_22[94]},
      {stage3_22[50]}
   );
   gpc1_1 gpc4074 (
      {stage2_24[66]},
      {stage3_24[37]}
   );
   gpc1_1 gpc4075 (
      {stage2_24[67]},
      {stage3_24[38]}
   );
   gpc1_1 gpc4076 (
      {stage2_24[68]},
      {stage3_24[39]}
   );
   gpc1_1 gpc4077 (
      {stage2_24[69]},
      {stage3_24[40]}
   );
   gpc1_1 gpc4078 (
      {stage2_24[70]},
      {stage3_24[41]}
   );
   gpc1_1 gpc4079 (
      {stage2_24[71]},
      {stage3_24[42]}
   );
   gpc1_1 gpc4080 (
      {stage2_24[72]},
      {stage3_24[43]}
   );
   gpc1_1 gpc4081 (
      {stage2_24[73]},
      {stage3_24[44]}
   );
   gpc1_1 gpc4082 (
      {stage2_24[74]},
      {stage3_24[45]}
   );
   gpc1_1 gpc4083 (
      {stage2_24[75]},
      {stage3_24[46]}
   );
   gpc1_1 gpc4084 (
      {stage2_24[76]},
      {stage3_24[47]}
   );
   gpc1_1 gpc4085 (
      {stage2_24[77]},
      {stage3_24[48]}
   );
   gpc1_1 gpc4086 (
      {stage2_24[78]},
      {stage3_24[49]}
   );
   gpc1_1 gpc4087 (
      {stage2_24[79]},
      {stage3_24[50]}
   );
   gpc1_1 gpc4088 (
      {stage2_24[80]},
      {stage3_24[51]}
   );
   gpc1_1 gpc4089 (
      {stage2_24[81]},
      {stage3_24[52]}
   );
   gpc1_1 gpc4090 (
      {stage2_24[82]},
      {stage3_24[53]}
   );
   gpc1_1 gpc4091 (
      {stage2_24[83]},
      {stage3_24[54]}
   );
   gpc1_1 gpc4092 (
      {stage2_24[84]},
      {stage3_24[55]}
   );
   gpc1_1 gpc4093 (
      {stage2_24[85]},
      {stage3_24[56]}
   );
   gpc1_1 gpc4094 (
      {stage2_24[86]},
      {stage3_24[57]}
   );
   gpc1_1 gpc4095 (
      {stage2_24[87]},
      {stage3_24[58]}
   );
   gpc1_1 gpc4096 (
      {stage2_24[88]},
      {stage3_24[59]}
   );
   gpc1_1 gpc4097 (
      {stage2_24[89]},
      {stage3_24[60]}
   );
   gpc1_1 gpc4098 (
      {stage2_25[84]},
      {stage3_25[30]}
   );
   gpc1_1 gpc4099 (
      {stage2_25[85]},
      {stage3_25[31]}
   );
   gpc1_1 gpc4100 (
      {stage2_25[86]},
      {stage3_25[32]}
   );
   gpc1_1 gpc4101 (
      {stage2_25[87]},
      {stage3_25[33]}
   );
   gpc1_1 gpc4102 (
      {stage2_25[88]},
      {stage3_25[34]}
   );
   gpc1_1 gpc4103 (
      {stage2_25[89]},
      {stage3_25[35]}
   );
   gpc1_1 gpc4104 (
      {stage2_25[90]},
      {stage3_25[36]}
   );
   gpc1_1 gpc4105 (
      {stage2_25[91]},
      {stage3_25[37]}
   );
   gpc1_1 gpc4106 (
      {stage2_25[92]},
      {stage3_25[38]}
   );
   gpc1_1 gpc4107 (
      {stage2_25[93]},
      {stage3_25[39]}
   );
   gpc1_1 gpc4108 (
      {stage2_25[94]},
      {stage3_25[40]}
   );
   gpc1_1 gpc4109 (
      {stage2_25[95]},
      {stage3_25[41]}
   );
   gpc1_1 gpc4110 (
      {stage2_25[96]},
      {stage3_25[42]}
   );
   gpc1_1 gpc4111 (
      {stage2_25[97]},
      {stage3_25[43]}
   );
   gpc1_1 gpc4112 (
      {stage2_25[98]},
      {stage3_25[44]}
   );
   gpc1_1 gpc4113 (
      {stage2_25[99]},
      {stage3_25[45]}
   );
   gpc1_1 gpc4114 (
      {stage2_25[100]},
      {stage3_25[46]}
   );
   gpc1_1 gpc4115 (
      {stage2_25[101]},
      {stage3_25[47]}
   );
   gpc1_1 gpc4116 (
      {stage2_25[102]},
      {stage3_25[48]}
   );
   gpc1_1 gpc4117 (
      {stage2_26[87]},
      {stage3_26[38]}
   );
   gpc1_1 gpc4118 (
      {stage2_26[88]},
      {stage3_26[39]}
   );
   gpc1_1 gpc4119 (
      {stage2_26[89]},
      {stage3_26[40]}
   );
   gpc1_1 gpc4120 (
      {stage2_26[90]},
      {stage3_26[41]}
   );
   gpc1_1 gpc4121 (
      {stage2_26[91]},
      {stage3_26[42]}
   );
   gpc1_1 gpc4122 (
      {stage2_26[92]},
      {stage3_26[43]}
   );
   gpc1_1 gpc4123 (
      {stage2_26[93]},
      {stage3_26[44]}
   );
   gpc1_1 gpc4124 (
      {stage2_26[94]},
      {stage3_26[45]}
   );
   gpc1_1 gpc4125 (
      {stage2_26[95]},
      {stage3_26[46]}
   );
   gpc1_1 gpc4126 (
      {stage2_26[96]},
      {stage3_26[47]}
   );
   gpc1_1 gpc4127 (
      {stage2_26[97]},
      {stage3_26[48]}
   );
   gpc1_1 gpc4128 (
      {stage2_26[98]},
      {stage3_26[49]}
   );
   gpc1_1 gpc4129 (
      {stage2_26[99]},
      {stage3_26[50]}
   );
   gpc1_1 gpc4130 (
      {stage2_27[72]},
      {stage3_27[42]}
   );
   gpc1_1 gpc4131 (
      {stage2_27[73]},
      {stage3_27[43]}
   );
   gpc1_1 gpc4132 (
      {stage2_27[74]},
      {stage3_27[44]}
   );
   gpc1_1 gpc4133 (
      {stage2_27[75]},
      {stage3_27[45]}
   );
   gpc1_1 gpc4134 (
      {stage2_27[76]},
      {stage3_27[46]}
   );
   gpc1_1 gpc4135 (
      {stage2_27[77]},
      {stage3_27[47]}
   );
   gpc1_1 gpc4136 (
      {stage2_27[78]},
      {stage3_27[48]}
   );
   gpc1_1 gpc4137 (
      {stage2_27[79]},
      {stage3_27[49]}
   );
   gpc1_1 gpc4138 (
      {stage2_27[80]},
      {stage3_27[50]}
   );
   gpc1_1 gpc4139 (
      {stage2_27[81]},
      {stage3_27[51]}
   );
   gpc1_1 gpc4140 (
      {stage2_27[82]},
      {stage3_27[52]}
   );
   gpc1_1 gpc4141 (
      {stage2_27[83]},
      {stage3_27[53]}
   );
   gpc1_1 gpc4142 (
      {stage2_27[84]},
      {stage3_27[54]}
   );
   gpc1_1 gpc4143 (
      {stage2_28[133]},
      {stage3_28[36]}
   );
   gpc1_1 gpc4144 (
      {stage2_28[134]},
      {stage3_28[37]}
   );
   gpc1_1 gpc4145 (
      {stage2_28[135]},
      {stage3_28[38]}
   );
   gpc1_1 gpc4146 (
      {stage2_28[136]},
      {stage3_28[39]}
   );
   gpc1_1 gpc4147 (
      {stage2_28[137]},
      {stage3_28[40]}
   );
   gpc1_1 gpc4148 (
      {stage2_28[138]},
      {stage3_28[41]}
   );
   gpc1_1 gpc4149 (
      {stage2_28[139]},
      {stage3_28[42]}
   );
   gpc1_1 gpc4150 (
      {stage2_28[140]},
      {stage3_28[43]}
   );
   gpc1_1 gpc4151 (
      {stage2_28[141]},
      {stage3_28[44]}
   );
   gpc1_1 gpc4152 (
      {stage2_28[142]},
      {stage3_28[45]}
   );
   gpc1_1 gpc4153 (
      {stage2_28[143]},
      {stage3_28[46]}
   );
   gpc1_1 gpc4154 (
      {stage2_28[144]},
      {stage3_28[47]}
   );
   gpc1_1 gpc4155 (
      {stage2_28[145]},
      {stage3_28[48]}
   );
   gpc1_1 gpc4156 (
      {stage2_28[146]},
      {stage3_28[49]}
   );
   gpc1_1 gpc4157 (
      {stage2_28[147]},
      {stage3_28[50]}
   );
   gpc1_1 gpc4158 (
      {stage2_28[148]},
      {stage3_28[51]}
   );
   gpc1_1 gpc4159 (
      {stage2_28[149]},
      {stage3_28[52]}
   );
   gpc1_1 gpc4160 (
      {stage2_28[150]},
      {stage3_28[53]}
   );
   gpc1_1 gpc4161 (
      {stage2_28[151]},
      {stage3_28[54]}
   );
   gpc1_1 gpc4162 (
      {stage2_28[152]},
      {stage3_28[55]}
   );
   gpc1_1 gpc4163 (
      {stage2_28[153]},
      {stage3_28[56]}
   );
   gpc1_1 gpc4164 (
      {stage2_28[154]},
      {stage3_28[57]}
   );
   gpc1_1 gpc4165 (
      {stage2_28[155]},
      {stage3_28[58]}
   );
   gpc1_1 gpc4166 (
      {stage2_28[156]},
      {stage3_28[59]}
   );
   gpc1_1 gpc4167 (
      {stage2_28[157]},
      {stage3_28[60]}
   );
   gpc1_1 gpc4168 (
      {stage2_28[158]},
      {stage3_28[61]}
   );
   gpc1_1 gpc4169 (
      {stage2_28[159]},
      {stage3_28[62]}
   );
   gpc1_1 gpc4170 (
      {stage2_28[160]},
      {stage3_28[63]}
   );
   gpc1_1 gpc4171 (
      {stage2_28[161]},
      {stage3_28[64]}
   );
   gpc1_1 gpc4172 (
      {stage2_28[162]},
      {stage3_28[65]}
   );
   gpc1_1 gpc4173 (
      {stage2_28[163]},
      {stage3_28[66]}
   );
   gpc1_1 gpc4174 (
      {stage2_28[164]},
      {stage3_28[67]}
   );
   gpc1_1 gpc4175 (
      {stage2_28[165]},
      {stage3_28[68]}
   );
   gpc1_1 gpc4176 (
      {stage2_28[166]},
      {stage3_28[69]}
   );
   gpc1_1 gpc4177 (
      {stage2_28[167]},
      {stage3_28[70]}
   );
   gpc1_1 gpc4178 (
      {stage2_28[168]},
      {stage3_28[71]}
   );
   gpc1_1 gpc4179 (
      {stage2_28[169]},
      {stage3_28[72]}
   );
   gpc1_1 gpc4180 (
      {stage2_28[170]},
      {stage3_28[73]}
   );
   gpc1_1 gpc4181 (
      {stage2_29[127]},
      {stage3_29[42]}
   );
   gpc1_1 gpc4182 (
      {stage2_29[128]},
      {stage3_29[43]}
   );
   gpc1_1 gpc4183 (
      {stage2_29[129]},
      {stage3_29[44]}
   );
   gpc1_1 gpc4184 (
      {stage2_29[130]},
      {stage3_29[45]}
   );
   gpc1_1 gpc4185 (
      {stage2_29[131]},
      {stage3_29[46]}
   );
   gpc1_1 gpc4186 (
      {stage2_29[132]},
      {stage3_29[47]}
   );
   gpc1_1 gpc4187 (
      {stage2_29[133]},
      {stage3_29[48]}
   );
   gpc1_1 gpc4188 (
      {stage2_29[134]},
      {stage3_29[49]}
   );
   gpc1_1 gpc4189 (
      {stage2_29[135]},
      {stage3_29[50]}
   );
   gpc1_1 gpc4190 (
      {stage2_29[136]},
      {stage3_29[51]}
   );
   gpc1_1 gpc4191 (
      {stage2_29[137]},
      {stage3_29[52]}
   );
   gpc1_1 gpc4192 (
      {stage2_29[138]},
      {stage3_29[53]}
   );
   gpc1_1 gpc4193 (
      {stage2_29[139]},
      {stage3_29[54]}
   );
   gpc1_1 gpc4194 (
      {stage2_29[140]},
      {stage3_29[55]}
   );
   gpc1_1 gpc4195 (
      {stage2_29[141]},
      {stage3_29[56]}
   );
   gpc1_1 gpc4196 (
      {stage2_29[142]},
      {stage3_29[57]}
   );
   gpc1_1 gpc4197 (
      {stage2_30[66]},
      {stage3_30[45]}
   );
   gpc1_1 gpc4198 (
      {stage2_30[67]},
      {stage3_30[46]}
   );
   gpc1_1 gpc4199 (
      {stage2_30[68]},
      {stage3_30[47]}
   );
   gpc1_1 gpc4200 (
      {stage2_30[69]},
      {stage3_30[48]}
   );
   gpc1_1 gpc4201 (
      {stage2_30[70]},
      {stage3_30[49]}
   );
   gpc1_1 gpc4202 (
      {stage2_30[71]},
      {stage3_30[50]}
   );
   gpc1_1 gpc4203 (
      {stage2_30[72]},
      {stage3_30[51]}
   );
   gpc1_1 gpc4204 (
      {stage2_30[73]},
      {stage3_30[52]}
   );
   gpc1_1 gpc4205 (
      {stage2_30[74]},
      {stage3_30[53]}
   );
   gpc1_1 gpc4206 (
      {stage2_30[75]},
      {stage3_30[54]}
   );
   gpc1_1 gpc4207 (
      {stage2_30[76]},
      {stage3_30[55]}
   );
   gpc1_1 gpc4208 (
      {stage2_30[77]},
      {stage3_30[56]}
   );
   gpc1_1 gpc4209 (
      {stage2_30[78]},
      {stage3_30[57]}
   );
   gpc1_1 gpc4210 (
      {stage2_30[79]},
      {stage3_30[58]}
   );
   gpc1_1 gpc4211 (
      {stage2_30[80]},
      {stage3_30[59]}
   );
   gpc1_1 gpc4212 (
      {stage2_30[81]},
      {stage3_30[60]}
   );
   gpc1_1 gpc4213 (
      {stage2_30[82]},
      {stage3_30[61]}
   );
   gpc1_1 gpc4214 (
      {stage2_30[83]},
      {stage3_30[62]}
   );
   gpc1_1 gpc4215 (
      {stage2_30[84]},
      {stage3_30[63]}
   );
   gpc1_1 gpc4216 (
      {stage2_30[85]},
      {stage3_30[64]}
   );
   gpc1_1 gpc4217 (
      {stage2_30[86]},
      {stage3_30[65]}
   );
   gpc1_1 gpc4218 (
      {stage2_30[87]},
      {stage3_30[66]}
   );
   gpc1_1 gpc4219 (
      {stage2_30[88]},
      {stage3_30[67]}
   );
   gpc1_1 gpc4220 (
      {stage2_30[89]},
      {stage3_30[68]}
   );
   gpc1_1 gpc4221 (
      {stage2_30[90]},
      {stage3_30[69]}
   );
   gpc1_1 gpc4222 (
      {stage2_30[91]},
      {stage3_30[70]}
   );
   gpc1_1 gpc4223 (
      {stage2_31[83]},
      {stage3_31[39]}
   );
   gpc1_1 gpc4224 (
      {stage2_31[84]},
      {stage3_31[40]}
   );
   gpc1_1 gpc4225 (
      {stage2_31[85]},
      {stage3_31[41]}
   );
   gpc1_1 gpc4226 (
      {stage2_31[86]},
      {stage3_31[42]}
   );
   gpc1_1 gpc4227 (
      {stage2_31[87]},
      {stage3_31[43]}
   );
   gpc1_1 gpc4228 (
      {stage2_31[88]},
      {stage3_31[44]}
   );
   gpc1_1 gpc4229 (
      {stage2_31[89]},
      {stage3_31[45]}
   );
   gpc1_1 gpc4230 (
      {stage2_31[90]},
      {stage3_31[46]}
   );
   gpc1_1 gpc4231 (
      {stage2_31[91]},
      {stage3_31[47]}
   );
   gpc1_1 gpc4232 (
      {stage2_31[92]},
      {stage3_31[48]}
   );
   gpc1_1 gpc4233 (
      {stage2_31[93]},
      {stage3_31[49]}
   );
   gpc1_1 gpc4234 (
      {stage2_31[94]},
      {stage3_31[50]}
   );
   gpc1_1 gpc4235 (
      {stage2_31[95]},
      {stage3_31[51]}
   );
   gpc1_1 gpc4236 (
      {stage2_31[96]},
      {stage3_31[52]}
   );
   gpc1_1 gpc4237 (
      {stage2_31[97]},
      {stage3_31[53]}
   );
   gpc1_1 gpc4238 (
      {stage2_31[98]},
      {stage3_31[54]}
   );
   gpc1_1 gpc4239 (
      {stage2_31[99]},
      {stage3_31[55]}
   );
   gpc1_1 gpc4240 (
      {stage2_31[100]},
      {stage3_31[56]}
   );
   gpc1_1 gpc4241 (
      {stage2_31[101]},
      {stage3_31[57]}
   );
   gpc1_1 gpc4242 (
      {stage2_32[46]},
      {stage3_32[30]}
   );
   gpc1_1 gpc4243 (
      {stage2_32[47]},
      {stage3_32[31]}
   );
   gpc1_1 gpc4244 (
      {stage2_32[48]},
      {stage3_32[32]}
   );
   gpc1_1 gpc4245 (
      {stage2_32[49]},
      {stage3_32[33]}
   );
   gpc1_1 gpc4246 (
      {stage2_32[50]},
      {stage3_32[34]}
   );
   gpc1_1 gpc4247 (
      {stage2_32[51]},
      {stage3_32[35]}
   );
   gpc1_1 gpc4248 (
      {stage2_32[52]},
      {stage3_32[36]}
   );
   gpc1_1 gpc4249 (
      {stage2_32[53]},
      {stage3_32[37]}
   );
   gpc1_1 gpc4250 (
      {stage2_32[54]},
      {stage3_32[38]}
   );
   gpc1_1 gpc4251 (
      {stage2_32[55]},
      {stage3_32[39]}
   );
   gpc1_1 gpc4252 (
      {stage2_32[56]},
      {stage3_32[40]}
   );
   gpc1_1 gpc4253 (
      {stage2_32[57]},
      {stage3_32[41]}
   );
   gpc1_1 gpc4254 (
      {stage2_32[58]},
      {stage3_32[42]}
   );
   gpc1_1 gpc4255 (
      {stage2_32[59]},
      {stage3_32[43]}
   );
   gpc1_1 gpc4256 (
      {stage2_32[60]},
      {stage3_32[44]}
   );
   gpc1_1 gpc4257 (
      {stage2_32[61]},
      {stage3_32[45]}
   );
   gpc1_1 gpc4258 (
      {stage2_32[62]},
      {stage3_32[46]}
   );
   gpc1_1 gpc4259 (
      {stage2_32[63]},
      {stage3_32[47]}
   );
   gpc1_1 gpc4260 (
      {stage2_32[64]},
      {stage3_32[48]}
   );
   gpc1_1 gpc4261 (
      {stage2_32[65]},
      {stage3_32[49]}
   );
   gpc1_1 gpc4262 (
      {stage2_32[66]},
      {stage3_32[50]}
   );
   gpc1_1 gpc4263 (
      {stage2_32[67]},
      {stage3_32[51]}
   );
   gpc1_1 gpc4264 (
      {stage2_32[68]},
      {stage3_32[52]}
   );
   gpc1_1 gpc4265 (
      {stage2_32[69]},
      {stage3_32[53]}
   );
   gpc1_1 gpc4266 (
      {stage2_32[70]},
      {stage3_32[54]}
   );
   gpc1_1 gpc4267 (
      {stage2_32[71]},
      {stage3_32[55]}
   );
   gpc1_1 gpc4268 (
      {stage2_32[72]},
      {stage3_32[56]}
   );
   gpc1_1 gpc4269 (
      {stage2_32[73]},
      {stage3_32[57]}
   );
   gpc1_1 gpc4270 (
      {stage2_33[57]},
      {stage3_33[24]}
   );
   gpc1_1 gpc4271 (
      {stage2_33[58]},
      {stage3_33[25]}
   );
   gpc1_1 gpc4272 (
      {stage2_33[59]},
      {stage3_33[26]}
   );
   gpc1_1 gpc4273 (
      {stage2_34[24]},
      {stage3_34[16]}
   );
   gpc1_1 gpc4274 (
      {stage2_34[25]},
      {stage3_34[17]}
   );
   gpc1_1 gpc4275 (
      {stage2_34[26]},
      {stage3_34[18]}
   );
   gpc1_1 gpc4276 (
      {stage2_34[27]},
      {stage3_34[19]}
   );
   gpc1_1 gpc4277 (
      {stage2_34[28]},
      {stage3_34[20]}
   );
   gpc1_1 gpc4278 (
      {stage2_34[29]},
      {stage3_34[21]}
   );
   gpc1_1 gpc4279 (
      {stage2_34[30]},
      {stage3_34[22]}
   );
   gpc1_1 gpc4280 (
      {stage2_34[31]},
      {stage3_34[23]}
   );
   gpc1_1 gpc4281 (
      {stage2_34[32]},
      {stage3_34[24]}
   );
   gpc1_1 gpc4282 (
      {stage2_34[33]},
      {stage3_34[25]}
   );
   gpc1_1 gpc4283 (
      {stage2_34[34]},
      {stage3_34[26]}
   );
   gpc606_5 gpc4284 (
      {stage3_1[0], stage3_1[1], stage3_1[2], stage3_1[3], stage3_1[4], stage3_1[5]},
      {stage3_3[0], stage3_3[1], stage3_3[2], stage3_3[3], stage3_3[4], stage3_3[5]},
      {stage4_5[0],stage4_4[0],stage4_3[0],stage4_2[0],stage4_1[0]}
   );
   gpc606_5 gpc4285 (
      {stage3_1[6], stage3_1[7], stage3_1[8], stage3_1[9], stage3_1[10], stage3_1[11]},
      {stage3_3[6], stage3_3[7], stage3_3[8], stage3_3[9], stage3_3[10], stage3_3[11]},
      {stage4_5[1],stage4_4[1],stage4_3[1],stage4_2[1],stage4_1[1]}
   );
   gpc606_5 gpc4286 (
      {stage3_2[0], stage3_2[1], stage3_2[2], stage3_2[3], stage3_2[4], stage3_2[5]},
      {stage3_4[0], stage3_4[1], stage3_4[2], stage3_4[3], stage3_4[4], stage3_4[5]},
      {stage4_6[0],stage4_5[2],stage4_4[2],stage4_3[2],stage4_2[2]}
   );
   gpc606_5 gpc4287 (
      {stage3_2[6], stage3_2[7], stage3_2[8], stage3_2[9], stage3_2[10], stage3_2[11]},
      {stage3_4[6], stage3_4[7], stage3_4[8], stage3_4[9], stage3_4[10], stage3_4[11]},
      {stage4_6[1],stage4_5[3],stage4_4[3],stage4_3[3],stage4_2[3]}
   );
   gpc606_5 gpc4288 (
      {stage3_2[12], stage3_2[13], stage3_2[14], stage3_2[15], stage3_2[16], stage3_2[17]},
      {stage3_4[12], stage3_4[13], stage3_4[14], stage3_4[15], stage3_4[16], stage3_4[17]},
      {stage4_6[2],stage4_5[4],stage4_4[4],stage4_3[4],stage4_2[4]}
   );
   gpc606_5 gpc4289 (
      {stage3_2[18], stage3_2[19], stage3_2[20], stage3_2[21], stage3_2[22], stage3_2[23]},
      {stage3_4[18], stage3_4[19], stage3_4[20], stage3_4[21], stage3_4[22], stage3_4[23]},
      {stage4_6[3],stage4_5[5],stage4_4[5],stage4_3[5],stage4_2[5]}
   );
   gpc606_5 gpc4290 (
      {stage3_2[24], stage3_2[25], stage3_2[26], stage3_2[27], stage3_2[28], stage3_2[29]},
      {stage3_4[24], stage3_4[25], stage3_4[26], stage3_4[27], stage3_4[28], stage3_4[29]},
      {stage4_6[4],stage4_5[6],stage4_4[6],stage4_3[6],stage4_2[6]}
   );
   gpc606_5 gpc4291 (
      {stage3_5[0], stage3_5[1], stage3_5[2], stage3_5[3], stage3_5[4], stage3_5[5]},
      {stage3_7[0], stage3_7[1], stage3_7[2], stage3_7[3], stage3_7[4], stage3_7[5]},
      {stage4_9[0],stage4_8[0],stage4_7[0],stage4_6[5],stage4_5[7]}
   );
   gpc606_5 gpc4292 (
      {stage3_5[6], stage3_5[7], stage3_5[8], stage3_5[9], stage3_5[10], stage3_5[11]},
      {stage3_7[6], stage3_7[7], stage3_7[8], stage3_7[9], stage3_7[10], stage3_7[11]},
      {stage4_9[1],stage4_8[1],stage4_7[1],stage4_6[6],stage4_5[8]}
   );
   gpc606_5 gpc4293 (
      {stage3_5[12], stage3_5[13], stage3_5[14], stage3_5[15], stage3_5[16], stage3_5[17]},
      {stage3_7[12], stage3_7[13], stage3_7[14], stage3_7[15], stage3_7[16], stage3_7[17]},
      {stage4_9[2],stage4_8[2],stage4_7[2],stage4_6[7],stage4_5[9]}
   );
   gpc606_5 gpc4294 (
      {stage3_5[18], stage3_5[19], stage3_5[20], stage3_5[21], stage3_5[22], stage3_5[23]},
      {stage3_7[18], stage3_7[19], stage3_7[20], stage3_7[21], stage3_7[22], stage3_7[23]},
      {stage4_9[3],stage4_8[3],stage4_7[3],stage4_6[8],stage4_5[10]}
   );
   gpc615_5 gpc4295 (
      {stage3_6[0], stage3_6[1], stage3_6[2], stage3_6[3], stage3_6[4]},
      {stage3_7[24]},
      {stage3_8[0], stage3_8[1], stage3_8[2], stage3_8[3], stage3_8[4], stage3_8[5]},
      {stage4_10[0],stage4_9[4],stage4_8[4],stage4_7[4],stage4_6[9]}
   );
   gpc615_5 gpc4296 (
      {stage3_6[5], stage3_6[6], stage3_6[7], stage3_6[8], stage3_6[9]},
      {stage3_7[25]},
      {stage3_8[6], stage3_8[7], stage3_8[8], stage3_8[9], stage3_8[10], stage3_8[11]},
      {stage4_10[1],stage4_9[5],stage4_8[5],stage4_7[5],stage4_6[10]}
   );
   gpc615_5 gpc4297 (
      {stage3_6[10], stage3_6[11], stage3_6[12], stage3_6[13], stage3_6[14]},
      {stage3_7[26]},
      {stage3_8[12], stage3_8[13], stage3_8[14], stage3_8[15], stage3_8[16], stage3_8[17]},
      {stage4_10[2],stage4_9[6],stage4_8[6],stage4_7[6],stage4_6[11]}
   );
   gpc615_5 gpc4298 (
      {stage3_6[15], stage3_6[16], stage3_6[17], stage3_6[18], stage3_6[19]},
      {stage3_7[27]},
      {stage3_8[18], stage3_8[19], stage3_8[20], stage3_8[21], stage3_8[22], stage3_8[23]},
      {stage4_10[3],stage4_9[7],stage4_8[7],stage4_7[7],stage4_6[12]}
   );
   gpc615_5 gpc4299 (
      {stage3_6[20], stage3_6[21], stage3_6[22], stage3_6[23], stage3_6[24]},
      {stage3_7[28]},
      {stage3_8[24], stage3_8[25], stage3_8[26], stage3_8[27], stage3_8[28], stage3_8[29]},
      {stage4_10[4],stage4_9[8],stage4_8[8],stage4_7[8],stage4_6[13]}
   );
   gpc615_5 gpc4300 (
      {stage3_6[25], stage3_6[26], stage3_6[27], stage3_6[28], stage3_6[29]},
      {stage3_7[29]},
      {stage3_8[30], stage3_8[31], stage3_8[32], stage3_8[33], stage3_8[34], stage3_8[35]},
      {stage4_10[5],stage4_9[9],stage4_8[9],stage4_7[9],stage4_6[14]}
   );
   gpc615_5 gpc4301 (
      {stage3_7[30], stage3_7[31], stage3_7[32], stage3_7[33], stage3_7[34]},
      {stage3_8[36]},
      {stage3_9[0], stage3_9[1], stage3_9[2], stage3_9[3], stage3_9[4], stage3_9[5]},
      {stage4_11[0],stage4_10[6],stage4_9[10],stage4_8[10],stage4_7[10]}
   );
   gpc615_5 gpc4302 (
      {stage3_7[35], stage3_7[36], stage3_7[37], stage3_7[38], stage3_7[39]},
      {stage3_8[37]},
      {stage3_9[6], stage3_9[7], stage3_9[8], stage3_9[9], stage3_9[10], stage3_9[11]},
      {stage4_11[1],stage4_10[7],stage4_9[11],stage4_8[11],stage4_7[11]}
   );
   gpc615_5 gpc4303 (
      {stage3_7[40], stage3_7[41], stage3_7[42], stage3_7[43], stage3_7[44]},
      {stage3_8[38]},
      {stage3_9[12], stage3_9[13], stage3_9[14], stage3_9[15], stage3_9[16], stage3_9[17]},
      {stage4_11[2],stage4_10[8],stage4_9[12],stage4_8[12],stage4_7[12]}
   );
   gpc117_4 gpc4304 (
      {stage3_8[39], stage3_8[40], stage3_8[41], stage3_8[42], stage3_8[43], stage3_8[44], stage3_8[45]},
      {stage3_9[18]},
      {stage3_10[0]},
      {stage4_11[3],stage4_10[9],stage4_9[13],stage4_8[13]}
   );
   gpc117_4 gpc4305 (
      {stage3_8[46], stage3_8[47], stage3_8[48], stage3_8[49], stage3_8[50], stage3_8[51], stage3_8[52]},
      {stage3_9[19]},
      {stage3_10[1]},
      {stage4_11[4],stage4_10[10],stage4_9[14],stage4_8[14]}
   );
   gpc606_5 gpc4306 (
      {stage3_8[53], stage3_8[54], stage3_8[55], stage3_8[56], stage3_8[57], stage3_8[58]},
      {stage3_10[2], stage3_10[3], stage3_10[4], stage3_10[5], stage3_10[6], stage3_10[7]},
      {stage4_12[0],stage4_11[5],stage4_10[11],stage4_9[15],stage4_8[15]}
   );
   gpc606_5 gpc4307 (
      {stage3_8[59], stage3_8[60], stage3_8[61], stage3_8[62], stage3_8[63], stage3_8[64]},
      {stage3_10[8], stage3_10[9], stage3_10[10], stage3_10[11], stage3_10[12], stage3_10[13]},
      {stage4_12[1],stage4_11[6],stage4_10[12],stage4_9[16],stage4_8[16]}
   );
   gpc615_5 gpc4308 (
      {stage3_8[65], stage3_8[66], stage3_8[67], stage3_8[68], stage3_8[69]},
      {stage3_9[20]},
      {stage3_10[14], stage3_10[15], stage3_10[16], stage3_10[17], stage3_10[18], stage3_10[19]},
      {stage4_12[2],stage4_11[7],stage4_10[13],stage4_9[17],stage4_8[17]}
   );
   gpc615_5 gpc4309 (
      {stage3_8[70], stage3_8[71], stage3_8[72], stage3_8[73], stage3_8[74]},
      {stage3_9[21]},
      {stage3_10[20], stage3_10[21], stage3_10[22], stage3_10[23], stage3_10[24], stage3_10[25]},
      {stage4_12[3],stage4_11[8],stage4_10[14],stage4_9[18],stage4_8[18]}
   );
   gpc615_5 gpc4310 (
      {stage3_8[75], stage3_8[76], stage3_8[77], stage3_8[78], stage3_8[79]},
      {stage3_9[22]},
      {stage3_10[26], stage3_10[27], stage3_10[28], stage3_10[29], stage3_10[30], stage3_10[31]},
      {stage4_12[4],stage4_11[9],stage4_10[15],stage4_9[19],stage4_8[19]}
   );
   gpc615_5 gpc4311 (
      {stage3_8[80], stage3_8[81], stage3_8[82], stage3_8[83], stage3_8[84]},
      {stage3_9[23]},
      {stage3_10[32], stage3_10[33], stage3_10[34], stage3_10[35], stage3_10[36], stage3_10[37]},
      {stage4_12[5],stage4_11[10],stage4_10[16],stage4_9[20],stage4_8[20]}
   );
   gpc606_5 gpc4312 (
      {stage3_9[24], stage3_9[25], stage3_9[26], stage3_9[27], stage3_9[28], stage3_9[29]},
      {stage3_11[0], stage3_11[1], stage3_11[2], stage3_11[3], stage3_11[4], stage3_11[5]},
      {stage4_13[0],stage4_12[6],stage4_11[11],stage4_10[17],stage4_9[21]}
   );
   gpc1163_5 gpc4313 (
      {stage3_11[6], stage3_11[7], stage3_11[8]},
      {stage3_12[0], stage3_12[1], stage3_12[2], stage3_12[3], stage3_12[4], stage3_12[5]},
      {stage3_13[0]},
      {stage3_14[0]},
      {stage4_15[0],stage4_14[0],stage4_13[1],stage4_12[7],stage4_11[12]}
   );
   gpc1163_5 gpc4314 (
      {stage3_11[9], stage3_11[10], stage3_11[11]},
      {stage3_12[6], stage3_12[7], stage3_12[8], stage3_12[9], stage3_12[10], stage3_12[11]},
      {stage3_13[1]},
      {stage3_14[1]},
      {stage4_15[1],stage4_14[1],stage4_13[2],stage4_12[8],stage4_11[13]}
   );
   gpc1163_5 gpc4315 (
      {stage3_11[12], stage3_11[13], stage3_11[14]},
      {stage3_12[12], stage3_12[13], stage3_12[14], stage3_12[15], stage3_12[16], stage3_12[17]},
      {stage3_13[2]},
      {stage3_14[2]},
      {stage4_15[2],stage4_14[2],stage4_13[3],stage4_12[9],stage4_11[14]}
   );
   gpc1163_5 gpc4316 (
      {stage3_11[15], stage3_11[16], stage3_11[17]},
      {stage3_12[18], stage3_12[19], stage3_12[20], stage3_12[21], stage3_12[22], stage3_12[23]},
      {stage3_13[3]},
      {stage3_14[3]},
      {stage4_15[3],stage4_14[3],stage4_13[4],stage4_12[10],stage4_11[15]}
   );
   gpc1163_5 gpc4317 (
      {stage3_11[18], stage3_11[19], stage3_11[20]},
      {stage3_12[24], stage3_12[25], stage3_12[26], stage3_12[27], stage3_12[28], stage3_12[29]},
      {stage3_13[4]},
      {stage3_14[4]},
      {stage4_15[4],stage4_14[4],stage4_13[5],stage4_12[11],stage4_11[16]}
   );
   gpc615_5 gpc4318 (
      {stage3_11[21], stage3_11[22], stage3_11[23], stage3_11[24], stage3_11[25]},
      {stage3_12[30]},
      {stage3_13[5], stage3_13[6], stage3_13[7], stage3_13[8], stage3_13[9], stage3_13[10]},
      {stage4_15[5],stage4_14[5],stage4_13[6],stage4_12[12],stage4_11[17]}
   );
   gpc615_5 gpc4319 (
      {stage3_11[26], stage3_11[27], stage3_11[28], stage3_11[29], stage3_11[30]},
      {stage3_12[31]},
      {stage3_13[11], stage3_13[12], stage3_13[13], stage3_13[14], stage3_13[15], stage3_13[16]},
      {stage4_15[6],stage4_14[6],stage4_13[7],stage4_12[13],stage4_11[18]}
   );
   gpc606_5 gpc4320 (
      {stage3_12[32], stage3_12[33], stage3_12[34], stage3_12[35], stage3_12[36], stage3_12[37]},
      {stage3_14[5], stage3_14[6], stage3_14[7], stage3_14[8], stage3_14[9], stage3_14[10]},
      {stage4_16[0],stage4_15[7],stage4_14[7],stage4_13[8],stage4_12[14]}
   );
   gpc606_5 gpc4321 (
      {stage3_13[17], stage3_13[18], stage3_13[19], stage3_13[20], stage3_13[21], stage3_13[22]},
      {stage3_15[0], stage3_15[1], stage3_15[2], stage3_15[3], stage3_15[4], stage3_15[5]},
      {stage4_17[0],stage4_16[1],stage4_15[8],stage4_14[8],stage4_13[9]}
   );
   gpc606_5 gpc4322 (
      {stage3_13[23], stage3_13[24], stage3_13[25], stage3_13[26], stage3_13[27], stage3_13[28]},
      {stage3_15[6], stage3_15[7], stage3_15[8], stage3_15[9], stage3_15[10], stage3_15[11]},
      {stage4_17[1],stage4_16[2],stage4_15[9],stage4_14[9],stage4_13[10]}
   );
   gpc615_5 gpc4323 (
      {stage3_14[11], stage3_14[12], stage3_14[13], stage3_14[14], stage3_14[15]},
      {stage3_15[12]},
      {stage3_16[0], stage3_16[1], stage3_16[2], stage3_16[3], stage3_16[4], stage3_16[5]},
      {stage4_18[0],stage4_17[2],stage4_16[3],stage4_15[10],stage4_14[10]}
   );
   gpc615_5 gpc4324 (
      {stage3_14[16], stage3_14[17], stage3_14[18], stage3_14[19], stage3_14[20]},
      {stage3_15[13]},
      {stage3_16[6], stage3_16[7], stage3_16[8], stage3_16[9], stage3_16[10], stage3_16[11]},
      {stage4_18[1],stage4_17[3],stage4_16[4],stage4_15[11],stage4_14[11]}
   );
   gpc615_5 gpc4325 (
      {stage3_14[21], stage3_14[22], stage3_14[23], stage3_14[24], stage3_14[25]},
      {stage3_15[14]},
      {stage3_16[12], stage3_16[13], stage3_16[14], stage3_16[15], stage3_16[16], stage3_16[17]},
      {stage4_18[2],stage4_17[4],stage4_16[5],stage4_15[12],stage4_14[12]}
   );
   gpc615_5 gpc4326 (
      {stage3_14[26], stage3_14[27], stage3_14[28], stage3_14[29], stage3_14[30]},
      {stage3_15[15]},
      {stage3_16[18], stage3_16[19], stage3_16[20], stage3_16[21], stage3_16[22], stage3_16[23]},
      {stage4_18[3],stage4_17[5],stage4_16[6],stage4_15[13],stage4_14[13]}
   );
   gpc615_5 gpc4327 (
      {stage3_14[31], stage3_14[32], stage3_14[33], stage3_14[34], stage3_14[35]},
      {stage3_15[16]},
      {stage3_16[24], stage3_16[25], stage3_16[26], stage3_16[27], stage3_16[28], stage3_16[29]},
      {stage4_18[4],stage4_17[6],stage4_16[7],stage4_15[14],stage4_14[14]}
   );
   gpc1163_5 gpc4328 (
      {stage3_15[17], stage3_15[18], stage3_15[19]},
      {stage3_16[30], stage3_16[31], stage3_16[32], stage3_16[33], stage3_16[34], stage3_16[35]},
      {stage3_17[0]},
      {stage3_18[0]},
      {stage4_19[0],stage4_18[5],stage4_17[7],stage4_16[8],stage4_15[15]}
   );
   gpc615_5 gpc4329 (
      {stage3_15[20], stage3_15[21], stage3_15[22], stage3_15[23], stage3_15[24]},
      {stage3_16[36]},
      {stage3_17[1], stage3_17[2], stage3_17[3], stage3_17[4], stage3_17[5], stage3_17[6]},
      {stage4_19[1],stage4_18[6],stage4_17[8],stage4_16[9],stage4_15[16]}
   );
   gpc615_5 gpc4330 (
      {stage3_15[25], stage3_15[26], stage3_15[27], stage3_15[28], stage3_15[29]},
      {stage3_16[37]},
      {stage3_17[7], stage3_17[8], stage3_17[9], stage3_17[10], stage3_17[11], stage3_17[12]},
      {stage4_19[2],stage4_18[7],stage4_17[9],stage4_16[10],stage4_15[17]}
   );
   gpc615_5 gpc4331 (
      {stage3_15[30], stage3_15[31], stage3_15[32], stage3_15[33], stage3_15[34]},
      {stage3_16[38]},
      {stage3_17[13], stage3_17[14], stage3_17[15], stage3_17[16], stage3_17[17], stage3_17[18]},
      {stage4_19[3],stage4_18[8],stage4_17[10],stage4_16[11],stage4_15[18]}
   );
   gpc615_5 gpc4332 (
      {stage3_15[35], stage3_15[36], stage3_15[37], stage3_15[38], stage3_15[39]},
      {stage3_16[39]},
      {stage3_17[19], stage3_17[20], stage3_17[21], stage3_17[22], stage3_17[23], stage3_17[24]},
      {stage4_19[4],stage4_18[9],stage4_17[11],stage4_16[12],stage4_15[19]}
   );
   gpc615_5 gpc4333 (
      {stage3_15[40], stage3_15[41], stage3_15[42], stage3_15[43], stage3_15[44]},
      {stage3_16[40]},
      {stage3_17[25], stage3_17[26], stage3_17[27], stage3_17[28], stage3_17[29], stage3_17[30]},
      {stage4_19[5],stage4_18[10],stage4_17[12],stage4_16[13],stage4_15[20]}
   );
   gpc615_5 gpc4334 (
      {stage3_15[45], stage3_15[46], stage3_15[47], stage3_15[48], stage3_15[49]},
      {stage3_16[41]},
      {stage3_17[31], stage3_17[32], stage3_17[33], stage3_17[34], stage3_17[35], stage3_17[36]},
      {stage4_19[6],stage4_18[11],stage4_17[13],stage4_16[14],stage4_15[21]}
   );
   gpc615_5 gpc4335 (
      {stage3_15[50], stage3_15[51], stage3_15[52], stage3_15[53], stage3_15[54]},
      {stage3_16[42]},
      {stage3_17[37], stage3_17[38], stage3_17[39], stage3_17[40], stage3_17[41], stage3_17[42]},
      {stage4_19[7],stage4_18[12],stage4_17[14],stage4_16[15],stage4_15[22]}
   );
   gpc606_5 gpc4336 (
      {stage3_16[43], stage3_16[44], stage3_16[45], stage3_16[46], stage3_16[47], stage3_16[48]},
      {stage3_18[1], stage3_18[2], stage3_18[3], stage3_18[4], stage3_18[5], stage3_18[6]},
      {stage4_20[0],stage4_19[8],stage4_18[13],stage4_17[15],stage4_16[16]}
   );
   gpc606_5 gpc4337 (
      {stage3_16[49], stage3_16[50], stage3_16[51], stage3_16[52], stage3_16[53], stage3_16[54]},
      {stage3_18[7], stage3_18[8], stage3_18[9], stage3_18[10], stage3_18[11], stage3_18[12]},
      {stage4_20[1],stage4_19[9],stage4_18[14],stage4_17[16],stage4_16[17]}
   );
   gpc606_5 gpc4338 (
      {stage3_16[55], stage3_16[56], stage3_16[57], stage3_16[58], stage3_16[59], stage3_16[60]},
      {stage3_18[13], stage3_18[14], stage3_18[15], stage3_18[16], stage3_18[17], stage3_18[18]},
      {stage4_20[2],stage4_19[10],stage4_18[15],stage4_17[17],stage4_16[18]}
   );
   gpc606_5 gpc4339 (
      {stage3_16[61], stage3_16[62], stage3_16[63], stage3_16[64], stage3_16[65], stage3_16[66]},
      {stage3_18[19], stage3_18[20], stage3_18[21], stage3_18[22], stage3_18[23], stage3_18[24]},
      {stage4_20[3],stage4_19[11],stage4_18[16],stage4_17[18],stage4_16[19]}
   );
   gpc606_5 gpc4340 (
      {stage3_17[43], stage3_17[44], stage3_17[45], stage3_17[46], stage3_17[47], stage3_17[48]},
      {stage3_19[0], stage3_19[1], stage3_19[2], stage3_19[3], stage3_19[4], stage3_19[5]},
      {stage4_21[0],stage4_20[4],stage4_19[12],stage4_18[17],stage4_17[19]}
   );
   gpc606_5 gpc4341 (
      {stage3_17[49], stage3_17[50], stage3_17[51], stage3_17[52], stage3_17[53], stage3_17[54]},
      {stage3_19[6], stage3_19[7], stage3_19[8], stage3_19[9], stage3_19[10], stage3_19[11]},
      {stage4_21[1],stage4_20[5],stage4_19[13],stage4_18[18],stage4_17[20]}
   );
   gpc615_5 gpc4342 (
      {stage3_19[12], stage3_19[13], stage3_19[14], stage3_19[15], stage3_19[16]},
      {stage3_20[0]},
      {stage3_21[0], stage3_21[1], stage3_21[2], stage3_21[3], stage3_21[4], stage3_21[5]},
      {stage4_23[0],stage4_22[0],stage4_21[2],stage4_20[6],stage4_19[14]}
   );
   gpc615_5 gpc4343 (
      {stage3_19[17], stage3_19[18], stage3_19[19], stage3_19[20], stage3_19[21]},
      {stage3_20[1]},
      {stage3_21[6], stage3_21[7], stage3_21[8], stage3_21[9], stage3_21[10], stage3_21[11]},
      {stage4_23[1],stage4_22[1],stage4_21[3],stage4_20[7],stage4_19[15]}
   );
   gpc615_5 gpc4344 (
      {stage3_19[22], stage3_19[23], stage3_19[24], stage3_19[25], stage3_19[26]},
      {stage3_20[2]},
      {stage3_21[12], stage3_21[13], stage3_21[14], stage3_21[15], stage3_21[16], stage3_21[17]},
      {stage4_23[2],stage4_22[2],stage4_21[4],stage4_20[8],stage4_19[16]}
   );
   gpc615_5 gpc4345 (
      {stage3_19[27], stage3_19[28], stage3_19[29], stage3_19[30], stage3_19[31]},
      {stage3_20[3]},
      {stage3_21[18], stage3_21[19], stage3_21[20], stage3_21[21], stage3_21[22], stage3_21[23]},
      {stage4_23[3],stage4_22[3],stage4_21[5],stage4_20[9],stage4_19[17]}
   );
   gpc615_5 gpc4346 (
      {stage3_19[32], stage3_19[33], stage3_19[34], stage3_19[35], stage3_19[36]},
      {stage3_20[4]},
      {stage3_21[24], stage3_21[25], stage3_21[26], stage3_21[27], stage3_21[28], stage3_21[29]},
      {stage4_23[4],stage4_22[4],stage4_21[6],stage4_20[10],stage4_19[18]}
   );
   gpc615_5 gpc4347 (
      {stage3_19[37], stage3_19[38], stage3_19[39], stage3_19[40], stage3_19[41]},
      {stage3_20[5]},
      {stage3_21[30], stage3_21[31], stage3_21[32], stage3_21[33], stage3_21[34], stage3_21[35]},
      {stage4_23[5],stage4_22[5],stage4_21[7],stage4_20[11],stage4_19[19]}
   );
   gpc615_5 gpc4348 (
      {stage3_19[42], stage3_19[43], stage3_19[44], stage3_19[45], stage3_19[46]},
      {stage3_20[6]},
      {stage3_21[36], stage3_21[37], stage3_21[38], stage3_21[39], stage3_21[40], stage3_21[41]},
      {stage4_23[6],stage4_22[6],stage4_21[8],stage4_20[12],stage4_19[20]}
   );
   gpc615_5 gpc4349 (
      {stage3_19[47], stage3_19[48], stage3_19[49], stage3_19[50], stage3_19[51]},
      {stage3_20[7]},
      {stage3_21[42], stage3_21[43], stage3_21[44], stage3_21[45], stage3_21[46], stage3_21[47]},
      {stage4_23[7],stage4_22[7],stage4_21[9],stage4_20[13],stage4_19[21]}
   );
   gpc1325_5 gpc4350 (
      {stage3_19[52], stage3_19[53], stage3_19[54], stage3_19[55], stage3_19[56]},
      {stage3_20[8], stage3_20[9]},
      {stage3_21[48], stage3_21[49], stage3_21[50]},
      {stage3_22[0]},
      {stage4_23[8],stage4_22[8],stage4_21[10],stage4_20[14],stage4_19[22]}
   );
   gpc1325_5 gpc4351 (
      {stage3_19[57], stage3_19[58], stage3_19[59], stage3_19[60], stage3_19[61]},
      {stage3_20[10], stage3_20[11]},
      {stage3_21[51], stage3_21[52], stage3_21[53]},
      {stage3_22[1]},
      {stage4_23[9],stage4_22[9],stage4_21[11],stage4_20[15],stage4_19[23]}
   );
   gpc606_5 gpc4352 (
      {stage3_20[12], stage3_20[13], stage3_20[14], stage3_20[15], stage3_20[16], stage3_20[17]},
      {stage3_22[2], stage3_22[3], stage3_22[4], stage3_22[5], stage3_22[6], stage3_22[7]},
      {stage4_24[0],stage4_23[10],stage4_22[10],stage4_21[12],stage4_20[16]}
   );
   gpc606_5 gpc4353 (
      {stage3_20[18], stage3_20[19], stage3_20[20], stage3_20[21], stage3_20[22], stage3_20[23]},
      {stage3_22[8], stage3_22[9], stage3_22[10], stage3_22[11], stage3_22[12], stage3_22[13]},
      {stage4_24[1],stage4_23[11],stage4_22[11],stage4_21[13],stage4_20[17]}
   );
   gpc606_5 gpc4354 (
      {stage3_20[24], stage3_20[25], stage3_20[26], stage3_20[27], stage3_20[28], stage3_20[29]},
      {stage3_22[14], stage3_22[15], stage3_22[16], stage3_22[17], stage3_22[18], stage3_22[19]},
      {stage4_24[2],stage4_23[12],stage4_22[12],stage4_21[14],stage4_20[18]}
   );
   gpc606_5 gpc4355 (
      {stage3_21[54], stage3_21[55], stage3_21[56], stage3_21[57], stage3_21[58], stage3_21[59]},
      {stage3_23[0], stage3_23[1], stage3_23[2], stage3_23[3], stage3_23[4], stage3_23[5]},
      {stage4_25[0],stage4_24[3],stage4_23[13],stage4_22[13],stage4_21[15]}
   );
   gpc207_4 gpc4356 (
      {stage3_22[20], stage3_22[21], stage3_22[22], stage3_22[23], stage3_22[24], stage3_22[25], stage3_22[26]},
      {stage3_24[0], stage3_24[1]},
      {stage4_25[1],stage4_24[4],stage4_23[14],stage4_22[14]}
   );
   gpc615_5 gpc4357 (
      {stage3_22[27], stage3_22[28], stage3_22[29], stage3_22[30], stage3_22[31]},
      {stage3_23[6]},
      {stage3_24[2], stage3_24[3], stage3_24[4], stage3_24[5], stage3_24[6], stage3_24[7]},
      {stage4_26[0],stage4_25[2],stage4_24[5],stage4_23[15],stage4_22[15]}
   );
   gpc615_5 gpc4358 (
      {stage3_22[32], stage3_22[33], stage3_22[34], stage3_22[35], stage3_22[36]},
      {stage3_23[7]},
      {stage3_24[8], stage3_24[9], stage3_24[10], stage3_24[11], stage3_24[12], stage3_24[13]},
      {stage4_26[1],stage4_25[3],stage4_24[6],stage4_23[16],stage4_22[16]}
   );
   gpc606_5 gpc4359 (
      {stage3_23[8], stage3_23[9], stage3_23[10], stage3_23[11], stage3_23[12], stage3_23[13]},
      {stage3_25[0], stage3_25[1], stage3_25[2], stage3_25[3], stage3_25[4], stage3_25[5]},
      {stage4_27[0],stage4_26[2],stage4_25[4],stage4_24[7],stage4_23[17]}
   );
   gpc615_5 gpc4360 (
      {stage3_23[14], stage3_23[15], stage3_23[16], stage3_23[17], stage3_23[18]},
      {stage3_24[14]},
      {stage3_25[6], stage3_25[7], stage3_25[8], stage3_25[9], stage3_25[10], stage3_25[11]},
      {stage4_27[1],stage4_26[3],stage4_25[5],stage4_24[8],stage4_23[18]}
   );
   gpc615_5 gpc4361 (
      {stage3_23[19], stage3_23[20], stage3_23[21], stage3_23[22], stage3_23[23]},
      {stage3_24[15]},
      {stage3_25[12], stage3_25[13], stage3_25[14], stage3_25[15], stage3_25[16], stage3_25[17]},
      {stage4_27[2],stage4_26[4],stage4_25[6],stage4_24[9],stage4_23[19]}
   );
   gpc615_5 gpc4362 (
      {stage3_23[24], stage3_23[25], stage3_23[26], stage3_23[27], stage3_23[28]},
      {stage3_24[16]},
      {stage3_25[18], stage3_25[19], stage3_25[20], stage3_25[21], stage3_25[22], stage3_25[23]},
      {stage4_27[3],stage4_26[5],stage4_25[7],stage4_24[10],stage4_23[20]}
   );
   gpc606_5 gpc4363 (
      {stage3_24[17], stage3_24[18], stage3_24[19], stage3_24[20], stage3_24[21], stage3_24[22]},
      {stage3_26[0], stage3_26[1], stage3_26[2], stage3_26[3], stage3_26[4], stage3_26[5]},
      {stage4_28[0],stage4_27[4],stage4_26[6],stage4_25[8],stage4_24[11]}
   );
   gpc606_5 gpc4364 (
      {stage3_24[23], stage3_24[24], stage3_24[25], stage3_24[26], stage3_24[27], stage3_24[28]},
      {stage3_26[6], stage3_26[7], stage3_26[8], stage3_26[9], stage3_26[10], stage3_26[11]},
      {stage4_28[1],stage4_27[5],stage4_26[7],stage4_25[9],stage4_24[12]}
   );
   gpc606_5 gpc4365 (
      {stage3_24[29], stage3_24[30], stage3_24[31], stage3_24[32], stage3_24[33], stage3_24[34]},
      {stage3_26[12], stage3_26[13], stage3_26[14], stage3_26[15], stage3_26[16], stage3_26[17]},
      {stage4_28[2],stage4_27[6],stage4_26[8],stage4_25[10],stage4_24[13]}
   );
   gpc606_5 gpc4366 (
      {stage3_24[35], stage3_24[36], stage3_24[37], stage3_24[38], stage3_24[39], stage3_24[40]},
      {stage3_26[18], stage3_26[19], stage3_26[20], stage3_26[21], stage3_26[22], stage3_26[23]},
      {stage4_28[3],stage4_27[7],stage4_26[9],stage4_25[11],stage4_24[14]}
   );
   gpc606_5 gpc4367 (
      {stage3_24[41], stage3_24[42], stage3_24[43], stage3_24[44], stage3_24[45], stage3_24[46]},
      {stage3_26[24], stage3_26[25], stage3_26[26], stage3_26[27], stage3_26[28], stage3_26[29]},
      {stage4_28[4],stage4_27[8],stage4_26[10],stage4_25[12],stage4_24[15]}
   );
   gpc606_5 gpc4368 (
      {stage3_25[24], stage3_25[25], stage3_25[26], stage3_25[27], stage3_25[28], stage3_25[29]},
      {stage3_27[0], stage3_27[1], stage3_27[2], stage3_27[3], stage3_27[4], stage3_27[5]},
      {stage4_29[0],stage4_28[5],stage4_27[9],stage4_26[11],stage4_25[13]}
   );
   gpc606_5 gpc4369 (
      {stage3_25[30], stage3_25[31], stage3_25[32], stage3_25[33], stage3_25[34], stage3_25[35]},
      {stage3_27[6], stage3_27[7], stage3_27[8], stage3_27[9], stage3_27[10], stage3_27[11]},
      {stage4_29[1],stage4_28[6],stage4_27[10],stage4_26[12],stage4_25[14]}
   );
   gpc606_5 gpc4370 (
      {stage3_25[36], stage3_25[37], stage3_25[38], stage3_25[39], stage3_25[40], stage3_25[41]},
      {stage3_27[12], stage3_27[13], stage3_27[14], stage3_27[15], stage3_27[16], stage3_27[17]},
      {stage4_29[2],stage4_28[7],stage4_27[11],stage4_26[13],stage4_25[15]}
   );
   gpc615_5 gpc4371 (
      {stage3_25[42], stage3_25[43], stage3_25[44], stage3_25[45], stage3_25[46]},
      {stage3_26[30]},
      {stage3_27[18], stage3_27[19], stage3_27[20], stage3_27[21], stage3_27[22], stage3_27[23]},
      {stage4_29[3],stage4_28[8],stage4_27[12],stage4_26[14],stage4_25[16]}
   );
   gpc615_5 gpc4372 (
      {stage3_26[31], stage3_26[32], stage3_26[33], stage3_26[34], stage3_26[35]},
      {stage3_27[24]},
      {stage3_28[0], stage3_28[1], stage3_28[2], stage3_28[3], stage3_28[4], stage3_28[5]},
      {stage4_30[0],stage4_29[4],stage4_28[9],stage4_27[13],stage4_26[15]}
   );
   gpc615_5 gpc4373 (
      {stage3_26[36], stage3_26[37], stage3_26[38], stage3_26[39], stage3_26[40]},
      {stage3_27[25]},
      {stage3_28[6], stage3_28[7], stage3_28[8], stage3_28[9], stage3_28[10], stage3_28[11]},
      {stage4_30[1],stage4_29[5],stage4_28[10],stage4_27[14],stage4_26[16]}
   );
   gpc615_5 gpc4374 (
      {stage3_26[41], stage3_26[42], stage3_26[43], stage3_26[44], stage3_26[45]},
      {stage3_27[26]},
      {stage3_28[12], stage3_28[13], stage3_28[14], stage3_28[15], stage3_28[16], stage3_28[17]},
      {stage4_30[2],stage4_29[6],stage4_28[11],stage4_27[15],stage4_26[17]}
   );
   gpc606_5 gpc4375 (
      {stage3_27[27], stage3_27[28], stage3_27[29], stage3_27[30], stage3_27[31], stage3_27[32]},
      {stage3_29[0], stage3_29[1], stage3_29[2], stage3_29[3], stage3_29[4], stage3_29[5]},
      {stage4_31[0],stage4_30[3],stage4_29[7],stage4_28[12],stage4_27[16]}
   );
   gpc615_5 gpc4376 (
      {stage3_27[33], stage3_27[34], stage3_27[35], stage3_27[36], stage3_27[37]},
      {stage3_28[18]},
      {stage3_29[6], stage3_29[7], stage3_29[8], stage3_29[9], stage3_29[10], stage3_29[11]},
      {stage4_31[1],stage4_30[4],stage4_29[8],stage4_28[13],stage4_27[17]}
   );
   gpc615_5 gpc4377 (
      {stage3_27[38], stage3_27[39], stage3_27[40], stage3_27[41], stage3_27[42]},
      {stage3_28[19]},
      {stage3_29[12], stage3_29[13], stage3_29[14], stage3_29[15], stage3_29[16], stage3_29[17]},
      {stage4_31[2],stage4_30[5],stage4_29[9],stage4_28[14],stage4_27[18]}
   );
   gpc615_5 gpc4378 (
      {stage3_27[43], stage3_27[44], stage3_27[45], stage3_27[46], stage3_27[47]},
      {stage3_28[20]},
      {stage3_29[18], stage3_29[19], stage3_29[20], stage3_29[21], stage3_29[22], stage3_29[23]},
      {stage4_31[3],stage4_30[6],stage4_29[10],stage4_28[15],stage4_27[19]}
   );
   gpc606_5 gpc4379 (
      {stage3_28[21], stage3_28[22], stage3_28[23], stage3_28[24], stage3_28[25], stage3_28[26]},
      {stage3_30[0], stage3_30[1], stage3_30[2], stage3_30[3], stage3_30[4], stage3_30[5]},
      {stage4_32[0],stage4_31[4],stage4_30[7],stage4_29[11],stage4_28[16]}
   );
   gpc606_5 gpc4380 (
      {stage3_28[27], stage3_28[28], stage3_28[29], stage3_28[30], stage3_28[31], stage3_28[32]},
      {stage3_30[6], stage3_30[7], stage3_30[8], stage3_30[9], stage3_30[10], stage3_30[11]},
      {stage4_32[1],stage4_31[5],stage4_30[8],stage4_29[12],stage4_28[17]}
   );
   gpc606_5 gpc4381 (
      {stage3_28[33], stage3_28[34], stage3_28[35], stage3_28[36], stage3_28[37], stage3_28[38]},
      {stage3_30[12], stage3_30[13], stage3_30[14], stage3_30[15], stage3_30[16], stage3_30[17]},
      {stage4_32[2],stage4_31[6],stage4_30[9],stage4_29[13],stage4_28[18]}
   );
   gpc606_5 gpc4382 (
      {stage3_28[39], stage3_28[40], stage3_28[41], stage3_28[42], stage3_28[43], stage3_28[44]},
      {stage3_30[18], stage3_30[19], stage3_30[20], stage3_30[21], stage3_30[22], stage3_30[23]},
      {stage4_32[3],stage4_31[7],stage4_30[10],stage4_29[14],stage4_28[19]}
   );
   gpc606_5 gpc4383 (
      {stage3_28[45], stage3_28[46], stage3_28[47], stage3_28[48], stage3_28[49], stage3_28[50]},
      {stage3_30[24], stage3_30[25], stage3_30[26], stage3_30[27], stage3_30[28], stage3_30[29]},
      {stage4_32[4],stage4_31[8],stage4_30[11],stage4_29[15],stage4_28[20]}
   );
   gpc606_5 gpc4384 (
      {stage3_28[51], stage3_28[52], stage3_28[53], stage3_28[54], stage3_28[55], stage3_28[56]},
      {stage3_30[30], stage3_30[31], stage3_30[32], stage3_30[33], stage3_30[34], stage3_30[35]},
      {stage4_32[5],stage4_31[9],stage4_30[12],stage4_29[16],stage4_28[21]}
   );
   gpc606_5 gpc4385 (
      {stage3_28[57], stage3_28[58], stage3_28[59], stage3_28[60], stage3_28[61], stage3_28[62]},
      {stage3_30[36], stage3_30[37], stage3_30[38], stage3_30[39], stage3_30[40], stage3_30[41]},
      {stage4_32[6],stage4_31[10],stage4_30[13],stage4_29[17],stage4_28[22]}
   );
   gpc606_5 gpc4386 (
      {stage3_28[63], stage3_28[64], stage3_28[65], stage3_28[66], stage3_28[67], stage3_28[68]},
      {stage3_30[42], stage3_30[43], stage3_30[44], stage3_30[45], stage3_30[46], stage3_30[47]},
      {stage4_32[7],stage4_31[11],stage4_30[14],stage4_29[18],stage4_28[23]}
   );
   gpc606_5 gpc4387 (
      {stage3_28[69], stage3_28[70], stage3_28[71], stage3_28[72], stage3_28[73], 1'b0},
      {stage3_30[48], stage3_30[49], stage3_30[50], stage3_30[51], stage3_30[52], stage3_30[53]},
      {stage4_32[8],stage4_31[12],stage4_30[15],stage4_29[19],stage4_28[24]}
   );
   gpc606_5 gpc4388 (
      {stage3_29[24], stage3_29[25], stage3_29[26], stage3_29[27], stage3_29[28], stage3_29[29]},
      {stage3_31[0], stage3_31[1], stage3_31[2], stage3_31[3], stage3_31[4], stage3_31[5]},
      {stage4_33[0],stage4_32[9],stage4_31[13],stage4_30[16],stage4_29[20]}
   );
   gpc606_5 gpc4389 (
      {stage3_29[30], stage3_29[31], stage3_29[32], stage3_29[33], stage3_29[34], stage3_29[35]},
      {stage3_31[6], stage3_31[7], stage3_31[8], stage3_31[9], stage3_31[10], stage3_31[11]},
      {stage4_33[1],stage4_32[10],stage4_31[14],stage4_30[17],stage4_29[21]}
   );
   gpc606_5 gpc4390 (
      {stage3_29[36], stage3_29[37], stage3_29[38], stage3_29[39], stage3_29[40], stage3_29[41]},
      {stage3_31[12], stage3_31[13], stage3_31[14], stage3_31[15], stage3_31[16], stage3_31[17]},
      {stage4_33[2],stage4_32[11],stage4_31[15],stage4_30[18],stage4_29[22]}
   );
   gpc606_5 gpc4391 (
      {stage3_29[42], stage3_29[43], stage3_29[44], stage3_29[45], stage3_29[46], stage3_29[47]},
      {stage3_31[18], stage3_31[19], stage3_31[20], stage3_31[21], stage3_31[22], stage3_31[23]},
      {stage4_33[3],stage4_32[12],stage4_31[16],stage4_30[19],stage4_29[23]}
   );
   gpc615_5 gpc4392 (
      {stage3_29[48], stage3_29[49], stage3_29[50], stage3_29[51], stage3_29[52]},
      {stage3_30[54]},
      {stage3_31[24], stage3_31[25], stage3_31[26], stage3_31[27], stage3_31[28], stage3_31[29]},
      {stage4_33[4],stage4_32[13],stage4_31[17],stage4_30[20],stage4_29[24]}
   );
   gpc615_5 gpc4393 (
      {stage3_29[53], stage3_29[54], stage3_29[55], stage3_29[56], stage3_29[57]},
      {stage3_30[55]},
      {stage3_31[30], stage3_31[31], stage3_31[32], stage3_31[33], stage3_31[34], stage3_31[35]},
      {stage4_33[5],stage4_32[14],stage4_31[18],stage4_30[21],stage4_29[25]}
   );
   gpc606_5 gpc4394 (
      {stage3_30[56], stage3_30[57], stage3_30[58], stage3_30[59], stage3_30[60], stage3_30[61]},
      {stage3_32[0], stage3_32[1], stage3_32[2], stage3_32[3], stage3_32[4], stage3_32[5]},
      {stage4_34[0],stage4_33[6],stage4_32[15],stage4_31[19],stage4_30[22]}
   );
   gpc606_5 gpc4395 (
      {stage3_30[62], stage3_30[63], stage3_30[64], stage3_30[65], stage3_30[66], stage3_30[67]},
      {stage3_32[6], stage3_32[7], stage3_32[8], stage3_32[9], stage3_32[10], stage3_32[11]},
      {stage4_34[1],stage4_33[7],stage4_32[16],stage4_31[20],stage4_30[23]}
   );
   gpc615_5 gpc4396 (
      {stage3_31[36], stage3_31[37], stage3_31[38], stage3_31[39], stage3_31[40]},
      {stage3_32[12]},
      {stage3_33[0], stage3_33[1], stage3_33[2], stage3_33[3], stage3_33[4], stage3_33[5]},
      {stage4_35[0],stage4_34[2],stage4_33[8],stage4_32[17],stage4_31[21]}
   );
   gpc615_5 gpc4397 (
      {stage3_31[41], stage3_31[42], stage3_31[43], stage3_31[44], stage3_31[45]},
      {stage3_32[13]},
      {stage3_33[6], stage3_33[7], stage3_33[8], stage3_33[9], stage3_33[10], stage3_33[11]},
      {stage4_35[1],stage4_34[3],stage4_33[9],stage4_32[18],stage4_31[22]}
   );
   gpc615_5 gpc4398 (
      {stage3_31[46], stage3_31[47], stage3_31[48], stage3_31[49], stage3_31[50]},
      {stage3_32[14]},
      {stage3_33[12], stage3_33[13], stage3_33[14], stage3_33[15], stage3_33[16], stage3_33[17]},
      {stage4_35[2],stage4_34[4],stage4_33[10],stage4_32[19],stage4_31[23]}
   );
   gpc606_5 gpc4399 (
      {stage3_32[15], stage3_32[16], stage3_32[17], stage3_32[18], stage3_32[19], stage3_32[20]},
      {stage3_34[0], stage3_34[1], stage3_34[2], stage3_34[3], stage3_34[4], stage3_34[5]},
      {stage4_36[0],stage4_35[3],stage4_34[5],stage4_33[11],stage4_32[20]}
   );
   gpc606_5 gpc4400 (
      {stage3_32[21], stage3_32[22], stage3_32[23], stage3_32[24], stage3_32[25], stage3_32[26]},
      {stage3_34[6], stage3_34[7], stage3_34[8], stage3_34[9], stage3_34[10], stage3_34[11]},
      {stage4_36[1],stage4_35[4],stage4_34[6],stage4_33[12],stage4_32[21]}
   );
   gpc606_5 gpc4401 (
      {stage3_32[27], stage3_32[28], stage3_32[29], stage3_32[30], stage3_32[31], stage3_32[32]},
      {stage3_34[12], stage3_34[13], stage3_34[14], stage3_34[15], stage3_34[16], stage3_34[17]},
      {stage4_36[2],stage4_35[5],stage4_34[7],stage4_33[13],stage4_32[22]}
   );
   gpc606_5 gpc4402 (
      {stage3_32[33], stage3_32[34], stage3_32[35], stage3_32[36], stage3_32[37], stage3_32[38]},
      {stage3_34[18], stage3_34[19], stage3_34[20], stage3_34[21], stage3_34[22], stage3_34[23]},
      {stage4_36[3],stage4_35[6],stage4_34[8],stage4_33[14],stage4_32[23]}
   );
   gpc606_5 gpc4403 (
      {stage3_33[18], stage3_33[19], stage3_33[20], stage3_33[21], stage3_33[22], stage3_33[23]},
      {stage3_35[0], stage3_35[1], stage3_35[2], stage3_35[3], stage3_35[4], stage3_35[5]},
      {stage4_37[0],stage4_36[4],stage4_35[7],stage4_34[9],stage4_33[15]}
   );
   gpc1_1 gpc4404 (
      {stage3_0[0]},
      {stage4_0[0]}
   );
   gpc1_1 gpc4405 (
      {stage3_0[1]},
      {stage4_0[1]}
   );
   gpc1_1 gpc4406 (
      {stage3_0[2]},
      {stage4_0[2]}
   );
   gpc1_1 gpc4407 (
      {stage3_0[3]},
      {stage4_0[3]}
   );
   gpc1_1 gpc4408 (
      {stage3_0[4]},
      {stage4_0[4]}
   );
   gpc1_1 gpc4409 (
      {stage3_0[5]},
      {stage4_0[5]}
   );
   gpc1_1 gpc4410 (
      {stage3_0[6]},
      {stage4_0[6]}
   );
   gpc1_1 gpc4411 (
      {stage3_0[7]},
      {stage4_0[7]}
   );
   gpc1_1 gpc4412 (
      {stage3_0[8]},
      {stage4_0[8]}
   );
   gpc1_1 gpc4413 (
      {stage3_0[9]},
      {stage4_0[9]}
   );
   gpc1_1 gpc4414 (
      {stage3_0[10]},
      {stage4_0[10]}
   );
   gpc1_1 gpc4415 (
      {stage3_1[12]},
      {stage4_1[2]}
   );
   gpc1_1 gpc4416 (
      {stage3_1[13]},
      {stage4_1[3]}
   );
   gpc1_1 gpc4417 (
      {stage3_1[14]},
      {stage4_1[4]}
   );
   gpc1_1 gpc4418 (
      {stage3_1[15]},
      {stage4_1[5]}
   );
   gpc1_1 gpc4419 (
      {stage3_1[16]},
      {stage4_1[6]}
   );
   gpc1_1 gpc4420 (
      {stage3_1[17]},
      {stage4_1[7]}
   );
   gpc1_1 gpc4421 (
      {stage3_1[18]},
      {stage4_1[8]}
   );
   gpc1_1 gpc4422 (
      {stage3_1[19]},
      {stage4_1[9]}
   );
   gpc1_1 gpc4423 (
      {stage3_1[20]},
      {stage4_1[10]}
   );
   gpc1_1 gpc4424 (
      {stage3_1[21]},
      {stage4_1[11]}
   );
   gpc1_1 gpc4425 (
      {stage3_1[22]},
      {stage4_1[12]}
   );
   gpc1_1 gpc4426 (
      {stage3_1[23]},
      {stage4_1[13]}
   );
   gpc1_1 gpc4427 (
      {stage3_1[24]},
      {stage4_1[14]}
   );
   gpc1_1 gpc4428 (
      {stage3_1[25]},
      {stage4_1[15]}
   );
   gpc1_1 gpc4429 (
      {stage3_2[30]},
      {stage4_2[7]}
   );
   gpc1_1 gpc4430 (
      {stage3_2[31]},
      {stage4_2[8]}
   );
   gpc1_1 gpc4431 (
      {stage3_2[32]},
      {stage4_2[9]}
   );
   gpc1_1 gpc4432 (
      {stage3_2[33]},
      {stage4_2[10]}
   );
   gpc1_1 gpc4433 (
      {stage3_2[34]},
      {stage4_2[11]}
   );
   gpc1_1 gpc4434 (
      {stage3_2[35]},
      {stage4_2[12]}
   );
   gpc1_1 gpc4435 (
      {stage3_3[12]},
      {stage4_3[7]}
   );
   gpc1_1 gpc4436 (
      {stage3_3[13]},
      {stage4_3[8]}
   );
   gpc1_1 gpc4437 (
      {stage3_3[14]},
      {stage4_3[9]}
   );
   gpc1_1 gpc4438 (
      {stage3_3[15]},
      {stage4_3[10]}
   );
   gpc1_1 gpc4439 (
      {stage3_3[16]},
      {stage4_3[11]}
   );
   gpc1_1 gpc4440 (
      {stage3_3[17]},
      {stage4_3[12]}
   );
   gpc1_1 gpc4441 (
      {stage3_3[18]},
      {stage4_3[13]}
   );
   gpc1_1 gpc4442 (
      {stage3_3[19]},
      {stage4_3[14]}
   );
   gpc1_1 gpc4443 (
      {stage3_3[20]},
      {stage4_3[15]}
   );
   gpc1_1 gpc4444 (
      {stage3_3[21]},
      {stage4_3[16]}
   );
   gpc1_1 gpc4445 (
      {stage3_3[22]},
      {stage4_3[17]}
   );
   gpc1_1 gpc4446 (
      {stage3_3[23]},
      {stage4_3[18]}
   );
   gpc1_1 gpc4447 (
      {stage3_3[24]},
      {stage4_3[19]}
   );
   gpc1_1 gpc4448 (
      {stage3_3[25]},
      {stage4_3[20]}
   );
   gpc1_1 gpc4449 (
      {stage3_3[26]},
      {stage4_3[21]}
   );
   gpc1_1 gpc4450 (
      {stage3_3[27]},
      {stage4_3[22]}
   );
   gpc1_1 gpc4451 (
      {stage3_4[30]},
      {stage4_4[7]}
   );
   gpc1_1 gpc4452 (
      {stage3_4[31]},
      {stage4_4[8]}
   );
   gpc1_1 gpc4453 (
      {stage3_4[32]},
      {stage4_4[9]}
   );
   gpc1_1 gpc4454 (
      {stage3_4[33]},
      {stage4_4[10]}
   );
   gpc1_1 gpc4455 (
      {stage3_4[34]},
      {stage4_4[11]}
   );
   gpc1_1 gpc4456 (
      {stage3_4[35]},
      {stage4_4[12]}
   );
   gpc1_1 gpc4457 (
      {stage3_4[36]},
      {stage4_4[13]}
   );
   gpc1_1 gpc4458 (
      {stage3_4[37]},
      {stage4_4[14]}
   );
   gpc1_1 gpc4459 (
      {stage3_4[38]},
      {stage4_4[15]}
   );
   gpc1_1 gpc4460 (
      {stage3_4[39]},
      {stage4_4[16]}
   );
   gpc1_1 gpc4461 (
      {stage3_4[40]},
      {stage4_4[17]}
   );
   gpc1_1 gpc4462 (
      {stage3_4[41]},
      {stage4_4[18]}
   );
   gpc1_1 gpc4463 (
      {stage3_4[42]},
      {stage4_4[19]}
   );
   gpc1_1 gpc4464 (
      {stage3_4[43]},
      {stage4_4[20]}
   );
   gpc1_1 gpc4465 (
      {stage3_4[44]},
      {stage4_4[21]}
   );
   gpc1_1 gpc4466 (
      {stage3_4[45]},
      {stage4_4[22]}
   );
   gpc1_1 gpc4467 (
      {stage3_4[46]},
      {stage4_4[23]}
   );
   gpc1_1 gpc4468 (
      {stage3_5[24]},
      {stage4_5[11]}
   );
   gpc1_1 gpc4469 (
      {stage3_5[25]},
      {stage4_5[12]}
   );
   gpc1_1 gpc4470 (
      {stage3_5[26]},
      {stage4_5[13]}
   );
   gpc1_1 gpc4471 (
      {stage3_5[27]},
      {stage4_5[14]}
   );
   gpc1_1 gpc4472 (
      {stage3_5[28]},
      {stage4_5[15]}
   );
   gpc1_1 gpc4473 (
      {stage3_5[29]},
      {stage4_5[16]}
   );
   gpc1_1 gpc4474 (
      {stage3_5[30]},
      {stage4_5[17]}
   );
   gpc1_1 gpc4475 (
      {stage3_5[31]},
      {stage4_5[18]}
   );
   gpc1_1 gpc4476 (
      {stage3_5[32]},
      {stage4_5[19]}
   );
   gpc1_1 gpc4477 (
      {stage3_5[33]},
      {stage4_5[20]}
   );
   gpc1_1 gpc4478 (
      {stage3_5[34]},
      {stage4_5[21]}
   );
   gpc1_1 gpc4479 (
      {stage3_5[35]},
      {stage4_5[22]}
   );
   gpc1_1 gpc4480 (
      {stage3_5[36]},
      {stage4_5[23]}
   );
   gpc1_1 gpc4481 (
      {stage3_5[37]},
      {stage4_5[24]}
   );
   gpc1_1 gpc4482 (
      {stage3_5[38]},
      {stage4_5[25]}
   );
   gpc1_1 gpc4483 (
      {stage3_5[39]},
      {stage4_5[26]}
   );
   gpc1_1 gpc4484 (
      {stage3_5[40]},
      {stage4_5[27]}
   );
   gpc1_1 gpc4485 (
      {stage3_5[41]},
      {stage4_5[28]}
   );
   gpc1_1 gpc4486 (
      {stage3_5[42]},
      {stage4_5[29]}
   );
   gpc1_1 gpc4487 (
      {stage3_5[43]},
      {stage4_5[30]}
   );
   gpc1_1 gpc4488 (
      {stage3_5[44]},
      {stage4_5[31]}
   );
   gpc1_1 gpc4489 (
      {stage3_5[45]},
      {stage4_5[32]}
   );
   gpc1_1 gpc4490 (
      {stage3_5[46]},
      {stage4_5[33]}
   );
   gpc1_1 gpc4491 (
      {stage3_5[47]},
      {stage4_5[34]}
   );
   gpc1_1 gpc4492 (
      {stage3_5[48]},
      {stage4_5[35]}
   );
   gpc1_1 gpc4493 (
      {stage3_5[49]},
      {stage4_5[36]}
   );
   gpc1_1 gpc4494 (
      {stage3_5[50]},
      {stage4_5[37]}
   );
   gpc1_1 gpc4495 (
      {stage3_5[51]},
      {stage4_5[38]}
   );
   gpc1_1 gpc4496 (
      {stage3_5[52]},
      {stage4_5[39]}
   );
   gpc1_1 gpc4497 (
      {stage3_5[53]},
      {stage4_5[40]}
   );
   gpc1_1 gpc4498 (
      {stage3_5[54]},
      {stage4_5[41]}
   );
   gpc1_1 gpc4499 (
      {stage3_5[55]},
      {stage4_5[42]}
   );
   gpc1_1 gpc4500 (
      {stage3_5[56]},
      {stage4_5[43]}
   );
   gpc1_1 gpc4501 (
      {stage3_5[57]},
      {stage4_5[44]}
   );
   gpc1_1 gpc4502 (
      {stage3_5[58]},
      {stage4_5[45]}
   );
   gpc1_1 gpc4503 (
      {stage3_6[30]},
      {stage4_6[15]}
   );
   gpc1_1 gpc4504 (
      {stage3_6[31]},
      {stage4_6[16]}
   );
   gpc1_1 gpc4505 (
      {stage3_6[32]},
      {stage4_6[17]}
   );
   gpc1_1 gpc4506 (
      {stage3_6[33]},
      {stage4_6[18]}
   );
   gpc1_1 gpc4507 (
      {stage3_6[34]},
      {stage4_6[19]}
   );
   gpc1_1 gpc4508 (
      {stage3_6[35]},
      {stage4_6[20]}
   );
   gpc1_1 gpc4509 (
      {stage3_6[36]},
      {stage4_6[21]}
   );
   gpc1_1 gpc4510 (
      {stage3_6[37]},
      {stage4_6[22]}
   );
   gpc1_1 gpc4511 (
      {stage3_7[45]},
      {stage4_7[13]}
   );
   gpc1_1 gpc4512 (
      {stage3_7[46]},
      {stage4_7[14]}
   );
   gpc1_1 gpc4513 (
      {stage3_8[85]},
      {stage4_8[21]}
   );
   gpc1_1 gpc4514 (
      {stage3_8[86]},
      {stage4_8[22]}
   );
   gpc1_1 gpc4515 (
      {stage3_8[87]},
      {stage4_8[23]}
   );
   gpc1_1 gpc4516 (
      {stage3_8[88]},
      {stage4_8[24]}
   );
   gpc1_1 gpc4517 (
      {stage3_8[89]},
      {stage4_8[25]}
   );
   gpc1_1 gpc4518 (
      {stage3_8[90]},
      {stage4_8[26]}
   );
   gpc1_1 gpc4519 (
      {stage3_8[91]},
      {stage4_8[27]}
   );
   gpc1_1 gpc4520 (
      {stage3_8[92]},
      {stage4_8[28]}
   );
   gpc1_1 gpc4521 (
      {stage3_9[30]},
      {stage4_9[22]}
   );
   gpc1_1 gpc4522 (
      {stage3_9[31]},
      {stage4_9[23]}
   );
   gpc1_1 gpc4523 (
      {stage3_9[32]},
      {stage4_9[24]}
   );
   gpc1_1 gpc4524 (
      {stage3_9[33]},
      {stage4_9[25]}
   );
   gpc1_1 gpc4525 (
      {stage3_9[34]},
      {stage4_9[26]}
   );
   gpc1_1 gpc4526 (
      {stage3_9[35]},
      {stage4_9[27]}
   );
   gpc1_1 gpc4527 (
      {stage3_9[36]},
      {stage4_9[28]}
   );
   gpc1_1 gpc4528 (
      {stage3_9[37]},
      {stage4_9[29]}
   );
   gpc1_1 gpc4529 (
      {stage3_9[38]},
      {stage4_9[30]}
   );
   gpc1_1 gpc4530 (
      {stage3_9[39]},
      {stage4_9[31]}
   );
   gpc1_1 gpc4531 (
      {stage3_9[40]},
      {stage4_9[32]}
   );
   gpc1_1 gpc4532 (
      {stage3_9[41]},
      {stage4_9[33]}
   );
   gpc1_1 gpc4533 (
      {stage3_9[42]},
      {stage4_9[34]}
   );
   gpc1_1 gpc4534 (
      {stage3_9[43]},
      {stage4_9[35]}
   );
   gpc1_1 gpc4535 (
      {stage3_9[44]},
      {stage4_9[36]}
   );
   gpc1_1 gpc4536 (
      {stage3_9[45]},
      {stage4_9[37]}
   );
   gpc1_1 gpc4537 (
      {stage3_9[46]},
      {stage4_9[38]}
   );
   gpc1_1 gpc4538 (
      {stage3_9[47]},
      {stage4_9[39]}
   );
   gpc1_1 gpc4539 (
      {stage3_9[48]},
      {stage4_9[40]}
   );
   gpc1_1 gpc4540 (
      {stage3_9[49]},
      {stage4_9[41]}
   );
   gpc1_1 gpc4541 (
      {stage3_11[31]},
      {stage4_11[19]}
   );
   gpc1_1 gpc4542 (
      {stage3_11[32]},
      {stage4_11[20]}
   );
   gpc1_1 gpc4543 (
      {stage3_11[33]},
      {stage4_11[21]}
   );
   gpc1_1 gpc4544 (
      {stage3_11[34]},
      {stage4_11[22]}
   );
   gpc1_1 gpc4545 (
      {stage3_11[35]},
      {stage4_11[23]}
   );
   gpc1_1 gpc4546 (
      {stage3_11[36]},
      {stage4_11[24]}
   );
   gpc1_1 gpc4547 (
      {stage3_11[37]},
      {stage4_11[25]}
   );
   gpc1_1 gpc4548 (
      {stage3_11[38]},
      {stage4_11[26]}
   );
   gpc1_1 gpc4549 (
      {stage3_11[39]},
      {stage4_11[27]}
   );
   gpc1_1 gpc4550 (
      {stage3_11[40]},
      {stage4_11[28]}
   );
   gpc1_1 gpc4551 (
      {stage3_11[41]},
      {stage4_11[29]}
   );
   gpc1_1 gpc4552 (
      {stage3_11[42]},
      {stage4_11[30]}
   );
   gpc1_1 gpc4553 (
      {stage3_11[43]},
      {stage4_11[31]}
   );
   gpc1_1 gpc4554 (
      {stage3_11[44]},
      {stage4_11[32]}
   );
   gpc1_1 gpc4555 (
      {stage3_11[45]},
      {stage4_11[33]}
   );
   gpc1_1 gpc4556 (
      {stage3_11[46]},
      {stage4_11[34]}
   );
   gpc1_1 gpc4557 (
      {stage3_11[47]},
      {stage4_11[35]}
   );
   gpc1_1 gpc4558 (
      {stage3_11[48]},
      {stage4_11[36]}
   );
   gpc1_1 gpc4559 (
      {stage3_11[49]},
      {stage4_11[37]}
   );
   gpc1_1 gpc4560 (
      {stage3_11[50]},
      {stage4_11[38]}
   );
   gpc1_1 gpc4561 (
      {stage3_11[51]},
      {stage4_11[39]}
   );
   gpc1_1 gpc4562 (
      {stage3_11[52]},
      {stage4_11[40]}
   );
   gpc1_1 gpc4563 (
      {stage3_11[53]},
      {stage4_11[41]}
   );
   gpc1_1 gpc4564 (
      {stage3_11[54]},
      {stage4_11[42]}
   );
   gpc1_1 gpc4565 (
      {stage3_12[38]},
      {stage4_12[15]}
   );
   gpc1_1 gpc4566 (
      {stage3_12[39]},
      {stage4_12[16]}
   );
   gpc1_1 gpc4567 (
      {stage3_12[40]},
      {stage4_12[17]}
   );
   gpc1_1 gpc4568 (
      {stage3_12[41]},
      {stage4_12[18]}
   );
   gpc1_1 gpc4569 (
      {stage3_12[42]},
      {stage4_12[19]}
   );
   gpc1_1 gpc4570 (
      {stage3_12[43]},
      {stage4_12[20]}
   );
   gpc1_1 gpc4571 (
      {stage3_12[44]},
      {stage4_12[21]}
   );
   gpc1_1 gpc4572 (
      {stage3_12[45]},
      {stage4_12[22]}
   );
   gpc1_1 gpc4573 (
      {stage3_12[46]},
      {stage4_12[23]}
   );
   gpc1_1 gpc4574 (
      {stage3_13[29]},
      {stage4_13[11]}
   );
   gpc1_1 gpc4575 (
      {stage3_13[30]},
      {stage4_13[12]}
   );
   gpc1_1 gpc4576 (
      {stage3_13[31]},
      {stage4_13[13]}
   );
   gpc1_1 gpc4577 (
      {stage3_13[32]},
      {stage4_13[14]}
   );
   gpc1_1 gpc4578 (
      {stage3_13[33]},
      {stage4_13[15]}
   );
   gpc1_1 gpc4579 (
      {stage3_13[34]},
      {stage4_13[16]}
   );
   gpc1_1 gpc4580 (
      {stage3_13[35]},
      {stage4_13[17]}
   );
   gpc1_1 gpc4581 (
      {stage3_13[36]},
      {stage4_13[18]}
   );
   gpc1_1 gpc4582 (
      {stage3_14[36]},
      {stage4_14[15]}
   );
   gpc1_1 gpc4583 (
      {stage3_14[37]},
      {stage4_14[16]}
   );
   gpc1_1 gpc4584 (
      {stage3_14[38]},
      {stage4_14[17]}
   );
   gpc1_1 gpc4585 (
      {stage3_14[39]},
      {stage4_14[18]}
   );
   gpc1_1 gpc4586 (
      {stage3_14[40]},
      {stage4_14[19]}
   );
   gpc1_1 gpc4587 (
      {stage3_14[41]},
      {stage4_14[20]}
   );
   gpc1_1 gpc4588 (
      {stage3_14[42]},
      {stage4_14[21]}
   );
   gpc1_1 gpc4589 (
      {stage3_14[43]},
      {stage4_14[22]}
   );
   gpc1_1 gpc4590 (
      {stage3_14[44]},
      {stage4_14[23]}
   );
   gpc1_1 gpc4591 (
      {stage3_14[45]},
      {stage4_14[24]}
   );
   gpc1_1 gpc4592 (
      {stage3_14[46]},
      {stage4_14[25]}
   );
   gpc1_1 gpc4593 (
      {stage3_14[47]},
      {stage4_14[26]}
   );
   gpc1_1 gpc4594 (
      {stage3_14[48]},
      {stage4_14[27]}
   );
   gpc1_1 gpc4595 (
      {stage3_14[49]},
      {stage4_14[28]}
   );
   gpc1_1 gpc4596 (
      {stage3_14[50]},
      {stage4_14[29]}
   );
   gpc1_1 gpc4597 (
      {stage3_14[51]},
      {stage4_14[30]}
   );
   gpc1_1 gpc4598 (
      {stage3_14[52]},
      {stage4_14[31]}
   );
   gpc1_1 gpc4599 (
      {stage3_14[53]},
      {stage4_14[32]}
   );
   gpc1_1 gpc4600 (
      {stage3_14[54]},
      {stage4_14[33]}
   );
   gpc1_1 gpc4601 (
      {stage3_14[55]},
      {stage4_14[34]}
   );
   gpc1_1 gpc4602 (
      {stage3_15[55]},
      {stage4_15[23]}
   );
   gpc1_1 gpc4603 (
      {stage3_15[56]},
      {stage4_15[24]}
   );
   gpc1_1 gpc4604 (
      {stage3_15[57]},
      {stage4_15[25]}
   );
   gpc1_1 gpc4605 (
      {stage3_15[58]},
      {stage4_15[26]}
   );
   gpc1_1 gpc4606 (
      {stage3_15[59]},
      {stage4_15[27]}
   );
   gpc1_1 gpc4607 (
      {stage3_15[60]},
      {stage4_15[28]}
   );
   gpc1_1 gpc4608 (
      {stage3_15[61]},
      {stage4_15[29]}
   );
   gpc1_1 gpc4609 (
      {stage3_15[62]},
      {stage4_15[30]}
   );
   gpc1_1 gpc4610 (
      {stage3_15[63]},
      {stage4_15[31]}
   );
   gpc1_1 gpc4611 (
      {stage3_15[64]},
      {stage4_15[32]}
   );
   gpc1_1 gpc4612 (
      {stage3_15[65]},
      {stage4_15[33]}
   );
   gpc1_1 gpc4613 (
      {stage3_15[66]},
      {stage4_15[34]}
   );
   gpc1_1 gpc4614 (
      {stage3_15[67]},
      {stage4_15[35]}
   );
   gpc1_1 gpc4615 (
      {stage3_15[68]},
      {stage4_15[36]}
   );
   gpc1_1 gpc4616 (
      {stage3_15[69]},
      {stage4_15[37]}
   );
   gpc1_1 gpc4617 (
      {stage3_15[70]},
      {stage4_15[38]}
   );
   gpc1_1 gpc4618 (
      {stage3_17[55]},
      {stage4_17[21]}
   );
   gpc1_1 gpc4619 (
      {stage3_17[56]},
      {stage4_17[22]}
   );
   gpc1_1 gpc4620 (
      {stage3_17[57]},
      {stage4_17[23]}
   );
   gpc1_1 gpc4621 (
      {stage3_17[58]},
      {stage4_17[24]}
   );
   gpc1_1 gpc4622 (
      {stage3_17[59]},
      {stage4_17[25]}
   );
   gpc1_1 gpc4623 (
      {stage3_17[60]},
      {stage4_17[26]}
   );
   gpc1_1 gpc4624 (
      {stage3_17[61]},
      {stage4_17[27]}
   );
   gpc1_1 gpc4625 (
      {stage3_17[62]},
      {stage4_17[28]}
   );
   gpc1_1 gpc4626 (
      {stage3_17[63]},
      {stage4_17[29]}
   );
   gpc1_1 gpc4627 (
      {stage3_17[64]},
      {stage4_17[30]}
   );
   gpc1_1 gpc4628 (
      {stage3_17[65]},
      {stage4_17[31]}
   );
   gpc1_1 gpc4629 (
      {stage3_17[66]},
      {stage4_17[32]}
   );
   gpc1_1 gpc4630 (
      {stage3_17[67]},
      {stage4_17[33]}
   );
   gpc1_1 gpc4631 (
      {stage3_17[68]},
      {stage4_17[34]}
   );
   gpc1_1 gpc4632 (
      {stage3_17[69]},
      {stage4_17[35]}
   );
   gpc1_1 gpc4633 (
      {stage3_17[70]},
      {stage4_17[36]}
   );
   gpc1_1 gpc4634 (
      {stage3_17[71]},
      {stage4_17[37]}
   );
   gpc1_1 gpc4635 (
      {stage3_17[72]},
      {stage4_17[38]}
   );
   gpc1_1 gpc4636 (
      {stage3_17[73]},
      {stage4_17[39]}
   );
   gpc1_1 gpc4637 (
      {stage3_17[74]},
      {stage4_17[40]}
   );
   gpc1_1 gpc4638 (
      {stage3_17[75]},
      {stage4_17[41]}
   );
   gpc1_1 gpc4639 (
      {stage3_17[76]},
      {stage4_17[42]}
   );
   gpc1_1 gpc4640 (
      {stage3_18[25]},
      {stage4_18[19]}
   );
   gpc1_1 gpc4641 (
      {stage3_18[26]},
      {stage4_18[20]}
   );
   gpc1_1 gpc4642 (
      {stage3_18[27]},
      {stage4_18[21]}
   );
   gpc1_1 gpc4643 (
      {stage3_18[28]},
      {stage4_18[22]}
   );
   gpc1_1 gpc4644 (
      {stage3_18[29]},
      {stage4_18[23]}
   );
   gpc1_1 gpc4645 (
      {stage3_18[30]},
      {stage4_18[24]}
   );
   gpc1_1 gpc4646 (
      {stage3_18[31]},
      {stage4_18[25]}
   );
   gpc1_1 gpc4647 (
      {stage3_18[32]},
      {stage4_18[26]}
   );
   gpc1_1 gpc4648 (
      {stage3_18[33]},
      {stage4_18[27]}
   );
   gpc1_1 gpc4649 (
      {stage3_18[34]},
      {stage4_18[28]}
   );
   gpc1_1 gpc4650 (
      {stage3_19[62]},
      {stage4_19[24]}
   );
   gpc1_1 gpc4651 (
      {stage3_19[63]},
      {stage4_19[25]}
   );
   gpc1_1 gpc4652 (
      {stage3_19[64]},
      {stage4_19[26]}
   );
   gpc1_1 gpc4653 (
      {stage3_19[65]},
      {stage4_19[27]}
   );
   gpc1_1 gpc4654 (
      {stage3_19[66]},
      {stage4_19[28]}
   );
   gpc1_1 gpc4655 (
      {stage3_19[67]},
      {stage4_19[29]}
   );
   gpc1_1 gpc4656 (
      {stage3_19[68]},
      {stage4_19[30]}
   );
   gpc1_1 gpc4657 (
      {stage3_19[69]},
      {stage4_19[31]}
   );
   gpc1_1 gpc4658 (
      {stage3_21[60]},
      {stage4_21[16]}
   );
   gpc1_1 gpc4659 (
      {stage3_21[61]},
      {stage4_21[17]}
   );
   gpc1_1 gpc4660 (
      {stage3_21[62]},
      {stage4_21[18]}
   );
   gpc1_1 gpc4661 (
      {stage3_22[37]},
      {stage4_22[17]}
   );
   gpc1_1 gpc4662 (
      {stage3_22[38]},
      {stage4_22[18]}
   );
   gpc1_1 gpc4663 (
      {stage3_22[39]},
      {stage4_22[19]}
   );
   gpc1_1 gpc4664 (
      {stage3_22[40]},
      {stage4_22[20]}
   );
   gpc1_1 gpc4665 (
      {stage3_22[41]},
      {stage4_22[21]}
   );
   gpc1_1 gpc4666 (
      {stage3_22[42]},
      {stage4_22[22]}
   );
   gpc1_1 gpc4667 (
      {stage3_22[43]},
      {stage4_22[23]}
   );
   gpc1_1 gpc4668 (
      {stage3_22[44]},
      {stage4_22[24]}
   );
   gpc1_1 gpc4669 (
      {stage3_22[45]},
      {stage4_22[25]}
   );
   gpc1_1 gpc4670 (
      {stage3_22[46]},
      {stage4_22[26]}
   );
   gpc1_1 gpc4671 (
      {stage3_22[47]},
      {stage4_22[27]}
   );
   gpc1_1 gpc4672 (
      {stage3_22[48]},
      {stage4_22[28]}
   );
   gpc1_1 gpc4673 (
      {stage3_22[49]},
      {stage4_22[29]}
   );
   gpc1_1 gpc4674 (
      {stage3_22[50]},
      {stage4_22[30]}
   );
   gpc1_1 gpc4675 (
      {stage3_23[29]},
      {stage4_23[21]}
   );
   gpc1_1 gpc4676 (
      {stage3_23[30]},
      {stage4_23[22]}
   );
   gpc1_1 gpc4677 (
      {stage3_23[31]},
      {stage4_23[23]}
   );
   gpc1_1 gpc4678 (
      {stage3_23[32]},
      {stage4_23[24]}
   );
   gpc1_1 gpc4679 (
      {stage3_23[33]},
      {stage4_23[25]}
   );
   gpc1_1 gpc4680 (
      {stage3_23[34]},
      {stage4_23[26]}
   );
   gpc1_1 gpc4681 (
      {stage3_23[35]},
      {stage4_23[27]}
   );
   gpc1_1 gpc4682 (
      {stage3_23[36]},
      {stage4_23[28]}
   );
   gpc1_1 gpc4683 (
      {stage3_23[37]},
      {stage4_23[29]}
   );
   gpc1_1 gpc4684 (
      {stage3_23[38]},
      {stage4_23[30]}
   );
   gpc1_1 gpc4685 (
      {stage3_23[39]},
      {stage4_23[31]}
   );
   gpc1_1 gpc4686 (
      {stage3_23[40]},
      {stage4_23[32]}
   );
   gpc1_1 gpc4687 (
      {stage3_23[41]},
      {stage4_23[33]}
   );
   gpc1_1 gpc4688 (
      {stage3_23[42]},
      {stage4_23[34]}
   );
   gpc1_1 gpc4689 (
      {stage3_23[43]},
      {stage4_23[35]}
   );
   gpc1_1 gpc4690 (
      {stage3_23[44]},
      {stage4_23[36]}
   );
   gpc1_1 gpc4691 (
      {stage3_23[45]},
      {stage4_23[37]}
   );
   gpc1_1 gpc4692 (
      {stage3_24[47]},
      {stage4_24[16]}
   );
   gpc1_1 gpc4693 (
      {stage3_24[48]},
      {stage4_24[17]}
   );
   gpc1_1 gpc4694 (
      {stage3_24[49]},
      {stage4_24[18]}
   );
   gpc1_1 gpc4695 (
      {stage3_24[50]},
      {stage4_24[19]}
   );
   gpc1_1 gpc4696 (
      {stage3_24[51]},
      {stage4_24[20]}
   );
   gpc1_1 gpc4697 (
      {stage3_24[52]},
      {stage4_24[21]}
   );
   gpc1_1 gpc4698 (
      {stage3_24[53]},
      {stage4_24[22]}
   );
   gpc1_1 gpc4699 (
      {stage3_24[54]},
      {stage4_24[23]}
   );
   gpc1_1 gpc4700 (
      {stage3_24[55]},
      {stage4_24[24]}
   );
   gpc1_1 gpc4701 (
      {stage3_24[56]},
      {stage4_24[25]}
   );
   gpc1_1 gpc4702 (
      {stage3_24[57]},
      {stage4_24[26]}
   );
   gpc1_1 gpc4703 (
      {stage3_24[58]},
      {stage4_24[27]}
   );
   gpc1_1 gpc4704 (
      {stage3_24[59]},
      {stage4_24[28]}
   );
   gpc1_1 gpc4705 (
      {stage3_24[60]},
      {stage4_24[29]}
   );
   gpc1_1 gpc4706 (
      {stage3_25[47]},
      {stage4_25[17]}
   );
   gpc1_1 gpc4707 (
      {stage3_25[48]},
      {stage4_25[18]}
   );
   gpc1_1 gpc4708 (
      {stage3_26[46]},
      {stage4_26[18]}
   );
   gpc1_1 gpc4709 (
      {stage3_26[47]},
      {stage4_26[19]}
   );
   gpc1_1 gpc4710 (
      {stage3_26[48]},
      {stage4_26[20]}
   );
   gpc1_1 gpc4711 (
      {stage3_26[49]},
      {stage4_26[21]}
   );
   gpc1_1 gpc4712 (
      {stage3_26[50]},
      {stage4_26[22]}
   );
   gpc1_1 gpc4713 (
      {stage3_27[48]},
      {stage4_27[20]}
   );
   gpc1_1 gpc4714 (
      {stage3_27[49]},
      {stage4_27[21]}
   );
   gpc1_1 gpc4715 (
      {stage3_27[50]},
      {stage4_27[22]}
   );
   gpc1_1 gpc4716 (
      {stage3_27[51]},
      {stage4_27[23]}
   );
   gpc1_1 gpc4717 (
      {stage3_27[52]},
      {stage4_27[24]}
   );
   gpc1_1 gpc4718 (
      {stage3_27[53]},
      {stage4_27[25]}
   );
   gpc1_1 gpc4719 (
      {stage3_27[54]},
      {stage4_27[26]}
   );
   gpc1_1 gpc4720 (
      {stage3_30[68]},
      {stage4_30[24]}
   );
   gpc1_1 gpc4721 (
      {stage3_30[69]},
      {stage4_30[25]}
   );
   gpc1_1 gpc4722 (
      {stage3_30[70]},
      {stage4_30[26]}
   );
   gpc1_1 gpc4723 (
      {stage3_31[51]},
      {stage4_31[24]}
   );
   gpc1_1 gpc4724 (
      {stage3_31[52]},
      {stage4_31[25]}
   );
   gpc1_1 gpc4725 (
      {stage3_31[53]},
      {stage4_31[26]}
   );
   gpc1_1 gpc4726 (
      {stage3_31[54]},
      {stage4_31[27]}
   );
   gpc1_1 gpc4727 (
      {stage3_31[55]},
      {stage4_31[28]}
   );
   gpc1_1 gpc4728 (
      {stage3_31[56]},
      {stage4_31[29]}
   );
   gpc1_1 gpc4729 (
      {stage3_31[57]},
      {stage4_31[30]}
   );
   gpc1_1 gpc4730 (
      {stage3_32[39]},
      {stage4_32[24]}
   );
   gpc1_1 gpc4731 (
      {stage3_32[40]},
      {stage4_32[25]}
   );
   gpc1_1 gpc4732 (
      {stage3_32[41]},
      {stage4_32[26]}
   );
   gpc1_1 gpc4733 (
      {stage3_32[42]},
      {stage4_32[27]}
   );
   gpc1_1 gpc4734 (
      {stage3_32[43]},
      {stage4_32[28]}
   );
   gpc1_1 gpc4735 (
      {stage3_32[44]},
      {stage4_32[29]}
   );
   gpc1_1 gpc4736 (
      {stage3_32[45]},
      {stage4_32[30]}
   );
   gpc1_1 gpc4737 (
      {stage3_32[46]},
      {stage4_32[31]}
   );
   gpc1_1 gpc4738 (
      {stage3_32[47]},
      {stage4_32[32]}
   );
   gpc1_1 gpc4739 (
      {stage3_32[48]},
      {stage4_32[33]}
   );
   gpc1_1 gpc4740 (
      {stage3_32[49]},
      {stage4_32[34]}
   );
   gpc1_1 gpc4741 (
      {stage3_32[50]},
      {stage4_32[35]}
   );
   gpc1_1 gpc4742 (
      {stage3_32[51]},
      {stage4_32[36]}
   );
   gpc1_1 gpc4743 (
      {stage3_32[52]},
      {stage4_32[37]}
   );
   gpc1_1 gpc4744 (
      {stage3_32[53]},
      {stage4_32[38]}
   );
   gpc1_1 gpc4745 (
      {stage3_32[54]},
      {stage4_32[39]}
   );
   gpc1_1 gpc4746 (
      {stage3_32[55]},
      {stage4_32[40]}
   );
   gpc1_1 gpc4747 (
      {stage3_32[56]},
      {stage4_32[41]}
   );
   gpc1_1 gpc4748 (
      {stage3_32[57]},
      {stage4_32[42]}
   );
   gpc1_1 gpc4749 (
      {stage3_33[24]},
      {stage4_33[16]}
   );
   gpc1_1 gpc4750 (
      {stage3_33[25]},
      {stage4_33[17]}
   );
   gpc1_1 gpc4751 (
      {stage3_33[26]},
      {stage4_33[18]}
   );
   gpc1_1 gpc4752 (
      {stage3_34[24]},
      {stage4_34[10]}
   );
   gpc1_1 gpc4753 (
      {stage3_34[25]},
      {stage4_34[11]}
   );
   gpc1_1 gpc4754 (
      {stage3_34[26]},
      {stage4_34[12]}
   );
   gpc1_1 gpc4755 (
      {stage3_35[6]},
      {stage4_35[8]}
   );
   gpc1_1 gpc4756 (
      {stage3_35[7]},
      {stage4_35[9]}
   );
   gpc1_1 gpc4757 (
      {stage3_35[8]},
      {stage4_35[10]}
   );
   gpc1_1 gpc4758 (
      {stage3_35[9]},
      {stage4_35[11]}
   );
   gpc1_1 gpc4759 (
      {stage3_35[10]},
      {stage4_35[12]}
   );
   gpc1_1 gpc4760 (
      {stage3_35[11]},
      {stage4_35[13]}
   );
   gpc1_1 gpc4761 (
      {stage3_35[12]},
      {stage4_35[14]}
   );
   gpc1_1 gpc4762 (
      {stage3_36[0]},
      {stage4_36[5]}
   );
   gpc1_1 gpc4763 (
      {stage3_36[1]},
      {stage4_36[6]}
   );
   gpc1_1 gpc4764 (
      {stage3_36[2]},
      {stage4_36[7]}
   );
   gpc1_1 gpc4765 (
      {stage3_36[3]},
      {stage4_36[8]}
   );
   gpc1_1 gpc4766 (
      {stage3_36[4]},
      {stage4_36[9]}
   );
   gpc1_1 gpc4767 (
      {stage3_36[5]},
      {stage4_36[10]}
   );
   gpc1_1 gpc4768 (
      {stage3_37[0]},
      {stage4_37[1]}
   );
   gpc1_1 gpc4769 (
      {stage3_37[1]},
      {stage4_37[2]}
   );
   gpc606_5 gpc4770 (
      {stage4_1[0], stage4_1[1], stage4_1[2], stage4_1[3], stage4_1[4], stage4_1[5]},
      {stage4_3[0], stage4_3[1], stage4_3[2], stage4_3[3], stage4_3[4], stage4_3[5]},
      {stage5_5[0],stage5_4[0],stage5_3[0],stage5_2[0],stage5_1[0]}
   );
   gpc615_5 gpc4771 (
      {stage4_2[0], stage4_2[1], stage4_2[2], stage4_2[3], stage4_2[4]},
      {stage4_3[6]},
      {stage4_4[0], stage4_4[1], stage4_4[2], stage4_4[3], stage4_4[4], stage4_4[5]},
      {stage5_6[0],stage5_5[1],stage5_4[1],stage5_3[1],stage5_2[1]}
   );
   gpc615_5 gpc4772 (
      {stage4_3[7], stage4_3[8], stage4_3[9], stage4_3[10], stage4_3[11]},
      {stage4_4[6]},
      {stage4_5[0], stage4_5[1], stage4_5[2], stage4_5[3], stage4_5[4], stage4_5[5]},
      {stage5_7[0],stage5_6[1],stage5_5[2],stage5_4[2],stage5_3[2]}
   );
   gpc615_5 gpc4773 (
      {stage4_3[12], stage4_3[13], stage4_3[14], stage4_3[15], stage4_3[16]},
      {stage4_4[7]},
      {stage4_5[6], stage4_5[7], stage4_5[8], stage4_5[9], stage4_5[10], stage4_5[11]},
      {stage5_7[1],stage5_6[2],stage5_5[3],stage5_4[3],stage5_3[3]}
   );
   gpc615_5 gpc4774 (
      {stage4_3[17], stage4_3[18], stage4_3[19], stage4_3[20], stage4_3[21]},
      {stage4_4[8]},
      {stage4_5[12], stage4_5[13], stage4_5[14], stage4_5[15], stage4_5[16], stage4_5[17]},
      {stage5_7[2],stage5_6[3],stage5_5[4],stage5_4[4],stage5_3[4]}
   );
   gpc606_5 gpc4775 (
      {stage4_4[9], stage4_4[10], stage4_4[11], stage4_4[12], stage4_4[13], stage4_4[14]},
      {stage4_6[0], stage4_6[1], stage4_6[2], stage4_6[3], stage4_6[4], stage4_6[5]},
      {stage5_8[0],stage5_7[3],stage5_6[4],stage5_5[5],stage5_4[5]}
   );
   gpc606_5 gpc4776 (
      {stage4_4[15], stage4_4[16], stage4_4[17], stage4_4[18], stage4_4[19], stage4_4[20]},
      {stage4_6[6], stage4_6[7], stage4_6[8], stage4_6[9], stage4_6[10], stage4_6[11]},
      {stage5_8[1],stage5_7[4],stage5_6[5],stage5_5[6],stage5_4[6]}
   );
   gpc7_3 gpc4777 (
      {stage4_5[18], stage4_5[19], stage4_5[20], stage4_5[21], stage4_5[22], stage4_5[23], stage4_5[24]},
      {stage5_7[5],stage5_6[6],stage5_5[7]}
   );
   gpc7_3 gpc4778 (
      {stage4_5[25], stage4_5[26], stage4_5[27], stage4_5[28], stage4_5[29], stage4_5[30], stage4_5[31]},
      {stage5_7[6],stage5_6[7],stage5_5[8]}
   );
   gpc7_3 gpc4779 (
      {stage4_5[32], stage4_5[33], stage4_5[34], stage4_5[35], stage4_5[36], stage4_5[37], stage4_5[38]},
      {stage5_7[7],stage5_6[8],stage5_5[9]}
   );
   gpc7_3 gpc4780 (
      {stage4_5[39], stage4_5[40], stage4_5[41], stage4_5[42], stage4_5[43], stage4_5[44], stage4_5[45]},
      {stage5_7[8],stage5_6[9],stage5_5[10]}
   );
   gpc615_5 gpc4781 (
      {stage4_6[12], stage4_6[13], stage4_6[14], stage4_6[15], stage4_6[16]},
      {stage4_7[0]},
      {stage4_8[0], stage4_8[1], stage4_8[2], stage4_8[3], stage4_8[4], stage4_8[5]},
      {stage5_10[0],stage5_9[0],stage5_8[2],stage5_7[9],stage5_6[10]}
   );
   gpc615_5 gpc4782 (
      {stage4_6[17], stage4_6[18], stage4_6[19], stage4_6[20], stage4_6[21]},
      {stage4_7[1]},
      {stage4_8[6], stage4_8[7], stage4_8[8], stage4_8[9], stage4_8[10], stage4_8[11]},
      {stage5_10[1],stage5_9[1],stage5_8[3],stage5_7[10],stage5_6[11]}
   );
   gpc1163_5 gpc4783 (
      {stage4_7[2], stage4_7[3], stage4_7[4]},
      {stage4_8[12], stage4_8[13], stage4_8[14], stage4_8[15], stage4_8[16], stage4_8[17]},
      {stage4_9[0]},
      {stage4_10[0]},
      {stage5_11[0],stage5_10[2],stage5_9[2],stage5_8[4],stage5_7[11]}
   );
   gpc623_5 gpc4784 (
      {stage4_7[5], stage4_7[6], stage4_7[7]},
      {stage4_8[18], stage4_8[19]},
      {stage4_9[1], stage4_9[2], stage4_9[3], stage4_9[4], stage4_9[5], stage4_9[6]},
      {stage5_11[1],stage5_10[3],stage5_9[3],stage5_8[5],stage5_7[12]}
   );
   gpc606_5 gpc4785 (
      {stage4_8[20], stage4_8[21], stage4_8[22], stage4_8[23], stage4_8[24], stage4_8[25]},
      {stage4_10[1], stage4_10[2], stage4_10[3], stage4_10[4], stage4_10[5], stage4_10[6]},
      {stage5_12[0],stage5_11[2],stage5_10[4],stage5_9[4],stage5_8[6]}
   );
   gpc606_5 gpc4786 (
      {stage4_9[7], stage4_9[8], stage4_9[9], stage4_9[10], stage4_9[11], stage4_9[12]},
      {stage4_11[0], stage4_11[1], stage4_11[2], stage4_11[3], stage4_11[4], stage4_11[5]},
      {stage5_13[0],stage5_12[1],stage5_11[3],stage5_10[5],stage5_9[5]}
   );
   gpc606_5 gpc4787 (
      {stage4_9[13], stage4_9[14], stage4_9[15], stage4_9[16], stage4_9[17], stage4_9[18]},
      {stage4_11[6], stage4_11[7], stage4_11[8], stage4_11[9], stage4_11[10], stage4_11[11]},
      {stage5_13[1],stage5_12[2],stage5_11[4],stage5_10[6],stage5_9[6]}
   );
   gpc606_5 gpc4788 (
      {stage4_9[19], stage4_9[20], stage4_9[21], stage4_9[22], stage4_9[23], stage4_9[24]},
      {stage4_11[12], stage4_11[13], stage4_11[14], stage4_11[15], stage4_11[16], stage4_11[17]},
      {stage5_13[2],stage5_12[3],stage5_11[5],stage5_10[7],stage5_9[7]}
   );
   gpc606_5 gpc4789 (
      {stage4_9[25], stage4_9[26], stage4_9[27], stage4_9[28], stage4_9[29], stage4_9[30]},
      {stage4_11[18], stage4_11[19], stage4_11[20], stage4_11[21], stage4_11[22], stage4_11[23]},
      {stage5_13[3],stage5_12[4],stage5_11[6],stage5_10[8],stage5_9[8]}
   );
   gpc606_5 gpc4790 (
      {stage4_9[31], stage4_9[32], stage4_9[33], stage4_9[34], stage4_9[35], stage4_9[36]},
      {stage4_11[24], stage4_11[25], stage4_11[26], stage4_11[27], stage4_11[28], stage4_11[29]},
      {stage5_13[4],stage5_12[5],stage5_11[7],stage5_10[9],stage5_9[9]}
   );
   gpc615_5 gpc4791 (
      {stage4_9[37], stage4_9[38], stage4_9[39], stage4_9[40], stage4_9[41]},
      {stage4_10[7]},
      {stage4_11[30], stage4_11[31], stage4_11[32], stage4_11[33], stage4_11[34], stage4_11[35]},
      {stage5_13[5],stage5_12[6],stage5_11[8],stage5_10[10],stage5_9[10]}
   );
   gpc615_5 gpc4792 (
      {stage4_10[8], stage4_10[9], stage4_10[10], stage4_10[11], stage4_10[12]},
      {stage4_11[36]},
      {stage4_12[0], stage4_12[1], stage4_12[2], stage4_12[3], stage4_12[4], stage4_12[5]},
      {stage5_14[0],stage5_13[6],stage5_12[7],stage5_11[9],stage5_10[11]}
   );
   gpc615_5 gpc4793 (
      {stage4_10[13], stage4_10[14], stage4_10[15], stage4_10[16], stage4_10[17]},
      {stage4_11[37]},
      {stage4_12[6], stage4_12[7], stage4_12[8], stage4_12[9], stage4_12[10], stage4_12[11]},
      {stage5_14[1],stage5_13[7],stage5_12[8],stage5_11[10],stage5_10[12]}
   );
   gpc606_5 gpc4794 (
      {stage4_12[12], stage4_12[13], stage4_12[14], stage4_12[15], stage4_12[16], stage4_12[17]},
      {stage4_14[0], stage4_14[1], stage4_14[2], stage4_14[3], stage4_14[4], stage4_14[5]},
      {stage5_16[0],stage5_15[0],stage5_14[2],stage5_13[8],stage5_12[9]}
   );
   gpc606_5 gpc4795 (
      {stage4_12[18], stage4_12[19], stage4_12[20], stage4_12[21], stage4_12[22], stage4_12[23]},
      {stage4_14[6], stage4_14[7], stage4_14[8], stage4_14[9], stage4_14[10], stage4_14[11]},
      {stage5_16[1],stage5_15[1],stage5_14[3],stage5_13[9],stage5_12[10]}
   );
   gpc1163_5 gpc4796 (
      {stage4_13[0], stage4_13[1], stage4_13[2]},
      {stage4_14[12], stage4_14[13], stage4_14[14], stage4_14[15], stage4_14[16], stage4_14[17]},
      {stage4_15[0]},
      {stage4_16[0]},
      {stage5_17[0],stage5_16[2],stage5_15[2],stage5_14[4],stage5_13[10]}
   );
   gpc1163_5 gpc4797 (
      {stage4_13[3], stage4_13[4], stage4_13[5]},
      {stage4_14[18], stage4_14[19], stage4_14[20], stage4_14[21], stage4_14[22], stage4_14[23]},
      {stage4_15[1]},
      {stage4_16[1]},
      {stage5_17[1],stage5_16[3],stage5_15[3],stage5_14[5],stage5_13[11]}
   );
   gpc1163_5 gpc4798 (
      {stage4_13[6], stage4_13[7], stage4_13[8]},
      {stage4_14[24], stage4_14[25], stage4_14[26], stage4_14[27], stage4_14[28], stage4_14[29]},
      {stage4_15[2]},
      {stage4_16[2]},
      {stage5_17[2],stage5_16[4],stage5_15[4],stage5_14[6],stage5_13[12]}
   );
   gpc606_5 gpc4799 (
      {stage4_13[9], stage4_13[10], stage4_13[11], stage4_13[12], stage4_13[13], stage4_13[14]},
      {stage4_15[3], stage4_15[4], stage4_15[5], stage4_15[6], stage4_15[7], stage4_15[8]},
      {stage5_17[3],stage5_16[5],stage5_15[5],stage5_14[7],stage5_13[13]}
   );
   gpc606_5 gpc4800 (
      {stage4_13[15], stage4_13[16], stage4_13[17], stage4_13[18], 1'b0, 1'b0},
      {stage4_15[9], stage4_15[10], stage4_15[11], stage4_15[12], stage4_15[13], stage4_15[14]},
      {stage5_17[4],stage5_16[6],stage5_15[6],stage5_14[8],stage5_13[14]}
   );
   gpc135_4 gpc4801 (
      {stage4_14[30], stage4_14[31], stage4_14[32], stage4_14[33], stage4_14[34]},
      {stage4_15[15], stage4_15[16], stage4_15[17]},
      {stage4_16[3]},
      {stage5_17[5],stage5_16[7],stage5_15[7],stage5_14[9]}
   );
   gpc615_5 gpc4802 (
      {stage4_15[18], stage4_15[19], stage4_15[20], stage4_15[21], stage4_15[22]},
      {stage4_16[4]},
      {stage4_17[0], stage4_17[1], stage4_17[2], stage4_17[3], stage4_17[4], stage4_17[5]},
      {stage5_19[0],stage5_18[0],stage5_17[6],stage5_16[8],stage5_15[8]}
   );
   gpc615_5 gpc4803 (
      {stage4_15[23], stage4_15[24], stage4_15[25], stage4_15[26], stage4_15[27]},
      {stage4_16[5]},
      {stage4_17[6], stage4_17[7], stage4_17[8], stage4_17[9], stage4_17[10], stage4_17[11]},
      {stage5_19[1],stage5_18[1],stage5_17[7],stage5_16[9],stage5_15[9]}
   );
   gpc615_5 gpc4804 (
      {stage4_15[28], stage4_15[29], stage4_15[30], stage4_15[31], stage4_15[32]},
      {stage4_16[6]},
      {stage4_17[12], stage4_17[13], stage4_17[14], stage4_17[15], stage4_17[16], stage4_17[17]},
      {stage5_19[2],stage5_18[2],stage5_17[8],stage5_16[10],stage5_15[10]}
   );
   gpc615_5 gpc4805 (
      {stage4_15[33], stage4_15[34], stage4_15[35], stage4_15[36], stage4_15[37]},
      {stage4_16[7]},
      {stage4_17[18], stage4_17[19], stage4_17[20], stage4_17[21], stage4_17[22], stage4_17[23]},
      {stage5_19[3],stage5_18[3],stage5_17[9],stage5_16[11],stage5_15[11]}
   );
   gpc606_5 gpc4806 (
      {stage4_16[8], stage4_16[9], stage4_16[10], stage4_16[11], stage4_16[12], stage4_16[13]},
      {stage4_18[0], stage4_18[1], stage4_18[2], stage4_18[3], stage4_18[4], stage4_18[5]},
      {stage5_20[0],stage5_19[4],stage5_18[4],stage5_17[10],stage5_16[12]}
   );
   gpc615_5 gpc4807 (
      {stage4_16[14], stage4_16[15], stage4_16[16], stage4_16[17], stage4_16[18]},
      {stage4_17[24]},
      {stage4_18[6], stage4_18[7], stage4_18[8], stage4_18[9], stage4_18[10], stage4_18[11]},
      {stage5_20[1],stage5_19[5],stage5_18[5],stage5_17[11],stage5_16[13]}
   );
   gpc606_5 gpc4808 (
      {stage4_17[25], stage4_17[26], stage4_17[27], stage4_17[28], stage4_17[29], stage4_17[30]},
      {stage4_19[0], stage4_19[1], stage4_19[2], stage4_19[3], stage4_19[4], stage4_19[5]},
      {stage5_21[0],stage5_20[2],stage5_19[6],stage5_18[6],stage5_17[12]}
   );
   gpc606_5 gpc4809 (
      {stage4_17[31], stage4_17[32], stage4_17[33], stage4_17[34], stage4_17[35], stage4_17[36]},
      {stage4_19[6], stage4_19[7], stage4_19[8], stage4_19[9], stage4_19[10], stage4_19[11]},
      {stage5_21[1],stage5_20[3],stage5_19[7],stage5_18[7],stage5_17[13]}
   );
   gpc606_5 gpc4810 (
      {stage4_17[37], stage4_17[38], stage4_17[39], stage4_17[40], stage4_17[41], stage4_17[42]},
      {stage4_19[12], stage4_19[13], stage4_19[14], stage4_19[15], stage4_19[16], stage4_19[17]},
      {stage5_21[2],stage5_20[4],stage5_19[8],stage5_18[8],stage5_17[14]}
   );
   gpc606_5 gpc4811 (
      {stage4_18[12], stage4_18[13], stage4_18[14], stage4_18[15], stage4_18[16], stage4_18[17]},
      {stage4_20[0], stage4_20[1], stage4_20[2], stage4_20[3], stage4_20[4], stage4_20[5]},
      {stage5_22[0],stage5_21[3],stage5_20[5],stage5_19[9],stage5_18[9]}
   );
   gpc615_5 gpc4812 (
      {stage4_18[18], stage4_18[19], stage4_18[20], stage4_18[21], stage4_18[22]},
      {stage4_19[18]},
      {stage4_20[6], stage4_20[7], stage4_20[8], stage4_20[9], stage4_20[10], stage4_20[11]},
      {stage5_22[1],stage5_21[4],stage5_20[6],stage5_19[10],stage5_18[10]}
   );
   gpc615_5 gpc4813 (
      {stage4_21[0], stage4_21[1], stage4_21[2], stage4_21[3], stage4_21[4]},
      {stage4_22[0]},
      {stage4_23[0], stage4_23[1], stage4_23[2], stage4_23[3], stage4_23[4], stage4_23[5]},
      {stage5_25[0],stage5_24[0],stage5_23[0],stage5_22[2],stage5_21[5]}
   );
   gpc615_5 gpc4814 (
      {stage4_21[5], stage4_21[6], stage4_21[7], stage4_21[8], stage4_21[9]},
      {stage4_22[1]},
      {stage4_23[6], stage4_23[7], stage4_23[8], stage4_23[9], stage4_23[10], stage4_23[11]},
      {stage5_25[1],stage5_24[1],stage5_23[1],stage5_22[3],stage5_21[6]}
   );
   gpc615_5 gpc4815 (
      {stage4_21[10], stage4_21[11], stage4_21[12], stage4_21[13], stage4_21[14]},
      {stage4_22[2]},
      {stage4_23[12], stage4_23[13], stage4_23[14], stage4_23[15], stage4_23[16], stage4_23[17]},
      {stage5_25[2],stage5_24[2],stage5_23[2],stage5_22[4],stage5_21[7]}
   );
   gpc615_5 gpc4816 (
      {stage4_21[15], stage4_21[16], stage4_21[17], stage4_21[18], 1'b0},
      {stage4_22[3]},
      {stage4_23[18], stage4_23[19], stage4_23[20], stage4_23[21], stage4_23[22], stage4_23[23]},
      {stage5_25[3],stage5_24[3],stage5_23[3],stage5_22[5],stage5_21[8]}
   );
   gpc615_5 gpc4817 (
      {stage4_22[4], stage4_22[5], stage4_22[6], stage4_22[7], stage4_22[8]},
      {stage4_23[24]},
      {stage4_24[0], stage4_24[1], stage4_24[2], stage4_24[3], stage4_24[4], stage4_24[5]},
      {stage5_26[0],stage5_25[4],stage5_24[4],stage5_23[4],stage5_22[6]}
   );
   gpc615_5 gpc4818 (
      {stage4_22[9], stage4_22[10], stage4_22[11], stage4_22[12], stage4_22[13]},
      {stage4_23[25]},
      {stage4_24[6], stage4_24[7], stage4_24[8], stage4_24[9], stage4_24[10], stage4_24[11]},
      {stage5_26[1],stage5_25[5],stage5_24[5],stage5_23[5],stage5_22[7]}
   );
   gpc615_5 gpc4819 (
      {stage4_22[14], stage4_22[15], stage4_22[16], stage4_22[17], stage4_22[18]},
      {stage4_23[26]},
      {stage4_24[12], stage4_24[13], stage4_24[14], stage4_24[15], stage4_24[16], stage4_24[17]},
      {stage5_26[2],stage5_25[6],stage5_24[6],stage5_23[6],stage5_22[8]}
   );
   gpc615_5 gpc4820 (
      {stage4_22[19], stage4_22[20], stage4_22[21], stage4_22[22], stage4_22[23]},
      {stage4_23[27]},
      {stage4_24[18], stage4_24[19], stage4_24[20], stage4_24[21], stage4_24[22], stage4_24[23]},
      {stage5_26[3],stage5_25[7],stage5_24[7],stage5_23[7],stage5_22[9]}
   );
   gpc615_5 gpc4821 (
      {stage4_23[28], stage4_23[29], stage4_23[30], stage4_23[31], stage4_23[32]},
      {stage4_24[24]},
      {stage4_25[0], stage4_25[1], stage4_25[2], stage4_25[3], stage4_25[4], stage4_25[5]},
      {stage5_27[0],stage5_26[4],stage5_25[8],stage5_24[8],stage5_23[8]}
   );
   gpc615_5 gpc4822 (
      {stage4_23[33], stage4_23[34], stage4_23[35], stage4_23[36], stage4_23[37]},
      {stage4_24[25]},
      {stage4_25[6], stage4_25[7], stage4_25[8], stage4_25[9], stage4_25[10], stage4_25[11]},
      {stage5_27[1],stage5_26[5],stage5_25[9],stage5_24[9],stage5_23[9]}
   );
   gpc606_5 gpc4823 (
      {stage4_25[12], stage4_25[13], stage4_25[14], stage4_25[15], stage4_25[16], stage4_25[17]},
      {stage4_27[0], stage4_27[1], stage4_27[2], stage4_27[3], stage4_27[4], stage4_27[5]},
      {stage5_29[0],stage5_28[0],stage5_27[2],stage5_26[6],stage5_25[10]}
   );
   gpc615_5 gpc4824 (
      {stage4_26[0], stage4_26[1], stage4_26[2], stage4_26[3], stage4_26[4]},
      {stage4_27[6]},
      {stage4_28[0], stage4_28[1], stage4_28[2], stage4_28[3], stage4_28[4], stage4_28[5]},
      {stage5_30[0],stage5_29[1],stage5_28[1],stage5_27[3],stage5_26[7]}
   );
   gpc615_5 gpc4825 (
      {stage4_26[5], stage4_26[6], stage4_26[7], stage4_26[8], stage4_26[9]},
      {stage4_27[7]},
      {stage4_28[6], stage4_28[7], stage4_28[8], stage4_28[9], stage4_28[10], stage4_28[11]},
      {stage5_30[1],stage5_29[2],stage5_28[2],stage5_27[4],stage5_26[8]}
   );
   gpc615_5 gpc4826 (
      {stage4_26[10], stage4_26[11], stage4_26[12], stage4_26[13], stage4_26[14]},
      {stage4_27[8]},
      {stage4_28[12], stage4_28[13], stage4_28[14], stage4_28[15], stage4_28[16], stage4_28[17]},
      {stage5_30[2],stage5_29[3],stage5_28[3],stage5_27[5],stage5_26[9]}
   );
   gpc615_5 gpc4827 (
      {stage4_26[15], stage4_26[16], stage4_26[17], stage4_26[18], stage4_26[19]},
      {stage4_27[9]},
      {stage4_28[18], stage4_28[19], stage4_28[20], stage4_28[21], stage4_28[22], stage4_28[23]},
      {stage5_30[3],stage5_29[4],stage5_28[4],stage5_27[6],stage5_26[10]}
   );
   gpc207_4 gpc4828 (
      {stage4_27[10], stage4_27[11], stage4_27[12], stage4_27[13], stage4_27[14], stage4_27[15], stage4_27[16]},
      {stage4_29[0], stage4_29[1]},
      {stage5_30[4],stage5_29[5],stage5_28[5],stage5_27[7]}
   );
   gpc615_5 gpc4829 (
      {stage4_27[17], stage4_27[18], stage4_27[19], stage4_27[20], stage4_27[21]},
      {stage4_28[24]},
      {stage4_29[2], stage4_29[3], stage4_29[4], stage4_29[5], stage4_29[6], stage4_29[7]},
      {stage5_31[0],stage5_30[5],stage5_29[6],stage5_28[6],stage5_27[8]}
   );
   gpc615_5 gpc4830 (
      {stage4_29[8], stage4_29[9], stage4_29[10], stage4_29[11], stage4_29[12]},
      {stage4_30[0]},
      {stage4_31[0], stage4_31[1], stage4_31[2], stage4_31[3], stage4_31[4], stage4_31[5]},
      {stage5_33[0],stage5_32[0],stage5_31[1],stage5_30[6],stage5_29[7]}
   );
   gpc615_5 gpc4831 (
      {stage4_29[13], stage4_29[14], stage4_29[15], stage4_29[16], stage4_29[17]},
      {stage4_30[1]},
      {stage4_31[6], stage4_31[7], stage4_31[8], stage4_31[9], stage4_31[10], stage4_31[11]},
      {stage5_33[1],stage5_32[1],stage5_31[2],stage5_30[7],stage5_29[8]}
   );
   gpc615_5 gpc4832 (
      {stage4_29[18], stage4_29[19], stage4_29[20], stage4_29[21], stage4_29[22]},
      {stage4_30[2]},
      {stage4_31[12], stage4_31[13], stage4_31[14], stage4_31[15], stage4_31[16], stage4_31[17]},
      {stage5_33[2],stage5_32[2],stage5_31[3],stage5_30[8],stage5_29[9]}
   );
   gpc615_5 gpc4833 (
      {stage4_30[3], stage4_30[4], stage4_30[5], stage4_30[6], stage4_30[7]},
      {stage4_31[18]},
      {stage4_32[0], stage4_32[1], stage4_32[2], stage4_32[3], stage4_32[4], stage4_32[5]},
      {stage5_34[0],stage5_33[3],stage5_32[3],stage5_31[4],stage5_30[9]}
   );
   gpc615_5 gpc4834 (
      {stage4_30[8], stage4_30[9], stage4_30[10], stage4_30[11], stage4_30[12]},
      {stage4_31[19]},
      {stage4_32[6], stage4_32[7], stage4_32[8], stage4_32[9], stage4_32[10], stage4_32[11]},
      {stage5_34[1],stage5_33[4],stage5_32[4],stage5_31[5],stage5_30[10]}
   );
   gpc615_5 gpc4835 (
      {stage4_30[13], stage4_30[14], stage4_30[15], stage4_30[16], stage4_30[17]},
      {stage4_31[20]},
      {stage4_32[12], stage4_32[13], stage4_32[14], stage4_32[15], stage4_32[16], stage4_32[17]},
      {stage5_34[2],stage5_33[5],stage5_32[5],stage5_31[6],stage5_30[11]}
   );
   gpc615_5 gpc4836 (
      {stage4_30[18], stage4_30[19], stage4_30[20], stage4_30[21], stage4_30[22]},
      {stage4_31[21]},
      {stage4_32[18], stage4_32[19], stage4_32[20], stage4_32[21], stage4_32[22], stage4_32[23]},
      {stage5_34[3],stage5_33[6],stage5_32[6],stage5_31[7],stage5_30[12]}
   );
   gpc615_5 gpc4837 (
      {stage4_31[22], stage4_31[23], stage4_31[24], stage4_31[25], stage4_31[26]},
      {stage4_32[24]},
      {stage4_33[0], stage4_33[1], stage4_33[2], stage4_33[3], stage4_33[4], stage4_33[5]},
      {stage5_35[0],stage5_34[4],stage5_33[7],stage5_32[7],stage5_31[8]}
   );
   gpc606_5 gpc4838 (
      {stage4_33[6], stage4_33[7], stage4_33[8], stage4_33[9], stage4_33[10], stage4_33[11]},
      {stage4_35[0], stage4_35[1], stage4_35[2], stage4_35[3], stage4_35[4], stage4_35[5]},
      {stage5_37[0],stage5_36[0],stage5_35[1],stage5_34[5],stage5_33[8]}
   );
   gpc606_5 gpc4839 (
      {stage4_33[12], stage4_33[13], stage4_33[14], stage4_33[15], stage4_33[16], stage4_33[17]},
      {stage4_35[6], stage4_35[7], stage4_35[8], stage4_35[9], stage4_35[10], stage4_35[11]},
      {stage5_37[1],stage5_36[1],stage5_35[2],stage5_34[6],stage5_33[9]}
   );
   gpc606_5 gpc4840 (
      {stage4_34[0], stage4_34[1], stage4_34[2], stage4_34[3], stage4_34[4], stage4_34[5]},
      {stage4_36[0], stage4_36[1], stage4_36[2], stage4_36[3], stage4_36[4], stage4_36[5]},
      {stage5_38[0],stage5_37[2],stage5_36[2],stage5_35[3],stage5_34[7]}
   );
   gpc606_5 gpc4841 (
      {stage4_34[6], stage4_34[7], stage4_34[8], stage4_34[9], stage4_34[10], stage4_34[11]},
      {stage4_36[6], stage4_36[7], stage4_36[8], stage4_36[9], stage4_36[10], 1'b0},
      {stage5_38[1],stage5_37[3],stage5_36[3],stage5_35[4],stage5_34[8]}
   );
   gpc1_1 gpc4842 (
      {stage4_0[0]},
      {stage5_0[0]}
   );
   gpc1_1 gpc4843 (
      {stage4_0[1]},
      {stage5_0[1]}
   );
   gpc1_1 gpc4844 (
      {stage4_0[2]},
      {stage5_0[2]}
   );
   gpc1_1 gpc4845 (
      {stage4_0[3]},
      {stage5_0[3]}
   );
   gpc1_1 gpc4846 (
      {stage4_0[4]},
      {stage5_0[4]}
   );
   gpc1_1 gpc4847 (
      {stage4_0[5]},
      {stage5_0[5]}
   );
   gpc1_1 gpc4848 (
      {stage4_0[6]},
      {stage5_0[6]}
   );
   gpc1_1 gpc4849 (
      {stage4_0[7]},
      {stage5_0[7]}
   );
   gpc1_1 gpc4850 (
      {stage4_0[8]},
      {stage5_0[8]}
   );
   gpc1_1 gpc4851 (
      {stage4_0[9]},
      {stage5_0[9]}
   );
   gpc1_1 gpc4852 (
      {stage4_0[10]},
      {stage5_0[10]}
   );
   gpc1_1 gpc4853 (
      {stage4_1[6]},
      {stage5_1[1]}
   );
   gpc1_1 gpc4854 (
      {stage4_1[7]},
      {stage5_1[2]}
   );
   gpc1_1 gpc4855 (
      {stage4_1[8]},
      {stage5_1[3]}
   );
   gpc1_1 gpc4856 (
      {stage4_1[9]},
      {stage5_1[4]}
   );
   gpc1_1 gpc4857 (
      {stage4_1[10]},
      {stage5_1[5]}
   );
   gpc1_1 gpc4858 (
      {stage4_1[11]},
      {stage5_1[6]}
   );
   gpc1_1 gpc4859 (
      {stage4_1[12]},
      {stage5_1[7]}
   );
   gpc1_1 gpc4860 (
      {stage4_1[13]},
      {stage5_1[8]}
   );
   gpc1_1 gpc4861 (
      {stage4_1[14]},
      {stage5_1[9]}
   );
   gpc1_1 gpc4862 (
      {stage4_1[15]},
      {stage5_1[10]}
   );
   gpc1_1 gpc4863 (
      {stage4_2[5]},
      {stage5_2[2]}
   );
   gpc1_1 gpc4864 (
      {stage4_2[6]},
      {stage5_2[3]}
   );
   gpc1_1 gpc4865 (
      {stage4_2[7]},
      {stage5_2[4]}
   );
   gpc1_1 gpc4866 (
      {stage4_2[8]},
      {stage5_2[5]}
   );
   gpc1_1 gpc4867 (
      {stage4_2[9]},
      {stage5_2[6]}
   );
   gpc1_1 gpc4868 (
      {stage4_2[10]},
      {stage5_2[7]}
   );
   gpc1_1 gpc4869 (
      {stage4_2[11]},
      {stage5_2[8]}
   );
   gpc1_1 gpc4870 (
      {stage4_2[12]},
      {stage5_2[9]}
   );
   gpc1_1 gpc4871 (
      {stage4_3[22]},
      {stage5_3[5]}
   );
   gpc1_1 gpc4872 (
      {stage4_4[21]},
      {stage5_4[7]}
   );
   gpc1_1 gpc4873 (
      {stage4_4[22]},
      {stage5_4[8]}
   );
   gpc1_1 gpc4874 (
      {stage4_4[23]},
      {stage5_4[9]}
   );
   gpc1_1 gpc4875 (
      {stage4_6[22]},
      {stage5_6[12]}
   );
   gpc1_1 gpc4876 (
      {stage4_7[8]},
      {stage5_7[13]}
   );
   gpc1_1 gpc4877 (
      {stage4_7[9]},
      {stage5_7[14]}
   );
   gpc1_1 gpc4878 (
      {stage4_7[10]},
      {stage5_7[15]}
   );
   gpc1_1 gpc4879 (
      {stage4_7[11]},
      {stage5_7[16]}
   );
   gpc1_1 gpc4880 (
      {stage4_7[12]},
      {stage5_7[17]}
   );
   gpc1_1 gpc4881 (
      {stage4_7[13]},
      {stage5_7[18]}
   );
   gpc1_1 gpc4882 (
      {stage4_7[14]},
      {stage5_7[19]}
   );
   gpc1_1 gpc4883 (
      {stage4_8[26]},
      {stage5_8[7]}
   );
   gpc1_1 gpc4884 (
      {stage4_8[27]},
      {stage5_8[8]}
   );
   gpc1_1 gpc4885 (
      {stage4_8[28]},
      {stage5_8[9]}
   );
   gpc1_1 gpc4886 (
      {stage4_11[38]},
      {stage5_11[11]}
   );
   gpc1_1 gpc4887 (
      {stage4_11[39]},
      {stage5_11[12]}
   );
   gpc1_1 gpc4888 (
      {stage4_11[40]},
      {stage5_11[13]}
   );
   gpc1_1 gpc4889 (
      {stage4_11[41]},
      {stage5_11[14]}
   );
   gpc1_1 gpc4890 (
      {stage4_11[42]},
      {stage5_11[15]}
   );
   gpc1_1 gpc4891 (
      {stage4_15[38]},
      {stage5_15[12]}
   );
   gpc1_1 gpc4892 (
      {stage4_16[19]},
      {stage5_16[14]}
   );
   gpc1_1 gpc4893 (
      {stage4_18[23]},
      {stage5_18[11]}
   );
   gpc1_1 gpc4894 (
      {stage4_18[24]},
      {stage5_18[12]}
   );
   gpc1_1 gpc4895 (
      {stage4_18[25]},
      {stage5_18[13]}
   );
   gpc1_1 gpc4896 (
      {stage4_18[26]},
      {stage5_18[14]}
   );
   gpc1_1 gpc4897 (
      {stage4_18[27]},
      {stage5_18[15]}
   );
   gpc1_1 gpc4898 (
      {stage4_18[28]},
      {stage5_18[16]}
   );
   gpc1_1 gpc4899 (
      {stage4_19[19]},
      {stage5_19[11]}
   );
   gpc1_1 gpc4900 (
      {stage4_19[20]},
      {stage5_19[12]}
   );
   gpc1_1 gpc4901 (
      {stage4_19[21]},
      {stage5_19[13]}
   );
   gpc1_1 gpc4902 (
      {stage4_19[22]},
      {stage5_19[14]}
   );
   gpc1_1 gpc4903 (
      {stage4_19[23]},
      {stage5_19[15]}
   );
   gpc1_1 gpc4904 (
      {stage4_19[24]},
      {stage5_19[16]}
   );
   gpc1_1 gpc4905 (
      {stage4_19[25]},
      {stage5_19[17]}
   );
   gpc1_1 gpc4906 (
      {stage4_19[26]},
      {stage5_19[18]}
   );
   gpc1_1 gpc4907 (
      {stage4_19[27]},
      {stage5_19[19]}
   );
   gpc1_1 gpc4908 (
      {stage4_19[28]},
      {stage5_19[20]}
   );
   gpc1_1 gpc4909 (
      {stage4_19[29]},
      {stage5_19[21]}
   );
   gpc1_1 gpc4910 (
      {stage4_19[30]},
      {stage5_19[22]}
   );
   gpc1_1 gpc4911 (
      {stage4_19[31]},
      {stage5_19[23]}
   );
   gpc1_1 gpc4912 (
      {stage4_20[12]},
      {stage5_20[7]}
   );
   gpc1_1 gpc4913 (
      {stage4_20[13]},
      {stage5_20[8]}
   );
   gpc1_1 gpc4914 (
      {stage4_20[14]},
      {stage5_20[9]}
   );
   gpc1_1 gpc4915 (
      {stage4_20[15]},
      {stage5_20[10]}
   );
   gpc1_1 gpc4916 (
      {stage4_20[16]},
      {stage5_20[11]}
   );
   gpc1_1 gpc4917 (
      {stage4_20[17]},
      {stage5_20[12]}
   );
   gpc1_1 gpc4918 (
      {stage4_20[18]},
      {stage5_20[13]}
   );
   gpc1_1 gpc4919 (
      {stage4_22[24]},
      {stage5_22[10]}
   );
   gpc1_1 gpc4920 (
      {stage4_22[25]},
      {stage5_22[11]}
   );
   gpc1_1 gpc4921 (
      {stage4_22[26]},
      {stage5_22[12]}
   );
   gpc1_1 gpc4922 (
      {stage4_22[27]},
      {stage5_22[13]}
   );
   gpc1_1 gpc4923 (
      {stage4_22[28]},
      {stage5_22[14]}
   );
   gpc1_1 gpc4924 (
      {stage4_22[29]},
      {stage5_22[15]}
   );
   gpc1_1 gpc4925 (
      {stage4_22[30]},
      {stage5_22[16]}
   );
   gpc1_1 gpc4926 (
      {stage4_24[26]},
      {stage5_24[10]}
   );
   gpc1_1 gpc4927 (
      {stage4_24[27]},
      {stage5_24[11]}
   );
   gpc1_1 gpc4928 (
      {stage4_24[28]},
      {stage5_24[12]}
   );
   gpc1_1 gpc4929 (
      {stage4_24[29]},
      {stage5_24[13]}
   );
   gpc1_1 gpc4930 (
      {stage4_25[18]},
      {stage5_25[11]}
   );
   gpc1_1 gpc4931 (
      {stage4_26[20]},
      {stage5_26[11]}
   );
   gpc1_1 gpc4932 (
      {stage4_26[21]},
      {stage5_26[12]}
   );
   gpc1_1 gpc4933 (
      {stage4_26[22]},
      {stage5_26[13]}
   );
   gpc1_1 gpc4934 (
      {stage4_27[22]},
      {stage5_27[9]}
   );
   gpc1_1 gpc4935 (
      {stage4_27[23]},
      {stage5_27[10]}
   );
   gpc1_1 gpc4936 (
      {stage4_27[24]},
      {stage5_27[11]}
   );
   gpc1_1 gpc4937 (
      {stage4_27[25]},
      {stage5_27[12]}
   );
   gpc1_1 gpc4938 (
      {stage4_27[26]},
      {stage5_27[13]}
   );
   gpc1_1 gpc4939 (
      {stage4_29[23]},
      {stage5_29[10]}
   );
   gpc1_1 gpc4940 (
      {stage4_29[24]},
      {stage5_29[11]}
   );
   gpc1_1 gpc4941 (
      {stage4_29[25]},
      {stage5_29[12]}
   );
   gpc1_1 gpc4942 (
      {stage4_30[23]},
      {stage5_30[13]}
   );
   gpc1_1 gpc4943 (
      {stage4_30[24]},
      {stage5_30[14]}
   );
   gpc1_1 gpc4944 (
      {stage4_30[25]},
      {stage5_30[15]}
   );
   gpc1_1 gpc4945 (
      {stage4_30[26]},
      {stage5_30[16]}
   );
   gpc1_1 gpc4946 (
      {stage4_31[27]},
      {stage5_31[9]}
   );
   gpc1_1 gpc4947 (
      {stage4_31[28]},
      {stage5_31[10]}
   );
   gpc1_1 gpc4948 (
      {stage4_31[29]},
      {stage5_31[11]}
   );
   gpc1_1 gpc4949 (
      {stage4_31[30]},
      {stage5_31[12]}
   );
   gpc1_1 gpc4950 (
      {stage4_32[25]},
      {stage5_32[8]}
   );
   gpc1_1 gpc4951 (
      {stage4_32[26]},
      {stage5_32[9]}
   );
   gpc1_1 gpc4952 (
      {stage4_32[27]},
      {stage5_32[10]}
   );
   gpc1_1 gpc4953 (
      {stage4_32[28]},
      {stage5_32[11]}
   );
   gpc1_1 gpc4954 (
      {stage4_32[29]},
      {stage5_32[12]}
   );
   gpc1_1 gpc4955 (
      {stage4_32[30]},
      {stage5_32[13]}
   );
   gpc1_1 gpc4956 (
      {stage4_32[31]},
      {stage5_32[14]}
   );
   gpc1_1 gpc4957 (
      {stage4_32[32]},
      {stage5_32[15]}
   );
   gpc1_1 gpc4958 (
      {stage4_32[33]},
      {stage5_32[16]}
   );
   gpc1_1 gpc4959 (
      {stage4_32[34]},
      {stage5_32[17]}
   );
   gpc1_1 gpc4960 (
      {stage4_32[35]},
      {stage5_32[18]}
   );
   gpc1_1 gpc4961 (
      {stage4_32[36]},
      {stage5_32[19]}
   );
   gpc1_1 gpc4962 (
      {stage4_32[37]},
      {stage5_32[20]}
   );
   gpc1_1 gpc4963 (
      {stage4_32[38]},
      {stage5_32[21]}
   );
   gpc1_1 gpc4964 (
      {stage4_32[39]},
      {stage5_32[22]}
   );
   gpc1_1 gpc4965 (
      {stage4_32[40]},
      {stage5_32[23]}
   );
   gpc1_1 gpc4966 (
      {stage4_32[41]},
      {stage5_32[24]}
   );
   gpc1_1 gpc4967 (
      {stage4_32[42]},
      {stage5_32[25]}
   );
   gpc1_1 gpc4968 (
      {stage4_33[18]},
      {stage5_33[10]}
   );
   gpc1_1 gpc4969 (
      {stage4_34[12]},
      {stage5_34[9]}
   );
   gpc1_1 gpc4970 (
      {stage4_35[12]},
      {stage5_35[5]}
   );
   gpc1_1 gpc4971 (
      {stage4_35[13]},
      {stage5_35[6]}
   );
   gpc1_1 gpc4972 (
      {stage4_35[14]},
      {stage5_35[7]}
   );
   gpc1_1 gpc4973 (
      {stage4_37[0]},
      {stage5_37[4]}
   );
   gpc1_1 gpc4974 (
      {stage4_37[1]},
      {stage5_37[5]}
   );
   gpc1_1 gpc4975 (
      {stage4_37[2]},
      {stage5_37[6]}
   );
   gpc1343_5 gpc4976 (
      {stage5_0[0], stage5_0[1], stage5_0[2]},
      {stage5_1[0], stage5_1[1], stage5_1[2], stage5_1[3]},
      {stage5_2[0], stage5_2[1], stage5_2[2]},
      {stage5_3[0]},
      {stage6_4[0],stage6_3[0],stage6_2[0],stage6_1[0],stage6_0[0]}
   );
   gpc1343_5 gpc4977 (
      {stage5_0[3], stage5_0[4], stage5_0[5]},
      {stage5_1[4], stage5_1[5], stage5_1[6], stage5_1[7]},
      {stage5_2[3], stage5_2[4], stage5_2[5]},
      {stage5_3[1]},
      {stage6_4[1],stage6_3[1],stage6_2[1],stage6_1[1],stage6_0[1]}
   );
   gpc117_4 gpc4978 (
      {stage5_4[0], stage5_4[1], stage5_4[2], stage5_4[3], stage5_4[4], stage5_4[5], stage5_4[6]},
      {stage5_5[0]},
      {stage5_6[0]},
      {stage6_7[0],stage6_6[0],stage6_5[0],stage6_4[2]}
   );
   gpc1343_5 gpc4979 (
      {stage5_5[1], stage5_5[2], stage5_5[3]},
      {stage5_6[1], stage5_6[2], stage5_6[3], stage5_6[4]},
      {stage5_7[0], stage5_7[1], stage5_7[2]},
      {stage5_8[0]},
      {stage6_9[0],stage6_8[0],stage6_7[1],stage6_6[1],stage6_5[1]}
   );
   gpc1343_5 gpc4980 (
      {stage5_5[4], stage5_5[5], stage5_5[6]},
      {stage5_6[5], stage5_6[6], stage5_6[7], stage5_6[8]},
      {stage5_7[3], stage5_7[4], stage5_7[5]},
      {stage5_8[1]},
      {stage6_9[1],stage6_8[1],stage6_7[2],stage6_6[2],stage6_5[2]}
   );
   gpc1343_5 gpc4981 (
      {stage5_5[7], stage5_5[8], stage5_5[9]},
      {stage5_6[9], stage5_6[10], stage5_6[11], stage5_6[12]},
      {stage5_7[6], stage5_7[7], stage5_7[8]},
      {stage5_8[2]},
      {stage6_9[2],stage6_8[2],stage6_7[3],stage6_6[3],stage6_5[3]}
   );
   gpc606_5 gpc4982 (
      {stage5_7[9], stage5_7[10], stage5_7[11], stage5_7[12], stage5_7[13], stage5_7[14]},
      {stage5_9[0], stage5_9[1], stage5_9[2], stage5_9[3], stage5_9[4], stage5_9[5]},
      {stage6_11[0],stage6_10[0],stage6_9[3],stage6_8[3],stage6_7[4]}
   );
   gpc615_5 gpc4983 (
      {stage5_7[15], stage5_7[16], stage5_7[17], stage5_7[18], stage5_7[19]},
      {stage5_8[3]},
      {stage5_9[6], stage5_9[7], stage5_9[8], stage5_9[9], stage5_9[10], 1'b0},
      {stage6_11[1],stage6_10[1],stage6_9[4],stage6_8[4],stage6_7[5]}
   );
   gpc606_5 gpc4984 (
      {stage5_8[4], stage5_8[5], stage5_8[6], stage5_8[7], stage5_8[8], stage5_8[9]},
      {stage5_10[0], stage5_10[1], stage5_10[2], stage5_10[3], stage5_10[4], stage5_10[5]},
      {stage6_12[0],stage6_11[2],stage6_10[2],stage6_9[5],stage6_8[5]}
   );
   gpc7_3 gpc4985 (
      {stage5_10[6], stage5_10[7], stage5_10[8], stage5_10[9], stage5_10[10], stage5_10[11], stage5_10[12]},
      {stage6_12[1],stage6_11[3],stage6_10[3]}
   );
   gpc207_4 gpc4986 (
      {stage5_11[0], stage5_11[1], stage5_11[2], stage5_11[3], stage5_11[4], stage5_11[5], stage5_11[6]},
      {stage5_13[0], stage5_13[1]},
      {stage6_14[0],stage6_13[0],stage6_12[2],stage6_11[4]}
   );
   gpc207_4 gpc4987 (
      {stage5_11[7], stage5_11[8], stage5_11[9], stage5_11[10], stage5_11[11], stage5_11[12], stage5_11[13]},
      {stage5_13[2], stage5_13[3]},
      {stage6_14[1],stage6_13[1],stage6_12[3],stage6_11[5]}
   );
   gpc7_3 gpc4988 (
      {stage5_12[0], stage5_12[1], stage5_12[2], stage5_12[3], stage5_12[4], stage5_12[5], stage5_12[6]},
      {stage6_14[2],stage6_13[2],stage6_12[4]}
   );
   gpc623_5 gpc4989 (
      {stage5_12[7], stage5_12[8], stage5_12[9]},
      {stage5_13[4], stage5_13[5]},
      {stage5_14[0], stage5_14[1], stage5_14[2], stage5_14[3], stage5_14[4], stage5_14[5]},
      {stage6_16[0],stage6_15[0],stage6_14[3],stage6_13[3],stage6_12[5]}
   );
   gpc623_5 gpc4990 (
      {stage5_13[6], stage5_13[7], stage5_13[8]},
      {stage5_14[6], stage5_14[7]},
      {stage5_15[0], stage5_15[1], stage5_15[2], stage5_15[3], stage5_15[4], stage5_15[5]},
      {stage6_17[0],stage6_16[1],stage6_15[1],stage6_14[4],stage6_13[4]}
   );
   gpc623_5 gpc4991 (
      {stage5_13[9], stage5_13[10], stage5_13[11]},
      {stage5_14[8], stage5_14[9]},
      {stage5_15[6], stage5_15[7], stage5_15[8], stage5_15[9], stage5_15[10], stage5_15[11]},
      {stage6_17[1],stage6_16[2],stage6_15[2],stage6_14[5],stage6_13[5]}
   );
   gpc207_4 gpc4992 (
      {stage5_16[0], stage5_16[1], stage5_16[2], stage5_16[3], stage5_16[4], stage5_16[5], stage5_16[6]},
      {stage5_18[0], stage5_18[1]},
      {stage6_19[0],stage6_18[0],stage6_17[2],stage6_16[3]}
   );
   gpc207_4 gpc4993 (
      {stage5_16[7], stage5_16[8], stage5_16[9], stage5_16[10], stage5_16[11], stage5_16[12], stage5_16[13]},
      {stage5_18[2], stage5_18[3]},
      {stage6_19[1],stage6_18[1],stage6_17[3],stage6_16[4]}
   );
   gpc1163_5 gpc4994 (
      {stage5_17[0], stage5_17[1], stage5_17[2]},
      {stage5_18[4], stage5_18[5], stage5_18[6], stage5_18[7], stage5_18[8], stage5_18[9]},
      {stage5_19[0]},
      {stage5_20[0]},
      {stage6_21[0],stage6_20[0],stage6_19[2],stage6_18[2],stage6_17[4]}
   );
   gpc1163_5 gpc4995 (
      {stage5_17[3], stage5_17[4], stage5_17[5]},
      {stage5_18[10], stage5_18[11], stage5_18[12], stage5_18[13], stage5_18[14], stage5_18[15]},
      {stage5_19[1]},
      {stage5_20[1]},
      {stage6_21[1],stage6_20[1],stage6_19[3],stage6_18[3],stage6_17[5]}
   );
   gpc606_5 gpc4996 (
      {stage5_17[6], stage5_17[7], stage5_17[8], stage5_17[9], stage5_17[10], stage5_17[11]},
      {stage5_19[2], stage5_19[3], stage5_19[4], stage5_19[5], stage5_19[6], stage5_19[7]},
      {stage6_21[2],stage6_20[2],stage6_19[4],stage6_18[4],stage6_17[6]}
   );
   gpc207_4 gpc4997 (
      {stage5_19[8], stage5_19[9], stage5_19[10], stage5_19[11], stage5_19[12], stage5_19[13], stage5_19[14]},
      {stage5_21[0], stage5_21[1]},
      {stage6_22[0],stage6_21[3],stage6_20[3],stage6_19[5]}
   );
   gpc606_5 gpc4998 (
      {stage5_20[2], stage5_20[3], stage5_20[4], stage5_20[5], stage5_20[6], stage5_20[7]},
      {stage5_22[0], stage5_22[1], stage5_22[2], stage5_22[3], stage5_22[4], stage5_22[5]},
      {stage6_24[0],stage6_23[0],stage6_22[1],stage6_21[4],stage6_20[4]}
   );
   gpc606_5 gpc4999 (
      {stage5_20[8], stage5_20[9], stage5_20[10], stage5_20[11], stage5_20[12], stage5_20[13]},
      {stage5_22[6], stage5_22[7], stage5_22[8], stage5_22[9], stage5_22[10], stage5_22[11]},
      {stage6_24[1],stage6_23[1],stage6_22[2],stage6_21[5],stage6_20[5]}
   );
   gpc1415_5 gpc5000 (
      {stage5_23[0], stage5_23[1], stage5_23[2], stage5_23[3], stage5_23[4]},
      {stage5_24[0]},
      {stage5_25[0], stage5_25[1], stage5_25[2], stage5_25[3]},
      {stage5_26[0]},
      {stage6_27[0],stage6_26[0],stage6_25[0],stage6_24[2],stage6_23[2]}
   );
   gpc615_5 gpc5001 (
      {stage5_23[5], stage5_23[6], stage5_23[7], stage5_23[8], stage5_23[9]},
      {stage5_24[1]},
      {stage5_25[4], stage5_25[5], stage5_25[6], stage5_25[7], stage5_25[8], stage5_25[9]},
      {stage6_27[1],stage6_26[1],stage6_25[1],stage6_24[3],stage6_23[3]}
   );
   gpc606_5 gpc5002 (
      {stage5_24[2], stage5_24[3], stage5_24[4], stage5_24[5], stage5_24[6], stage5_24[7]},
      {stage5_26[1], stage5_26[2], stage5_26[3], stage5_26[4], stage5_26[5], stage5_26[6]},
      {stage6_28[0],stage6_27[2],stage6_26[2],stage6_25[2],stage6_24[4]}
   );
   gpc606_5 gpc5003 (
      {stage5_24[8], stage5_24[9], stage5_24[10], stage5_24[11], stage5_24[12], stage5_24[13]},
      {stage5_26[7], stage5_26[8], stage5_26[9], stage5_26[10], stage5_26[11], stage5_26[12]},
      {stage6_28[1],stage6_27[3],stage6_26[3],stage6_25[3],stage6_24[5]}
   );
   gpc606_5 gpc5004 (
      {stage5_27[0], stage5_27[1], stage5_27[2], stage5_27[3], stage5_27[4], stage5_27[5]},
      {stage5_29[0], stage5_29[1], stage5_29[2], stage5_29[3], stage5_29[4], stage5_29[5]},
      {stage6_31[0],stage6_30[0],stage6_29[0],stage6_28[2],stage6_27[4]}
   );
   gpc606_5 gpc5005 (
      {stage5_27[6], stage5_27[7], stage5_27[8], stage5_27[9], stage5_27[10], stage5_27[11]},
      {stage5_29[6], stage5_29[7], stage5_29[8], stage5_29[9], stage5_29[10], stage5_29[11]},
      {stage6_31[1],stage6_30[1],stage6_29[1],stage6_28[3],stage6_27[5]}
   );
   gpc207_4 gpc5006 (
      {stage5_28[0], stage5_28[1], stage5_28[2], stage5_28[3], stage5_28[4], stage5_28[5], stage5_28[6]},
      {stage5_30[0], stage5_30[1]},
      {stage6_31[2],stage6_30[2],stage6_29[2],stage6_28[4]}
   );
   gpc615_5 gpc5007 (
      {stage5_30[2], stage5_30[3], stage5_30[4], stage5_30[5], stage5_30[6]},
      {stage5_31[0]},
      {stage5_32[0], stage5_32[1], stage5_32[2], stage5_32[3], stage5_32[4], stage5_32[5]},
      {stage6_34[0],stage6_33[0],stage6_32[0],stage6_31[3],stage6_30[3]}
   );
   gpc615_5 gpc5008 (
      {stage5_30[7], stage5_30[8], stage5_30[9], stage5_30[10], stage5_30[11]},
      {stage5_31[1]},
      {stage5_32[6], stage5_32[7], stage5_32[8], stage5_32[9], stage5_32[10], stage5_32[11]},
      {stage6_34[1],stage6_33[1],stage6_32[1],stage6_31[4],stage6_30[4]}
   );
   gpc615_5 gpc5009 (
      {stage5_30[12], stage5_30[13], stage5_30[14], stage5_30[15], stage5_30[16]},
      {stage5_31[2]},
      {stage5_32[12], stage5_32[13], stage5_32[14], stage5_32[15], stage5_32[16], stage5_32[17]},
      {stage6_34[2],stage6_33[2],stage6_32[2],stage6_31[5],stage6_30[5]}
   );
   gpc615_5 gpc5010 (
      {stage5_31[3], stage5_31[4], stage5_31[5], stage5_31[6], stage5_31[7]},
      {stage5_32[18]},
      {stage5_33[0], stage5_33[1], stage5_33[2], stage5_33[3], stage5_33[4], stage5_33[5]},
      {stage6_35[0],stage6_34[3],stage6_33[3],stage6_32[3],stage6_31[6]}
   );
   gpc615_5 gpc5011 (
      {stage5_31[8], stage5_31[9], stage5_31[10], stage5_31[11], stage5_31[12]},
      {stage5_32[19]},
      {stage5_33[6], stage5_33[7], stage5_33[8], stage5_33[9], stage5_33[10], 1'b0},
      {stage6_35[1],stage6_34[4],stage6_33[4],stage6_32[4],stage6_31[7]}
   );
   gpc606_5 gpc5012 (
      {stage5_32[20], stage5_32[21], stage5_32[22], stage5_32[23], stage5_32[24], stage5_32[25]},
      {stage5_34[0], stage5_34[1], stage5_34[2], stage5_34[3], stage5_34[4], stage5_34[5]},
      {stage6_36[0],stage6_35[2],stage6_34[5],stage6_33[5],stage6_32[5]}
   );
   gpc606_5 gpc5013 (
      {stage5_35[0], stage5_35[1], stage5_35[2], stage5_35[3], stage5_35[4], stage5_35[5]},
      {stage5_37[0], stage5_37[1], stage5_37[2], stage5_37[3], stage5_37[4], stage5_37[5]},
      {stage6_39[0],stage6_38[0],stage6_37[0],stage6_36[1],stage6_35[3]}
   );
   gpc1325_5 gpc5014 (
      {stage5_36[0], stage5_36[1], stage5_36[2], stage5_36[3], 1'b0},
      {stage5_37[6], 1'b0},
      {stage5_38[0], stage5_38[1], 1'b0},
      {1'b0},
      {stage6_40[0],stage6_39[1],stage6_38[1],stage6_37[1],stage6_36[2]}
   );
   gpc1_1 gpc5015 (
      {stage5_0[6]},
      {stage6_0[2]}
   );
   gpc1_1 gpc5016 (
      {stage5_0[7]},
      {stage6_0[3]}
   );
   gpc1_1 gpc5017 (
      {stage5_0[8]},
      {stage6_0[4]}
   );
   gpc1_1 gpc5018 (
      {stage5_0[9]},
      {stage6_0[5]}
   );
   gpc1_1 gpc5019 (
      {stage5_0[10]},
      {stage6_0[6]}
   );
   gpc1_1 gpc5020 (
      {stage5_1[8]},
      {stage6_1[2]}
   );
   gpc1_1 gpc5021 (
      {stage5_1[9]},
      {stage6_1[3]}
   );
   gpc1_1 gpc5022 (
      {stage5_1[10]},
      {stage6_1[4]}
   );
   gpc1_1 gpc5023 (
      {stage5_2[6]},
      {stage6_2[2]}
   );
   gpc1_1 gpc5024 (
      {stage5_2[7]},
      {stage6_2[3]}
   );
   gpc1_1 gpc5025 (
      {stage5_2[8]},
      {stage6_2[4]}
   );
   gpc1_1 gpc5026 (
      {stage5_2[9]},
      {stage6_2[5]}
   );
   gpc1_1 gpc5027 (
      {stage5_3[2]},
      {stage6_3[2]}
   );
   gpc1_1 gpc5028 (
      {stage5_3[3]},
      {stage6_3[3]}
   );
   gpc1_1 gpc5029 (
      {stage5_3[4]},
      {stage6_3[4]}
   );
   gpc1_1 gpc5030 (
      {stage5_3[5]},
      {stage6_3[5]}
   );
   gpc1_1 gpc5031 (
      {stage5_4[7]},
      {stage6_4[3]}
   );
   gpc1_1 gpc5032 (
      {stage5_4[8]},
      {stage6_4[4]}
   );
   gpc1_1 gpc5033 (
      {stage5_4[9]},
      {stage6_4[5]}
   );
   gpc1_1 gpc5034 (
      {stage5_5[10]},
      {stage6_5[4]}
   );
   gpc1_1 gpc5035 (
      {stage5_11[14]},
      {stage6_11[6]}
   );
   gpc1_1 gpc5036 (
      {stage5_11[15]},
      {stage6_11[7]}
   );
   gpc1_1 gpc5037 (
      {stage5_12[10]},
      {stage6_12[6]}
   );
   gpc1_1 gpc5038 (
      {stage5_13[12]},
      {stage6_13[6]}
   );
   gpc1_1 gpc5039 (
      {stage5_13[13]},
      {stage6_13[7]}
   );
   gpc1_1 gpc5040 (
      {stage5_13[14]},
      {stage6_13[8]}
   );
   gpc1_1 gpc5041 (
      {stage5_15[12]},
      {stage6_15[3]}
   );
   gpc1_1 gpc5042 (
      {stage5_16[14]},
      {stage6_16[5]}
   );
   gpc1_1 gpc5043 (
      {stage5_17[12]},
      {stage6_17[7]}
   );
   gpc1_1 gpc5044 (
      {stage5_17[13]},
      {stage6_17[8]}
   );
   gpc1_1 gpc5045 (
      {stage5_17[14]},
      {stage6_17[9]}
   );
   gpc1_1 gpc5046 (
      {stage5_18[16]},
      {stage6_18[5]}
   );
   gpc1_1 gpc5047 (
      {stage5_19[15]},
      {stage6_19[6]}
   );
   gpc1_1 gpc5048 (
      {stage5_19[16]},
      {stage6_19[7]}
   );
   gpc1_1 gpc5049 (
      {stage5_19[17]},
      {stage6_19[8]}
   );
   gpc1_1 gpc5050 (
      {stage5_19[18]},
      {stage6_19[9]}
   );
   gpc1_1 gpc5051 (
      {stage5_19[19]},
      {stage6_19[10]}
   );
   gpc1_1 gpc5052 (
      {stage5_19[20]},
      {stage6_19[11]}
   );
   gpc1_1 gpc5053 (
      {stage5_19[21]},
      {stage6_19[12]}
   );
   gpc1_1 gpc5054 (
      {stage5_19[22]},
      {stage6_19[13]}
   );
   gpc1_1 gpc5055 (
      {stage5_19[23]},
      {stage6_19[14]}
   );
   gpc1_1 gpc5056 (
      {stage5_21[2]},
      {stage6_21[6]}
   );
   gpc1_1 gpc5057 (
      {stage5_21[3]},
      {stage6_21[7]}
   );
   gpc1_1 gpc5058 (
      {stage5_21[4]},
      {stage6_21[8]}
   );
   gpc1_1 gpc5059 (
      {stage5_21[5]},
      {stage6_21[9]}
   );
   gpc1_1 gpc5060 (
      {stage5_21[6]},
      {stage6_21[10]}
   );
   gpc1_1 gpc5061 (
      {stage5_21[7]},
      {stage6_21[11]}
   );
   gpc1_1 gpc5062 (
      {stage5_21[8]},
      {stage6_21[12]}
   );
   gpc1_1 gpc5063 (
      {stage5_22[12]},
      {stage6_22[3]}
   );
   gpc1_1 gpc5064 (
      {stage5_22[13]},
      {stage6_22[4]}
   );
   gpc1_1 gpc5065 (
      {stage5_22[14]},
      {stage6_22[5]}
   );
   gpc1_1 gpc5066 (
      {stage5_22[15]},
      {stage6_22[6]}
   );
   gpc1_1 gpc5067 (
      {stage5_22[16]},
      {stage6_22[7]}
   );
   gpc1_1 gpc5068 (
      {stage5_25[10]},
      {stage6_25[4]}
   );
   gpc1_1 gpc5069 (
      {stage5_25[11]},
      {stage6_25[5]}
   );
   gpc1_1 gpc5070 (
      {stage5_26[13]},
      {stage6_26[4]}
   );
   gpc1_1 gpc5071 (
      {stage5_27[12]},
      {stage6_27[6]}
   );
   gpc1_1 gpc5072 (
      {stage5_27[13]},
      {stage6_27[7]}
   );
   gpc1_1 gpc5073 (
      {stage5_29[12]},
      {stage6_29[3]}
   );
   gpc1_1 gpc5074 (
      {stage5_34[6]},
      {stage6_34[6]}
   );
   gpc1_1 gpc5075 (
      {stage5_34[7]},
      {stage6_34[7]}
   );
   gpc1_1 gpc5076 (
      {stage5_34[8]},
      {stage6_34[8]}
   );
   gpc1_1 gpc5077 (
      {stage5_34[9]},
      {stage6_34[9]}
   );
   gpc1_1 gpc5078 (
      {stage5_35[6]},
      {stage6_35[4]}
   );
   gpc1_1 gpc5079 (
      {stage5_35[7]},
      {stage6_35[5]}
   );
   gpc606_5 gpc5080 (
      {stage6_1[0], stage6_1[1], stage6_1[2], stage6_1[3], stage6_1[4], 1'b0},
      {stage6_3[0], stage6_3[1], stage6_3[2], stage6_3[3], stage6_3[4], stage6_3[5]},
      {stage7_5[0],stage7_4[0],stage7_3[0],stage7_2[0],stage7_1[0]}
   );
   gpc15_3 gpc5081 (
      {stage6_5[0], stage6_5[1], stage6_5[2], stage6_5[3], stage6_5[4]},
      {stage6_6[0]},
      {stage7_7[0],stage7_6[0],stage7_5[1]}
   );
   gpc606_5 gpc5082 (
      {stage6_7[0], stage6_7[1], stage6_7[2], stage6_7[3], stage6_7[4], stage6_7[5]},
      {stage6_9[0], stage6_9[1], stage6_9[2], stage6_9[3], stage6_9[4], stage6_9[5]},
      {stage7_11[0],stage7_10[0],stage7_9[0],stage7_8[0],stage7_7[1]}
   );
   gpc1343_5 gpc5083 (
      {stage6_11[0], stage6_11[1], stage6_11[2]},
      {stage6_12[0], stage6_12[1], stage6_12[2], stage6_12[3]},
      {stage6_13[0], stage6_13[1], stage6_13[2]},
      {stage6_14[0]},
      {stage7_15[0],stage7_14[0],stage7_13[0],stage7_12[0],stage7_11[1]}
   );
   gpc615_5 gpc5084 (
      {stage6_11[3], stage6_11[4], stage6_11[5], stage6_11[6], stage6_11[7]},
      {stage6_12[4]},
      {stage6_13[3], stage6_13[4], stage6_13[5], stage6_13[6], stage6_13[7], stage6_13[8]},
      {stage7_15[1],stage7_14[1],stage7_13[1],stage7_12[1],stage7_11[2]}
   );
   gpc1343_5 gpc5085 (
      {stage6_16[0], stage6_16[1], stage6_16[2]},
      {stage6_17[0], stage6_17[1], stage6_17[2], stage6_17[3]},
      {stage6_18[0], stage6_18[1], stage6_18[2]},
      {stage6_19[0]},
      {stage7_20[0],stage7_19[0],stage7_18[0],stage7_17[0],stage7_16[0]}
   );
   gpc1343_5 gpc5086 (
      {stage6_16[3], stage6_16[4], stage6_16[5]},
      {stage6_17[4], stage6_17[5], stage6_17[6], stage6_17[7]},
      {stage6_18[3], stage6_18[4], stage6_18[5]},
      {stage6_19[1]},
      {stage7_20[1],stage7_19[1],stage7_18[1],stage7_17[1],stage7_16[1]}
   );
   gpc606_5 gpc5087 (
      {stage6_19[2], stage6_19[3], stage6_19[4], stage6_19[5], stage6_19[6], stage6_19[7]},
      {stage6_21[0], stage6_21[1], stage6_21[2], stage6_21[3], stage6_21[4], stage6_21[5]},
      {stage7_23[0],stage7_22[0],stage7_21[0],stage7_20[2],stage7_19[2]}
   );
   gpc606_5 gpc5088 (
      {stage6_19[8], stage6_19[9], stage6_19[10], stage6_19[11], stage6_19[12], stage6_19[13]},
      {stage6_21[6], stage6_21[7], stage6_21[8], stage6_21[9], stage6_21[10], stage6_21[11]},
      {stage7_23[1],stage7_22[1],stage7_21[1],stage7_20[3],stage7_19[3]}
   );
   gpc15_3 gpc5089 (
      {stage6_20[0], stage6_20[1], stage6_20[2], stage6_20[3], stage6_20[4]},
      {stage6_21[12]},
      {stage7_22[2],stage7_21[2],stage7_20[4]}
   );
   gpc606_5 gpc5090 (
      {stage6_22[0], stage6_22[1], stage6_22[2], stage6_22[3], stage6_22[4], stage6_22[5]},
      {stage6_24[0], stage6_24[1], stage6_24[2], stage6_24[3], stage6_24[4], stage6_24[5]},
      {stage7_26[0],stage7_25[0],stage7_24[0],stage7_23[2],stage7_22[3]}
   );
   gpc606_5 gpc5091 (
      {stage6_25[0], stage6_25[1], stage6_25[2], stage6_25[3], stage6_25[4], stage6_25[5]},
      {stage6_27[0], stage6_27[1], stage6_27[2], stage6_27[3], stage6_27[4], stage6_27[5]},
      {stage7_29[0],stage7_28[0],stage7_27[0],stage7_26[1],stage7_25[1]}
   );
   gpc15_3 gpc5092 (
      {stage6_26[0], stage6_26[1], stage6_26[2], stage6_26[3], stage6_26[4]},
      {stage6_27[6]},
      {stage7_28[1],stage7_27[1],stage7_26[2]}
   );
   gpc606_5 gpc5093 (
      {stage6_30[0], stage6_30[1], stage6_30[2], stage6_30[3], stage6_30[4], stage6_30[5]},
      {stage6_32[0], stage6_32[1], stage6_32[2], stage6_32[3], stage6_32[4], stage6_32[5]},
      {stage7_34[0],stage7_33[0],stage7_32[0],stage7_31[0],stage7_30[0]}
   );
   gpc606_5 gpc5094 (
      {stage6_33[0], stage6_33[1], stage6_33[2], stage6_33[3], stage6_33[4], stage6_33[5]},
      {stage6_35[0], stage6_35[1], stage6_35[2], stage6_35[3], stage6_35[4], stage6_35[5]},
      {stage7_37[0],stage7_36[0],stage7_35[0],stage7_34[1],stage7_33[1]}
   );
   gpc606_5 gpc5095 (
      {stage6_34[0], stage6_34[1], stage6_34[2], stage6_34[3], stage6_34[4], stage6_34[5]},
      {stage6_36[0], stage6_36[1], stage6_36[2], 1'b0, 1'b0, 1'b0},
      {stage7_38[0],stage7_37[1],stage7_36[1],stage7_35[1],stage7_34[2]}
   );
   gpc1_1 gpc5096 (
      {stage6_0[0]},
      {stage7_0[0]}
   );
   gpc1_1 gpc5097 (
      {stage6_0[1]},
      {stage7_0[1]}
   );
   gpc1_1 gpc5098 (
      {stage6_0[2]},
      {stage7_0[2]}
   );
   gpc1_1 gpc5099 (
      {stage6_0[3]},
      {stage7_0[3]}
   );
   gpc1_1 gpc5100 (
      {stage6_0[4]},
      {stage7_0[4]}
   );
   gpc1_1 gpc5101 (
      {stage6_0[5]},
      {stage7_0[5]}
   );
   gpc1_1 gpc5102 (
      {stage6_0[6]},
      {stage7_0[6]}
   );
   gpc1_1 gpc5103 (
      {stage6_2[0]},
      {stage7_2[1]}
   );
   gpc1_1 gpc5104 (
      {stage6_2[1]},
      {stage7_2[2]}
   );
   gpc1_1 gpc5105 (
      {stage6_2[2]},
      {stage7_2[3]}
   );
   gpc1_1 gpc5106 (
      {stage6_2[3]},
      {stage7_2[4]}
   );
   gpc1_1 gpc5107 (
      {stage6_2[4]},
      {stage7_2[5]}
   );
   gpc1_1 gpc5108 (
      {stage6_2[5]},
      {stage7_2[6]}
   );
   gpc1_1 gpc5109 (
      {stage6_4[0]},
      {stage7_4[1]}
   );
   gpc1_1 gpc5110 (
      {stage6_4[1]},
      {stage7_4[2]}
   );
   gpc1_1 gpc5111 (
      {stage6_4[2]},
      {stage7_4[3]}
   );
   gpc1_1 gpc5112 (
      {stage6_4[3]},
      {stage7_4[4]}
   );
   gpc1_1 gpc5113 (
      {stage6_4[4]},
      {stage7_4[5]}
   );
   gpc1_1 gpc5114 (
      {stage6_4[5]},
      {stage7_4[6]}
   );
   gpc1_1 gpc5115 (
      {stage6_6[1]},
      {stage7_6[1]}
   );
   gpc1_1 gpc5116 (
      {stage6_6[2]},
      {stage7_6[2]}
   );
   gpc1_1 gpc5117 (
      {stage6_6[3]},
      {stage7_6[3]}
   );
   gpc1_1 gpc5118 (
      {stage6_8[0]},
      {stage7_8[1]}
   );
   gpc1_1 gpc5119 (
      {stage6_8[1]},
      {stage7_8[2]}
   );
   gpc1_1 gpc5120 (
      {stage6_8[2]},
      {stage7_8[3]}
   );
   gpc1_1 gpc5121 (
      {stage6_8[3]},
      {stage7_8[4]}
   );
   gpc1_1 gpc5122 (
      {stage6_8[4]},
      {stage7_8[5]}
   );
   gpc1_1 gpc5123 (
      {stage6_8[5]},
      {stage7_8[6]}
   );
   gpc1_1 gpc5124 (
      {stage6_10[0]},
      {stage7_10[1]}
   );
   gpc1_1 gpc5125 (
      {stage6_10[1]},
      {stage7_10[2]}
   );
   gpc1_1 gpc5126 (
      {stage6_10[2]},
      {stage7_10[3]}
   );
   gpc1_1 gpc5127 (
      {stage6_10[3]},
      {stage7_10[4]}
   );
   gpc1_1 gpc5128 (
      {stage6_12[5]},
      {stage7_12[2]}
   );
   gpc1_1 gpc5129 (
      {stage6_12[6]},
      {stage7_12[3]}
   );
   gpc1_1 gpc5130 (
      {stage6_14[1]},
      {stage7_14[2]}
   );
   gpc1_1 gpc5131 (
      {stage6_14[2]},
      {stage7_14[3]}
   );
   gpc1_1 gpc5132 (
      {stage6_14[3]},
      {stage7_14[4]}
   );
   gpc1_1 gpc5133 (
      {stage6_14[4]},
      {stage7_14[5]}
   );
   gpc1_1 gpc5134 (
      {stage6_14[5]},
      {stage7_14[6]}
   );
   gpc1_1 gpc5135 (
      {stage6_15[0]},
      {stage7_15[2]}
   );
   gpc1_1 gpc5136 (
      {stage6_15[1]},
      {stage7_15[3]}
   );
   gpc1_1 gpc5137 (
      {stage6_15[2]},
      {stage7_15[4]}
   );
   gpc1_1 gpc5138 (
      {stage6_15[3]},
      {stage7_15[5]}
   );
   gpc1_1 gpc5139 (
      {stage6_17[8]},
      {stage7_17[2]}
   );
   gpc1_1 gpc5140 (
      {stage6_17[9]},
      {stage7_17[3]}
   );
   gpc1_1 gpc5141 (
      {stage6_19[14]},
      {stage7_19[4]}
   );
   gpc1_1 gpc5142 (
      {stage6_20[5]},
      {stage7_20[5]}
   );
   gpc1_1 gpc5143 (
      {stage6_22[6]},
      {stage7_22[4]}
   );
   gpc1_1 gpc5144 (
      {stage6_22[7]},
      {stage7_22[5]}
   );
   gpc1_1 gpc5145 (
      {stage6_23[0]},
      {stage7_23[3]}
   );
   gpc1_1 gpc5146 (
      {stage6_23[1]},
      {stage7_23[4]}
   );
   gpc1_1 gpc5147 (
      {stage6_23[2]},
      {stage7_23[5]}
   );
   gpc1_1 gpc5148 (
      {stage6_23[3]},
      {stage7_23[6]}
   );
   gpc1_1 gpc5149 (
      {stage6_27[7]},
      {stage7_27[2]}
   );
   gpc1_1 gpc5150 (
      {stage6_28[0]},
      {stage7_28[2]}
   );
   gpc1_1 gpc5151 (
      {stage6_28[1]},
      {stage7_28[3]}
   );
   gpc1_1 gpc5152 (
      {stage6_28[2]},
      {stage7_28[4]}
   );
   gpc1_1 gpc5153 (
      {stage6_28[3]},
      {stage7_28[5]}
   );
   gpc1_1 gpc5154 (
      {stage6_28[4]},
      {stage7_28[6]}
   );
   gpc1_1 gpc5155 (
      {stage6_29[0]},
      {stage7_29[1]}
   );
   gpc1_1 gpc5156 (
      {stage6_29[1]},
      {stage7_29[2]}
   );
   gpc1_1 gpc5157 (
      {stage6_29[2]},
      {stage7_29[3]}
   );
   gpc1_1 gpc5158 (
      {stage6_29[3]},
      {stage7_29[4]}
   );
   gpc1_1 gpc5159 (
      {stage6_31[0]},
      {stage7_31[1]}
   );
   gpc1_1 gpc5160 (
      {stage6_31[1]},
      {stage7_31[2]}
   );
   gpc1_1 gpc5161 (
      {stage6_31[2]},
      {stage7_31[3]}
   );
   gpc1_1 gpc5162 (
      {stage6_31[3]},
      {stage7_31[4]}
   );
   gpc1_1 gpc5163 (
      {stage6_31[4]},
      {stage7_31[5]}
   );
   gpc1_1 gpc5164 (
      {stage6_31[5]},
      {stage7_31[6]}
   );
   gpc1_1 gpc5165 (
      {stage6_31[6]},
      {stage7_31[7]}
   );
   gpc1_1 gpc5166 (
      {stage6_31[7]},
      {stage7_31[8]}
   );
   gpc1_1 gpc5167 (
      {stage6_34[6]},
      {stage7_34[3]}
   );
   gpc1_1 gpc5168 (
      {stage6_34[7]},
      {stage7_34[4]}
   );
   gpc1_1 gpc5169 (
      {stage6_34[8]},
      {stage7_34[5]}
   );
   gpc1_1 gpc5170 (
      {stage6_34[9]},
      {stage7_34[6]}
   );
   gpc1_1 gpc5171 (
      {stage6_37[0]},
      {stage7_37[2]}
   );
   gpc1_1 gpc5172 (
      {stage6_37[1]},
      {stage7_37[3]}
   );
   gpc1_1 gpc5173 (
      {stage6_38[0]},
      {stage7_38[1]}
   );
   gpc1_1 gpc5174 (
      {stage6_38[1]},
      {stage7_38[2]}
   );
   gpc1_1 gpc5175 (
      {stage6_39[0]},
      {stage7_39[0]}
   );
   gpc1_1 gpc5176 (
      {stage6_39[1]},
      {stage7_39[1]}
   );
   gpc1_1 gpc5177 (
      {stage6_40[0]},
      {stage7_40[0]}
   );
   gpc606_5 gpc5178 (
      {stage7_0[0], stage7_0[1], stage7_0[2], stage7_0[3], stage7_0[4], stage7_0[5]},
      {stage7_2[0], stage7_2[1], stage7_2[2], stage7_2[3], stage7_2[4], stage7_2[5]},
      {stage8_4[0],stage8_3[0],stage8_2[0],stage8_1[0],stage8_0[0]}
   );
   gpc117_4 gpc5179 (
      {stage7_4[0], stage7_4[1], stage7_4[2], stage7_4[3], stage7_4[4], stage7_4[5], stage7_4[6]},
      {stage7_5[0]},
      {stage7_6[0]},
      {stage8_7[0],stage8_6[0],stage8_5[0],stage8_4[1]}
   );
   gpc623_5 gpc5180 (
      {stage7_6[1], stage7_6[2], stage7_6[3]},
      {stage7_7[0], stage7_7[1]},
      {stage7_8[0], stage7_8[1], stage7_8[2], stage7_8[3], stage7_8[4], stage7_8[5]},
      {stage8_10[0],stage8_9[0],stage8_8[0],stage8_7[1],stage8_6[1]}
   );
   gpc1325_5 gpc5181 (
      {stage7_10[0], stage7_10[1], stage7_10[2], stage7_10[3], stage7_10[4]},
      {stage7_11[0], stage7_11[1]},
      {stage7_12[0], stage7_12[1], stage7_12[2]},
      {stage7_13[0]},
      {stage8_14[0],stage8_13[0],stage8_12[0],stage8_11[0],stage8_10[1]}
   );
   gpc117_4 gpc5182 (
      {stage7_14[0], stage7_14[1], stage7_14[2], stage7_14[3], stage7_14[4], stage7_14[5], stage7_14[6]},
      {stage7_15[0]},
      {stage7_16[0]},
      {stage8_17[0],stage8_16[0],stage8_15[0],stage8_14[1]}
   );
   gpc1415_5 gpc5183 (
      {stage7_15[1], stage7_15[2], stage7_15[3], stage7_15[4], stage7_15[5]},
      {stage7_16[1]},
      {stage7_17[0], stage7_17[1], stage7_17[2], stage7_17[3]},
      {stage7_18[0]},
      {stage8_19[0],stage8_18[0],stage8_17[1],stage8_16[1],stage8_15[1]}
   );
   gpc135_4 gpc5184 (
      {stage7_19[0], stage7_19[1], stage7_19[2], stage7_19[3], stage7_19[4]},
      {stage7_20[0], stage7_20[1], stage7_20[2]},
      {stage7_21[0]},
      {stage8_22[0],stage8_21[0],stage8_20[0],stage8_19[1]}
   );
   gpc623_5 gpc5185 (
      {stage7_20[3], stage7_20[4], stage7_20[5]},
      {stage7_21[1], stage7_21[2]},
      {stage7_22[0], stage7_22[1], stage7_22[2], stage7_22[3], stage7_22[4], stage7_22[5]},
      {stage8_24[0],stage8_23[0],stage8_22[1],stage8_21[1],stage8_20[1]}
   );
   gpc117_4 gpc5186 (
      {stage7_23[0], stage7_23[1], stage7_23[2], stage7_23[3], stage7_23[4], stage7_23[5], stage7_23[6]},
      {stage7_24[0]},
      {stage7_25[0]},
      {stage8_26[0],stage8_25[0],stage8_24[1],stage8_23[1]}
   );
   gpc2223_5 gpc5187 (
      {stage7_26[0], stage7_26[1], stage7_26[2]},
      {stage7_27[0], stage7_27[1]},
      {stage7_28[0], stage7_28[1]},
      {stage7_29[0], stage7_29[1]},
      {stage8_30[0],stage8_29[0],stage8_28[0],stage8_27[0],stage8_26[1]}
   );
   gpc2135_5 gpc5188 (
      {stage7_28[2], stage7_28[3], stage7_28[4], stage7_28[5], stage7_28[6]},
      {stage7_29[2], stage7_29[3], stage7_29[4]},
      {stage7_30[0]},
      {stage7_31[0], stage7_31[1]},
      {stage8_32[0],stage8_31[0],stage8_30[1],stage8_29[1],stage8_28[1]}
   );
   gpc117_4 gpc5189 (
      {stage7_31[2], stage7_31[3], stage7_31[4], stage7_31[5], stage7_31[6], stage7_31[7], stage7_31[8]},
      {stage7_32[0]},
      {stage7_33[0]},
      {stage8_34[0],stage8_33[0],stage8_32[1],stage8_31[1]}
   );
   gpc117_4 gpc5190 (
      {stage7_34[0], stage7_34[1], stage7_34[2], stage7_34[3], stage7_34[4], stage7_34[5], stage7_34[6]},
      {stage7_35[0]},
      {stage7_36[0]},
      {stage8_37[0],stage8_36[0],stage8_35[0],stage8_34[1]}
   );
   gpc615_5 gpc5191 (
      {stage7_35[1], 1'b0, 1'b0, 1'b0, 1'b0},
      {stage7_36[1]},
      {stage7_37[0], stage7_37[1], stage7_37[2], stage7_37[3], 1'b0, 1'b0},
      {stage8_39[0],stage8_38[0],stage8_37[1],stage8_36[1],stage8_35[1]}
   );
   gpc1163_5 gpc5192 (
      {stage7_38[0], stage7_38[1], stage7_38[2]},
      {stage7_39[0], stage7_39[1], 1'b0, 1'b0, 1'b0, 1'b0},
      {stage7_40[0]},
      {1'b0},
      {stage8_40[0],stage8_39[1],stage8_38[1]}
   );
   gpc1_1 gpc5193 (
      {stage7_0[6]},
      {stage8_0[1]}
   );
   gpc1_1 gpc5194 (
      {stage7_1[0]},
      {stage8_1[1]}
   );
   gpc1_1 gpc5195 (
      {stage7_2[6]},
      {stage8_2[1]}
   );
   gpc1_1 gpc5196 (
      {stage7_3[0]},
      {stage8_3[1]}
   );
   gpc1_1 gpc5197 (
      {stage7_5[1]},
      {stage8_5[1]}
   );
   gpc1_1 gpc5198 (
      {stage7_8[6]},
      {stage8_8[1]}
   );
   gpc1_1 gpc5199 (
      {stage7_9[0]},
      {stage8_9[1]}
   );
   gpc1_1 gpc5200 (
      {stage7_11[2]},
      {stage8_11[1]}
   );
   gpc1_1 gpc5201 (
      {stage7_12[3]},
      {stage8_12[1]}
   );
   gpc1_1 gpc5202 (
      {stage7_13[1]},
      {stage8_13[1]}
   );
   gpc1_1 gpc5203 (
      {stage7_18[1]},
      {stage8_18[1]}
   );
   gpc1_1 gpc5204 (
      {stage7_25[1]},
      {stage8_25[1]}
   );
   gpc1_1 gpc5205 (
      {stage7_27[2]},
      {stage8_27[1]}
   );
   gpc1_1 gpc5206 (
      {stage7_33[1]},
      {stage8_33[1]}
   );
endmodule
module rowadder2_1_41(input [40:0] src0, input [40:0] src1, output [41:0] dst0);
    wire [40:0] gene;
    wire [40:0] prop;
    wire [43:0] out;
    wire [43:0] carryout;
    LUT2 #(
        .INIT(4'h8)
    ) lut_0_gene (
        .I0(src0[0]),
        .I1(src1[0]),
        .O(gene[0])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_0_prop (
        .I0(src0[0]),
        .I1(src1[0]),
        .O(prop[0])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_1_gene (
        .I0(src0[1]),
        .I1(src1[1]),
        .O(gene[1])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_1_prop (
        .I0(src0[1]),
        .I1(src1[1]),
        .O(prop[1])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_2_gene (
        .I0(src0[2]),
        .I1(src1[2]),
        .O(gene[2])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_2_prop (
        .I0(src0[2]),
        .I1(src1[2]),
        .O(prop[2])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_3_gene (
        .I0(src0[3]),
        .I1(src1[3]),
        .O(gene[3])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_3_prop (
        .I0(src0[3]),
        .I1(src1[3]),
        .O(prop[3])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_4_gene (
        .I0(src0[4]),
        .I1(src1[4]),
        .O(gene[4])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_4_prop (
        .I0(src0[4]),
        .I1(src1[4]),
        .O(prop[4])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_5_gene (
        .I0(src0[5]),
        .I1(src1[5]),
        .O(gene[5])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_5_prop (
        .I0(src0[5]),
        .I1(src1[5]),
        .O(prop[5])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_6_gene (
        .I0(src0[6]),
        .I1(src1[6]),
        .O(gene[6])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_6_prop (
        .I0(src0[6]),
        .I1(src1[6]),
        .O(prop[6])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_7_gene (
        .I0(src0[7]),
        .I1(src1[7]),
        .O(gene[7])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_7_prop (
        .I0(src0[7]),
        .I1(src1[7]),
        .O(prop[7])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_8_gene (
        .I0(src0[8]),
        .I1(src1[8]),
        .O(gene[8])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_8_prop (
        .I0(src0[8]),
        .I1(src1[8]),
        .O(prop[8])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_9_gene (
        .I0(src0[9]),
        .I1(src1[9]),
        .O(gene[9])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_9_prop (
        .I0(src0[9]),
        .I1(src1[9]),
        .O(prop[9])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_10_gene (
        .I0(src0[10]),
        .I1(src1[10]),
        .O(gene[10])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_10_prop (
        .I0(src0[10]),
        .I1(src1[10]),
        .O(prop[10])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_11_gene (
        .I0(src0[11]),
        .I1(src1[11]),
        .O(gene[11])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_11_prop (
        .I0(src0[11]),
        .I1(src1[11]),
        .O(prop[11])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_12_gene (
        .I0(src0[12]),
        .I1(src1[12]),
        .O(gene[12])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_12_prop (
        .I0(src0[12]),
        .I1(src1[12]),
        .O(prop[12])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_13_gene (
        .I0(src0[13]),
        .I1(src1[13]),
        .O(gene[13])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_13_prop (
        .I0(src0[13]),
        .I1(src1[13]),
        .O(prop[13])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_14_gene (
        .I0(src0[14]),
        .I1(src1[14]),
        .O(gene[14])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_14_prop (
        .I0(src0[14]),
        .I1(src1[14]),
        .O(prop[14])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_15_gene (
        .I0(src0[15]),
        .I1(src1[15]),
        .O(gene[15])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_15_prop (
        .I0(src0[15]),
        .I1(src1[15]),
        .O(prop[15])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_16_gene (
        .I0(src0[16]),
        .I1(src1[16]),
        .O(gene[16])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_16_prop (
        .I0(src0[16]),
        .I1(src1[16]),
        .O(prop[16])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_17_gene (
        .I0(src0[17]),
        .I1(src1[17]),
        .O(gene[17])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_17_prop (
        .I0(src0[17]),
        .I1(src1[17]),
        .O(prop[17])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_18_gene (
        .I0(src0[18]),
        .I1(src1[18]),
        .O(gene[18])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_18_prop (
        .I0(src0[18]),
        .I1(src1[18]),
        .O(prop[18])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_19_gene (
        .I0(src0[19]),
        .I1(src1[19]),
        .O(gene[19])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_19_prop (
        .I0(src0[19]),
        .I1(src1[19]),
        .O(prop[19])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_20_gene (
        .I0(src0[20]),
        .I1(src1[20]),
        .O(gene[20])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_20_prop (
        .I0(src0[20]),
        .I1(src1[20]),
        .O(prop[20])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_21_gene (
        .I0(src0[21]),
        .I1(src1[21]),
        .O(gene[21])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_21_prop (
        .I0(src0[21]),
        .I1(src1[21]),
        .O(prop[21])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_22_gene (
        .I0(src0[22]),
        .I1(src1[22]),
        .O(gene[22])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_22_prop (
        .I0(src0[22]),
        .I1(src1[22]),
        .O(prop[22])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_23_gene (
        .I0(src0[23]),
        .I1(src1[23]),
        .O(gene[23])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_23_prop (
        .I0(src0[23]),
        .I1(src1[23]),
        .O(prop[23])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_24_gene (
        .I0(src0[24]),
        .I1(src1[24]),
        .O(gene[24])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_24_prop (
        .I0(src0[24]),
        .I1(src1[24]),
        .O(prop[24])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_25_gene (
        .I0(src0[25]),
        .I1(src1[25]),
        .O(gene[25])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_25_prop (
        .I0(src0[25]),
        .I1(src1[25]),
        .O(prop[25])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_26_gene (
        .I0(src0[26]),
        .I1(src1[26]),
        .O(gene[26])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_26_prop (
        .I0(src0[26]),
        .I1(src1[26]),
        .O(prop[26])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_27_gene (
        .I0(src0[27]),
        .I1(src1[27]),
        .O(gene[27])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_27_prop (
        .I0(src0[27]),
        .I1(src1[27]),
        .O(prop[27])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_28_gene (
        .I0(src0[28]),
        .I1(src1[28]),
        .O(gene[28])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_28_prop (
        .I0(src0[28]),
        .I1(src1[28]),
        .O(prop[28])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_29_gene (
        .I0(src0[29]),
        .I1(src1[29]),
        .O(gene[29])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_29_prop (
        .I0(src0[29]),
        .I1(src1[29]),
        .O(prop[29])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_30_gene (
        .I0(src0[30]),
        .I1(src1[30]),
        .O(gene[30])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_30_prop (
        .I0(src0[30]),
        .I1(src1[30]),
        .O(prop[30])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_31_gene (
        .I0(src0[31]),
        .I1(src1[31]),
        .O(gene[31])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_31_prop (
        .I0(src0[31]),
        .I1(src1[31]),
        .O(prop[31])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_32_gene (
        .I0(src0[32]),
        .I1(src1[32]),
        .O(gene[32])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_32_prop (
        .I0(src0[32]),
        .I1(src1[32]),
        .O(prop[32])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_33_gene (
        .I0(src0[33]),
        .I1(src1[33]),
        .O(gene[33])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_33_prop (
        .I0(src0[33]),
        .I1(src1[33]),
        .O(prop[33])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_34_gene (
        .I0(src0[34]),
        .I1(src1[34]),
        .O(gene[34])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_34_prop (
        .I0(src0[34]),
        .I1(src1[34]),
        .O(prop[34])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_35_gene (
        .I0(src0[35]),
        .I1(src1[35]),
        .O(gene[35])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_35_prop (
        .I0(src0[35]),
        .I1(src1[35]),
        .O(prop[35])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_36_gene (
        .I0(src0[36]),
        .I1(src1[36]),
        .O(gene[36])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_36_prop (
        .I0(src0[36]),
        .I1(src1[36]),
        .O(prop[36])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_37_gene (
        .I0(src0[37]),
        .I1(src1[37]),
        .O(gene[37])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_37_prop (
        .I0(src0[37]),
        .I1(src1[37]),
        .O(prop[37])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_38_gene (
        .I0(src0[38]),
        .I1(src1[38]),
        .O(gene[38])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_38_prop (
        .I0(src0[38]),
        .I1(src1[38]),
        .O(prop[38])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_39_gene (
        .I0(src0[39]),
        .I1(src1[39]),
        .O(gene[39])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_39_prop (
        .I0(src0[39]),
        .I1(src1[39]),
        .O(prop[39])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_40_gene (
        .I0(src0[40]),
        .I1(src1[40]),
        .O(gene[40])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_40_prop (
        .I0(src0[40]),
        .I1(src1[40]),
        .O(prop[40])
    );
    CARRY4 carry4_3_0 (
        .CO(carryout[3:0]),
        .O(out[3:0]),
        .CI(1'h0),
        .CYINIT(1'h0),
        .DI(gene[3:0]),
        .S(prop[3:0])
    );
    CARRY4 carry4_7_4 (
        .CO(carryout[7:4]),
        .O(out[7:4]),
        .CI(carryout[3]),
        .CYINIT(1'h0),
        .DI(gene[7:4]),
        .S(prop[7:4])
    );
    CARRY4 carry4_11_8 (
        .CO(carryout[11:8]),
        .O(out[11:8]),
        .CI(carryout[7]),
        .CYINIT(1'h0),
        .DI(gene[11:8]),
        .S(prop[11:8])
    );
    CARRY4 carry4_15_12 (
        .CO(carryout[15:12]),
        .O(out[15:12]),
        .CI(carryout[11]),
        .CYINIT(1'h0),
        .DI(gene[15:12]),
        .S(prop[15:12])
    );
    CARRY4 carry4_19_16 (
        .CO(carryout[19:16]),
        .O(out[19:16]),
        .CI(carryout[15]),
        .CYINIT(1'h0),
        .DI(gene[19:16]),
        .S(prop[19:16])
    );
    CARRY4 carry4_23_20 (
        .CO(carryout[23:20]),
        .O(out[23:20]),
        .CI(carryout[19]),
        .CYINIT(1'h0),
        .DI(gene[23:20]),
        .S(prop[23:20])
    );
    CARRY4 carry4_27_24 (
        .CO(carryout[27:24]),
        .O(out[27:24]),
        .CI(carryout[23]),
        .CYINIT(1'h0),
        .DI(gene[27:24]),
        .S(prop[27:24])
    );
    CARRY4 carry4_31_28 (
        .CO(carryout[31:28]),
        .O(out[31:28]),
        .CI(carryout[27]),
        .CYINIT(1'h0),
        .DI(gene[31:28]),
        .S(prop[31:28])
    );
    CARRY4 carry4_35_32 (
        .CO(carryout[35:32]),
        .O(out[35:32]),
        .CI(carryout[31]),
        .CYINIT(1'h0),
        .DI(gene[35:32]),
        .S(prop[35:32])
    );
    CARRY4 carry4_39_36 (
        .CO(carryout[39:36]),
        .O(out[39:36]),
        .CI(carryout[35]),
        .CYINIT(1'h0),
        .DI(gene[39:36]),
        .S(prop[39:36])
    );
    CARRY4 carry4_43_40 (
        .CO(carryout[43:40]),
        .O(out[43:40]),
        .CI(carryout[39]),
        .CYINIT(1'h0),
        .DI({3'h0, gene[40:40]}),
        .S({3'h0, prop[40:40]})
    );
    assign dst0 = {carryout[40], out[40:0]};
endmodule


module testbench();
    reg [511:0] src0;
    reg [511:0] src1;
    reg [511:0] src2;
    reg [511:0] src3;
    reg [511:0] src4;
    reg [511:0] src5;
    reg [511:0] src6;
    reg [511:0] src7;
    reg [511:0] src8;
    reg [511:0] src9;
    reg [511:0] src10;
    reg [511:0] src11;
    reg [511:0] src12;
    reg [511:0] src13;
    reg [511:0] src14;
    reg [511:0] src15;
    reg [511:0] src16;
    reg [511:0] src17;
    reg [511:0] src18;
    reg [511:0] src19;
    reg [511:0] src20;
    reg [511:0] src21;
    reg [511:0] src22;
    reg [511:0] src23;
    reg [511:0] src24;
    reg [511:0] src25;
    reg [511:0] src26;
    reg [511:0] src27;
    reg [511:0] src28;
    reg [511:0] src29;
    reg [511:0] src30;
    reg [511:0] src31;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [0:0] dst26;
    wire [0:0] dst27;
    wire [0:0] dst28;
    wire [0:0] dst29;
    wire [0:0] dst30;
    wire [0:0] dst31;
    wire [0:0] dst32;
    wire [0:0] dst33;
    wire [0:0] dst34;
    wire [0:0] dst35;
    wire [0:0] dst36;
    wire [0:0] dst37;
    wire [0:0] dst38;
    wire [0:0] dst39;
    wire [0:0] dst40;
    wire [40:0] srcsum;
    wire [40:0] dstsum;
    wire test;
    compressor2_1_512_32 compressor2_1_512_32(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .src31(src31),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25),
        .dst26(dst26),
        .dst27(dst27),
        .dst28(dst28),
        .dst29(dst29),
        .dst30(dst30),
        .dst31(dst31),
        .dst32(dst32),
        .dst33(dst33),
        .dst34(dst34),
        .dst35(dst35),
        .dst36(dst36),
        .dst37(dst37),
        .dst38(dst38),
        .dst39(dst39),
        .dst40(dst40));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13] + src0[14] + src0[15] + src0[16] + src0[17] + src0[18] + src0[19] + src0[20] + src0[21] + src0[22] + src0[23] + src0[24] + src0[25] + src0[26] + src0[27] + src0[28] + src0[29] + src0[30] + src0[31] + src0[32] + src0[33] + src0[34] + src0[35] + src0[36] + src0[37] + src0[38] + src0[39] + src0[40] + src0[41] + src0[42] + src0[43] + src0[44] + src0[45] + src0[46] + src0[47] + src0[48] + src0[49] + src0[50] + src0[51] + src0[52] + src0[53] + src0[54] + src0[55] + src0[56] + src0[57] + src0[58] + src0[59] + src0[60] + src0[61] + src0[62] + src0[63] + src0[64] + src0[65] + src0[66] + src0[67] + src0[68] + src0[69] + src0[70] + src0[71] + src0[72] + src0[73] + src0[74] + src0[75] + src0[76] + src0[77] + src0[78] + src0[79] + src0[80] + src0[81] + src0[82] + src0[83] + src0[84] + src0[85] + src0[86] + src0[87] + src0[88] + src0[89] + src0[90] + src0[91] + src0[92] + src0[93] + src0[94] + src0[95] + src0[96] + src0[97] + src0[98] + src0[99] + src0[100] + src0[101] + src0[102] + src0[103] + src0[104] + src0[105] + src0[106] + src0[107] + src0[108] + src0[109] + src0[110] + src0[111] + src0[112] + src0[113] + src0[114] + src0[115] + src0[116] + src0[117] + src0[118] + src0[119] + src0[120] + src0[121] + src0[122] + src0[123] + src0[124] + src0[125] + src0[126] + src0[127] + src0[128] + src0[129] + src0[130] + src0[131] + src0[132] + src0[133] + src0[134] + src0[135] + src0[136] + src0[137] + src0[138] + src0[139] + src0[140] + src0[141] + src0[142] + src0[143] + src0[144] + src0[145] + src0[146] + src0[147] + src0[148] + src0[149] + src0[150] + src0[151] + src0[152] + src0[153] + src0[154] + src0[155] + src0[156] + src0[157] + src0[158] + src0[159] + src0[160] + src0[161] + src0[162] + src0[163] + src0[164] + src0[165] + src0[166] + src0[167] + src0[168] + src0[169] + src0[170] + src0[171] + src0[172] + src0[173] + src0[174] + src0[175] + src0[176] + src0[177] + src0[178] + src0[179] + src0[180] + src0[181] + src0[182] + src0[183] + src0[184] + src0[185] + src0[186] + src0[187] + src0[188] + src0[189] + src0[190] + src0[191] + src0[192] + src0[193] + src0[194] + src0[195] + src0[196] + src0[197] + src0[198] + src0[199] + src0[200] + src0[201] + src0[202] + src0[203] + src0[204] + src0[205] + src0[206] + src0[207] + src0[208] + src0[209] + src0[210] + src0[211] + src0[212] + src0[213] + src0[214] + src0[215] + src0[216] + src0[217] + src0[218] + src0[219] + src0[220] + src0[221] + src0[222] + src0[223] + src0[224] + src0[225] + src0[226] + src0[227] + src0[228] + src0[229] + src0[230] + src0[231] + src0[232] + src0[233] + src0[234] + src0[235] + src0[236] + src0[237] + src0[238] + src0[239] + src0[240] + src0[241] + src0[242] + src0[243] + src0[244] + src0[245] + src0[246] + src0[247] + src0[248] + src0[249] + src0[250] + src0[251] + src0[252] + src0[253] + src0[254] + src0[255] + src0[256] + src0[257] + src0[258] + src0[259] + src0[260] + src0[261] + src0[262] + src0[263] + src0[264] + src0[265] + src0[266] + src0[267] + src0[268] + src0[269] + src0[270] + src0[271] + src0[272] + src0[273] + src0[274] + src0[275] + src0[276] + src0[277] + src0[278] + src0[279] + src0[280] + src0[281] + src0[282] + src0[283] + src0[284] + src0[285] + src0[286] + src0[287] + src0[288] + src0[289] + src0[290] + src0[291] + src0[292] + src0[293] + src0[294] + src0[295] + src0[296] + src0[297] + src0[298] + src0[299] + src0[300] + src0[301] + src0[302] + src0[303] + src0[304] + src0[305] + src0[306] + src0[307] + src0[308] + src0[309] + src0[310] + src0[311] + src0[312] + src0[313] + src0[314] + src0[315] + src0[316] + src0[317] + src0[318] + src0[319] + src0[320] + src0[321] + src0[322] + src0[323] + src0[324] + src0[325] + src0[326] + src0[327] + src0[328] + src0[329] + src0[330] + src0[331] + src0[332] + src0[333] + src0[334] + src0[335] + src0[336] + src0[337] + src0[338] + src0[339] + src0[340] + src0[341] + src0[342] + src0[343] + src0[344] + src0[345] + src0[346] + src0[347] + src0[348] + src0[349] + src0[350] + src0[351] + src0[352] + src0[353] + src0[354] + src0[355] + src0[356] + src0[357] + src0[358] + src0[359] + src0[360] + src0[361] + src0[362] + src0[363] + src0[364] + src0[365] + src0[366] + src0[367] + src0[368] + src0[369] + src0[370] + src0[371] + src0[372] + src0[373] + src0[374] + src0[375] + src0[376] + src0[377] + src0[378] + src0[379] + src0[380] + src0[381] + src0[382] + src0[383] + src0[384] + src0[385] + src0[386] + src0[387] + src0[388] + src0[389] + src0[390] + src0[391] + src0[392] + src0[393] + src0[394] + src0[395] + src0[396] + src0[397] + src0[398] + src0[399] + src0[400] + src0[401] + src0[402] + src0[403] + src0[404] + src0[405] + src0[406] + src0[407] + src0[408] + src0[409] + src0[410] + src0[411] + src0[412] + src0[413] + src0[414] + src0[415] + src0[416] + src0[417] + src0[418] + src0[419] + src0[420] + src0[421] + src0[422] + src0[423] + src0[424] + src0[425] + src0[426] + src0[427] + src0[428] + src0[429] + src0[430] + src0[431] + src0[432] + src0[433] + src0[434] + src0[435] + src0[436] + src0[437] + src0[438] + src0[439] + src0[440] + src0[441] + src0[442] + src0[443] + src0[444] + src0[445] + src0[446] + src0[447] + src0[448] + src0[449] + src0[450] + src0[451] + src0[452] + src0[453] + src0[454] + src0[455] + src0[456] + src0[457] + src0[458] + src0[459] + src0[460] + src0[461] + src0[462] + src0[463] + src0[464] + src0[465] + src0[466] + src0[467] + src0[468] + src0[469] + src0[470] + src0[471] + src0[472] + src0[473] + src0[474] + src0[475] + src0[476] + src0[477] + src0[478] + src0[479] + src0[480] + src0[481] + src0[482] + src0[483] + src0[484] + src0[485] + src0[486] + src0[487] + src0[488] + src0[489] + src0[490] + src0[491] + src0[492] + src0[493] + src0[494] + src0[495] + src0[496] + src0[497] + src0[498] + src0[499] + src0[500] + src0[501] + src0[502] + src0[503] + src0[504] + src0[505] + src0[506] + src0[507] + src0[508] + src0[509] + src0[510] + src0[511])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13] + src1[14] + src1[15] + src1[16] + src1[17] + src1[18] + src1[19] + src1[20] + src1[21] + src1[22] + src1[23] + src1[24] + src1[25] + src1[26] + src1[27] + src1[28] + src1[29] + src1[30] + src1[31] + src1[32] + src1[33] + src1[34] + src1[35] + src1[36] + src1[37] + src1[38] + src1[39] + src1[40] + src1[41] + src1[42] + src1[43] + src1[44] + src1[45] + src1[46] + src1[47] + src1[48] + src1[49] + src1[50] + src1[51] + src1[52] + src1[53] + src1[54] + src1[55] + src1[56] + src1[57] + src1[58] + src1[59] + src1[60] + src1[61] + src1[62] + src1[63] + src1[64] + src1[65] + src1[66] + src1[67] + src1[68] + src1[69] + src1[70] + src1[71] + src1[72] + src1[73] + src1[74] + src1[75] + src1[76] + src1[77] + src1[78] + src1[79] + src1[80] + src1[81] + src1[82] + src1[83] + src1[84] + src1[85] + src1[86] + src1[87] + src1[88] + src1[89] + src1[90] + src1[91] + src1[92] + src1[93] + src1[94] + src1[95] + src1[96] + src1[97] + src1[98] + src1[99] + src1[100] + src1[101] + src1[102] + src1[103] + src1[104] + src1[105] + src1[106] + src1[107] + src1[108] + src1[109] + src1[110] + src1[111] + src1[112] + src1[113] + src1[114] + src1[115] + src1[116] + src1[117] + src1[118] + src1[119] + src1[120] + src1[121] + src1[122] + src1[123] + src1[124] + src1[125] + src1[126] + src1[127] + src1[128] + src1[129] + src1[130] + src1[131] + src1[132] + src1[133] + src1[134] + src1[135] + src1[136] + src1[137] + src1[138] + src1[139] + src1[140] + src1[141] + src1[142] + src1[143] + src1[144] + src1[145] + src1[146] + src1[147] + src1[148] + src1[149] + src1[150] + src1[151] + src1[152] + src1[153] + src1[154] + src1[155] + src1[156] + src1[157] + src1[158] + src1[159] + src1[160] + src1[161] + src1[162] + src1[163] + src1[164] + src1[165] + src1[166] + src1[167] + src1[168] + src1[169] + src1[170] + src1[171] + src1[172] + src1[173] + src1[174] + src1[175] + src1[176] + src1[177] + src1[178] + src1[179] + src1[180] + src1[181] + src1[182] + src1[183] + src1[184] + src1[185] + src1[186] + src1[187] + src1[188] + src1[189] + src1[190] + src1[191] + src1[192] + src1[193] + src1[194] + src1[195] + src1[196] + src1[197] + src1[198] + src1[199] + src1[200] + src1[201] + src1[202] + src1[203] + src1[204] + src1[205] + src1[206] + src1[207] + src1[208] + src1[209] + src1[210] + src1[211] + src1[212] + src1[213] + src1[214] + src1[215] + src1[216] + src1[217] + src1[218] + src1[219] + src1[220] + src1[221] + src1[222] + src1[223] + src1[224] + src1[225] + src1[226] + src1[227] + src1[228] + src1[229] + src1[230] + src1[231] + src1[232] + src1[233] + src1[234] + src1[235] + src1[236] + src1[237] + src1[238] + src1[239] + src1[240] + src1[241] + src1[242] + src1[243] + src1[244] + src1[245] + src1[246] + src1[247] + src1[248] + src1[249] + src1[250] + src1[251] + src1[252] + src1[253] + src1[254] + src1[255] + src1[256] + src1[257] + src1[258] + src1[259] + src1[260] + src1[261] + src1[262] + src1[263] + src1[264] + src1[265] + src1[266] + src1[267] + src1[268] + src1[269] + src1[270] + src1[271] + src1[272] + src1[273] + src1[274] + src1[275] + src1[276] + src1[277] + src1[278] + src1[279] + src1[280] + src1[281] + src1[282] + src1[283] + src1[284] + src1[285] + src1[286] + src1[287] + src1[288] + src1[289] + src1[290] + src1[291] + src1[292] + src1[293] + src1[294] + src1[295] + src1[296] + src1[297] + src1[298] + src1[299] + src1[300] + src1[301] + src1[302] + src1[303] + src1[304] + src1[305] + src1[306] + src1[307] + src1[308] + src1[309] + src1[310] + src1[311] + src1[312] + src1[313] + src1[314] + src1[315] + src1[316] + src1[317] + src1[318] + src1[319] + src1[320] + src1[321] + src1[322] + src1[323] + src1[324] + src1[325] + src1[326] + src1[327] + src1[328] + src1[329] + src1[330] + src1[331] + src1[332] + src1[333] + src1[334] + src1[335] + src1[336] + src1[337] + src1[338] + src1[339] + src1[340] + src1[341] + src1[342] + src1[343] + src1[344] + src1[345] + src1[346] + src1[347] + src1[348] + src1[349] + src1[350] + src1[351] + src1[352] + src1[353] + src1[354] + src1[355] + src1[356] + src1[357] + src1[358] + src1[359] + src1[360] + src1[361] + src1[362] + src1[363] + src1[364] + src1[365] + src1[366] + src1[367] + src1[368] + src1[369] + src1[370] + src1[371] + src1[372] + src1[373] + src1[374] + src1[375] + src1[376] + src1[377] + src1[378] + src1[379] + src1[380] + src1[381] + src1[382] + src1[383] + src1[384] + src1[385] + src1[386] + src1[387] + src1[388] + src1[389] + src1[390] + src1[391] + src1[392] + src1[393] + src1[394] + src1[395] + src1[396] + src1[397] + src1[398] + src1[399] + src1[400] + src1[401] + src1[402] + src1[403] + src1[404] + src1[405] + src1[406] + src1[407] + src1[408] + src1[409] + src1[410] + src1[411] + src1[412] + src1[413] + src1[414] + src1[415] + src1[416] + src1[417] + src1[418] + src1[419] + src1[420] + src1[421] + src1[422] + src1[423] + src1[424] + src1[425] + src1[426] + src1[427] + src1[428] + src1[429] + src1[430] + src1[431] + src1[432] + src1[433] + src1[434] + src1[435] + src1[436] + src1[437] + src1[438] + src1[439] + src1[440] + src1[441] + src1[442] + src1[443] + src1[444] + src1[445] + src1[446] + src1[447] + src1[448] + src1[449] + src1[450] + src1[451] + src1[452] + src1[453] + src1[454] + src1[455] + src1[456] + src1[457] + src1[458] + src1[459] + src1[460] + src1[461] + src1[462] + src1[463] + src1[464] + src1[465] + src1[466] + src1[467] + src1[468] + src1[469] + src1[470] + src1[471] + src1[472] + src1[473] + src1[474] + src1[475] + src1[476] + src1[477] + src1[478] + src1[479] + src1[480] + src1[481] + src1[482] + src1[483] + src1[484] + src1[485] + src1[486] + src1[487] + src1[488] + src1[489] + src1[490] + src1[491] + src1[492] + src1[493] + src1[494] + src1[495] + src1[496] + src1[497] + src1[498] + src1[499] + src1[500] + src1[501] + src1[502] + src1[503] + src1[504] + src1[505] + src1[506] + src1[507] + src1[508] + src1[509] + src1[510] + src1[511])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13] + src2[14] + src2[15] + src2[16] + src2[17] + src2[18] + src2[19] + src2[20] + src2[21] + src2[22] + src2[23] + src2[24] + src2[25] + src2[26] + src2[27] + src2[28] + src2[29] + src2[30] + src2[31] + src2[32] + src2[33] + src2[34] + src2[35] + src2[36] + src2[37] + src2[38] + src2[39] + src2[40] + src2[41] + src2[42] + src2[43] + src2[44] + src2[45] + src2[46] + src2[47] + src2[48] + src2[49] + src2[50] + src2[51] + src2[52] + src2[53] + src2[54] + src2[55] + src2[56] + src2[57] + src2[58] + src2[59] + src2[60] + src2[61] + src2[62] + src2[63] + src2[64] + src2[65] + src2[66] + src2[67] + src2[68] + src2[69] + src2[70] + src2[71] + src2[72] + src2[73] + src2[74] + src2[75] + src2[76] + src2[77] + src2[78] + src2[79] + src2[80] + src2[81] + src2[82] + src2[83] + src2[84] + src2[85] + src2[86] + src2[87] + src2[88] + src2[89] + src2[90] + src2[91] + src2[92] + src2[93] + src2[94] + src2[95] + src2[96] + src2[97] + src2[98] + src2[99] + src2[100] + src2[101] + src2[102] + src2[103] + src2[104] + src2[105] + src2[106] + src2[107] + src2[108] + src2[109] + src2[110] + src2[111] + src2[112] + src2[113] + src2[114] + src2[115] + src2[116] + src2[117] + src2[118] + src2[119] + src2[120] + src2[121] + src2[122] + src2[123] + src2[124] + src2[125] + src2[126] + src2[127] + src2[128] + src2[129] + src2[130] + src2[131] + src2[132] + src2[133] + src2[134] + src2[135] + src2[136] + src2[137] + src2[138] + src2[139] + src2[140] + src2[141] + src2[142] + src2[143] + src2[144] + src2[145] + src2[146] + src2[147] + src2[148] + src2[149] + src2[150] + src2[151] + src2[152] + src2[153] + src2[154] + src2[155] + src2[156] + src2[157] + src2[158] + src2[159] + src2[160] + src2[161] + src2[162] + src2[163] + src2[164] + src2[165] + src2[166] + src2[167] + src2[168] + src2[169] + src2[170] + src2[171] + src2[172] + src2[173] + src2[174] + src2[175] + src2[176] + src2[177] + src2[178] + src2[179] + src2[180] + src2[181] + src2[182] + src2[183] + src2[184] + src2[185] + src2[186] + src2[187] + src2[188] + src2[189] + src2[190] + src2[191] + src2[192] + src2[193] + src2[194] + src2[195] + src2[196] + src2[197] + src2[198] + src2[199] + src2[200] + src2[201] + src2[202] + src2[203] + src2[204] + src2[205] + src2[206] + src2[207] + src2[208] + src2[209] + src2[210] + src2[211] + src2[212] + src2[213] + src2[214] + src2[215] + src2[216] + src2[217] + src2[218] + src2[219] + src2[220] + src2[221] + src2[222] + src2[223] + src2[224] + src2[225] + src2[226] + src2[227] + src2[228] + src2[229] + src2[230] + src2[231] + src2[232] + src2[233] + src2[234] + src2[235] + src2[236] + src2[237] + src2[238] + src2[239] + src2[240] + src2[241] + src2[242] + src2[243] + src2[244] + src2[245] + src2[246] + src2[247] + src2[248] + src2[249] + src2[250] + src2[251] + src2[252] + src2[253] + src2[254] + src2[255] + src2[256] + src2[257] + src2[258] + src2[259] + src2[260] + src2[261] + src2[262] + src2[263] + src2[264] + src2[265] + src2[266] + src2[267] + src2[268] + src2[269] + src2[270] + src2[271] + src2[272] + src2[273] + src2[274] + src2[275] + src2[276] + src2[277] + src2[278] + src2[279] + src2[280] + src2[281] + src2[282] + src2[283] + src2[284] + src2[285] + src2[286] + src2[287] + src2[288] + src2[289] + src2[290] + src2[291] + src2[292] + src2[293] + src2[294] + src2[295] + src2[296] + src2[297] + src2[298] + src2[299] + src2[300] + src2[301] + src2[302] + src2[303] + src2[304] + src2[305] + src2[306] + src2[307] + src2[308] + src2[309] + src2[310] + src2[311] + src2[312] + src2[313] + src2[314] + src2[315] + src2[316] + src2[317] + src2[318] + src2[319] + src2[320] + src2[321] + src2[322] + src2[323] + src2[324] + src2[325] + src2[326] + src2[327] + src2[328] + src2[329] + src2[330] + src2[331] + src2[332] + src2[333] + src2[334] + src2[335] + src2[336] + src2[337] + src2[338] + src2[339] + src2[340] + src2[341] + src2[342] + src2[343] + src2[344] + src2[345] + src2[346] + src2[347] + src2[348] + src2[349] + src2[350] + src2[351] + src2[352] + src2[353] + src2[354] + src2[355] + src2[356] + src2[357] + src2[358] + src2[359] + src2[360] + src2[361] + src2[362] + src2[363] + src2[364] + src2[365] + src2[366] + src2[367] + src2[368] + src2[369] + src2[370] + src2[371] + src2[372] + src2[373] + src2[374] + src2[375] + src2[376] + src2[377] + src2[378] + src2[379] + src2[380] + src2[381] + src2[382] + src2[383] + src2[384] + src2[385] + src2[386] + src2[387] + src2[388] + src2[389] + src2[390] + src2[391] + src2[392] + src2[393] + src2[394] + src2[395] + src2[396] + src2[397] + src2[398] + src2[399] + src2[400] + src2[401] + src2[402] + src2[403] + src2[404] + src2[405] + src2[406] + src2[407] + src2[408] + src2[409] + src2[410] + src2[411] + src2[412] + src2[413] + src2[414] + src2[415] + src2[416] + src2[417] + src2[418] + src2[419] + src2[420] + src2[421] + src2[422] + src2[423] + src2[424] + src2[425] + src2[426] + src2[427] + src2[428] + src2[429] + src2[430] + src2[431] + src2[432] + src2[433] + src2[434] + src2[435] + src2[436] + src2[437] + src2[438] + src2[439] + src2[440] + src2[441] + src2[442] + src2[443] + src2[444] + src2[445] + src2[446] + src2[447] + src2[448] + src2[449] + src2[450] + src2[451] + src2[452] + src2[453] + src2[454] + src2[455] + src2[456] + src2[457] + src2[458] + src2[459] + src2[460] + src2[461] + src2[462] + src2[463] + src2[464] + src2[465] + src2[466] + src2[467] + src2[468] + src2[469] + src2[470] + src2[471] + src2[472] + src2[473] + src2[474] + src2[475] + src2[476] + src2[477] + src2[478] + src2[479] + src2[480] + src2[481] + src2[482] + src2[483] + src2[484] + src2[485] + src2[486] + src2[487] + src2[488] + src2[489] + src2[490] + src2[491] + src2[492] + src2[493] + src2[494] + src2[495] + src2[496] + src2[497] + src2[498] + src2[499] + src2[500] + src2[501] + src2[502] + src2[503] + src2[504] + src2[505] + src2[506] + src2[507] + src2[508] + src2[509] + src2[510] + src2[511])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13] + src3[14] + src3[15] + src3[16] + src3[17] + src3[18] + src3[19] + src3[20] + src3[21] + src3[22] + src3[23] + src3[24] + src3[25] + src3[26] + src3[27] + src3[28] + src3[29] + src3[30] + src3[31] + src3[32] + src3[33] + src3[34] + src3[35] + src3[36] + src3[37] + src3[38] + src3[39] + src3[40] + src3[41] + src3[42] + src3[43] + src3[44] + src3[45] + src3[46] + src3[47] + src3[48] + src3[49] + src3[50] + src3[51] + src3[52] + src3[53] + src3[54] + src3[55] + src3[56] + src3[57] + src3[58] + src3[59] + src3[60] + src3[61] + src3[62] + src3[63] + src3[64] + src3[65] + src3[66] + src3[67] + src3[68] + src3[69] + src3[70] + src3[71] + src3[72] + src3[73] + src3[74] + src3[75] + src3[76] + src3[77] + src3[78] + src3[79] + src3[80] + src3[81] + src3[82] + src3[83] + src3[84] + src3[85] + src3[86] + src3[87] + src3[88] + src3[89] + src3[90] + src3[91] + src3[92] + src3[93] + src3[94] + src3[95] + src3[96] + src3[97] + src3[98] + src3[99] + src3[100] + src3[101] + src3[102] + src3[103] + src3[104] + src3[105] + src3[106] + src3[107] + src3[108] + src3[109] + src3[110] + src3[111] + src3[112] + src3[113] + src3[114] + src3[115] + src3[116] + src3[117] + src3[118] + src3[119] + src3[120] + src3[121] + src3[122] + src3[123] + src3[124] + src3[125] + src3[126] + src3[127] + src3[128] + src3[129] + src3[130] + src3[131] + src3[132] + src3[133] + src3[134] + src3[135] + src3[136] + src3[137] + src3[138] + src3[139] + src3[140] + src3[141] + src3[142] + src3[143] + src3[144] + src3[145] + src3[146] + src3[147] + src3[148] + src3[149] + src3[150] + src3[151] + src3[152] + src3[153] + src3[154] + src3[155] + src3[156] + src3[157] + src3[158] + src3[159] + src3[160] + src3[161] + src3[162] + src3[163] + src3[164] + src3[165] + src3[166] + src3[167] + src3[168] + src3[169] + src3[170] + src3[171] + src3[172] + src3[173] + src3[174] + src3[175] + src3[176] + src3[177] + src3[178] + src3[179] + src3[180] + src3[181] + src3[182] + src3[183] + src3[184] + src3[185] + src3[186] + src3[187] + src3[188] + src3[189] + src3[190] + src3[191] + src3[192] + src3[193] + src3[194] + src3[195] + src3[196] + src3[197] + src3[198] + src3[199] + src3[200] + src3[201] + src3[202] + src3[203] + src3[204] + src3[205] + src3[206] + src3[207] + src3[208] + src3[209] + src3[210] + src3[211] + src3[212] + src3[213] + src3[214] + src3[215] + src3[216] + src3[217] + src3[218] + src3[219] + src3[220] + src3[221] + src3[222] + src3[223] + src3[224] + src3[225] + src3[226] + src3[227] + src3[228] + src3[229] + src3[230] + src3[231] + src3[232] + src3[233] + src3[234] + src3[235] + src3[236] + src3[237] + src3[238] + src3[239] + src3[240] + src3[241] + src3[242] + src3[243] + src3[244] + src3[245] + src3[246] + src3[247] + src3[248] + src3[249] + src3[250] + src3[251] + src3[252] + src3[253] + src3[254] + src3[255] + src3[256] + src3[257] + src3[258] + src3[259] + src3[260] + src3[261] + src3[262] + src3[263] + src3[264] + src3[265] + src3[266] + src3[267] + src3[268] + src3[269] + src3[270] + src3[271] + src3[272] + src3[273] + src3[274] + src3[275] + src3[276] + src3[277] + src3[278] + src3[279] + src3[280] + src3[281] + src3[282] + src3[283] + src3[284] + src3[285] + src3[286] + src3[287] + src3[288] + src3[289] + src3[290] + src3[291] + src3[292] + src3[293] + src3[294] + src3[295] + src3[296] + src3[297] + src3[298] + src3[299] + src3[300] + src3[301] + src3[302] + src3[303] + src3[304] + src3[305] + src3[306] + src3[307] + src3[308] + src3[309] + src3[310] + src3[311] + src3[312] + src3[313] + src3[314] + src3[315] + src3[316] + src3[317] + src3[318] + src3[319] + src3[320] + src3[321] + src3[322] + src3[323] + src3[324] + src3[325] + src3[326] + src3[327] + src3[328] + src3[329] + src3[330] + src3[331] + src3[332] + src3[333] + src3[334] + src3[335] + src3[336] + src3[337] + src3[338] + src3[339] + src3[340] + src3[341] + src3[342] + src3[343] + src3[344] + src3[345] + src3[346] + src3[347] + src3[348] + src3[349] + src3[350] + src3[351] + src3[352] + src3[353] + src3[354] + src3[355] + src3[356] + src3[357] + src3[358] + src3[359] + src3[360] + src3[361] + src3[362] + src3[363] + src3[364] + src3[365] + src3[366] + src3[367] + src3[368] + src3[369] + src3[370] + src3[371] + src3[372] + src3[373] + src3[374] + src3[375] + src3[376] + src3[377] + src3[378] + src3[379] + src3[380] + src3[381] + src3[382] + src3[383] + src3[384] + src3[385] + src3[386] + src3[387] + src3[388] + src3[389] + src3[390] + src3[391] + src3[392] + src3[393] + src3[394] + src3[395] + src3[396] + src3[397] + src3[398] + src3[399] + src3[400] + src3[401] + src3[402] + src3[403] + src3[404] + src3[405] + src3[406] + src3[407] + src3[408] + src3[409] + src3[410] + src3[411] + src3[412] + src3[413] + src3[414] + src3[415] + src3[416] + src3[417] + src3[418] + src3[419] + src3[420] + src3[421] + src3[422] + src3[423] + src3[424] + src3[425] + src3[426] + src3[427] + src3[428] + src3[429] + src3[430] + src3[431] + src3[432] + src3[433] + src3[434] + src3[435] + src3[436] + src3[437] + src3[438] + src3[439] + src3[440] + src3[441] + src3[442] + src3[443] + src3[444] + src3[445] + src3[446] + src3[447] + src3[448] + src3[449] + src3[450] + src3[451] + src3[452] + src3[453] + src3[454] + src3[455] + src3[456] + src3[457] + src3[458] + src3[459] + src3[460] + src3[461] + src3[462] + src3[463] + src3[464] + src3[465] + src3[466] + src3[467] + src3[468] + src3[469] + src3[470] + src3[471] + src3[472] + src3[473] + src3[474] + src3[475] + src3[476] + src3[477] + src3[478] + src3[479] + src3[480] + src3[481] + src3[482] + src3[483] + src3[484] + src3[485] + src3[486] + src3[487] + src3[488] + src3[489] + src3[490] + src3[491] + src3[492] + src3[493] + src3[494] + src3[495] + src3[496] + src3[497] + src3[498] + src3[499] + src3[500] + src3[501] + src3[502] + src3[503] + src3[504] + src3[505] + src3[506] + src3[507] + src3[508] + src3[509] + src3[510] + src3[511])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13] + src4[14] + src4[15] + src4[16] + src4[17] + src4[18] + src4[19] + src4[20] + src4[21] + src4[22] + src4[23] + src4[24] + src4[25] + src4[26] + src4[27] + src4[28] + src4[29] + src4[30] + src4[31] + src4[32] + src4[33] + src4[34] + src4[35] + src4[36] + src4[37] + src4[38] + src4[39] + src4[40] + src4[41] + src4[42] + src4[43] + src4[44] + src4[45] + src4[46] + src4[47] + src4[48] + src4[49] + src4[50] + src4[51] + src4[52] + src4[53] + src4[54] + src4[55] + src4[56] + src4[57] + src4[58] + src4[59] + src4[60] + src4[61] + src4[62] + src4[63] + src4[64] + src4[65] + src4[66] + src4[67] + src4[68] + src4[69] + src4[70] + src4[71] + src4[72] + src4[73] + src4[74] + src4[75] + src4[76] + src4[77] + src4[78] + src4[79] + src4[80] + src4[81] + src4[82] + src4[83] + src4[84] + src4[85] + src4[86] + src4[87] + src4[88] + src4[89] + src4[90] + src4[91] + src4[92] + src4[93] + src4[94] + src4[95] + src4[96] + src4[97] + src4[98] + src4[99] + src4[100] + src4[101] + src4[102] + src4[103] + src4[104] + src4[105] + src4[106] + src4[107] + src4[108] + src4[109] + src4[110] + src4[111] + src4[112] + src4[113] + src4[114] + src4[115] + src4[116] + src4[117] + src4[118] + src4[119] + src4[120] + src4[121] + src4[122] + src4[123] + src4[124] + src4[125] + src4[126] + src4[127] + src4[128] + src4[129] + src4[130] + src4[131] + src4[132] + src4[133] + src4[134] + src4[135] + src4[136] + src4[137] + src4[138] + src4[139] + src4[140] + src4[141] + src4[142] + src4[143] + src4[144] + src4[145] + src4[146] + src4[147] + src4[148] + src4[149] + src4[150] + src4[151] + src4[152] + src4[153] + src4[154] + src4[155] + src4[156] + src4[157] + src4[158] + src4[159] + src4[160] + src4[161] + src4[162] + src4[163] + src4[164] + src4[165] + src4[166] + src4[167] + src4[168] + src4[169] + src4[170] + src4[171] + src4[172] + src4[173] + src4[174] + src4[175] + src4[176] + src4[177] + src4[178] + src4[179] + src4[180] + src4[181] + src4[182] + src4[183] + src4[184] + src4[185] + src4[186] + src4[187] + src4[188] + src4[189] + src4[190] + src4[191] + src4[192] + src4[193] + src4[194] + src4[195] + src4[196] + src4[197] + src4[198] + src4[199] + src4[200] + src4[201] + src4[202] + src4[203] + src4[204] + src4[205] + src4[206] + src4[207] + src4[208] + src4[209] + src4[210] + src4[211] + src4[212] + src4[213] + src4[214] + src4[215] + src4[216] + src4[217] + src4[218] + src4[219] + src4[220] + src4[221] + src4[222] + src4[223] + src4[224] + src4[225] + src4[226] + src4[227] + src4[228] + src4[229] + src4[230] + src4[231] + src4[232] + src4[233] + src4[234] + src4[235] + src4[236] + src4[237] + src4[238] + src4[239] + src4[240] + src4[241] + src4[242] + src4[243] + src4[244] + src4[245] + src4[246] + src4[247] + src4[248] + src4[249] + src4[250] + src4[251] + src4[252] + src4[253] + src4[254] + src4[255] + src4[256] + src4[257] + src4[258] + src4[259] + src4[260] + src4[261] + src4[262] + src4[263] + src4[264] + src4[265] + src4[266] + src4[267] + src4[268] + src4[269] + src4[270] + src4[271] + src4[272] + src4[273] + src4[274] + src4[275] + src4[276] + src4[277] + src4[278] + src4[279] + src4[280] + src4[281] + src4[282] + src4[283] + src4[284] + src4[285] + src4[286] + src4[287] + src4[288] + src4[289] + src4[290] + src4[291] + src4[292] + src4[293] + src4[294] + src4[295] + src4[296] + src4[297] + src4[298] + src4[299] + src4[300] + src4[301] + src4[302] + src4[303] + src4[304] + src4[305] + src4[306] + src4[307] + src4[308] + src4[309] + src4[310] + src4[311] + src4[312] + src4[313] + src4[314] + src4[315] + src4[316] + src4[317] + src4[318] + src4[319] + src4[320] + src4[321] + src4[322] + src4[323] + src4[324] + src4[325] + src4[326] + src4[327] + src4[328] + src4[329] + src4[330] + src4[331] + src4[332] + src4[333] + src4[334] + src4[335] + src4[336] + src4[337] + src4[338] + src4[339] + src4[340] + src4[341] + src4[342] + src4[343] + src4[344] + src4[345] + src4[346] + src4[347] + src4[348] + src4[349] + src4[350] + src4[351] + src4[352] + src4[353] + src4[354] + src4[355] + src4[356] + src4[357] + src4[358] + src4[359] + src4[360] + src4[361] + src4[362] + src4[363] + src4[364] + src4[365] + src4[366] + src4[367] + src4[368] + src4[369] + src4[370] + src4[371] + src4[372] + src4[373] + src4[374] + src4[375] + src4[376] + src4[377] + src4[378] + src4[379] + src4[380] + src4[381] + src4[382] + src4[383] + src4[384] + src4[385] + src4[386] + src4[387] + src4[388] + src4[389] + src4[390] + src4[391] + src4[392] + src4[393] + src4[394] + src4[395] + src4[396] + src4[397] + src4[398] + src4[399] + src4[400] + src4[401] + src4[402] + src4[403] + src4[404] + src4[405] + src4[406] + src4[407] + src4[408] + src4[409] + src4[410] + src4[411] + src4[412] + src4[413] + src4[414] + src4[415] + src4[416] + src4[417] + src4[418] + src4[419] + src4[420] + src4[421] + src4[422] + src4[423] + src4[424] + src4[425] + src4[426] + src4[427] + src4[428] + src4[429] + src4[430] + src4[431] + src4[432] + src4[433] + src4[434] + src4[435] + src4[436] + src4[437] + src4[438] + src4[439] + src4[440] + src4[441] + src4[442] + src4[443] + src4[444] + src4[445] + src4[446] + src4[447] + src4[448] + src4[449] + src4[450] + src4[451] + src4[452] + src4[453] + src4[454] + src4[455] + src4[456] + src4[457] + src4[458] + src4[459] + src4[460] + src4[461] + src4[462] + src4[463] + src4[464] + src4[465] + src4[466] + src4[467] + src4[468] + src4[469] + src4[470] + src4[471] + src4[472] + src4[473] + src4[474] + src4[475] + src4[476] + src4[477] + src4[478] + src4[479] + src4[480] + src4[481] + src4[482] + src4[483] + src4[484] + src4[485] + src4[486] + src4[487] + src4[488] + src4[489] + src4[490] + src4[491] + src4[492] + src4[493] + src4[494] + src4[495] + src4[496] + src4[497] + src4[498] + src4[499] + src4[500] + src4[501] + src4[502] + src4[503] + src4[504] + src4[505] + src4[506] + src4[507] + src4[508] + src4[509] + src4[510] + src4[511])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13] + src5[14] + src5[15] + src5[16] + src5[17] + src5[18] + src5[19] + src5[20] + src5[21] + src5[22] + src5[23] + src5[24] + src5[25] + src5[26] + src5[27] + src5[28] + src5[29] + src5[30] + src5[31] + src5[32] + src5[33] + src5[34] + src5[35] + src5[36] + src5[37] + src5[38] + src5[39] + src5[40] + src5[41] + src5[42] + src5[43] + src5[44] + src5[45] + src5[46] + src5[47] + src5[48] + src5[49] + src5[50] + src5[51] + src5[52] + src5[53] + src5[54] + src5[55] + src5[56] + src5[57] + src5[58] + src5[59] + src5[60] + src5[61] + src5[62] + src5[63] + src5[64] + src5[65] + src5[66] + src5[67] + src5[68] + src5[69] + src5[70] + src5[71] + src5[72] + src5[73] + src5[74] + src5[75] + src5[76] + src5[77] + src5[78] + src5[79] + src5[80] + src5[81] + src5[82] + src5[83] + src5[84] + src5[85] + src5[86] + src5[87] + src5[88] + src5[89] + src5[90] + src5[91] + src5[92] + src5[93] + src5[94] + src5[95] + src5[96] + src5[97] + src5[98] + src5[99] + src5[100] + src5[101] + src5[102] + src5[103] + src5[104] + src5[105] + src5[106] + src5[107] + src5[108] + src5[109] + src5[110] + src5[111] + src5[112] + src5[113] + src5[114] + src5[115] + src5[116] + src5[117] + src5[118] + src5[119] + src5[120] + src5[121] + src5[122] + src5[123] + src5[124] + src5[125] + src5[126] + src5[127] + src5[128] + src5[129] + src5[130] + src5[131] + src5[132] + src5[133] + src5[134] + src5[135] + src5[136] + src5[137] + src5[138] + src5[139] + src5[140] + src5[141] + src5[142] + src5[143] + src5[144] + src5[145] + src5[146] + src5[147] + src5[148] + src5[149] + src5[150] + src5[151] + src5[152] + src5[153] + src5[154] + src5[155] + src5[156] + src5[157] + src5[158] + src5[159] + src5[160] + src5[161] + src5[162] + src5[163] + src5[164] + src5[165] + src5[166] + src5[167] + src5[168] + src5[169] + src5[170] + src5[171] + src5[172] + src5[173] + src5[174] + src5[175] + src5[176] + src5[177] + src5[178] + src5[179] + src5[180] + src5[181] + src5[182] + src5[183] + src5[184] + src5[185] + src5[186] + src5[187] + src5[188] + src5[189] + src5[190] + src5[191] + src5[192] + src5[193] + src5[194] + src5[195] + src5[196] + src5[197] + src5[198] + src5[199] + src5[200] + src5[201] + src5[202] + src5[203] + src5[204] + src5[205] + src5[206] + src5[207] + src5[208] + src5[209] + src5[210] + src5[211] + src5[212] + src5[213] + src5[214] + src5[215] + src5[216] + src5[217] + src5[218] + src5[219] + src5[220] + src5[221] + src5[222] + src5[223] + src5[224] + src5[225] + src5[226] + src5[227] + src5[228] + src5[229] + src5[230] + src5[231] + src5[232] + src5[233] + src5[234] + src5[235] + src5[236] + src5[237] + src5[238] + src5[239] + src5[240] + src5[241] + src5[242] + src5[243] + src5[244] + src5[245] + src5[246] + src5[247] + src5[248] + src5[249] + src5[250] + src5[251] + src5[252] + src5[253] + src5[254] + src5[255] + src5[256] + src5[257] + src5[258] + src5[259] + src5[260] + src5[261] + src5[262] + src5[263] + src5[264] + src5[265] + src5[266] + src5[267] + src5[268] + src5[269] + src5[270] + src5[271] + src5[272] + src5[273] + src5[274] + src5[275] + src5[276] + src5[277] + src5[278] + src5[279] + src5[280] + src5[281] + src5[282] + src5[283] + src5[284] + src5[285] + src5[286] + src5[287] + src5[288] + src5[289] + src5[290] + src5[291] + src5[292] + src5[293] + src5[294] + src5[295] + src5[296] + src5[297] + src5[298] + src5[299] + src5[300] + src5[301] + src5[302] + src5[303] + src5[304] + src5[305] + src5[306] + src5[307] + src5[308] + src5[309] + src5[310] + src5[311] + src5[312] + src5[313] + src5[314] + src5[315] + src5[316] + src5[317] + src5[318] + src5[319] + src5[320] + src5[321] + src5[322] + src5[323] + src5[324] + src5[325] + src5[326] + src5[327] + src5[328] + src5[329] + src5[330] + src5[331] + src5[332] + src5[333] + src5[334] + src5[335] + src5[336] + src5[337] + src5[338] + src5[339] + src5[340] + src5[341] + src5[342] + src5[343] + src5[344] + src5[345] + src5[346] + src5[347] + src5[348] + src5[349] + src5[350] + src5[351] + src5[352] + src5[353] + src5[354] + src5[355] + src5[356] + src5[357] + src5[358] + src5[359] + src5[360] + src5[361] + src5[362] + src5[363] + src5[364] + src5[365] + src5[366] + src5[367] + src5[368] + src5[369] + src5[370] + src5[371] + src5[372] + src5[373] + src5[374] + src5[375] + src5[376] + src5[377] + src5[378] + src5[379] + src5[380] + src5[381] + src5[382] + src5[383] + src5[384] + src5[385] + src5[386] + src5[387] + src5[388] + src5[389] + src5[390] + src5[391] + src5[392] + src5[393] + src5[394] + src5[395] + src5[396] + src5[397] + src5[398] + src5[399] + src5[400] + src5[401] + src5[402] + src5[403] + src5[404] + src5[405] + src5[406] + src5[407] + src5[408] + src5[409] + src5[410] + src5[411] + src5[412] + src5[413] + src5[414] + src5[415] + src5[416] + src5[417] + src5[418] + src5[419] + src5[420] + src5[421] + src5[422] + src5[423] + src5[424] + src5[425] + src5[426] + src5[427] + src5[428] + src5[429] + src5[430] + src5[431] + src5[432] + src5[433] + src5[434] + src5[435] + src5[436] + src5[437] + src5[438] + src5[439] + src5[440] + src5[441] + src5[442] + src5[443] + src5[444] + src5[445] + src5[446] + src5[447] + src5[448] + src5[449] + src5[450] + src5[451] + src5[452] + src5[453] + src5[454] + src5[455] + src5[456] + src5[457] + src5[458] + src5[459] + src5[460] + src5[461] + src5[462] + src5[463] + src5[464] + src5[465] + src5[466] + src5[467] + src5[468] + src5[469] + src5[470] + src5[471] + src5[472] + src5[473] + src5[474] + src5[475] + src5[476] + src5[477] + src5[478] + src5[479] + src5[480] + src5[481] + src5[482] + src5[483] + src5[484] + src5[485] + src5[486] + src5[487] + src5[488] + src5[489] + src5[490] + src5[491] + src5[492] + src5[493] + src5[494] + src5[495] + src5[496] + src5[497] + src5[498] + src5[499] + src5[500] + src5[501] + src5[502] + src5[503] + src5[504] + src5[505] + src5[506] + src5[507] + src5[508] + src5[509] + src5[510] + src5[511])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13] + src6[14] + src6[15] + src6[16] + src6[17] + src6[18] + src6[19] + src6[20] + src6[21] + src6[22] + src6[23] + src6[24] + src6[25] + src6[26] + src6[27] + src6[28] + src6[29] + src6[30] + src6[31] + src6[32] + src6[33] + src6[34] + src6[35] + src6[36] + src6[37] + src6[38] + src6[39] + src6[40] + src6[41] + src6[42] + src6[43] + src6[44] + src6[45] + src6[46] + src6[47] + src6[48] + src6[49] + src6[50] + src6[51] + src6[52] + src6[53] + src6[54] + src6[55] + src6[56] + src6[57] + src6[58] + src6[59] + src6[60] + src6[61] + src6[62] + src6[63] + src6[64] + src6[65] + src6[66] + src6[67] + src6[68] + src6[69] + src6[70] + src6[71] + src6[72] + src6[73] + src6[74] + src6[75] + src6[76] + src6[77] + src6[78] + src6[79] + src6[80] + src6[81] + src6[82] + src6[83] + src6[84] + src6[85] + src6[86] + src6[87] + src6[88] + src6[89] + src6[90] + src6[91] + src6[92] + src6[93] + src6[94] + src6[95] + src6[96] + src6[97] + src6[98] + src6[99] + src6[100] + src6[101] + src6[102] + src6[103] + src6[104] + src6[105] + src6[106] + src6[107] + src6[108] + src6[109] + src6[110] + src6[111] + src6[112] + src6[113] + src6[114] + src6[115] + src6[116] + src6[117] + src6[118] + src6[119] + src6[120] + src6[121] + src6[122] + src6[123] + src6[124] + src6[125] + src6[126] + src6[127] + src6[128] + src6[129] + src6[130] + src6[131] + src6[132] + src6[133] + src6[134] + src6[135] + src6[136] + src6[137] + src6[138] + src6[139] + src6[140] + src6[141] + src6[142] + src6[143] + src6[144] + src6[145] + src6[146] + src6[147] + src6[148] + src6[149] + src6[150] + src6[151] + src6[152] + src6[153] + src6[154] + src6[155] + src6[156] + src6[157] + src6[158] + src6[159] + src6[160] + src6[161] + src6[162] + src6[163] + src6[164] + src6[165] + src6[166] + src6[167] + src6[168] + src6[169] + src6[170] + src6[171] + src6[172] + src6[173] + src6[174] + src6[175] + src6[176] + src6[177] + src6[178] + src6[179] + src6[180] + src6[181] + src6[182] + src6[183] + src6[184] + src6[185] + src6[186] + src6[187] + src6[188] + src6[189] + src6[190] + src6[191] + src6[192] + src6[193] + src6[194] + src6[195] + src6[196] + src6[197] + src6[198] + src6[199] + src6[200] + src6[201] + src6[202] + src6[203] + src6[204] + src6[205] + src6[206] + src6[207] + src6[208] + src6[209] + src6[210] + src6[211] + src6[212] + src6[213] + src6[214] + src6[215] + src6[216] + src6[217] + src6[218] + src6[219] + src6[220] + src6[221] + src6[222] + src6[223] + src6[224] + src6[225] + src6[226] + src6[227] + src6[228] + src6[229] + src6[230] + src6[231] + src6[232] + src6[233] + src6[234] + src6[235] + src6[236] + src6[237] + src6[238] + src6[239] + src6[240] + src6[241] + src6[242] + src6[243] + src6[244] + src6[245] + src6[246] + src6[247] + src6[248] + src6[249] + src6[250] + src6[251] + src6[252] + src6[253] + src6[254] + src6[255] + src6[256] + src6[257] + src6[258] + src6[259] + src6[260] + src6[261] + src6[262] + src6[263] + src6[264] + src6[265] + src6[266] + src6[267] + src6[268] + src6[269] + src6[270] + src6[271] + src6[272] + src6[273] + src6[274] + src6[275] + src6[276] + src6[277] + src6[278] + src6[279] + src6[280] + src6[281] + src6[282] + src6[283] + src6[284] + src6[285] + src6[286] + src6[287] + src6[288] + src6[289] + src6[290] + src6[291] + src6[292] + src6[293] + src6[294] + src6[295] + src6[296] + src6[297] + src6[298] + src6[299] + src6[300] + src6[301] + src6[302] + src6[303] + src6[304] + src6[305] + src6[306] + src6[307] + src6[308] + src6[309] + src6[310] + src6[311] + src6[312] + src6[313] + src6[314] + src6[315] + src6[316] + src6[317] + src6[318] + src6[319] + src6[320] + src6[321] + src6[322] + src6[323] + src6[324] + src6[325] + src6[326] + src6[327] + src6[328] + src6[329] + src6[330] + src6[331] + src6[332] + src6[333] + src6[334] + src6[335] + src6[336] + src6[337] + src6[338] + src6[339] + src6[340] + src6[341] + src6[342] + src6[343] + src6[344] + src6[345] + src6[346] + src6[347] + src6[348] + src6[349] + src6[350] + src6[351] + src6[352] + src6[353] + src6[354] + src6[355] + src6[356] + src6[357] + src6[358] + src6[359] + src6[360] + src6[361] + src6[362] + src6[363] + src6[364] + src6[365] + src6[366] + src6[367] + src6[368] + src6[369] + src6[370] + src6[371] + src6[372] + src6[373] + src6[374] + src6[375] + src6[376] + src6[377] + src6[378] + src6[379] + src6[380] + src6[381] + src6[382] + src6[383] + src6[384] + src6[385] + src6[386] + src6[387] + src6[388] + src6[389] + src6[390] + src6[391] + src6[392] + src6[393] + src6[394] + src6[395] + src6[396] + src6[397] + src6[398] + src6[399] + src6[400] + src6[401] + src6[402] + src6[403] + src6[404] + src6[405] + src6[406] + src6[407] + src6[408] + src6[409] + src6[410] + src6[411] + src6[412] + src6[413] + src6[414] + src6[415] + src6[416] + src6[417] + src6[418] + src6[419] + src6[420] + src6[421] + src6[422] + src6[423] + src6[424] + src6[425] + src6[426] + src6[427] + src6[428] + src6[429] + src6[430] + src6[431] + src6[432] + src6[433] + src6[434] + src6[435] + src6[436] + src6[437] + src6[438] + src6[439] + src6[440] + src6[441] + src6[442] + src6[443] + src6[444] + src6[445] + src6[446] + src6[447] + src6[448] + src6[449] + src6[450] + src6[451] + src6[452] + src6[453] + src6[454] + src6[455] + src6[456] + src6[457] + src6[458] + src6[459] + src6[460] + src6[461] + src6[462] + src6[463] + src6[464] + src6[465] + src6[466] + src6[467] + src6[468] + src6[469] + src6[470] + src6[471] + src6[472] + src6[473] + src6[474] + src6[475] + src6[476] + src6[477] + src6[478] + src6[479] + src6[480] + src6[481] + src6[482] + src6[483] + src6[484] + src6[485] + src6[486] + src6[487] + src6[488] + src6[489] + src6[490] + src6[491] + src6[492] + src6[493] + src6[494] + src6[495] + src6[496] + src6[497] + src6[498] + src6[499] + src6[500] + src6[501] + src6[502] + src6[503] + src6[504] + src6[505] + src6[506] + src6[507] + src6[508] + src6[509] + src6[510] + src6[511])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13] + src7[14] + src7[15] + src7[16] + src7[17] + src7[18] + src7[19] + src7[20] + src7[21] + src7[22] + src7[23] + src7[24] + src7[25] + src7[26] + src7[27] + src7[28] + src7[29] + src7[30] + src7[31] + src7[32] + src7[33] + src7[34] + src7[35] + src7[36] + src7[37] + src7[38] + src7[39] + src7[40] + src7[41] + src7[42] + src7[43] + src7[44] + src7[45] + src7[46] + src7[47] + src7[48] + src7[49] + src7[50] + src7[51] + src7[52] + src7[53] + src7[54] + src7[55] + src7[56] + src7[57] + src7[58] + src7[59] + src7[60] + src7[61] + src7[62] + src7[63] + src7[64] + src7[65] + src7[66] + src7[67] + src7[68] + src7[69] + src7[70] + src7[71] + src7[72] + src7[73] + src7[74] + src7[75] + src7[76] + src7[77] + src7[78] + src7[79] + src7[80] + src7[81] + src7[82] + src7[83] + src7[84] + src7[85] + src7[86] + src7[87] + src7[88] + src7[89] + src7[90] + src7[91] + src7[92] + src7[93] + src7[94] + src7[95] + src7[96] + src7[97] + src7[98] + src7[99] + src7[100] + src7[101] + src7[102] + src7[103] + src7[104] + src7[105] + src7[106] + src7[107] + src7[108] + src7[109] + src7[110] + src7[111] + src7[112] + src7[113] + src7[114] + src7[115] + src7[116] + src7[117] + src7[118] + src7[119] + src7[120] + src7[121] + src7[122] + src7[123] + src7[124] + src7[125] + src7[126] + src7[127] + src7[128] + src7[129] + src7[130] + src7[131] + src7[132] + src7[133] + src7[134] + src7[135] + src7[136] + src7[137] + src7[138] + src7[139] + src7[140] + src7[141] + src7[142] + src7[143] + src7[144] + src7[145] + src7[146] + src7[147] + src7[148] + src7[149] + src7[150] + src7[151] + src7[152] + src7[153] + src7[154] + src7[155] + src7[156] + src7[157] + src7[158] + src7[159] + src7[160] + src7[161] + src7[162] + src7[163] + src7[164] + src7[165] + src7[166] + src7[167] + src7[168] + src7[169] + src7[170] + src7[171] + src7[172] + src7[173] + src7[174] + src7[175] + src7[176] + src7[177] + src7[178] + src7[179] + src7[180] + src7[181] + src7[182] + src7[183] + src7[184] + src7[185] + src7[186] + src7[187] + src7[188] + src7[189] + src7[190] + src7[191] + src7[192] + src7[193] + src7[194] + src7[195] + src7[196] + src7[197] + src7[198] + src7[199] + src7[200] + src7[201] + src7[202] + src7[203] + src7[204] + src7[205] + src7[206] + src7[207] + src7[208] + src7[209] + src7[210] + src7[211] + src7[212] + src7[213] + src7[214] + src7[215] + src7[216] + src7[217] + src7[218] + src7[219] + src7[220] + src7[221] + src7[222] + src7[223] + src7[224] + src7[225] + src7[226] + src7[227] + src7[228] + src7[229] + src7[230] + src7[231] + src7[232] + src7[233] + src7[234] + src7[235] + src7[236] + src7[237] + src7[238] + src7[239] + src7[240] + src7[241] + src7[242] + src7[243] + src7[244] + src7[245] + src7[246] + src7[247] + src7[248] + src7[249] + src7[250] + src7[251] + src7[252] + src7[253] + src7[254] + src7[255] + src7[256] + src7[257] + src7[258] + src7[259] + src7[260] + src7[261] + src7[262] + src7[263] + src7[264] + src7[265] + src7[266] + src7[267] + src7[268] + src7[269] + src7[270] + src7[271] + src7[272] + src7[273] + src7[274] + src7[275] + src7[276] + src7[277] + src7[278] + src7[279] + src7[280] + src7[281] + src7[282] + src7[283] + src7[284] + src7[285] + src7[286] + src7[287] + src7[288] + src7[289] + src7[290] + src7[291] + src7[292] + src7[293] + src7[294] + src7[295] + src7[296] + src7[297] + src7[298] + src7[299] + src7[300] + src7[301] + src7[302] + src7[303] + src7[304] + src7[305] + src7[306] + src7[307] + src7[308] + src7[309] + src7[310] + src7[311] + src7[312] + src7[313] + src7[314] + src7[315] + src7[316] + src7[317] + src7[318] + src7[319] + src7[320] + src7[321] + src7[322] + src7[323] + src7[324] + src7[325] + src7[326] + src7[327] + src7[328] + src7[329] + src7[330] + src7[331] + src7[332] + src7[333] + src7[334] + src7[335] + src7[336] + src7[337] + src7[338] + src7[339] + src7[340] + src7[341] + src7[342] + src7[343] + src7[344] + src7[345] + src7[346] + src7[347] + src7[348] + src7[349] + src7[350] + src7[351] + src7[352] + src7[353] + src7[354] + src7[355] + src7[356] + src7[357] + src7[358] + src7[359] + src7[360] + src7[361] + src7[362] + src7[363] + src7[364] + src7[365] + src7[366] + src7[367] + src7[368] + src7[369] + src7[370] + src7[371] + src7[372] + src7[373] + src7[374] + src7[375] + src7[376] + src7[377] + src7[378] + src7[379] + src7[380] + src7[381] + src7[382] + src7[383] + src7[384] + src7[385] + src7[386] + src7[387] + src7[388] + src7[389] + src7[390] + src7[391] + src7[392] + src7[393] + src7[394] + src7[395] + src7[396] + src7[397] + src7[398] + src7[399] + src7[400] + src7[401] + src7[402] + src7[403] + src7[404] + src7[405] + src7[406] + src7[407] + src7[408] + src7[409] + src7[410] + src7[411] + src7[412] + src7[413] + src7[414] + src7[415] + src7[416] + src7[417] + src7[418] + src7[419] + src7[420] + src7[421] + src7[422] + src7[423] + src7[424] + src7[425] + src7[426] + src7[427] + src7[428] + src7[429] + src7[430] + src7[431] + src7[432] + src7[433] + src7[434] + src7[435] + src7[436] + src7[437] + src7[438] + src7[439] + src7[440] + src7[441] + src7[442] + src7[443] + src7[444] + src7[445] + src7[446] + src7[447] + src7[448] + src7[449] + src7[450] + src7[451] + src7[452] + src7[453] + src7[454] + src7[455] + src7[456] + src7[457] + src7[458] + src7[459] + src7[460] + src7[461] + src7[462] + src7[463] + src7[464] + src7[465] + src7[466] + src7[467] + src7[468] + src7[469] + src7[470] + src7[471] + src7[472] + src7[473] + src7[474] + src7[475] + src7[476] + src7[477] + src7[478] + src7[479] + src7[480] + src7[481] + src7[482] + src7[483] + src7[484] + src7[485] + src7[486] + src7[487] + src7[488] + src7[489] + src7[490] + src7[491] + src7[492] + src7[493] + src7[494] + src7[495] + src7[496] + src7[497] + src7[498] + src7[499] + src7[500] + src7[501] + src7[502] + src7[503] + src7[504] + src7[505] + src7[506] + src7[507] + src7[508] + src7[509] + src7[510] + src7[511])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13] + src8[14] + src8[15] + src8[16] + src8[17] + src8[18] + src8[19] + src8[20] + src8[21] + src8[22] + src8[23] + src8[24] + src8[25] + src8[26] + src8[27] + src8[28] + src8[29] + src8[30] + src8[31] + src8[32] + src8[33] + src8[34] + src8[35] + src8[36] + src8[37] + src8[38] + src8[39] + src8[40] + src8[41] + src8[42] + src8[43] + src8[44] + src8[45] + src8[46] + src8[47] + src8[48] + src8[49] + src8[50] + src8[51] + src8[52] + src8[53] + src8[54] + src8[55] + src8[56] + src8[57] + src8[58] + src8[59] + src8[60] + src8[61] + src8[62] + src8[63] + src8[64] + src8[65] + src8[66] + src8[67] + src8[68] + src8[69] + src8[70] + src8[71] + src8[72] + src8[73] + src8[74] + src8[75] + src8[76] + src8[77] + src8[78] + src8[79] + src8[80] + src8[81] + src8[82] + src8[83] + src8[84] + src8[85] + src8[86] + src8[87] + src8[88] + src8[89] + src8[90] + src8[91] + src8[92] + src8[93] + src8[94] + src8[95] + src8[96] + src8[97] + src8[98] + src8[99] + src8[100] + src8[101] + src8[102] + src8[103] + src8[104] + src8[105] + src8[106] + src8[107] + src8[108] + src8[109] + src8[110] + src8[111] + src8[112] + src8[113] + src8[114] + src8[115] + src8[116] + src8[117] + src8[118] + src8[119] + src8[120] + src8[121] + src8[122] + src8[123] + src8[124] + src8[125] + src8[126] + src8[127] + src8[128] + src8[129] + src8[130] + src8[131] + src8[132] + src8[133] + src8[134] + src8[135] + src8[136] + src8[137] + src8[138] + src8[139] + src8[140] + src8[141] + src8[142] + src8[143] + src8[144] + src8[145] + src8[146] + src8[147] + src8[148] + src8[149] + src8[150] + src8[151] + src8[152] + src8[153] + src8[154] + src8[155] + src8[156] + src8[157] + src8[158] + src8[159] + src8[160] + src8[161] + src8[162] + src8[163] + src8[164] + src8[165] + src8[166] + src8[167] + src8[168] + src8[169] + src8[170] + src8[171] + src8[172] + src8[173] + src8[174] + src8[175] + src8[176] + src8[177] + src8[178] + src8[179] + src8[180] + src8[181] + src8[182] + src8[183] + src8[184] + src8[185] + src8[186] + src8[187] + src8[188] + src8[189] + src8[190] + src8[191] + src8[192] + src8[193] + src8[194] + src8[195] + src8[196] + src8[197] + src8[198] + src8[199] + src8[200] + src8[201] + src8[202] + src8[203] + src8[204] + src8[205] + src8[206] + src8[207] + src8[208] + src8[209] + src8[210] + src8[211] + src8[212] + src8[213] + src8[214] + src8[215] + src8[216] + src8[217] + src8[218] + src8[219] + src8[220] + src8[221] + src8[222] + src8[223] + src8[224] + src8[225] + src8[226] + src8[227] + src8[228] + src8[229] + src8[230] + src8[231] + src8[232] + src8[233] + src8[234] + src8[235] + src8[236] + src8[237] + src8[238] + src8[239] + src8[240] + src8[241] + src8[242] + src8[243] + src8[244] + src8[245] + src8[246] + src8[247] + src8[248] + src8[249] + src8[250] + src8[251] + src8[252] + src8[253] + src8[254] + src8[255] + src8[256] + src8[257] + src8[258] + src8[259] + src8[260] + src8[261] + src8[262] + src8[263] + src8[264] + src8[265] + src8[266] + src8[267] + src8[268] + src8[269] + src8[270] + src8[271] + src8[272] + src8[273] + src8[274] + src8[275] + src8[276] + src8[277] + src8[278] + src8[279] + src8[280] + src8[281] + src8[282] + src8[283] + src8[284] + src8[285] + src8[286] + src8[287] + src8[288] + src8[289] + src8[290] + src8[291] + src8[292] + src8[293] + src8[294] + src8[295] + src8[296] + src8[297] + src8[298] + src8[299] + src8[300] + src8[301] + src8[302] + src8[303] + src8[304] + src8[305] + src8[306] + src8[307] + src8[308] + src8[309] + src8[310] + src8[311] + src8[312] + src8[313] + src8[314] + src8[315] + src8[316] + src8[317] + src8[318] + src8[319] + src8[320] + src8[321] + src8[322] + src8[323] + src8[324] + src8[325] + src8[326] + src8[327] + src8[328] + src8[329] + src8[330] + src8[331] + src8[332] + src8[333] + src8[334] + src8[335] + src8[336] + src8[337] + src8[338] + src8[339] + src8[340] + src8[341] + src8[342] + src8[343] + src8[344] + src8[345] + src8[346] + src8[347] + src8[348] + src8[349] + src8[350] + src8[351] + src8[352] + src8[353] + src8[354] + src8[355] + src8[356] + src8[357] + src8[358] + src8[359] + src8[360] + src8[361] + src8[362] + src8[363] + src8[364] + src8[365] + src8[366] + src8[367] + src8[368] + src8[369] + src8[370] + src8[371] + src8[372] + src8[373] + src8[374] + src8[375] + src8[376] + src8[377] + src8[378] + src8[379] + src8[380] + src8[381] + src8[382] + src8[383] + src8[384] + src8[385] + src8[386] + src8[387] + src8[388] + src8[389] + src8[390] + src8[391] + src8[392] + src8[393] + src8[394] + src8[395] + src8[396] + src8[397] + src8[398] + src8[399] + src8[400] + src8[401] + src8[402] + src8[403] + src8[404] + src8[405] + src8[406] + src8[407] + src8[408] + src8[409] + src8[410] + src8[411] + src8[412] + src8[413] + src8[414] + src8[415] + src8[416] + src8[417] + src8[418] + src8[419] + src8[420] + src8[421] + src8[422] + src8[423] + src8[424] + src8[425] + src8[426] + src8[427] + src8[428] + src8[429] + src8[430] + src8[431] + src8[432] + src8[433] + src8[434] + src8[435] + src8[436] + src8[437] + src8[438] + src8[439] + src8[440] + src8[441] + src8[442] + src8[443] + src8[444] + src8[445] + src8[446] + src8[447] + src8[448] + src8[449] + src8[450] + src8[451] + src8[452] + src8[453] + src8[454] + src8[455] + src8[456] + src8[457] + src8[458] + src8[459] + src8[460] + src8[461] + src8[462] + src8[463] + src8[464] + src8[465] + src8[466] + src8[467] + src8[468] + src8[469] + src8[470] + src8[471] + src8[472] + src8[473] + src8[474] + src8[475] + src8[476] + src8[477] + src8[478] + src8[479] + src8[480] + src8[481] + src8[482] + src8[483] + src8[484] + src8[485] + src8[486] + src8[487] + src8[488] + src8[489] + src8[490] + src8[491] + src8[492] + src8[493] + src8[494] + src8[495] + src8[496] + src8[497] + src8[498] + src8[499] + src8[500] + src8[501] + src8[502] + src8[503] + src8[504] + src8[505] + src8[506] + src8[507] + src8[508] + src8[509] + src8[510] + src8[511])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13] + src9[14] + src9[15] + src9[16] + src9[17] + src9[18] + src9[19] + src9[20] + src9[21] + src9[22] + src9[23] + src9[24] + src9[25] + src9[26] + src9[27] + src9[28] + src9[29] + src9[30] + src9[31] + src9[32] + src9[33] + src9[34] + src9[35] + src9[36] + src9[37] + src9[38] + src9[39] + src9[40] + src9[41] + src9[42] + src9[43] + src9[44] + src9[45] + src9[46] + src9[47] + src9[48] + src9[49] + src9[50] + src9[51] + src9[52] + src9[53] + src9[54] + src9[55] + src9[56] + src9[57] + src9[58] + src9[59] + src9[60] + src9[61] + src9[62] + src9[63] + src9[64] + src9[65] + src9[66] + src9[67] + src9[68] + src9[69] + src9[70] + src9[71] + src9[72] + src9[73] + src9[74] + src9[75] + src9[76] + src9[77] + src9[78] + src9[79] + src9[80] + src9[81] + src9[82] + src9[83] + src9[84] + src9[85] + src9[86] + src9[87] + src9[88] + src9[89] + src9[90] + src9[91] + src9[92] + src9[93] + src9[94] + src9[95] + src9[96] + src9[97] + src9[98] + src9[99] + src9[100] + src9[101] + src9[102] + src9[103] + src9[104] + src9[105] + src9[106] + src9[107] + src9[108] + src9[109] + src9[110] + src9[111] + src9[112] + src9[113] + src9[114] + src9[115] + src9[116] + src9[117] + src9[118] + src9[119] + src9[120] + src9[121] + src9[122] + src9[123] + src9[124] + src9[125] + src9[126] + src9[127] + src9[128] + src9[129] + src9[130] + src9[131] + src9[132] + src9[133] + src9[134] + src9[135] + src9[136] + src9[137] + src9[138] + src9[139] + src9[140] + src9[141] + src9[142] + src9[143] + src9[144] + src9[145] + src9[146] + src9[147] + src9[148] + src9[149] + src9[150] + src9[151] + src9[152] + src9[153] + src9[154] + src9[155] + src9[156] + src9[157] + src9[158] + src9[159] + src9[160] + src9[161] + src9[162] + src9[163] + src9[164] + src9[165] + src9[166] + src9[167] + src9[168] + src9[169] + src9[170] + src9[171] + src9[172] + src9[173] + src9[174] + src9[175] + src9[176] + src9[177] + src9[178] + src9[179] + src9[180] + src9[181] + src9[182] + src9[183] + src9[184] + src9[185] + src9[186] + src9[187] + src9[188] + src9[189] + src9[190] + src9[191] + src9[192] + src9[193] + src9[194] + src9[195] + src9[196] + src9[197] + src9[198] + src9[199] + src9[200] + src9[201] + src9[202] + src9[203] + src9[204] + src9[205] + src9[206] + src9[207] + src9[208] + src9[209] + src9[210] + src9[211] + src9[212] + src9[213] + src9[214] + src9[215] + src9[216] + src9[217] + src9[218] + src9[219] + src9[220] + src9[221] + src9[222] + src9[223] + src9[224] + src9[225] + src9[226] + src9[227] + src9[228] + src9[229] + src9[230] + src9[231] + src9[232] + src9[233] + src9[234] + src9[235] + src9[236] + src9[237] + src9[238] + src9[239] + src9[240] + src9[241] + src9[242] + src9[243] + src9[244] + src9[245] + src9[246] + src9[247] + src9[248] + src9[249] + src9[250] + src9[251] + src9[252] + src9[253] + src9[254] + src9[255] + src9[256] + src9[257] + src9[258] + src9[259] + src9[260] + src9[261] + src9[262] + src9[263] + src9[264] + src9[265] + src9[266] + src9[267] + src9[268] + src9[269] + src9[270] + src9[271] + src9[272] + src9[273] + src9[274] + src9[275] + src9[276] + src9[277] + src9[278] + src9[279] + src9[280] + src9[281] + src9[282] + src9[283] + src9[284] + src9[285] + src9[286] + src9[287] + src9[288] + src9[289] + src9[290] + src9[291] + src9[292] + src9[293] + src9[294] + src9[295] + src9[296] + src9[297] + src9[298] + src9[299] + src9[300] + src9[301] + src9[302] + src9[303] + src9[304] + src9[305] + src9[306] + src9[307] + src9[308] + src9[309] + src9[310] + src9[311] + src9[312] + src9[313] + src9[314] + src9[315] + src9[316] + src9[317] + src9[318] + src9[319] + src9[320] + src9[321] + src9[322] + src9[323] + src9[324] + src9[325] + src9[326] + src9[327] + src9[328] + src9[329] + src9[330] + src9[331] + src9[332] + src9[333] + src9[334] + src9[335] + src9[336] + src9[337] + src9[338] + src9[339] + src9[340] + src9[341] + src9[342] + src9[343] + src9[344] + src9[345] + src9[346] + src9[347] + src9[348] + src9[349] + src9[350] + src9[351] + src9[352] + src9[353] + src9[354] + src9[355] + src9[356] + src9[357] + src9[358] + src9[359] + src9[360] + src9[361] + src9[362] + src9[363] + src9[364] + src9[365] + src9[366] + src9[367] + src9[368] + src9[369] + src9[370] + src9[371] + src9[372] + src9[373] + src9[374] + src9[375] + src9[376] + src9[377] + src9[378] + src9[379] + src9[380] + src9[381] + src9[382] + src9[383] + src9[384] + src9[385] + src9[386] + src9[387] + src9[388] + src9[389] + src9[390] + src9[391] + src9[392] + src9[393] + src9[394] + src9[395] + src9[396] + src9[397] + src9[398] + src9[399] + src9[400] + src9[401] + src9[402] + src9[403] + src9[404] + src9[405] + src9[406] + src9[407] + src9[408] + src9[409] + src9[410] + src9[411] + src9[412] + src9[413] + src9[414] + src9[415] + src9[416] + src9[417] + src9[418] + src9[419] + src9[420] + src9[421] + src9[422] + src9[423] + src9[424] + src9[425] + src9[426] + src9[427] + src9[428] + src9[429] + src9[430] + src9[431] + src9[432] + src9[433] + src9[434] + src9[435] + src9[436] + src9[437] + src9[438] + src9[439] + src9[440] + src9[441] + src9[442] + src9[443] + src9[444] + src9[445] + src9[446] + src9[447] + src9[448] + src9[449] + src9[450] + src9[451] + src9[452] + src9[453] + src9[454] + src9[455] + src9[456] + src9[457] + src9[458] + src9[459] + src9[460] + src9[461] + src9[462] + src9[463] + src9[464] + src9[465] + src9[466] + src9[467] + src9[468] + src9[469] + src9[470] + src9[471] + src9[472] + src9[473] + src9[474] + src9[475] + src9[476] + src9[477] + src9[478] + src9[479] + src9[480] + src9[481] + src9[482] + src9[483] + src9[484] + src9[485] + src9[486] + src9[487] + src9[488] + src9[489] + src9[490] + src9[491] + src9[492] + src9[493] + src9[494] + src9[495] + src9[496] + src9[497] + src9[498] + src9[499] + src9[500] + src9[501] + src9[502] + src9[503] + src9[504] + src9[505] + src9[506] + src9[507] + src9[508] + src9[509] + src9[510] + src9[511])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13] + src10[14] + src10[15] + src10[16] + src10[17] + src10[18] + src10[19] + src10[20] + src10[21] + src10[22] + src10[23] + src10[24] + src10[25] + src10[26] + src10[27] + src10[28] + src10[29] + src10[30] + src10[31] + src10[32] + src10[33] + src10[34] + src10[35] + src10[36] + src10[37] + src10[38] + src10[39] + src10[40] + src10[41] + src10[42] + src10[43] + src10[44] + src10[45] + src10[46] + src10[47] + src10[48] + src10[49] + src10[50] + src10[51] + src10[52] + src10[53] + src10[54] + src10[55] + src10[56] + src10[57] + src10[58] + src10[59] + src10[60] + src10[61] + src10[62] + src10[63] + src10[64] + src10[65] + src10[66] + src10[67] + src10[68] + src10[69] + src10[70] + src10[71] + src10[72] + src10[73] + src10[74] + src10[75] + src10[76] + src10[77] + src10[78] + src10[79] + src10[80] + src10[81] + src10[82] + src10[83] + src10[84] + src10[85] + src10[86] + src10[87] + src10[88] + src10[89] + src10[90] + src10[91] + src10[92] + src10[93] + src10[94] + src10[95] + src10[96] + src10[97] + src10[98] + src10[99] + src10[100] + src10[101] + src10[102] + src10[103] + src10[104] + src10[105] + src10[106] + src10[107] + src10[108] + src10[109] + src10[110] + src10[111] + src10[112] + src10[113] + src10[114] + src10[115] + src10[116] + src10[117] + src10[118] + src10[119] + src10[120] + src10[121] + src10[122] + src10[123] + src10[124] + src10[125] + src10[126] + src10[127] + src10[128] + src10[129] + src10[130] + src10[131] + src10[132] + src10[133] + src10[134] + src10[135] + src10[136] + src10[137] + src10[138] + src10[139] + src10[140] + src10[141] + src10[142] + src10[143] + src10[144] + src10[145] + src10[146] + src10[147] + src10[148] + src10[149] + src10[150] + src10[151] + src10[152] + src10[153] + src10[154] + src10[155] + src10[156] + src10[157] + src10[158] + src10[159] + src10[160] + src10[161] + src10[162] + src10[163] + src10[164] + src10[165] + src10[166] + src10[167] + src10[168] + src10[169] + src10[170] + src10[171] + src10[172] + src10[173] + src10[174] + src10[175] + src10[176] + src10[177] + src10[178] + src10[179] + src10[180] + src10[181] + src10[182] + src10[183] + src10[184] + src10[185] + src10[186] + src10[187] + src10[188] + src10[189] + src10[190] + src10[191] + src10[192] + src10[193] + src10[194] + src10[195] + src10[196] + src10[197] + src10[198] + src10[199] + src10[200] + src10[201] + src10[202] + src10[203] + src10[204] + src10[205] + src10[206] + src10[207] + src10[208] + src10[209] + src10[210] + src10[211] + src10[212] + src10[213] + src10[214] + src10[215] + src10[216] + src10[217] + src10[218] + src10[219] + src10[220] + src10[221] + src10[222] + src10[223] + src10[224] + src10[225] + src10[226] + src10[227] + src10[228] + src10[229] + src10[230] + src10[231] + src10[232] + src10[233] + src10[234] + src10[235] + src10[236] + src10[237] + src10[238] + src10[239] + src10[240] + src10[241] + src10[242] + src10[243] + src10[244] + src10[245] + src10[246] + src10[247] + src10[248] + src10[249] + src10[250] + src10[251] + src10[252] + src10[253] + src10[254] + src10[255] + src10[256] + src10[257] + src10[258] + src10[259] + src10[260] + src10[261] + src10[262] + src10[263] + src10[264] + src10[265] + src10[266] + src10[267] + src10[268] + src10[269] + src10[270] + src10[271] + src10[272] + src10[273] + src10[274] + src10[275] + src10[276] + src10[277] + src10[278] + src10[279] + src10[280] + src10[281] + src10[282] + src10[283] + src10[284] + src10[285] + src10[286] + src10[287] + src10[288] + src10[289] + src10[290] + src10[291] + src10[292] + src10[293] + src10[294] + src10[295] + src10[296] + src10[297] + src10[298] + src10[299] + src10[300] + src10[301] + src10[302] + src10[303] + src10[304] + src10[305] + src10[306] + src10[307] + src10[308] + src10[309] + src10[310] + src10[311] + src10[312] + src10[313] + src10[314] + src10[315] + src10[316] + src10[317] + src10[318] + src10[319] + src10[320] + src10[321] + src10[322] + src10[323] + src10[324] + src10[325] + src10[326] + src10[327] + src10[328] + src10[329] + src10[330] + src10[331] + src10[332] + src10[333] + src10[334] + src10[335] + src10[336] + src10[337] + src10[338] + src10[339] + src10[340] + src10[341] + src10[342] + src10[343] + src10[344] + src10[345] + src10[346] + src10[347] + src10[348] + src10[349] + src10[350] + src10[351] + src10[352] + src10[353] + src10[354] + src10[355] + src10[356] + src10[357] + src10[358] + src10[359] + src10[360] + src10[361] + src10[362] + src10[363] + src10[364] + src10[365] + src10[366] + src10[367] + src10[368] + src10[369] + src10[370] + src10[371] + src10[372] + src10[373] + src10[374] + src10[375] + src10[376] + src10[377] + src10[378] + src10[379] + src10[380] + src10[381] + src10[382] + src10[383] + src10[384] + src10[385] + src10[386] + src10[387] + src10[388] + src10[389] + src10[390] + src10[391] + src10[392] + src10[393] + src10[394] + src10[395] + src10[396] + src10[397] + src10[398] + src10[399] + src10[400] + src10[401] + src10[402] + src10[403] + src10[404] + src10[405] + src10[406] + src10[407] + src10[408] + src10[409] + src10[410] + src10[411] + src10[412] + src10[413] + src10[414] + src10[415] + src10[416] + src10[417] + src10[418] + src10[419] + src10[420] + src10[421] + src10[422] + src10[423] + src10[424] + src10[425] + src10[426] + src10[427] + src10[428] + src10[429] + src10[430] + src10[431] + src10[432] + src10[433] + src10[434] + src10[435] + src10[436] + src10[437] + src10[438] + src10[439] + src10[440] + src10[441] + src10[442] + src10[443] + src10[444] + src10[445] + src10[446] + src10[447] + src10[448] + src10[449] + src10[450] + src10[451] + src10[452] + src10[453] + src10[454] + src10[455] + src10[456] + src10[457] + src10[458] + src10[459] + src10[460] + src10[461] + src10[462] + src10[463] + src10[464] + src10[465] + src10[466] + src10[467] + src10[468] + src10[469] + src10[470] + src10[471] + src10[472] + src10[473] + src10[474] + src10[475] + src10[476] + src10[477] + src10[478] + src10[479] + src10[480] + src10[481] + src10[482] + src10[483] + src10[484] + src10[485] + src10[486] + src10[487] + src10[488] + src10[489] + src10[490] + src10[491] + src10[492] + src10[493] + src10[494] + src10[495] + src10[496] + src10[497] + src10[498] + src10[499] + src10[500] + src10[501] + src10[502] + src10[503] + src10[504] + src10[505] + src10[506] + src10[507] + src10[508] + src10[509] + src10[510] + src10[511])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13] + src11[14] + src11[15] + src11[16] + src11[17] + src11[18] + src11[19] + src11[20] + src11[21] + src11[22] + src11[23] + src11[24] + src11[25] + src11[26] + src11[27] + src11[28] + src11[29] + src11[30] + src11[31] + src11[32] + src11[33] + src11[34] + src11[35] + src11[36] + src11[37] + src11[38] + src11[39] + src11[40] + src11[41] + src11[42] + src11[43] + src11[44] + src11[45] + src11[46] + src11[47] + src11[48] + src11[49] + src11[50] + src11[51] + src11[52] + src11[53] + src11[54] + src11[55] + src11[56] + src11[57] + src11[58] + src11[59] + src11[60] + src11[61] + src11[62] + src11[63] + src11[64] + src11[65] + src11[66] + src11[67] + src11[68] + src11[69] + src11[70] + src11[71] + src11[72] + src11[73] + src11[74] + src11[75] + src11[76] + src11[77] + src11[78] + src11[79] + src11[80] + src11[81] + src11[82] + src11[83] + src11[84] + src11[85] + src11[86] + src11[87] + src11[88] + src11[89] + src11[90] + src11[91] + src11[92] + src11[93] + src11[94] + src11[95] + src11[96] + src11[97] + src11[98] + src11[99] + src11[100] + src11[101] + src11[102] + src11[103] + src11[104] + src11[105] + src11[106] + src11[107] + src11[108] + src11[109] + src11[110] + src11[111] + src11[112] + src11[113] + src11[114] + src11[115] + src11[116] + src11[117] + src11[118] + src11[119] + src11[120] + src11[121] + src11[122] + src11[123] + src11[124] + src11[125] + src11[126] + src11[127] + src11[128] + src11[129] + src11[130] + src11[131] + src11[132] + src11[133] + src11[134] + src11[135] + src11[136] + src11[137] + src11[138] + src11[139] + src11[140] + src11[141] + src11[142] + src11[143] + src11[144] + src11[145] + src11[146] + src11[147] + src11[148] + src11[149] + src11[150] + src11[151] + src11[152] + src11[153] + src11[154] + src11[155] + src11[156] + src11[157] + src11[158] + src11[159] + src11[160] + src11[161] + src11[162] + src11[163] + src11[164] + src11[165] + src11[166] + src11[167] + src11[168] + src11[169] + src11[170] + src11[171] + src11[172] + src11[173] + src11[174] + src11[175] + src11[176] + src11[177] + src11[178] + src11[179] + src11[180] + src11[181] + src11[182] + src11[183] + src11[184] + src11[185] + src11[186] + src11[187] + src11[188] + src11[189] + src11[190] + src11[191] + src11[192] + src11[193] + src11[194] + src11[195] + src11[196] + src11[197] + src11[198] + src11[199] + src11[200] + src11[201] + src11[202] + src11[203] + src11[204] + src11[205] + src11[206] + src11[207] + src11[208] + src11[209] + src11[210] + src11[211] + src11[212] + src11[213] + src11[214] + src11[215] + src11[216] + src11[217] + src11[218] + src11[219] + src11[220] + src11[221] + src11[222] + src11[223] + src11[224] + src11[225] + src11[226] + src11[227] + src11[228] + src11[229] + src11[230] + src11[231] + src11[232] + src11[233] + src11[234] + src11[235] + src11[236] + src11[237] + src11[238] + src11[239] + src11[240] + src11[241] + src11[242] + src11[243] + src11[244] + src11[245] + src11[246] + src11[247] + src11[248] + src11[249] + src11[250] + src11[251] + src11[252] + src11[253] + src11[254] + src11[255] + src11[256] + src11[257] + src11[258] + src11[259] + src11[260] + src11[261] + src11[262] + src11[263] + src11[264] + src11[265] + src11[266] + src11[267] + src11[268] + src11[269] + src11[270] + src11[271] + src11[272] + src11[273] + src11[274] + src11[275] + src11[276] + src11[277] + src11[278] + src11[279] + src11[280] + src11[281] + src11[282] + src11[283] + src11[284] + src11[285] + src11[286] + src11[287] + src11[288] + src11[289] + src11[290] + src11[291] + src11[292] + src11[293] + src11[294] + src11[295] + src11[296] + src11[297] + src11[298] + src11[299] + src11[300] + src11[301] + src11[302] + src11[303] + src11[304] + src11[305] + src11[306] + src11[307] + src11[308] + src11[309] + src11[310] + src11[311] + src11[312] + src11[313] + src11[314] + src11[315] + src11[316] + src11[317] + src11[318] + src11[319] + src11[320] + src11[321] + src11[322] + src11[323] + src11[324] + src11[325] + src11[326] + src11[327] + src11[328] + src11[329] + src11[330] + src11[331] + src11[332] + src11[333] + src11[334] + src11[335] + src11[336] + src11[337] + src11[338] + src11[339] + src11[340] + src11[341] + src11[342] + src11[343] + src11[344] + src11[345] + src11[346] + src11[347] + src11[348] + src11[349] + src11[350] + src11[351] + src11[352] + src11[353] + src11[354] + src11[355] + src11[356] + src11[357] + src11[358] + src11[359] + src11[360] + src11[361] + src11[362] + src11[363] + src11[364] + src11[365] + src11[366] + src11[367] + src11[368] + src11[369] + src11[370] + src11[371] + src11[372] + src11[373] + src11[374] + src11[375] + src11[376] + src11[377] + src11[378] + src11[379] + src11[380] + src11[381] + src11[382] + src11[383] + src11[384] + src11[385] + src11[386] + src11[387] + src11[388] + src11[389] + src11[390] + src11[391] + src11[392] + src11[393] + src11[394] + src11[395] + src11[396] + src11[397] + src11[398] + src11[399] + src11[400] + src11[401] + src11[402] + src11[403] + src11[404] + src11[405] + src11[406] + src11[407] + src11[408] + src11[409] + src11[410] + src11[411] + src11[412] + src11[413] + src11[414] + src11[415] + src11[416] + src11[417] + src11[418] + src11[419] + src11[420] + src11[421] + src11[422] + src11[423] + src11[424] + src11[425] + src11[426] + src11[427] + src11[428] + src11[429] + src11[430] + src11[431] + src11[432] + src11[433] + src11[434] + src11[435] + src11[436] + src11[437] + src11[438] + src11[439] + src11[440] + src11[441] + src11[442] + src11[443] + src11[444] + src11[445] + src11[446] + src11[447] + src11[448] + src11[449] + src11[450] + src11[451] + src11[452] + src11[453] + src11[454] + src11[455] + src11[456] + src11[457] + src11[458] + src11[459] + src11[460] + src11[461] + src11[462] + src11[463] + src11[464] + src11[465] + src11[466] + src11[467] + src11[468] + src11[469] + src11[470] + src11[471] + src11[472] + src11[473] + src11[474] + src11[475] + src11[476] + src11[477] + src11[478] + src11[479] + src11[480] + src11[481] + src11[482] + src11[483] + src11[484] + src11[485] + src11[486] + src11[487] + src11[488] + src11[489] + src11[490] + src11[491] + src11[492] + src11[493] + src11[494] + src11[495] + src11[496] + src11[497] + src11[498] + src11[499] + src11[500] + src11[501] + src11[502] + src11[503] + src11[504] + src11[505] + src11[506] + src11[507] + src11[508] + src11[509] + src11[510] + src11[511])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12] + src12[13] + src12[14] + src12[15] + src12[16] + src12[17] + src12[18] + src12[19] + src12[20] + src12[21] + src12[22] + src12[23] + src12[24] + src12[25] + src12[26] + src12[27] + src12[28] + src12[29] + src12[30] + src12[31] + src12[32] + src12[33] + src12[34] + src12[35] + src12[36] + src12[37] + src12[38] + src12[39] + src12[40] + src12[41] + src12[42] + src12[43] + src12[44] + src12[45] + src12[46] + src12[47] + src12[48] + src12[49] + src12[50] + src12[51] + src12[52] + src12[53] + src12[54] + src12[55] + src12[56] + src12[57] + src12[58] + src12[59] + src12[60] + src12[61] + src12[62] + src12[63] + src12[64] + src12[65] + src12[66] + src12[67] + src12[68] + src12[69] + src12[70] + src12[71] + src12[72] + src12[73] + src12[74] + src12[75] + src12[76] + src12[77] + src12[78] + src12[79] + src12[80] + src12[81] + src12[82] + src12[83] + src12[84] + src12[85] + src12[86] + src12[87] + src12[88] + src12[89] + src12[90] + src12[91] + src12[92] + src12[93] + src12[94] + src12[95] + src12[96] + src12[97] + src12[98] + src12[99] + src12[100] + src12[101] + src12[102] + src12[103] + src12[104] + src12[105] + src12[106] + src12[107] + src12[108] + src12[109] + src12[110] + src12[111] + src12[112] + src12[113] + src12[114] + src12[115] + src12[116] + src12[117] + src12[118] + src12[119] + src12[120] + src12[121] + src12[122] + src12[123] + src12[124] + src12[125] + src12[126] + src12[127] + src12[128] + src12[129] + src12[130] + src12[131] + src12[132] + src12[133] + src12[134] + src12[135] + src12[136] + src12[137] + src12[138] + src12[139] + src12[140] + src12[141] + src12[142] + src12[143] + src12[144] + src12[145] + src12[146] + src12[147] + src12[148] + src12[149] + src12[150] + src12[151] + src12[152] + src12[153] + src12[154] + src12[155] + src12[156] + src12[157] + src12[158] + src12[159] + src12[160] + src12[161] + src12[162] + src12[163] + src12[164] + src12[165] + src12[166] + src12[167] + src12[168] + src12[169] + src12[170] + src12[171] + src12[172] + src12[173] + src12[174] + src12[175] + src12[176] + src12[177] + src12[178] + src12[179] + src12[180] + src12[181] + src12[182] + src12[183] + src12[184] + src12[185] + src12[186] + src12[187] + src12[188] + src12[189] + src12[190] + src12[191] + src12[192] + src12[193] + src12[194] + src12[195] + src12[196] + src12[197] + src12[198] + src12[199] + src12[200] + src12[201] + src12[202] + src12[203] + src12[204] + src12[205] + src12[206] + src12[207] + src12[208] + src12[209] + src12[210] + src12[211] + src12[212] + src12[213] + src12[214] + src12[215] + src12[216] + src12[217] + src12[218] + src12[219] + src12[220] + src12[221] + src12[222] + src12[223] + src12[224] + src12[225] + src12[226] + src12[227] + src12[228] + src12[229] + src12[230] + src12[231] + src12[232] + src12[233] + src12[234] + src12[235] + src12[236] + src12[237] + src12[238] + src12[239] + src12[240] + src12[241] + src12[242] + src12[243] + src12[244] + src12[245] + src12[246] + src12[247] + src12[248] + src12[249] + src12[250] + src12[251] + src12[252] + src12[253] + src12[254] + src12[255] + src12[256] + src12[257] + src12[258] + src12[259] + src12[260] + src12[261] + src12[262] + src12[263] + src12[264] + src12[265] + src12[266] + src12[267] + src12[268] + src12[269] + src12[270] + src12[271] + src12[272] + src12[273] + src12[274] + src12[275] + src12[276] + src12[277] + src12[278] + src12[279] + src12[280] + src12[281] + src12[282] + src12[283] + src12[284] + src12[285] + src12[286] + src12[287] + src12[288] + src12[289] + src12[290] + src12[291] + src12[292] + src12[293] + src12[294] + src12[295] + src12[296] + src12[297] + src12[298] + src12[299] + src12[300] + src12[301] + src12[302] + src12[303] + src12[304] + src12[305] + src12[306] + src12[307] + src12[308] + src12[309] + src12[310] + src12[311] + src12[312] + src12[313] + src12[314] + src12[315] + src12[316] + src12[317] + src12[318] + src12[319] + src12[320] + src12[321] + src12[322] + src12[323] + src12[324] + src12[325] + src12[326] + src12[327] + src12[328] + src12[329] + src12[330] + src12[331] + src12[332] + src12[333] + src12[334] + src12[335] + src12[336] + src12[337] + src12[338] + src12[339] + src12[340] + src12[341] + src12[342] + src12[343] + src12[344] + src12[345] + src12[346] + src12[347] + src12[348] + src12[349] + src12[350] + src12[351] + src12[352] + src12[353] + src12[354] + src12[355] + src12[356] + src12[357] + src12[358] + src12[359] + src12[360] + src12[361] + src12[362] + src12[363] + src12[364] + src12[365] + src12[366] + src12[367] + src12[368] + src12[369] + src12[370] + src12[371] + src12[372] + src12[373] + src12[374] + src12[375] + src12[376] + src12[377] + src12[378] + src12[379] + src12[380] + src12[381] + src12[382] + src12[383] + src12[384] + src12[385] + src12[386] + src12[387] + src12[388] + src12[389] + src12[390] + src12[391] + src12[392] + src12[393] + src12[394] + src12[395] + src12[396] + src12[397] + src12[398] + src12[399] + src12[400] + src12[401] + src12[402] + src12[403] + src12[404] + src12[405] + src12[406] + src12[407] + src12[408] + src12[409] + src12[410] + src12[411] + src12[412] + src12[413] + src12[414] + src12[415] + src12[416] + src12[417] + src12[418] + src12[419] + src12[420] + src12[421] + src12[422] + src12[423] + src12[424] + src12[425] + src12[426] + src12[427] + src12[428] + src12[429] + src12[430] + src12[431] + src12[432] + src12[433] + src12[434] + src12[435] + src12[436] + src12[437] + src12[438] + src12[439] + src12[440] + src12[441] + src12[442] + src12[443] + src12[444] + src12[445] + src12[446] + src12[447] + src12[448] + src12[449] + src12[450] + src12[451] + src12[452] + src12[453] + src12[454] + src12[455] + src12[456] + src12[457] + src12[458] + src12[459] + src12[460] + src12[461] + src12[462] + src12[463] + src12[464] + src12[465] + src12[466] + src12[467] + src12[468] + src12[469] + src12[470] + src12[471] + src12[472] + src12[473] + src12[474] + src12[475] + src12[476] + src12[477] + src12[478] + src12[479] + src12[480] + src12[481] + src12[482] + src12[483] + src12[484] + src12[485] + src12[486] + src12[487] + src12[488] + src12[489] + src12[490] + src12[491] + src12[492] + src12[493] + src12[494] + src12[495] + src12[496] + src12[497] + src12[498] + src12[499] + src12[500] + src12[501] + src12[502] + src12[503] + src12[504] + src12[505] + src12[506] + src12[507] + src12[508] + src12[509] + src12[510] + src12[511])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13] + src13[14] + src13[15] + src13[16] + src13[17] + src13[18] + src13[19] + src13[20] + src13[21] + src13[22] + src13[23] + src13[24] + src13[25] + src13[26] + src13[27] + src13[28] + src13[29] + src13[30] + src13[31] + src13[32] + src13[33] + src13[34] + src13[35] + src13[36] + src13[37] + src13[38] + src13[39] + src13[40] + src13[41] + src13[42] + src13[43] + src13[44] + src13[45] + src13[46] + src13[47] + src13[48] + src13[49] + src13[50] + src13[51] + src13[52] + src13[53] + src13[54] + src13[55] + src13[56] + src13[57] + src13[58] + src13[59] + src13[60] + src13[61] + src13[62] + src13[63] + src13[64] + src13[65] + src13[66] + src13[67] + src13[68] + src13[69] + src13[70] + src13[71] + src13[72] + src13[73] + src13[74] + src13[75] + src13[76] + src13[77] + src13[78] + src13[79] + src13[80] + src13[81] + src13[82] + src13[83] + src13[84] + src13[85] + src13[86] + src13[87] + src13[88] + src13[89] + src13[90] + src13[91] + src13[92] + src13[93] + src13[94] + src13[95] + src13[96] + src13[97] + src13[98] + src13[99] + src13[100] + src13[101] + src13[102] + src13[103] + src13[104] + src13[105] + src13[106] + src13[107] + src13[108] + src13[109] + src13[110] + src13[111] + src13[112] + src13[113] + src13[114] + src13[115] + src13[116] + src13[117] + src13[118] + src13[119] + src13[120] + src13[121] + src13[122] + src13[123] + src13[124] + src13[125] + src13[126] + src13[127] + src13[128] + src13[129] + src13[130] + src13[131] + src13[132] + src13[133] + src13[134] + src13[135] + src13[136] + src13[137] + src13[138] + src13[139] + src13[140] + src13[141] + src13[142] + src13[143] + src13[144] + src13[145] + src13[146] + src13[147] + src13[148] + src13[149] + src13[150] + src13[151] + src13[152] + src13[153] + src13[154] + src13[155] + src13[156] + src13[157] + src13[158] + src13[159] + src13[160] + src13[161] + src13[162] + src13[163] + src13[164] + src13[165] + src13[166] + src13[167] + src13[168] + src13[169] + src13[170] + src13[171] + src13[172] + src13[173] + src13[174] + src13[175] + src13[176] + src13[177] + src13[178] + src13[179] + src13[180] + src13[181] + src13[182] + src13[183] + src13[184] + src13[185] + src13[186] + src13[187] + src13[188] + src13[189] + src13[190] + src13[191] + src13[192] + src13[193] + src13[194] + src13[195] + src13[196] + src13[197] + src13[198] + src13[199] + src13[200] + src13[201] + src13[202] + src13[203] + src13[204] + src13[205] + src13[206] + src13[207] + src13[208] + src13[209] + src13[210] + src13[211] + src13[212] + src13[213] + src13[214] + src13[215] + src13[216] + src13[217] + src13[218] + src13[219] + src13[220] + src13[221] + src13[222] + src13[223] + src13[224] + src13[225] + src13[226] + src13[227] + src13[228] + src13[229] + src13[230] + src13[231] + src13[232] + src13[233] + src13[234] + src13[235] + src13[236] + src13[237] + src13[238] + src13[239] + src13[240] + src13[241] + src13[242] + src13[243] + src13[244] + src13[245] + src13[246] + src13[247] + src13[248] + src13[249] + src13[250] + src13[251] + src13[252] + src13[253] + src13[254] + src13[255] + src13[256] + src13[257] + src13[258] + src13[259] + src13[260] + src13[261] + src13[262] + src13[263] + src13[264] + src13[265] + src13[266] + src13[267] + src13[268] + src13[269] + src13[270] + src13[271] + src13[272] + src13[273] + src13[274] + src13[275] + src13[276] + src13[277] + src13[278] + src13[279] + src13[280] + src13[281] + src13[282] + src13[283] + src13[284] + src13[285] + src13[286] + src13[287] + src13[288] + src13[289] + src13[290] + src13[291] + src13[292] + src13[293] + src13[294] + src13[295] + src13[296] + src13[297] + src13[298] + src13[299] + src13[300] + src13[301] + src13[302] + src13[303] + src13[304] + src13[305] + src13[306] + src13[307] + src13[308] + src13[309] + src13[310] + src13[311] + src13[312] + src13[313] + src13[314] + src13[315] + src13[316] + src13[317] + src13[318] + src13[319] + src13[320] + src13[321] + src13[322] + src13[323] + src13[324] + src13[325] + src13[326] + src13[327] + src13[328] + src13[329] + src13[330] + src13[331] + src13[332] + src13[333] + src13[334] + src13[335] + src13[336] + src13[337] + src13[338] + src13[339] + src13[340] + src13[341] + src13[342] + src13[343] + src13[344] + src13[345] + src13[346] + src13[347] + src13[348] + src13[349] + src13[350] + src13[351] + src13[352] + src13[353] + src13[354] + src13[355] + src13[356] + src13[357] + src13[358] + src13[359] + src13[360] + src13[361] + src13[362] + src13[363] + src13[364] + src13[365] + src13[366] + src13[367] + src13[368] + src13[369] + src13[370] + src13[371] + src13[372] + src13[373] + src13[374] + src13[375] + src13[376] + src13[377] + src13[378] + src13[379] + src13[380] + src13[381] + src13[382] + src13[383] + src13[384] + src13[385] + src13[386] + src13[387] + src13[388] + src13[389] + src13[390] + src13[391] + src13[392] + src13[393] + src13[394] + src13[395] + src13[396] + src13[397] + src13[398] + src13[399] + src13[400] + src13[401] + src13[402] + src13[403] + src13[404] + src13[405] + src13[406] + src13[407] + src13[408] + src13[409] + src13[410] + src13[411] + src13[412] + src13[413] + src13[414] + src13[415] + src13[416] + src13[417] + src13[418] + src13[419] + src13[420] + src13[421] + src13[422] + src13[423] + src13[424] + src13[425] + src13[426] + src13[427] + src13[428] + src13[429] + src13[430] + src13[431] + src13[432] + src13[433] + src13[434] + src13[435] + src13[436] + src13[437] + src13[438] + src13[439] + src13[440] + src13[441] + src13[442] + src13[443] + src13[444] + src13[445] + src13[446] + src13[447] + src13[448] + src13[449] + src13[450] + src13[451] + src13[452] + src13[453] + src13[454] + src13[455] + src13[456] + src13[457] + src13[458] + src13[459] + src13[460] + src13[461] + src13[462] + src13[463] + src13[464] + src13[465] + src13[466] + src13[467] + src13[468] + src13[469] + src13[470] + src13[471] + src13[472] + src13[473] + src13[474] + src13[475] + src13[476] + src13[477] + src13[478] + src13[479] + src13[480] + src13[481] + src13[482] + src13[483] + src13[484] + src13[485] + src13[486] + src13[487] + src13[488] + src13[489] + src13[490] + src13[491] + src13[492] + src13[493] + src13[494] + src13[495] + src13[496] + src13[497] + src13[498] + src13[499] + src13[500] + src13[501] + src13[502] + src13[503] + src13[504] + src13[505] + src13[506] + src13[507] + src13[508] + src13[509] + src13[510] + src13[511])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14] + src14[15] + src14[16] + src14[17] + src14[18] + src14[19] + src14[20] + src14[21] + src14[22] + src14[23] + src14[24] + src14[25] + src14[26] + src14[27] + src14[28] + src14[29] + src14[30] + src14[31] + src14[32] + src14[33] + src14[34] + src14[35] + src14[36] + src14[37] + src14[38] + src14[39] + src14[40] + src14[41] + src14[42] + src14[43] + src14[44] + src14[45] + src14[46] + src14[47] + src14[48] + src14[49] + src14[50] + src14[51] + src14[52] + src14[53] + src14[54] + src14[55] + src14[56] + src14[57] + src14[58] + src14[59] + src14[60] + src14[61] + src14[62] + src14[63] + src14[64] + src14[65] + src14[66] + src14[67] + src14[68] + src14[69] + src14[70] + src14[71] + src14[72] + src14[73] + src14[74] + src14[75] + src14[76] + src14[77] + src14[78] + src14[79] + src14[80] + src14[81] + src14[82] + src14[83] + src14[84] + src14[85] + src14[86] + src14[87] + src14[88] + src14[89] + src14[90] + src14[91] + src14[92] + src14[93] + src14[94] + src14[95] + src14[96] + src14[97] + src14[98] + src14[99] + src14[100] + src14[101] + src14[102] + src14[103] + src14[104] + src14[105] + src14[106] + src14[107] + src14[108] + src14[109] + src14[110] + src14[111] + src14[112] + src14[113] + src14[114] + src14[115] + src14[116] + src14[117] + src14[118] + src14[119] + src14[120] + src14[121] + src14[122] + src14[123] + src14[124] + src14[125] + src14[126] + src14[127] + src14[128] + src14[129] + src14[130] + src14[131] + src14[132] + src14[133] + src14[134] + src14[135] + src14[136] + src14[137] + src14[138] + src14[139] + src14[140] + src14[141] + src14[142] + src14[143] + src14[144] + src14[145] + src14[146] + src14[147] + src14[148] + src14[149] + src14[150] + src14[151] + src14[152] + src14[153] + src14[154] + src14[155] + src14[156] + src14[157] + src14[158] + src14[159] + src14[160] + src14[161] + src14[162] + src14[163] + src14[164] + src14[165] + src14[166] + src14[167] + src14[168] + src14[169] + src14[170] + src14[171] + src14[172] + src14[173] + src14[174] + src14[175] + src14[176] + src14[177] + src14[178] + src14[179] + src14[180] + src14[181] + src14[182] + src14[183] + src14[184] + src14[185] + src14[186] + src14[187] + src14[188] + src14[189] + src14[190] + src14[191] + src14[192] + src14[193] + src14[194] + src14[195] + src14[196] + src14[197] + src14[198] + src14[199] + src14[200] + src14[201] + src14[202] + src14[203] + src14[204] + src14[205] + src14[206] + src14[207] + src14[208] + src14[209] + src14[210] + src14[211] + src14[212] + src14[213] + src14[214] + src14[215] + src14[216] + src14[217] + src14[218] + src14[219] + src14[220] + src14[221] + src14[222] + src14[223] + src14[224] + src14[225] + src14[226] + src14[227] + src14[228] + src14[229] + src14[230] + src14[231] + src14[232] + src14[233] + src14[234] + src14[235] + src14[236] + src14[237] + src14[238] + src14[239] + src14[240] + src14[241] + src14[242] + src14[243] + src14[244] + src14[245] + src14[246] + src14[247] + src14[248] + src14[249] + src14[250] + src14[251] + src14[252] + src14[253] + src14[254] + src14[255] + src14[256] + src14[257] + src14[258] + src14[259] + src14[260] + src14[261] + src14[262] + src14[263] + src14[264] + src14[265] + src14[266] + src14[267] + src14[268] + src14[269] + src14[270] + src14[271] + src14[272] + src14[273] + src14[274] + src14[275] + src14[276] + src14[277] + src14[278] + src14[279] + src14[280] + src14[281] + src14[282] + src14[283] + src14[284] + src14[285] + src14[286] + src14[287] + src14[288] + src14[289] + src14[290] + src14[291] + src14[292] + src14[293] + src14[294] + src14[295] + src14[296] + src14[297] + src14[298] + src14[299] + src14[300] + src14[301] + src14[302] + src14[303] + src14[304] + src14[305] + src14[306] + src14[307] + src14[308] + src14[309] + src14[310] + src14[311] + src14[312] + src14[313] + src14[314] + src14[315] + src14[316] + src14[317] + src14[318] + src14[319] + src14[320] + src14[321] + src14[322] + src14[323] + src14[324] + src14[325] + src14[326] + src14[327] + src14[328] + src14[329] + src14[330] + src14[331] + src14[332] + src14[333] + src14[334] + src14[335] + src14[336] + src14[337] + src14[338] + src14[339] + src14[340] + src14[341] + src14[342] + src14[343] + src14[344] + src14[345] + src14[346] + src14[347] + src14[348] + src14[349] + src14[350] + src14[351] + src14[352] + src14[353] + src14[354] + src14[355] + src14[356] + src14[357] + src14[358] + src14[359] + src14[360] + src14[361] + src14[362] + src14[363] + src14[364] + src14[365] + src14[366] + src14[367] + src14[368] + src14[369] + src14[370] + src14[371] + src14[372] + src14[373] + src14[374] + src14[375] + src14[376] + src14[377] + src14[378] + src14[379] + src14[380] + src14[381] + src14[382] + src14[383] + src14[384] + src14[385] + src14[386] + src14[387] + src14[388] + src14[389] + src14[390] + src14[391] + src14[392] + src14[393] + src14[394] + src14[395] + src14[396] + src14[397] + src14[398] + src14[399] + src14[400] + src14[401] + src14[402] + src14[403] + src14[404] + src14[405] + src14[406] + src14[407] + src14[408] + src14[409] + src14[410] + src14[411] + src14[412] + src14[413] + src14[414] + src14[415] + src14[416] + src14[417] + src14[418] + src14[419] + src14[420] + src14[421] + src14[422] + src14[423] + src14[424] + src14[425] + src14[426] + src14[427] + src14[428] + src14[429] + src14[430] + src14[431] + src14[432] + src14[433] + src14[434] + src14[435] + src14[436] + src14[437] + src14[438] + src14[439] + src14[440] + src14[441] + src14[442] + src14[443] + src14[444] + src14[445] + src14[446] + src14[447] + src14[448] + src14[449] + src14[450] + src14[451] + src14[452] + src14[453] + src14[454] + src14[455] + src14[456] + src14[457] + src14[458] + src14[459] + src14[460] + src14[461] + src14[462] + src14[463] + src14[464] + src14[465] + src14[466] + src14[467] + src14[468] + src14[469] + src14[470] + src14[471] + src14[472] + src14[473] + src14[474] + src14[475] + src14[476] + src14[477] + src14[478] + src14[479] + src14[480] + src14[481] + src14[482] + src14[483] + src14[484] + src14[485] + src14[486] + src14[487] + src14[488] + src14[489] + src14[490] + src14[491] + src14[492] + src14[493] + src14[494] + src14[495] + src14[496] + src14[497] + src14[498] + src14[499] + src14[500] + src14[501] + src14[502] + src14[503] + src14[504] + src14[505] + src14[506] + src14[507] + src14[508] + src14[509] + src14[510] + src14[511])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15] + src15[16] + src15[17] + src15[18] + src15[19] + src15[20] + src15[21] + src15[22] + src15[23] + src15[24] + src15[25] + src15[26] + src15[27] + src15[28] + src15[29] + src15[30] + src15[31] + src15[32] + src15[33] + src15[34] + src15[35] + src15[36] + src15[37] + src15[38] + src15[39] + src15[40] + src15[41] + src15[42] + src15[43] + src15[44] + src15[45] + src15[46] + src15[47] + src15[48] + src15[49] + src15[50] + src15[51] + src15[52] + src15[53] + src15[54] + src15[55] + src15[56] + src15[57] + src15[58] + src15[59] + src15[60] + src15[61] + src15[62] + src15[63] + src15[64] + src15[65] + src15[66] + src15[67] + src15[68] + src15[69] + src15[70] + src15[71] + src15[72] + src15[73] + src15[74] + src15[75] + src15[76] + src15[77] + src15[78] + src15[79] + src15[80] + src15[81] + src15[82] + src15[83] + src15[84] + src15[85] + src15[86] + src15[87] + src15[88] + src15[89] + src15[90] + src15[91] + src15[92] + src15[93] + src15[94] + src15[95] + src15[96] + src15[97] + src15[98] + src15[99] + src15[100] + src15[101] + src15[102] + src15[103] + src15[104] + src15[105] + src15[106] + src15[107] + src15[108] + src15[109] + src15[110] + src15[111] + src15[112] + src15[113] + src15[114] + src15[115] + src15[116] + src15[117] + src15[118] + src15[119] + src15[120] + src15[121] + src15[122] + src15[123] + src15[124] + src15[125] + src15[126] + src15[127] + src15[128] + src15[129] + src15[130] + src15[131] + src15[132] + src15[133] + src15[134] + src15[135] + src15[136] + src15[137] + src15[138] + src15[139] + src15[140] + src15[141] + src15[142] + src15[143] + src15[144] + src15[145] + src15[146] + src15[147] + src15[148] + src15[149] + src15[150] + src15[151] + src15[152] + src15[153] + src15[154] + src15[155] + src15[156] + src15[157] + src15[158] + src15[159] + src15[160] + src15[161] + src15[162] + src15[163] + src15[164] + src15[165] + src15[166] + src15[167] + src15[168] + src15[169] + src15[170] + src15[171] + src15[172] + src15[173] + src15[174] + src15[175] + src15[176] + src15[177] + src15[178] + src15[179] + src15[180] + src15[181] + src15[182] + src15[183] + src15[184] + src15[185] + src15[186] + src15[187] + src15[188] + src15[189] + src15[190] + src15[191] + src15[192] + src15[193] + src15[194] + src15[195] + src15[196] + src15[197] + src15[198] + src15[199] + src15[200] + src15[201] + src15[202] + src15[203] + src15[204] + src15[205] + src15[206] + src15[207] + src15[208] + src15[209] + src15[210] + src15[211] + src15[212] + src15[213] + src15[214] + src15[215] + src15[216] + src15[217] + src15[218] + src15[219] + src15[220] + src15[221] + src15[222] + src15[223] + src15[224] + src15[225] + src15[226] + src15[227] + src15[228] + src15[229] + src15[230] + src15[231] + src15[232] + src15[233] + src15[234] + src15[235] + src15[236] + src15[237] + src15[238] + src15[239] + src15[240] + src15[241] + src15[242] + src15[243] + src15[244] + src15[245] + src15[246] + src15[247] + src15[248] + src15[249] + src15[250] + src15[251] + src15[252] + src15[253] + src15[254] + src15[255] + src15[256] + src15[257] + src15[258] + src15[259] + src15[260] + src15[261] + src15[262] + src15[263] + src15[264] + src15[265] + src15[266] + src15[267] + src15[268] + src15[269] + src15[270] + src15[271] + src15[272] + src15[273] + src15[274] + src15[275] + src15[276] + src15[277] + src15[278] + src15[279] + src15[280] + src15[281] + src15[282] + src15[283] + src15[284] + src15[285] + src15[286] + src15[287] + src15[288] + src15[289] + src15[290] + src15[291] + src15[292] + src15[293] + src15[294] + src15[295] + src15[296] + src15[297] + src15[298] + src15[299] + src15[300] + src15[301] + src15[302] + src15[303] + src15[304] + src15[305] + src15[306] + src15[307] + src15[308] + src15[309] + src15[310] + src15[311] + src15[312] + src15[313] + src15[314] + src15[315] + src15[316] + src15[317] + src15[318] + src15[319] + src15[320] + src15[321] + src15[322] + src15[323] + src15[324] + src15[325] + src15[326] + src15[327] + src15[328] + src15[329] + src15[330] + src15[331] + src15[332] + src15[333] + src15[334] + src15[335] + src15[336] + src15[337] + src15[338] + src15[339] + src15[340] + src15[341] + src15[342] + src15[343] + src15[344] + src15[345] + src15[346] + src15[347] + src15[348] + src15[349] + src15[350] + src15[351] + src15[352] + src15[353] + src15[354] + src15[355] + src15[356] + src15[357] + src15[358] + src15[359] + src15[360] + src15[361] + src15[362] + src15[363] + src15[364] + src15[365] + src15[366] + src15[367] + src15[368] + src15[369] + src15[370] + src15[371] + src15[372] + src15[373] + src15[374] + src15[375] + src15[376] + src15[377] + src15[378] + src15[379] + src15[380] + src15[381] + src15[382] + src15[383] + src15[384] + src15[385] + src15[386] + src15[387] + src15[388] + src15[389] + src15[390] + src15[391] + src15[392] + src15[393] + src15[394] + src15[395] + src15[396] + src15[397] + src15[398] + src15[399] + src15[400] + src15[401] + src15[402] + src15[403] + src15[404] + src15[405] + src15[406] + src15[407] + src15[408] + src15[409] + src15[410] + src15[411] + src15[412] + src15[413] + src15[414] + src15[415] + src15[416] + src15[417] + src15[418] + src15[419] + src15[420] + src15[421] + src15[422] + src15[423] + src15[424] + src15[425] + src15[426] + src15[427] + src15[428] + src15[429] + src15[430] + src15[431] + src15[432] + src15[433] + src15[434] + src15[435] + src15[436] + src15[437] + src15[438] + src15[439] + src15[440] + src15[441] + src15[442] + src15[443] + src15[444] + src15[445] + src15[446] + src15[447] + src15[448] + src15[449] + src15[450] + src15[451] + src15[452] + src15[453] + src15[454] + src15[455] + src15[456] + src15[457] + src15[458] + src15[459] + src15[460] + src15[461] + src15[462] + src15[463] + src15[464] + src15[465] + src15[466] + src15[467] + src15[468] + src15[469] + src15[470] + src15[471] + src15[472] + src15[473] + src15[474] + src15[475] + src15[476] + src15[477] + src15[478] + src15[479] + src15[480] + src15[481] + src15[482] + src15[483] + src15[484] + src15[485] + src15[486] + src15[487] + src15[488] + src15[489] + src15[490] + src15[491] + src15[492] + src15[493] + src15[494] + src15[495] + src15[496] + src15[497] + src15[498] + src15[499] + src15[500] + src15[501] + src15[502] + src15[503] + src15[504] + src15[505] + src15[506] + src15[507] + src15[508] + src15[509] + src15[510] + src15[511])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16] + src16[17] + src16[18] + src16[19] + src16[20] + src16[21] + src16[22] + src16[23] + src16[24] + src16[25] + src16[26] + src16[27] + src16[28] + src16[29] + src16[30] + src16[31] + src16[32] + src16[33] + src16[34] + src16[35] + src16[36] + src16[37] + src16[38] + src16[39] + src16[40] + src16[41] + src16[42] + src16[43] + src16[44] + src16[45] + src16[46] + src16[47] + src16[48] + src16[49] + src16[50] + src16[51] + src16[52] + src16[53] + src16[54] + src16[55] + src16[56] + src16[57] + src16[58] + src16[59] + src16[60] + src16[61] + src16[62] + src16[63] + src16[64] + src16[65] + src16[66] + src16[67] + src16[68] + src16[69] + src16[70] + src16[71] + src16[72] + src16[73] + src16[74] + src16[75] + src16[76] + src16[77] + src16[78] + src16[79] + src16[80] + src16[81] + src16[82] + src16[83] + src16[84] + src16[85] + src16[86] + src16[87] + src16[88] + src16[89] + src16[90] + src16[91] + src16[92] + src16[93] + src16[94] + src16[95] + src16[96] + src16[97] + src16[98] + src16[99] + src16[100] + src16[101] + src16[102] + src16[103] + src16[104] + src16[105] + src16[106] + src16[107] + src16[108] + src16[109] + src16[110] + src16[111] + src16[112] + src16[113] + src16[114] + src16[115] + src16[116] + src16[117] + src16[118] + src16[119] + src16[120] + src16[121] + src16[122] + src16[123] + src16[124] + src16[125] + src16[126] + src16[127] + src16[128] + src16[129] + src16[130] + src16[131] + src16[132] + src16[133] + src16[134] + src16[135] + src16[136] + src16[137] + src16[138] + src16[139] + src16[140] + src16[141] + src16[142] + src16[143] + src16[144] + src16[145] + src16[146] + src16[147] + src16[148] + src16[149] + src16[150] + src16[151] + src16[152] + src16[153] + src16[154] + src16[155] + src16[156] + src16[157] + src16[158] + src16[159] + src16[160] + src16[161] + src16[162] + src16[163] + src16[164] + src16[165] + src16[166] + src16[167] + src16[168] + src16[169] + src16[170] + src16[171] + src16[172] + src16[173] + src16[174] + src16[175] + src16[176] + src16[177] + src16[178] + src16[179] + src16[180] + src16[181] + src16[182] + src16[183] + src16[184] + src16[185] + src16[186] + src16[187] + src16[188] + src16[189] + src16[190] + src16[191] + src16[192] + src16[193] + src16[194] + src16[195] + src16[196] + src16[197] + src16[198] + src16[199] + src16[200] + src16[201] + src16[202] + src16[203] + src16[204] + src16[205] + src16[206] + src16[207] + src16[208] + src16[209] + src16[210] + src16[211] + src16[212] + src16[213] + src16[214] + src16[215] + src16[216] + src16[217] + src16[218] + src16[219] + src16[220] + src16[221] + src16[222] + src16[223] + src16[224] + src16[225] + src16[226] + src16[227] + src16[228] + src16[229] + src16[230] + src16[231] + src16[232] + src16[233] + src16[234] + src16[235] + src16[236] + src16[237] + src16[238] + src16[239] + src16[240] + src16[241] + src16[242] + src16[243] + src16[244] + src16[245] + src16[246] + src16[247] + src16[248] + src16[249] + src16[250] + src16[251] + src16[252] + src16[253] + src16[254] + src16[255] + src16[256] + src16[257] + src16[258] + src16[259] + src16[260] + src16[261] + src16[262] + src16[263] + src16[264] + src16[265] + src16[266] + src16[267] + src16[268] + src16[269] + src16[270] + src16[271] + src16[272] + src16[273] + src16[274] + src16[275] + src16[276] + src16[277] + src16[278] + src16[279] + src16[280] + src16[281] + src16[282] + src16[283] + src16[284] + src16[285] + src16[286] + src16[287] + src16[288] + src16[289] + src16[290] + src16[291] + src16[292] + src16[293] + src16[294] + src16[295] + src16[296] + src16[297] + src16[298] + src16[299] + src16[300] + src16[301] + src16[302] + src16[303] + src16[304] + src16[305] + src16[306] + src16[307] + src16[308] + src16[309] + src16[310] + src16[311] + src16[312] + src16[313] + src16[314] + src16[315] + src16[316] + src16[317] + src16[318] + src16[319] + src16[320] + src16[321] + src16[322] + src16[323] + src16[324] + src16[325] + src16[326] + src16[327] + src16[328] + src16[329] + src16[330] + src16[331] + src16[332] + src16[333] + src16[334] + src16[335] + src16[336] + src16[337] + src16[338] + src16[339] + src16[340] + src16[341] + src16[342] + src16[343] + src16[344] + src16[345] + src16[346] + src16[347] + src16[348] + src16[349] + src16[350] + src16[351] + src16[352] + src16[353] + src16[354] + src16[355] + src16[356] + src16[357] + src16[358] + src16[359] + src16[360] + src16[361] + src16[362] + src16[363] + src16[364] + src16[365] + src16[366] + src16[367] + src16[368] + src16[369] + src16[370] + src16[371] + src16[372] + src16[373] + src16[374] + src16[375] + src16[376] + src16[377] + src16[378] + src16[379] + src16[380] + src16[381] + src16[382] + src16[383] + src16[384] + src16[385] + src16[386] + src16[387] + src16[388] + src16[389] + src16[390] + src16[391] + src16[392] + src16[393] + src16[394] + src16[395] + src16[396] + src16[397] + src16[398] + src16[399] + src16[400] + src16[401] + src16[402] + src16[403] + src16[404] + src16[405] + src16[406] + src16[407] + src16[408] + src16[409] + src16[410] + src16[411] + src16[412] + src16[413] + src16[414] + src16[415] + src16[416] + src16[417] + src16[418] + src16[419] + src16[420] + src16[421] + src16[422] + src16[423] + src16[424] + src16[425] + src16[426] + src16[427] + src16[428] + src16[429] + src16[430] + src16[431] + src16[432] + src16[433] + src16[434] + src16[435] + src16[436] + src16[437] + src16[438] + src16[439] + src16[440] + src16[441] + src16[442] + src16[443] + src16[444] + src16[445] + src16[446] + src16[447] + src16[448] + src16[449] + src16[450] + src16[451] + src16[452] + src16[453] + src16[454] + src16[455] + src16[456] + src16[457] + src16[458] + src16[459] + src16[460] + src16[461] + src16[462] + src16[463] + src16[464] + src16[465] + src16[466] + src16[467] + src16[468] + src16[469] + src16[470] + src16[471] + src16[472] + src16[473] + src16[474] + src16[475] + src16[476] + src16[477] + src16[478] + src16[479] + src16[480] + src16[481] + src16[482] + src16[483] + src16[484] + src16[485] + src16[486] + src16[487] + src16[488] + src16[489] + src16[490] + src16[491] + src16[492] + src16[493] + src16[494] + src16[495] + src16[496] + src16[497] + src16[498] + src16[499] + src16[500] + src16[501] + src16[502] + src16[503] + src16[504] + src16[505] + src16[506] + src16[507] + src16[508] + src16[509] + src16[510] + src16[511])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17] + src17[18] + src17[19] + src17[20] + src17[21] + src17[22] + src17[23] + src17[24] + src17[25] + src17[26] + src17[27] + src17[28] + src17[29] + src17[30] + src17[31] + src17[32] + src17[33] + src17[34] + src17[35] + src17[36] + src17[37] + src17[38] + src17[39] + src17[40] + src17[41] + src17[42] + src17[43] + src17[44] + src17[45] + src17[46] + src17[47] + src17[48] + src17[49] + src17[50] + src17[51] + src17[52] + src17[53] + src17[54] + src17[55] + src17[56] + src17[57] + src17[58] + src17[59] + src17[60] + src17[61] + src17[62] + src17[63] + src17[64] + src17[65] + src17[66] + src17[67] + src17[68] + src17[69] + src17[70] + src17[71] + src17[72] + src17[73] + src17[74] + src17[75] + src17[76] + src17[77] + src17[78] + src17[79] + src17[80] + src17[81] + src17[82] + src17[83] + src17[84] + src17[85] + src17[86] + src17[87] + src17[88] + src17[89] + src17[90] + src17[91] + src17[92] + src17[93] + src17[94] + src17[95] + src17[96] + src17[97] + src17[98] + src17[99] + src17[100] + src17[101] + src17[102] + src17[103] + src17[104] + src17[105] + src17[106] + src17[107] + src17[108] + src17[109] + src17[110] + src17[111] + src17[112] + src17[113] + src17[114] + src17[115] + src17[116] + src17[117] + src17[118] + src17[119] + src17[120] + src17[121] + src17[122] + src17[123] + src17[124] + src17[125] + src17[126] + src17[127] + src17[128] + src17[129] + src17[130] + src17[131] + src17[132] + src17[133] + src17[134] + src17[135] + src17[136] + src17[137] + src17[138] + src17[139] + src17[140] + src17[141] + src17[142] + src17[143] + src17[144] + src17[145] + src17[146] + src17[147] + src17[148] + src17[149] + src17[150] + src17[151] + src17[152] + src17[153] + src17[154] + src17[155] + src17[156] + src17[157] + src17[158] + src17[159] + src17[160] + src17[161] + src17[162] + src17[163] + src17[164] + src17[165] + src17[166] + src17[167] + src17[168] + src17[169] + src17[170] + src17[171] + src17[172] + src17[173] + src17[174] + src17[175] + src17[176] + src17[177] + src17[178] + src17[179] + src17[180] + src17[181] + src17[182] + src17[183] + src17[184] + src17[185] + src17[186] + src17[187] + src17[188] + src17[189] + src17[190] + src17[191] + src17[192] + src17[193] + src17[194] + src17[195] + src17[196] + src17[197] + src17[198] + src17[199] + src17[200] + src17[201] + src17[202] + src17[203] + src17[204] + src17[205] + src17[206] + src17[207] + src17[208] + src17[209] + src17[210] + src17[211] + src17[212] + src17[213] + src17[214] + src17[215] + src17[216] + src17[217] + src17[218] + src17[219] + src17[220] + src17[221] + src17[222] + src17[223] + src17[224] + src17[225] + src17[226] + src17[227] + src17[228] + src17[229] + src17[230] + src17[231] + src17[232] + src17[233] + src17[234] + src17[235] + src17[236] + src17[237] + src17[238] + src17[239] + src17[240] + src17[241] + src17[242] + src17[243] + src17[244] + src17[245] + src17[246] + src17[247] + src17[248] + src17[249] + src17[250] + src17[251] + src17[252] + src17[253] + src17[254] + src17[255] + src17[256] + src17[257] + src17[258] + src17[259] + src17[260] + src17[261] + src17[262] + src17[263] + src17[264] + src17[265] + src17[266] + src17[267] + src17[268] + src17[269] + src17[270] + src17[271] + src17[272] + src17[273] + src17[274] + src17[275] + src17[276] + src17[277] + src17[278] + src17[279] + src17[280] + src17[281] + src17[282] + src17[283] + src17[284] + src17[285] + src17[286] + src17[287] + src17[288] + src17[289] + src17[290] + src17[291] + src17[292] + src17[293] + src17[294] + src17[295] + src17[296] + src17[297] + src17[298] + src17[299] + src17[300] + src17[301] + src17[302] + src17[303] + src17[304] + src17[305] + src17[306] + src17[307] + src17[308] + src17[309] + src17[310] + src17[311] + src17[312] + src17[313] + src17[314] + src17[315] + src17[316] + src17[317] + src17[318] + src17[319] + src17[320] + src17[321] + src17[322] + src17[323] + src17[324] + src17[325] + src17[326] + src17[327] + src17[328] + src17[329] + src17[330] + src17[331] + src17[332] + src17[333] + src17[334] + src17[335] + src17[336] + src17[337] + src17[338] + src17[339] + src17[340] + src17[341] + src17[342] + src17[343] + src17[344] + src17[345] + src17[346] + src17[347] + src17[348] + src17[349] + src17[350] + src17[351] + src17[352] + src17[353] + src17[354] + src17[355] + src17[356] + src17[357] + src17[358] + src17[359] + src17[360] + src17[361] + src17[362] + src17[363] + src17[364] + src17[365] + src17[366] + src17[367] + src17[368] + src17[369] + src17[370] + src17[371] + src17[372] + src17[373] + src17[374] + src17[375] + src17[376] + src17[377] + src17[378] + src17[379] + src17[380] + src17[381] + src17[382] + src17[383] + src17[384] + src17[385] + src17[386] + src17[387] + src17[388] + src17[389] + src17[390] + src17[391] + src17[392] + src17[393] + src17[394] + src17[395] + src17[396] + src17[397] + src17[398] + src17[399] + src17[400] + src17[401] + src17[402] + src17[403] + src17[404] + src17[405] + src17[406] + src17[407] + src17[408] + src17[409] + src17[410] + src17[411] + src17[412] + src17[413] + src17[414] + src17[415] + src17[416] + src17[417] + src17[418] + src17[419] + src17[420] + src17[421] + src17[422] + src17[423] + src17[424] + src17[425] + src17[426] + src17[427] + src17[428] + src17[429] + src17[430] + src17[431] + src17[432] + src17[433] + src17[434] + src17[435] + src17[436] + src17[437] + src17[438] + src17[439] + src17[440] + src17[441] + src17[442] + src17[443] + src17[444] + src17[445] + src17[446] + src17[447] + src17[448] + src17[449] + src17[450] + src17[451] + src17[452] + src17[453] + src17[454] + src17[455] + src17[456] + src17[457] + src17[458] + src17[459] + src17[460] + src17[461] + src17[462] + src17[463] + src17[464] + src17[465] + src17[466] + src17[467] + src17[468] + src17[469] + src17[470] + src17[471] + src17[472] + src17[473] + src17[474] + src17[475] + src17[476] + src17[477] + src17[478] + src17[479] + src17[480] + src17[481] + src17[482] + src17[483] + src17[484] + src17[485] + src17[486] + src17[487] + src17[488] + src17[489] + src17[490] + src17[491] + src17[492] + src17[493] + src17[494] + src17[495] + src17[496] + src17[497] + src17[498] + src17[499] + src17[500] + src17[501] + src17[502] + src17[503] + src17[504] + src17[505] + src17[506] + src17[507] + src17[508] + src17[509] + src17[510] + src17[511])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15] + src18[16] + src18[17] + src18[18] + src18[19] + src18[20] + src18[21] + src18[22] + src18[23] + src18[24] + src18[25] + src18[26] + src18[27] + src18[28] + src18[29] + src18[30] + src18[31] + src18[32] + src18[33] + src18[34] + src18[35] + src18[36] + src18[37] + src18[38] + src18[39] + src18[40] + src18[41] + src18[42] + src18[43] + src18[44] + src18[45] + src18[46] + src18[47] + src18[48] + src18[49] + src18[50] + src18[51] + src18[52] + src18[53] + src18[54] + src18[55] + src18[56] + src18[57] + src18[58] + src18[59] + src18[60] + src18[61] + src18[62] + src18[63] + src18[64] + src18[65] + src18[66] + src18[67] + src18[68] + src18[69] + src18[70] + src18[71] + src18[72] + src18[73] + src18[74] + src18[75] + src18[76] + src18[77] + src18[78] + src18[79] + src18[80] + src18[81] + src18[82] + src18[83] + src18[84] + src18[85] + src18[86] + src18[87] + src18[88] + src18[89] + src18[90] + src18[91] + src18[92] + src18[93] + src18[94] + src18[95] + src18[96] + src18[97] + src18[98] + src18[99] + src18[100] + src18[101] + src18[102] + src18[103] + src18[104] + src18[105] + src18[106] + src18[107] + src18[108] + src18[109] + src18[110] + src18[111] + src18[112] + src18[113] + src18[114] + src18[115] + src18[116] + src18[117] + src18[118] + src18[119] + src18[120] + src18[121] + src18[122] + src18[123] + src18[124] + src18[125] + src18[126] + src18[127] + src18[128] + src18[129] + src18[130] + src18[131] + src18[132] + src18[133] + src18[134] + src18[135] + src18[136] + src18[137] + src18[138] + src18[139] + src18[140] + src18[141] + src18[142] + src18[143] + src18[144] + src18[145] + src18[146] + src18[147] + src18[148] + src18[149] + src18[150] + src18[151] + src18[152] + src18[153] + src18[154] + src18[155] + src18[156] + src18[157] + src18[158] + src18[159] + src18[160] + src18[161] + src18[162] + src18[163] + src18[164] + src18[165] + src18[166] + src18[167] + src18[168] + src18[169] + src18[170] + src18[171] + src18[172] + src18[173] + src18[174] + src18[175] + src18[176] + src18[177] + src18[178] + src18[179] + src18[180] + src18[181] + src18[182] + src18[183] + src18[184] + src18[185] + src18[186] + src18[187] + src18[188] + src18[189] + src18[190] + src18[191] + src18[192] + src18[193] + src18[194] + src18[195] + src18[196] + src18[197] + src18[198] + src18[199] + src18[200] + src18[201] + src18[202] + src18[203] + src18[204] + src18[205] + src18[206] + src18[207] + src18[208] + src18[209] + src18[210] + src18[211] + src18[212] + src18[213] + src18[214] + src18[215] + src18[216] + src18[217] + src18[218] + src18[219] + src18[220] + src18[221] + src18[222] + src18[223] + src18[224] + src18[225] + src18[226] + src18[227] + src18[228] + src18[229] + src18[230] + src18[231] + src18[232] + src18[233] + src18[234] + src18[235] + src18[236] + src18[237] + src18[238] + src18[239] + src18[240] + src18[241] + src18[242] + src18[243] + src18[244] + src18[245] + src18[246] + src18[247] + src18[248] + src18[249] + src18[250] + src18[251] + src18[252] + src18[253] + src18[254] + src18[255] + src18[256] + src18[257] + src18[258] + src18[259] + src18[260] + src18[261] + src18[262] + src18[263] + src18[264] + src18[265] + src18[266] + src18[267] + src18[268] + src18[269] + src18[270] + src18[271] + src18[272] + src18[273] + src18[274] + src18[275] + src18[276] + src18[277] + src18[278] + src18[279] + src18[280] + src18[281] + src18[282] + src18[283] + src18[284] + src18[285] + src18[286] + src18[287] + src18[288] + src18[289] + src18[290] + src18[291] + src18[292] + src18[293] + src18[294] + src18[295] + src18[296] + src18[297] + src18[298] + src18[299] + src18[300] + src18[301] + src18[302] + src18[303] + src18[304] + src18[305] + src18[306] + src18[307] + src18[308] + src18[309] + src18[310] + src18[311] + src18[312] + src18[313] + src18[314] + src18[315] + src18[316] + src18[317] + src18[318] + src18[319] + src18[320] + src18[321] + src18[322] + src18[323] + src18[324] + src18[325] + src18[326] + src18[327] + src18[328] + src18[329] + src18[330] + src18[331] + src18[332] + src18[333] + src18[334] + src18[335] + src18[336] + src18[337] + src18[338] + src18[339] + src18[340] + src18[341] + src18[342] + src18[343] + src18[344] + src18[345] + src18[346] + src18[347] + src18[348] + src18[349] + src18[350] + src18[351] + src18[352] + src18[353] + src18[354] + src18[355] + src18[356] + src18[357] + src18[358] + src18[359] + src18[360] + src18[361] + src18[362] + src18[363] + src18[364] + src18[365] + src18[366] + src18[367] + src18[368] + src18[369] + src18[370] + src18[371] + src18[372] + src18[373] + src18[374] + src18[375] + src18[376] + src18[377] + src18[378] + src18[379] + src18[380] + src18[381] + src18[382] + src18[383] + src18[384] + src18[385] + src18[386] + src18[387] + src18[388] + src18[389] + src18[390] + src18[391] + src18[392] + src18[393] + src18[394] + src18[395] + src18[396] + src18[397] + src18[398] + src18[399] + src18[400] + src18[401] + src18[402] + src18[403] + src18[404] + src18[405] + src18[406] + src18[407] + src18[408] + src18[409] + src18[410] + src18[411] + src18[412] + src18[413] + src18[414] + src18[415] + src18[416] + src18[417] + src18[418] + src18[419] + src18[420] + src18[421] + src18[422] + src18[423] + src18[424] + src18[425] + src18[426] + src18[427] + src18[428] + src18[429] + src18[430] + src18[431] + src18[432] + src18[433] + src18[434] + src18[435] + src18[436] + src18[437] + src18[438] + src18[439] + src18[440] + src18[441] + src18[442] + src18[443] + src18[444] + src18[445] + src18[446] + src18[447] + src18[448] + src18[449] + src18[450] + src18[451] + src18[452] + src18[453] + src18[454] + src18[455] + src18[456] + src18[457] + src18[458] + src18[459] + src18[460] + src18[461] + src18[462] + src18[463] + src18[464] + src18[465] + src18[466] + src18[467] + src18[468] + src18[469] + src18[470] + src18[471] + src18[472] + src18[473] + src18[474] + src18[475] + src18[476] + src18[477] + src18[478] + src18[479] + src18[480] + src18[481] + src18[482] + src18[483] + src18[484] + src18[485] + src18[486] + src18[487] + src18[488] + src18[489] + src18[490] + src18[491] + src18[492] + src18[493] + src18[494] + src18[495] + src18[496] + src18[497] + src18[498] + src18[499] + src18[500] + src18[501] + src18[502] + src18[503] + src18[504] + src18[505] + src18[506] + src18[507] + src18[508] + src18[509] + src18[510] + src18[511])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13] + src19[14] + src19[15] + src19[16] + src19[17] + src19[18] + src19[19] + src19[20] + src19[21] + src19[22] + src19[23] + src19[24] + src19[25] + src19[26] + src19[27] + src19[28] + src19[29] + src19[30] + src19[31] + src19[32] + src19[33] + src19[34] + src19[35] + src19[36] + src19[37] + src19[38] + src19[39] + src19[40] + src19[41] + src19[42] + src19[43] + src19[44] + src19[45] + src19[46] + src19[47] + src19[48] + src19[49] + src19[50] + src19[51] + src19[52] + src19[53] + src19[54] + src19[55] + src19[56] + src19[57] + src19[58] + src19[59] + src19[60] + src19[61] + src19[62] + src19[63] + src19[64] + src19[65] + src19[66] + src19[67] + src19[68] + src19[69] + src19[70] + src19[71] + src19[72] + src19[73] + src19[74] + src19[75] + src19[76] + src19[77] + src19[78] + src19[79] + src19[80] + src19[81] + src19[82] + src19[83] + src19[84] + src19[85] + src19[86] + src19[87] + src19[88] + src19[89] + src19[90] + src19[91] + src19[92] + src19[93] + src19[94] + src19[95] + src19[96] + src19[97] + src19[98] + src19[99] + src19[100] + src19[101] + src19[102] + src19[103] + src19[104] + src19[105] + src19[106] + src19[107] + src19[108] + src19[109] + src19[110] + src19[111] + src19[112] + src19[113] + src19[114] + src19[115] + src19[116] + src19[117] + src19[118] + src19[119] + src19[120] + src19[121] + src19[122] + src19[123] + src19[124] + src19[125] + src19[126] + src19[127] + src19[128] + src19[129] + src19[130] + src19[131] + src19[132] + src19[133] + src19[134] + src19[135] + src19[136] + src19[137] + src19[138] + src19[139] + src19[140] + src19[141] + src19[142] + src19[143] + src19[144] + src19[145] + src19[146] + src19[147] + src19[148] + src19[149] + src19[150] + src19[151] + src19[152] + src19[153] + src19[154] + src19[155] + src19[156] + src19[157] + src19[158] + src19[159] + src19[160] + src19[161] + src19[162] + src19[163] + src19[164] + src19[165] + src19[166] + src19[167] + src19[168] + src19[169] + src19[170] + src19[171] + src19[172] + src19[173] + src19[174] + src19[175] + src19[176] + src19[177] + src19[178] + src19[179] + src19[180] + src19[181] + src19[182] + src19[183] + src19[184] + src19[185] + src19[186] + src19[187] + src19[188] + src19[189] + src19[190] + src19[191] + src19[192] + src19[193] + src19[194] + src19[195] + src19[196] + src19[197] + src19[198] + src19[199] + src19[200] + src19[201] + src19[202] + src19[203] + src19[204] + src19[205] + src19[206] + src19[207] + src19[208] + src19[209] + src19[210] + src19[211] + src19[212] + src19[213] + src19[214] + src19[215] + src19[216] + src19[217] + src19[218] + src19[219] + src19[220] + src19[221] + src19[222] + src19[223] + src19[224] + src19[225] + src19[226] + src19[227] + src19[228] + src19[229] + src19[230] + src19[231] + src19[232] + src19[233] + src19[234] + src19[235] + src19[236] + src19[237] + src19[238] + src19[239] + src19[240] + src19[241] + src19[242] + src19[243] + src19[244] + src19[245] + src19[246] + src19[247] + src19[248] + src19[249] + src19[250] + src19[251] + src19[252] + src19[253] + src19[254] + src19[255] + src19[256] + src19[257] + src19[258] + src19[259] + src19[260] + src19[261] + src19[262] + src19[263] + src19[264] + src19[265] + src19[266] + src19[267] + src19[268] + src19[269] + src19[270] + src19[271] + src19[272] + src19[273] + src19[274] + src19[275] + src19[276] + src19[277] + src19[278] + src19[279] + src19[280] + src19[281] + src19[282] + src19[283] + src19[284] + src19[285] + src19[286] + src19[287] + src19[288] + src19[289] + src19[290] + src19[291] + src19[292] + src19[293] + src19[294] + src19[295] + src19[296] + src19[297] + src19[298] + src19[299] + src19[300] + src19[301] + src19[302] + src19[303] + src19[304] + src19[305] + src19[306] + src19[307] + src19[308] + src19[309] + src19[310] + src19[311] + src19[312] + src19[313] + src19[314] + src19[315] + src19[316] + src19[317] + src19[318] + src19[319] + src19[320] + src19[321] + src19[322] + src19[323] + src19[324] + src19[325] + src19[326] + src19[327] + src19[328] + src19[329] + src19[330] + src19[331] + src19[332] + src19[333] + src19[334] + src19[335] + src19[336] + src19[337] + src19[338] + src19[339] + src19[340] + src19[341] + src19[342] + src19[343] + src19[344] + src19[345] + src19[346] + src19[347] + src19[348] + src19[349] + src19[350] + src19[351] + src19[352] + src19[353] + src19[354] + src19[355] + src19[356] + src19[357] + src19[358] + src19[359] + src19[360] + src19[361] + src19[362] + src19[363] + src19[364] + src19[365] + src19[366] + src19[367] + src19[368] + src19[369] + src19[370] + src19[371] + src19[372] + src19[373] + src19[374] + src19[375] + src19[376] + src19[377] + src19[378] + src19[379] + src19[380] + src19[381] + src19[382] + src19[383] + src19[384] + src19[385] + src19[386] + src19[387] + src19[388] + src19[389] + src19[390] + src19[391] + src19[392] + src19[393] + src19[394] + src19[395] + src19[396] + src19[397] + src19[398] + src19[399] + src19[400] + src19[401] + src19[402] + src19[403] + src19[404] + src19[405] + src19[406] + src19[407] + src19[408] + src19[409] + src19[410] + src19[411] + src19[412] + src19[413] + src19[414] + src19[415] + src19[416] + src19[417] + src19[418] + src19[419] + src19[420] + src19[421] + src19[422] + src19[423] + src19[424] + src19[425] + src19[426] + src19[427] + src19[428] + src19[429] + src19[430] + src19[431] + src19[432] + src19[433] + src19[434] + src19[435] + src19[436] + src19[437] + src19[438] + src19[439] + src19[440] + src19[441] + src19[442] + src19[443] + src19[444] + src19[445] + src19[446] + src19[447] + src19[448] + src19[449] + src19[450] + src19[451] + src19[452] + src19[453] + src19[454] + src19[455] + src19[456] + src19[457] + src19[458] + src19[459] + src19[460] + src19[461] + src19[462] + src19[463] + src19[464] + src19[465] + src19[466] + src19[467] + src19[468] + src19[469] + src19[470] + src19[471] + src19[472] + src19[473] + src19[474] + src19[475] + src19[476] + src19[477] + src19[478] + src19[479] + src19[480] + src19[481] + src19[482] + src19[483] + src19[484] + src19[485] + src19[486] + src19[487] + src19[488] + src19[489] + src19[490] + src19[491] + src19[492] + src19[493] + src19[494] + src19[495] + src19[496] + src19[497] + src19[498] + src19[499] + src19[500] + src19[501] + src19[502] + src19[503] + src19[504] + src19[505] + src19[506] + src19[507] + src19[508] + src19[509] + src19[510] + src19[511])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6] + src20[7] + src20[8] + src20[9] + src20[10] + src20[11] + src20[12] + src20[13] + src20[14] + src20[15] + src20[16] + src20[17] + src20[18] + src20[19] + src20[20] + src20[21] + src20[22] + src20[23] + src20[24] + src20[25] + src20[26] + src20[27] + src20[28] + src20[29] + src20[30] + src20[31] + src20[32] + src20[33] + src20[34] + src20[35] + src20[36] + src20[37] + src20[38] + src20[39] + src20[40] + src20[41] + src20[42] + src20[43] + src20[44] + src20[45] + src20[46] + src20[47] + src20[48] + src20[49] + src20[50] + src20[51] + src20[52] + src20[53] + src20[54] + src20[55] + src20[56] + src20[57] + src20[58] + src20[59] + src20[60] + src20[61] + src20[62] + src20[63] + src20[64] + src20[65] + src20[66] + src20[67] + src20[68] + src20[69] + src20[70] + src20[71] + src20[72] + src20[73] + src20[74] + src20[75] + src20[76] + src20[77] + src20[78] + src20[79] + src20[80] + src20[81] + src20[82] + src20[83] + src20[84] + src20[85] + src20[86] + src20[87] + src20[88] + src20[89] + src20[90] + src20[91] + src20[92] + src20[93] + src20[94] + src20[95] + src20[96] + src20[97] + src20[98] + src20[99] + src20[100] + src20[101] + src20[102] + src20[103] + src20[104] + src20[105] + src20[106] + src20[107] + src20[108] + src20[109] + src20[110] + src20[111] + src20[112] + src20[113] + src20[114] + src20[115] + src20[116] + src20[117] + src20[118] + src20[119] + src20[120] + src20[121] + src20[122] + src20[123] + src20[124] + src20[125] + src20[126] + src20[127] + src20[128] + src20[129] + src20[130] + src20[131] + src20[132] + src20[133] + src20[134] + src20[135] + src20[136] + src20[137] + src20[138] + src20[139] + src20[140] + src20[141] + src20[142] + src20[143] + src20[144] + src20[145] + src20[146] + src20[147] + src20[148] + src20[149] + src20[150] + src20[151] + src20[152] + src20[153] + src20[154] + src20[155] + src20[156] + src20[157] + src20[158] + src20[159] + src20[160] + src20[161] + src20[162] + src20[163] + src20[164] + src20[165] + src20[166] + src20[167] + src20[168] + src20[169] + src20[170] + src20[171] + src20[172] + src20[173] + src20[174] + src20[175] + src20[176] + src20[177] + src20[178] + src20[179] + src20[180] + src20[181] + src20[182] + src20[183] + src20[184] + src20[185] + src20[186] + src20[187] + src20[188] + src20[189] + src20[190] + src20[191] + src20[192] + src20[193] + src20[194] + src20[195] + src20[196] + src20[197] + src20[198] + src20[199] + src20[200] + src20[201] + src20[202] + src20[203] + src20[204] + src20[205] + src20[206] + src20[207] + src20[208] + src20[209] + src20[210] + src20[211] + src20[212] + src20[213] + src20[214] + src20[215] + src20[216] + src20[217] + src20[218] + src20[219] + src20[220] + src20[221] + src20[222] + src20[223] + src20[224] + src20[225] + src20[226] + src20[227] + src20[228] + src20[229] + src20[230] + src20[231] + src20[232] + src20[233] + src20[234] + src20[235] + src20[236] + src20[237] + src20[238] + src20[239] + src20[240] + src20[241] + src20[242] + src20[243] + src20[244] + src20[245] + src20[246] + src20[247] + src20[248] + src20[249] + src20[250] + src20[251] + src20[252] + src20[253] + src20[254] + src20[255] + src20[256] + src20[257] + src20[258] + src20[259] + src20[260] + src20[261] + src20[262] + src20[263] + src20[264] + src20[265] + src20[266] + src20[267] + src20[268] + src20[269] + src20[270] + src20[271] + src20[272] + src20[273] + src20[274] + src20[275] + src20[276] + src20[277] + src20[278] + src20[279] + src20[280] + src20[281] + src20[282] + src20[283] + src20[284] + src20[285] + src20[286] + src20[287] + src20[288] + src20[289] + src20[290] + src20[291] + src20[292] + src20[293] + src20[294] + src20[295] + src20[296] + src20[297] + src20[298] + src20[299] + src20[300] + src20[301] + src20[302] + src20[303] + src20[304] + src20[305] + src20[306] + src20[307] + src20[308] + src20[309] + src20[310] + src20[311] + src20[312] + src20[313] + src20[314] + src20[315] + src20[316] + src20[317] + src20[318] + src20[319] + src20[320] + src20[321] + src20[322] + src20[323] + src20[324] + src20[325] + src20[326] + src20[327] + src20[328] + src20[329] + src20[330] + src20[331] + src20[332] + src20[333] + src20[334] + src20[335] + src20[336] + src20[337] + src20[338] + src20[339] + src20[340] + src20[341] + src20[342] + src20[343] + src20[344] + src20[345] + src20[346] + src20[347] + src20[348] + src20[349] + src20[350] + src20[351] + src20[352] + src20[353] + src20[354] + src20[355] + src20[356] + src20[357] + src20[358] + src20[359] + src20[360] + src20[361] + src20[362] + src20[363] + src20[364] + src20[365] + src20[366] + src20[367] + src20[368] + src20[369] + src20[370] + src20[371] + src20[372] + src20[373] + src20[374] + src20[375] + src20[376] + src20[377] + src20[378] + src20[379] + src20[380] + src20[381] + src20[382] + src20[383] + src20[384] + src20[385] + src20[386] + src20[387] + src20[388] + src20[389] + src20[390] + src20[391] + src20[392] + src20[393] + src20[394] + src20[395] + src20[396] + src20[397] + src20[398] + src20[399] + src20[400] + src20[401] + src20[402] + src20[403] + src20[404] + src20[405] + src20[406] + src20[407] + src20[408] + src20[409] + src20[410] + src20[411] + src20[412] + src20[413] + src20[414] + src20[415] + src20[416] + src20[417] + src20[418] + src20[419] + src20[420] + src20[421] + src20[422] + src20[423] + src20[424] + src20[425] + src20[426] + src20[427] + src20[428] + src20[429] + src20[430] + src20[431] + src20[432] + src20[433] + src20[434] + src20[435] + src20[436] + src20[437] + src20[438] + src20[439] + src20[440] + src20[441] + src20[442] + src20[443] + src20[444] + src20[445] + src20[446] + src20[447] + src20[448] + src20[449] + src20[450] + src20[451] + src20[452] + src20[453] + src20[454] + src20[455] + src20[456] + src20[457] + src20[458] + src20[459] + src20[460] + src20[461] + src20[462] + src20[463] + src20[464] + src20[465] + src20[466] + src20[467] + src20[468] + src20[469] + src20[470] + src20[471] + src20[472] + src20[473] + src20[474] + src20[475] + src20[476] + src20[477] + src20[478] + src20[479] + src20[480] + src20[481] + src20[482] + src20[483] + src20[484] + src20[485] + src20[486] + src20[487] + src20[488] + src20[489] + src20[490] + src20[491] + src20[492] + src20[493] + src20[494] + src20[495] + src20[496] + src20[497] + src20[498] + src20[499] + src20[500] + src20[501] + src20[502] + src20[503] + src20[504] + src20[505] + src20[506] + src20[507] + src20[508] + src20[509] + src20[510] + src20[511])<<20) + ((src21[0] + src21[1] + src21[2] + src21[3] + src21[4] + src21[5] + src21[6] + src21[7] + src21[8] + src21[9] + src21[10] + src21[11] + src21[12] + src21[13] + src21[14] + src21[15] + src21[16] + src21[17] + src21[18] + src21[19] + src21[20] + src21[21] + src21[22] + src21[23] + src21[24] + src21[25] + src21[26] + src21[27] + src21[28] + src21[29] + src21[30] + src21[31] + src21[32] + src21[33] + src21[34] + src21[35] + src21[36] + src21[37] + src21[38] + src21[39] + src21[40] + src21[41] + src21[42] + src21[43] + src21[44] + src21[45] + src21[46] + src21[47] + src21[48] + src21[49] + src21[50] + src21[51] + src21[52] + src21[53] + src21[54] + src21[55] + src21[56] + src21[57] + src21[58] + src21[59] + src21[60] + src21[61] + src21[62] + src21[63] + src21[64] + src21[65] + src21[66] + src21[67] + src21[68] + src21[69] + src21[70] + src21[71] + src21[72] + src21[73] + src21[74] + src21[75] + src21[76] + src21[77] + src21[78] + src21[79] + src21[80] + src21[81] + src21[82] + src21[83] + src21[84] + src21[85] + src21[86] + src21[87] + src21[88] + src21[89] + src21[90] + src21[91] + src21[92] + src21[93] + src21[94] + src21[95] + src21[96] + src21[97] + src21[98] + src21[99] + src21[100] + src21[101] + src21[102] + src21[103] + src21[104] + src21[105] + src21[106] + src21[107] + src21[108] + src21[109] + src21[110] + src21[111] + src21[112] + src21[113] + src21[114] + src21[115] + src21[116] + src21[117] + src21[118] + src21[119] + src21[120] + src21[121] + src21[122] + src21[123] + src21[124] + src21[125] + src21[126] + src21[127] + src21[128] + src21[129] + src21[130] + src21[131] + src21[132] + src21[133] + src21[134] + src21[135] + src21[136] + src21[137] + src21[138] + src21[139] + src21[140] + src21[141] + src21[142] + src21[143] + src21[144] + src21[145] + src21[146] + src21[147] + src21[148] + src21[149] + src21[150] + src21[151] + src21[152] + src21[153] + src21[154] + src21[155] + src21[156] + src21[157] + src21[158] + src21[159] + src21[160] + src21[161] + src21[162] + src21[163] + src21[164] + src21[165] + src21[166] + src21[167] + src21[168] + src21[169] + src21[170] + src21[171] + src21[172] + src21[173] + src21[174] + src21[175] + src21[176] + src21[177] + src21[178] + src21[179] + src21[180] + src21[181] + src21[182] + src21[183] + src21[184] + src21[185] + src21[186] + src21[187] + src21[188] + src21[189] + src21[190] + src21[191] + src21[192] + src21[193] + src21[194] + src21[195] + src21[196] + src21[197] + src21[198] + src21[199] + src21[200] + src21[201] + src21[202] + src21[203] + src21[204] + src21[205] + src21[206] + src21[207] + src21[208] + src21[209] + src21[210] + src21[211] + src21[212] + src21[213] + src21[214] + src21[215] + src21[216] + src21[217] + src21[218] + src21[219] + src21[220] + src21[221] + src21[222] + src21[223] + src21[224] + src21[225] + src21[226] + src21[227] + src21[228] + src21[229] + src21[230] + src21[231] + src21[232] + src21[233] + src21[234] + src21[235] + src21[236] + src21[237] + src21[238] + src21[239] + src21[240] + src21[241] + src21[242] + src21[243] + src21[244] + src21[245] + src21[246] + src21[247] + src21[248] + src21[249] + src21[250] + src21[251] + src21[252] + src21[253] + src21[254] + src21[255] + src21[256] + src21[257] + src21[258] + src21[259] + src21[260] + src21[261] + src21[262] + src21[263] + src21[264] + src21[265] + src21[266] + src21[267] + src21[268] + src21[269] + src21[270] + src21[271] + src21[272] + src21[273] + src21[274] + src21[275] + src21[276] + src21[277] + src21[278] + src21[279] + src21[280] + src21[281] + src21[282] + src21[283] + src21[284] + src21[285] + src21[286] + src21[287] + src21[288] + src21[289] + src21[290] + src21[291] + src21[292] + src21[293] + src21[294] + src21[295] + src21[296] + src21[297] + src21[298] + src21[299] + src21[300] + src21[301] + src21[302] + src21[303] + src21[304] + src21[305] + src21[306] + src21[307] + src21[308] + src21[309] + src21[310] + src21[311] + src21[312] + src21[313] + src21[314] + src21[315] + src21[316] + src21[317] + src21[318] + src21[319] + src21[320] + src21[321] + src21[322] + src21[323] + src21[324] + src21[325] + src21[326] + src21[327] + src21[328] + src21[329] + src21[330] + src21[331] + src21[332] + src21[333] + src21[334] + src21[335] + src21[336] + src21[337] + src21[338] + src21[339] + src21[340] + src21[341] + src21[342] + src21[343] + src21[344] + src21[345] + src21[346] + src21[347] + src21[348] + src21[349] + src21[350] + src21[351] + src21[352] + src21[353] + src21[354] + src21[355] + src21[356] + src21[357] + src21[358] + src21[359] + src21[360] + src21[361] + src21[362] + src21[363] + src21[364] + src21[365] + src21[366] + src21[367] + src21[368] + src21[369] + src21[370] + src21[371] + src21[372] + src21[373] + src21[374] + src21[375] + src21[376] + src21[377] + src21[378] + src21[379] + src21[380] + src21[381] + src21[382] + src21[383] + src21[384] + src21[385] + src21[386] + src21[387] + src21[388] + src21[389] + src21[390] + src21[391] + src21[392] + src21[393] + src21[394] + src21[395] + src21[396] + src21[397] + src21[398] + src21[399] + src21[400] + src21[401] + src21[402] + src21[403] + src21[404] + src21[405] + src21[406] + src21[407] + src21[408] + src21[409] + src21[410] + src21[411] + src21[412] + src21[413] + src21[414] + src21[415] + src21[416] + src21[417] + src21[418] + src21[419] + src21[420] + src21[421] + src21[422] + src21[423] + src21[424] + src21[425] + src21[426] + src21[427] + src21[428] + src21[429] + src21[430] + src21[431] + src21[432] + src21[433] + src21[434] + src21[435] + src21[436] + src21[437] + src21[438] + src21[439] + src21[440] + src21[441] + src21[442] + src21[443] + src21[444] + src21[445] + src21[446] + src21[447] + src21[448] + src21[449] + src21[450] + src21[451] + src21[452] + src21[453] + src21[454] + src21[455] + src21[456] + src21[457] + src21[458] + src21[459] + src21[460] + src21[461] + src21[462] + src21[463] + src21[464] + src21[465] + src21[466] + src21[467] + src21[468] + src21[469] + src21[470] + src21[471] + src21[472] + src21[473] + src21[474] + src21[475] + src21[476] + src21[477] + src21[478] + src21[479] + src21[480] + src21[481] + src21[482] + src21[483] + src21[484] + src21[485] + src21[486] + src21[487] + src21[488] + src21[489] + src21[490] + src21[491] + src21[492] + src21[493] + src21[494] + src21[495] + src21[496] + src21[497] + src21[498] + src21[499] + src21[500] + src21[501] + src21[502] + src21[503] + src21[504] + src21[505] + src21[506] + src21[507] + src21[508] + src21[509] + src21[510] + src21[511])<<21) + ((src22[0] + src22[1] + src22[2] + src22[3] + src22[4] + src22[5] + src22[6] + src22[7] + src22[8] + src22[9] + src22[10] + src22[11] + src22[12] + src22[13] + src22[14] + src22[15] + src22[16] + src22[17] + src22[18] + src22[19] + src22[20] + src22[21] + src22[22] + src22[23] + src22[24] + src22[25] + src22[26] + src22[27] + src22[28] + src22[29] + src22[30] + src22[31] + src22[32] + src22[33] + src22[34] + src22[35] + src22[36] + src22[37] + src22[38] + src22[39] + src22[40] + src22[41] + src22[42] + src22[43] + src22[44] + src22[45] + src22[46] + src22[47] + src22[48] + src22[49] + src22[50] + src22[51] + src22[52] + src22[53] + src22[54] + src22[55] + src22[56] + src22[57] + src22[58] + src22[59] + src22[60] + src22[61] + src22[62] + src22[63] + src22[64] + src22[65] + src22[66] + src22[67] + src22[68] + src22[69] + src22[70] + src22[71] + src22[72] + src22[73] + src22[74] + src22[75] + src22[76] + src22[77] + src22[78] + src22[79] + src22[80] + src22[81] + src22[82] + src22[83] + src22[84] + src22[85] + src22[86] + src22[87] + src22[88] + src22[89] + src22[90] + src22[91] + src22[92] + src22[93] + src22[94] + src22[95] + src22[96] + src22[97] + src22[98] + src22[99] + src22[100] + src22[101] + src22[102] + src22[103] + src22[104] + src22[105] + src22[106] + src22[107] + src22[108] + src22[109] + src22[110] + src22[111] + src22[112] + src22[113] + src22[114] + src22[115] + src22[116] + src22[117] + src22[118] + src22[119] + src22[120] + src22[121] + src22[122] + src22[123] + src22[124] + src22[125] + src22[126] + src22[127] + src22[128] + src22[129] + src22[130] + src22[131] + src22[132] + src22[133] + src22[134] + src22[135] + src22[136] + src22[137] + src22[138] + src22[139] + src22[140] + src22[141] + src22[142] + src22[143] + src22[144] + src22[145] + src22[146] + src22[147] + src22[148] + src22[149] + src22[150] + src22[151] + src22[152] + src22[153] + src22[154] + src22[155] + src22[156] + src22[157] + src22[158] + src22[159] + src22[160] + src22[161] + src22[162] + src22[163] + src22[164] + src22[165] + src22[166] + src22[167] + src22[168] + src22[169] + src22[170] + src22[171] + src22[172] + src22[173] + src22[174] + src22[175] + src22[176] + src22[177] + src22[178] + src22[179] + src22[180] + src22[181] + src22[182] + src22[183] + src22[184] + src22[185] + src22[186] + src22[187] + src22[188] + src22[189] + src22[190] + src22[191] + src22[192] + src22[193] + src22[194] + src22[195] + src22[196] + src22[197] + src22[198] + src22[199] + src22[200] + src22[201] + src22[202] + src22[203] + src22[204] + src22[205] + src22[206] + src22[207] + src22[208] + src22[209] + src22[210] + src22[211] + src22[212] + src22[213] + src22[214] + src22[215] + src22[216] + src22[217] + src22[218] + src22[219] + src22[220] + src22[221] + src22[222] + src22[223] + src22[224] + src22[225] + src22[226] + src22[227] + src22[228] + src22[229] + src22[230] + src22[231] + src22[232] + src22[233] + src22[234] + src22[235] + src22[236] + src22[237] + src22[238] + src22[239] + src22[240] + src22[241] + src22[242] + src22[243] + src22[244] + src22[245] + src22[246] + src22[247] + src22[248] + src22[249] + src22[250] + src22[251] + src22[252] + src22[253] + src22[254] + src22[255] + src22[256] + src22[257] + src22[258] + src22[259] + src22[260] + src22[261] + src22[262] + src22[263] + src22[264] + src22[265] + src22[266] + src22[267] + src22[268] + src22[269] + src22[270] + src22[271] + src22[272] + src22[273] + src22[274] + src22[275] + src22[276] + src22[277] + src22[278] + src22[279] + src22[280] + src22[281] + src22[282] + src22[283] + src22[284] + src22[285] + src22[286] + src22[287] + src22[288] + src22[289] + src22[290] + src22[291] + src22[292] + src22[293] + src22[294] + src22[295] + src22[296] + src22[297] + src22[298] + src22[299] + src22[300] + src22[301] + src22[302] + src22[303] + src22[304] + src22[305] + src22[306] + src22[307] + src22[308] + src22[309] + src22[310] + src22[311] + src22[312] + src22[313] + src22[314] + src22[315] + src22[316] + src22[317] + src22[318] + src22[319] + src22[320] + src22[321] + src22[322] + src22[323] + src22[324] + src22[325] + src22[326] + src22[327] + src22[328] + src22[329] + src22[330] + src22[331] + src22[332] + src22[333] + src22[334] + src22[335] + src22[336] + src22[337] + src22[338] + src22[339] + src22[340] + src22[341] + src22[342] + src22[343] + src22[344] + src22[345] + src22[346] + src22[347] + src22[348] + src22[349] + src22[350] + src22[351] + src22[352] + src22[353] + src22[354] + src22[355] + src22[356] + src22[357] + src22[358] + src22[359] + src22[360] + src22[361] + src22[362] + src22[363] + src22[364] + src22[365] + src22[366] + src22[367] + src22[368] + src22[369] + src22[370] + src22[371] + src22[372] + src22[373] + src22[374] + src22[375] + src22[376] + src22[377] + src22[378] + src22[379] + src22[380] + src22[381] + src22[382] + src22[383] + src22[384] + src22[385] + src22[386] + src22[387] + src22[388] + src22[389] + src22[390] + src22[391] + src22[392] + src22[393] + src22[394] + src22[395] + src22[396] + src22[397] + src22[398] + src22[399] + src22[400] + src22[401] + src22[402] + src22[403] + src22[404] + src22[405] + src22[406] + src22[407] + src22[408] + src22[409] + src22[410] + src22[411] + src22[412] + src22[413] + src22[414] + src22[415] + src22[416] + src22[417] + src22[418] + src22[419] + src22[420] + src22[421] + src22[422] + src22[423] + src22[424] + src22[425] + src22[426] + src22[427] + src22[428] + src22[429] + src22[430] + src22[431] + src22[432] + src22[433] + src22[434] + src22[435] + src22[436] + src22[437] + src22[438] + src22[439] + src22[440] + src22[441] + src22[442] + src22[443] + src22[444] + src22[445] + src22[446] + src22[447] + src22[448] + src22[449] + src22[450] + src22[451] + src22[452] + src22[453] + src22[454] + src22[455] + src22[456] + src22[457] + src22[458] + src22[459] + src22[460] + src22[461] + src22[462] + src22[463] + src22[464] + src22[465] + src22[466] + src22[467] + src22[468] + src22[469] + src22[470] + src22[471] + src22[472] + src22[473] + src22[474] + src22[475] + src22[476] + src22[477] + src22[478] + src22[479] + src22[480] + src22[481] + src22[482] + src22[483] + src22[484] + src22[485] + src22[486] + src22[487] + src22[488] + src22[489] + src22[490] + src22[491] + src22[492] + src22[493] + src22[494] + src22[495] + src22[496] + src22[497] + src22[498] + src22[499] + src22[500] + src22[501] + src22[502] + src22[503] + src22[504] + src22[505] + src22[506] + src22[507] + src22[508] + src22[509] + src22[510] + src22[511])<<22) + ((src23[0] + src23[1] + src23[2] + src23[3] + src23[4] + src23[5] + src23[6] + src23[7] + src23[8] + src23[9] + src23[10] + src23[11] + src23[12] + src23[13] + src23[14] + src23[15] + src23[16] + src23[17] + src23[18] + src23[19] + src23[20] + src23[21] + src23[22] + src23[23] + src23[24] + src23[25] + src23[26] + src23[27] + src23[28] + src23[29] + src23[30] + src23[31] + src23[32] + src23[33] + src23[34] + src23[35] + src23[36] + src23[37] + src23[38] + src23[39] + src23[40] + src23[41] + src23[42] + src23[43] + src23[44] + src23[45] + src23[46] + src23[47] + src23[48] + src23[49] + src23[50] + src23[51] + src23[52] + src23[53] + src23[54] + src23[55] + src23[56] + src23[57] + src23[58] + src23[59] + src23[60] + src23[61] + src23[62] + src23[63] + src23[64] + src23[65] + src23[66] + src23[67] + src23[68] + src23[69] + src23[70] + src23[71] + src23[72] + src23[73] + src23[74] + src23[75] + src23[76] + src23[77] + src23[78] + src23[79] + src23[80] + src23[81] + src23[82] + src23[83] + src23[84] + src23[85] + src23[86] + src23[87] + src23[88] + src23[89] + src23[90] + src23[91] + src23[92] + src23[93] + src23[94] + src23[95] + src23[96] + src23[97] + src23[98] + src23[99] + src23[100] + src23[101] + src23[102] + src23[103] + src23[104] + src23[105] + src23[106] + src23[107] + src23[108] + src23[109] + src23[110] + src23[111] + src23[112] + src23[113] + src23[114] + src23[115] + src23[116] + src23[117] + src23[118] + src23[119] + src23[120] + src23[121] + src23[122] + src23[123] + src23[124] + src23[125] + src23[126] + src23[127] + src23[128] + src23[129] + src23[130] + src23[131] + src23[132] + src23[133] + src23[134] + src23[135] + src23[136] + src23[137] + src23[138] + src23[139] + src23[140] + src23[141] + src23[142] + src23[143] + src23[144] + src23[145] + src23[146] + src23[147] + src23[148] + src23[149] + src23[150] + src23[151] + src23[152] + src23[153] + src23[154] + src23[155] + src23[156] + src23[157] + src23[158] + src23[159] + src23[160] + src23[161] + src23[162] + src23[163] + src23[164] + src23[165] + src23[166] + src23[167] + src23[168] + src23[169] + src23[170] + src23[171] + src23[172] + src23[173] + src23[174] + src23[175] + src23[176] + src23[177] + src23[178] + src23[179] + src23[180] + src23[181] + src23[182] + src23[183] + src23[184] + src23[185] + src23[186] + src23[187] + src23[188] + src23[189] + src23[190] + src23[191] + src23[192] + src23[193] + src23[194] + src23[195] + src23[196] + src23[197] + src23[198] + src23[199] + src23[200] + src23[201] + src23[202] + src23[203] + src23[204] + src23[205] + src23[206] + src23[207] + src23[208] + src23[209] + src23[210] + src23[211] + src23[212] + src23[213] + src23[214] + src23[215] + src23[216] + src23[217] + src23[218] + src23[219] + src23[220] + src23[221] + src23[222] + src23[223] + src23[224] + src23[225] + src23[226] + src23[227] + src23[228] + src23[229] + src23[230] + src23[231] + src23[232] + src23[233] + src23[234] + src23[235] + src23[236] + src23[237] + src23[238] + src23[239] + src23[240] + src23[241] + src23[242] + src23[243] + src23[244] + src23[245] + src23[246] + src23[247] + src23[248] + src23[249] + src23[250] + src23[251] + src23[252] + src23[253] + src23[254] + src23[255] + src23[256] + src23[257] + src23[258] + src23[259] + src23[260] + src23[261] + src23[262] + src23[263] + src23[264] + src23[265] + src23[266] + src23[267] + src23[268] + src23[269] + src23[270] + src23[271] + src23[272] + src23[273] + src23[274] + src23[275] + src23[276] + src23[277] + src23[278] + src23[279] + src23[280] + src23[281] + src23[282] + src23[283] + src23[284] + src23[285] + src23[286] + src23[287] + src23[288] + src23[289] + src23[290] + src23[291] + src23[292] + src23[293] + src23[294] + src23[295] + src23[296] + src23[297] + src23[298] + src23[299] + src23[300] + src23[301] + src23[302] + src23[303] + src23[304] + src23[305] + src23[306] + src23[307] + src23[308] + src23[309] + src23[310] + src23[311] + src23[312] + src23[313] + src23[314] + src23[315] + src23[316] + src23[317] + src23[318] + src23[319] + src23[320] + src23[321] + src23[322] + src23[323] + src23[324] + src23[325] + src23[326] + src23[327] + src23[328] + src23[329] + src23[330] + src23[331] + src23[332] + src23[333] + src23[334] + src23[335] + src23[336] + src23[337] + src23[338] + src23[339] + src23[340] + src23[341] + src23[342] + src23[343] + src23[344] + src23[345] + src23[346] + src23[347] + src23[348] + src23[349] + src23[350] + src23[351] + src23[352] + src23[353] + src23[354] + src23[355] + src23[356] + src23[357] + src23[358] + src23[359] + src23[360] + src23[361] + src23[362] + src23[363] + src23[364] + src23[365] + src23[366] + src23[367] + src23[368] + src23[369] + src23[370] + src23[371] + src23[372] + src23[373] + src23[374] + src23[375] + src23[376] + src23[377] + src23[378] + src23[379] + src23[380] + src23[381] + src23[382] + src23[383] + src23[384] + src23[385] + src23[386] + src23[387] + src23[388] + src23[389] + src23[390] + src23[391] + src23[392] + src23[393] + src23[394] + src23[395] + src23[396] + src23[397] + src23[398] + src23[399] + src23[400] + src23[401] + src23[402] + src23[403] + src23[404] + src23[405] + src23[406] + src23[407] + src23[408] + src23[409] + src23[410] + src23[411] + src23[412] + src23[413] + src23[414] + src23[415] + src23[416] + src23[417] + src23[418] + src23[419] + src23[420] + src23[421] + src23[422] + src23[423] + src23[424] + src23[425] + src23[426] + src23[427] + src23[428] + src23[429] + src23[430] + src23[431] + src23[432] + src23[433] + src23[434] + src23[435] + src23[436] + src23[437] + src23[438] + src23[439] + src23[440] + src23[441] + src23[442] + src23[443] + src23[444] + src23[445] + src23[446] + src23[447] + src23[448] + src23[449] + src23[450] + src23[451] + src23[452] + src23[453] + src23[454] + src23[455] + src23[456] + src23[457] + src23[458] + src23[459] + src23[460] + src23[461] + src23[462] + src23[463] + src23[464] + src23[465] + src23[466] + src23[467] + src23[468] + src23[469] + src23[470] + src23[471] + src23[472] + src23[473] + src23[474] + src23[475] + src23[476] + src23[477] + src23[478] + src23[479] + src23[480] + src23[481] + src23[482] + src23[483] + src23[484] + src23[485] + src23[486] + src23[487] + src23[488] + src23[489] + src23[490] + src23[491] + src23[492] + src23[493] + src23[494] + src23[495] + src23[496] + src23[497] + src23[498] + src23[499] + src23[500] + src23[501] + src23[502] + src23[503] + src23[504] + src23[505] + src23[506] + src23[507] + src23[508] + src23[509] + src23[510] + src23[511])<<23) + ((src24[0] + src24[1] + src24[2] + src24[3] + src24[4] + src24[5] + src24[6] + src24[7] + src24[8] + src24[9] + src24[10] + src24[11] + src24[12] + src24[13] + src24[14] + src24[15] + src24[16] + src24[17] + src24[18] + src24[19] + src24[20] + src24[21] + src24[22] + src24[23] + src24[24] + src24[25] + src24[26] + src24[27] + src24[28] + src24[29] + src24[30] + src24[31] + src24[32] + src24[33] + src24[34] + src24[35] + src24[36] + src24[37] + src24[38] + src24[39] + src24[40] + src24[41] + src24[42] + src24[43] + src24[44] + src24[45] + src24[46] + src24[47] + src24[48] + src24[49] + src24[50] + src24[51] + src24[52] + src24[53] + src24[54] + src24[55] + src24[56] + src24[57] + src24[58] + src24[59] + src24[60] + src24[61] + src24[62] + src24[63] + src24[64] + src24[65] + src24[66] + src24[67] + src24[68] + src24[69] + src24[70] + src24[71] + src24[72] + src24[73] + src24[74] + src24[75] + src24[76] + src24[77] + src24[78] + src24[79] + src24[80] + src24[81] + src24[82] + src24[83] + src24[84] + src24[85] + src24[86] + src24[87] + src24[88] + src24[89] + src24[90] + src24[91] + src24[92] + src24[93] + src24[94] + src24[95] + src24[96] + src24[97] + src24[98] + src24[99] + src24[100] + src24[101] + src24[102] + src24[103] + src24[104] + src24[105] + src24[106] + src24[107] + src24[108] + src24[109] + src24[110] + src24[111] + src24[112] + src24[113] + src24[114] + src24[115] + src24[116] + src24[117] + src24[118] + src24[119] + src24[120] + src24[121] + src24[122] + src24[123] + src24[124] + src24[125] + src24[126] + src24[127] + src24[128] + src24[129] + src24[130] + src24[131] + src24[132] + src24[133] + src24[134] + src24[135] + src24[136] + src24[137] + src24[138] + src24[139] + src24[140] + src24[141] + src24[142] + src24[143] + src24[144] + src24[145] + src24[146] + src24[147] + src24[148] + src24[149] + src24[150] + src24[151] + src24[152] + src24[153] + src24[154] + src24[155] + src24[156] + src24[157] + src24[158] + src24[159] + src24[160] + src24[161] + src24[162] + src24[163] + src24[164] + src24[165] + src24[166] + src24[167] + src24[168] + src24[169] + src24[170] + src24[171] + src24[172] + src24[173] + src24[174] + src24[175] + src24[176] + src24[177] + src24[178] + src24[179] + src24[180] + src24[181] + src24[182] + src24[183] + src24[184] + src24[185] + src24[186] + src24[187] + src24[188] + src24[189] + src24[190] + src24[191] + src24[192] + src24[193] + src24[194] + src24[195] + src24[196] + src24[197] + src24[198] + src24[199] + src24[200] + src24[201] + src24[202] + src24[203] + src24[204] + src24[205] + src24[206] + src24[207] + src24[208] + src24[209] + src24[210] + src24[211] + src24[212] + src24[213] + src24[214] + src24[215] + src24[216] + src24[217] + src24[218] + src24[219] + src24[220] + src24[221] + src24[222] + src24[223] + src24[224] + src24[225] + src24[226] + src24[227] + src24[228] + src24[229] + src24[230] + src24[231] + src24[232] + src24[233] + src24[234] + src24[235] + src24[236] + src24[237] + src24[238] + src24[239] + src24[240] + src24[241] + src24[242] + src24[243] + src24[244] + src24[245] + src24[246] + src24[247] + src24[248] + src24[249] + src24[250] + src24[251] + src24[252] + src24[253] + src24[254] + src24[255] + src24[256] + src24[257] + src24[258] + src24[259] + src24[260] + src24[261] + src24[262] + src24[263] + src24[264] + src24[265] + src24[266] + src24[267] + src24[268] + src24[269] + src24[270] + src24[271] + src24[272] + src24[273] + src24[274] + src24[275] + src24[276] + src24[277] + src24[278] + src24[279] + src24[280] + src24[281] + src24[282] + src24[283] + src24[284] + src24[285] + src24[286] + src24[287] + src24[288] + src24[289] + src24[290] + src24[291] + src24[292] + src24[293] + src24[294] + src24[295] + src24[296] + src24[297] + src24[298] + src24[299] + src24[300] + src24[301] + src24[302] + src24[303] + src24[304] + src24[305] + src24[306] + src24[307] + src24[308] + src24[309] + src24[310] + src24[311] + src24[312] + src24[313] + src24[314] + src24[315] + src24[316] + src24[317] + src24[318] + src24[319] + src24[320] + src24[321] + src24[322] + src24[323] + src24[324] + src24[325] + src24[326] + src24[327] + src24[328] + src24[329] + src24[330] + src24[331] + src24[332] + src24[333] + src24[334] + src24[335] + src24[336] + src24[337] + src24[338] + src24[339] + src24[340] + src24[341] + src24[342] + src24[343] + src24[344] + src24[345] + src24[346] + src24[347] + src24[348] + src24[349] + src24[350] + src24[351] + src24[352] + src24[353] + src24[354] + src24[355] + src24[356] + src24[357] + src24[358] + src24[359] + src24[360] + src24[361] + src24[362] + src24[363] + src24[364] + src24[365] + src24[366] + src24[367] + src24[368] + src24[369] + src24[370] + src24[371] + src24[372] + src24[373] + src24[374] + src24[375] + src24[376] + src24[377] + src24[378] + src24[379] + src24[380] + src24[381] + src24[382] + src24[383] + src24[384] + src24[385] + src24[386] + src24[387] + src24[388] + src24[389] + src24[390] + src24[391] + src24[392] + src24[393] + src24[394] + src24[395] + src24[396] + src24[397] + src24[398] + src24[399] + src24[400] + src24[401] + src24[402] + src24[403] + src24[404] + src24[405] + src24[406] + src24[407] + src24[408] + src24[409] + src24[410] + src24[411] + src24[412] + src24[413] + src24[414] + src24[415] + src24[416] + src24[417] + src24[418] + src24[419] + src24[420] + src24[421] + src24[422] + src24[423] + src24[424] + src24[425] + src24[426] + src24[427] + src24[428] + src24[429] + src24[430] + src24[431] + src24[432] + src24[433] + src24[434] + src24[435] + src24[436] + src24[437] + src24[438] + src24[439] + src24[440] + src24[441] + src24[442] + src24[443] + src24[444] + src24[445] + src24[446] + src24[447] + src24[448] + src24[449] + src24[450] + src24[451] + src24[452] + src24[453] + src24[454] + src24[455] + src24[456] + src24[457] + src24[458] + src24[459] + src24[460] + src24[461] + src24[462] + src24[463] + src24[464] + src24[465] + src24[466] + src24[467] + src24[468] + src24[469] + src24[470] + src24[471] + src24[472] + src24[473] + src24[474] + src24[475] + src24[476] + src24[477] + src24[478] + src24[479] + src24[480] + src24[481] + src24[482] + src24[483] + src24[484] + src24[485] + src24[486] + src24[487] + src24[488] + src24[489] + src24[490] + src24[491] + src24[492] + src24[493] + src24[494] + src24[495] + src24[496] + src24[497] + src24[498] + src24[499] + src24[500] + src24[501] + src24[502] + src24[503] + src24[504] + src24[505] + src24[506] + src24[507] + src24[508] + src24[509] + src24[510] + src24[511])<<24) + ((src25[0] + src25[1] + src25[2] + src25[3] + src25[4] + src25[5] + src25[6] + src25[7] + src25[8] + src25[9] + src25[10] + src25[11] + src25[12] + src25[13] + src25[14] + src25[15] + src25[16] + src25[17] + src25[18] + src25[19] + src25[20] + src25[21] + src25[22] + src25[23] + src25[24] + src25[25] + src25[26] + src25[27] + src25[28] + src25[29] + src25[30] + src25[31] + src25[32] + src25[33] + src25[34] + src25[35] + src25[36] + src25[37] + src25[38] + src25[39] + src25[40] + src25[41] + src25[42] + src25[43] + src25[44] + src25[45] + src25[46] + src25[47] + src25[48] + src25[49] + src25[50] + src25[51] + src25[52] + src25[53] + src25[54] + src25[55] + src25[56] + src25[57] + src25[58] + src25[59] + src25[60] + src25[61] + src25[62] + src25[63] + src25[64] + src25[65] + src25[66] + src25[67] + src25[68] + src25[69] + src25[70] + src25[71] + src25[72] + src25[73] + src25[74] + src25[75] + src25[76] + src25[77] + src25[78] + src25[79] + src25[80] + src25[81] + src25[82] + src25[83] + src25[84] + src25[85] + src25[86] + src25[87] + src25[88] + src25[89] + src25[90] + src25[91] + src25[92] + src25[93] + src25[94] + src25[95] + src25[96] + src25[97] + src25[98] + src25[99] + src25[100] + src25[101] + src25[102] + src25[103] + src25[104] + src25[105] + src25[106] + src25[107] + src25[108] + src25[109] + src25[110] + src25[111] + src25[112] + src25[113] + src25[114] + src25[115] + src25[116] + src25[117] + src25[118] + src25[119] + src25[120] + src25[121] + src25[122] + src25[123] + src25[124] + src25[125] + src25[126] + src25[127] + src25[128] + src25[129] + src25[130] + src25[131] + src25[132] + src25[133] + src25[134] + src25[135] + src25[136] + src25[137] + src25[138] + src25[139] + src25[140] + src25[141] + src25[142] + src25[143] + src25[144] + src25[145] + src25[146] + src25[147] + src25[148] + src25[149] + src25[150] + src25[151] + src25[152] + src25[153] + src25[154] + src25[155] + src25[156] + src25[157] + src25[158] + src25[159] + src25[160] + src25[161] + src25[162] + src25[163] + src25[164] + src25[165] + src25[166] + src25[167] + src25[168] + src25[169] + src25[170] + src25[171] + src25[172] + src25[173] + src25[174] + src25[175] + src25[176] + src25[177] + src25[178] + src25[179] + src25[180] + src25[181] + src25[182] + src25[183] + src25[184] + src25[185] + src25[186] + src25[187] + src25[188] + src25[189] + src25[190] + src25[191] + src25[192] + src25[193] + src25[194] + src25[195] + src25[196] + src25[197] + src25[198] + src25[199] + src25[200] + src25[201] + src25[202] + src25[203] + src25[204] + src25[205] + src25[206] + src25[207] + src25[208] + src25[209] + src25[210] + src25[211] + src25[212] + src25[213] + src25[214] + src25[215] + src25[216] + src25[217] + src25[218] + src25[219] + src25[220] + src25[221] + src25[222] + src25[223] + src25[224] + src25[225] + src25[226] + src25[227] + src25[228] + src25[229] + src25[230] + src25[231] + src25[232] + src25[233] + src25[234] + src25[235] + src25[236] + src25[237] + src25[238] + src25[239] + src25[240] + src25[241] + src25[242] + src25[243] + src25[244] + src25[245] + src25[246] + src25[247] + src25[248] + src25[249] + src25[250] + src25[251] + src25[252] + src25[253] + src25[254] + src25[255] + src25[256] + src25[257] + src25[258] + src25[259] + src25[260] + src25[261] + src25[262] + src25[263] + src25[264] + src25[265] + src25[266] + src25[267] + src25[268] + src25[269] + src25[270] + src25[271] + src25[272] + src25[273] + src25[274] + src25[275] + src25[276] + src25[277] + src25[278] + src25[279] + src25[280] + src25[281] + src25[282] + src25[283] + src25[284] + src25[285] + src25[286] + src25[287] + src25[288] + src25[289] + src25[290] + src25[291] + src25[292] + src25[293] + src25[294] + src25[295] + src25[296] + src25[297] + src25[298] + src25[299] + src25[300] + src25[301] + src25[302] + src25[303] + src25[304] + src25[305] + src25[306] + src25[307] + src25[308] + src25[309] + src25[310] + src25[311] + src25[312] + src25[313] + src25[314] + src25[315] + src25[316] + src25[317] + src25[318] + src25[319] + src25[320] + src25[321] + src25[322] + src25[323] + src25[324] + src25[325] + src25[326] + src25[327] + src25[328] + src25[329] + src25[330] + src25[331] + src25[332] + src25[333] + src25[334] + src25[335] + src25[336] + src25[337] + src25[338] + src25[339] + src25[340] + src25[341] + src25[342] + src25[343] + src25[344] + src25[345] + src25[346] + src25[347] + src25[348] + src25[349] + src25[350] + src25[351] + src25[352] + src25[353] + src25[354] + src25[355] + src25[356] + src25[357] + src25[358] + src25[359] + src25[360] + src25[361] + src25[362] + src25[363] + src25[364] + src25[365] + src25[366] + src25[367] + src25[368] + src25[369] + src25[370] + src25[371] + src25[372] + src25[373] + src25[374] + src25[375] + src25[376] + src25[377] + src25[378] + src25[379] + src25[380] + src25[381] + src25[382] + src25[383] + src25[384] + src25[385] + src25[386] + src25[387] + src25[388] + src25[389] + src25[390] + src25[391] + src25[392] + src25[393] + src25[394] + src25[395] + src25[396] + src25[397] + src25[398] + src25[399] + src25[400] + src25[401] + src25[402] + src25[403] + src25[404] + src25[405] + src25[406] + src25[407] + src25[408] + src25[409] + src25[410] + src25[411] + src25[412] + src25[413] + src25[414] + src25[415] + src25[416] + src25[417] + src25[418] + src25[419] + src25[420] + src25[421] + src25[422] + src25[423] + src25[424] + src25[425] + src25[426] + src25[427] + src25[428] + src25[429] + src25[430] + src25[431] + src25[432] + src25[433] + src25[434] + src25[435] + src25[436] + src25[437] + src25[438] + src25[439] + src25[440] + src25[441] + src25[442] + src25[443] + src25[444] + src25[445] + src25[446] + src25[447] + src25[448] + src25[449] + src25[450] + src25[451] + src25[452] + src25[453] + src25[454] + src25[455] + src25[456] + src25[457] + src25[458] + src25[459] + src25[460] + src25[461] + src25[462] + src25[463] + src25[464] + src25[465] + src25[466] + src25[467] + src25[468] + src25[469] + src25[470] + src25[471] + src25[472] + src25[473] + src25[474] + src25[475] + src25[476] + src25[477] + src25[478] + src25[479] + src25[480] + src25[481] + src25[482] + src25[483] + src25[484] + src25[485] + src25[486] + src25[487] + src25[488] + src25[489] + src25[490] + src25[491] + src25[492] + src25[493] + src25[494] + src25[495] + src25[496] + src25[497] + src25[498] + src25[499] + src25[500] + src25[501] + src25[502] + src25[503] + src25[504] + src25[505] + src25[506] + src25[507] + src25[508] + src25[509] + src25[510] + src25[511])<<25) + ((src26[0] + src26[1] + src26[2] + src26[3] + src26[4] + src26[5] + src26[6] + src26[7] + src26[8] + src26[9] + src26[10] + src26[11] + src26[12] + src26[13] + src26[14] + src26[15] + src26[16] + src26[17] + src26[18] + src26[19] + src26[20] + src26[21] + src26[22] + src26[23] + src26[24] + src26[25] + src26[26] + src26[27] + src26[28] + src26[29] + src26[30] + src26[31] + src26[32] + src26[33] + src26[34] + src26[35] + src26[36] + src26[37] + src26[38] + src26[39] + src26[40] + src26[41] + src26[42] + src26[43] + src26[44] + src26[45] + src26[46] + src26[47] + src26[48] + src26[49] + src26[50] + src26[51] + src26[52] + src26[53] + src26[54] + src26[55] + src26[56] + src26[57] + src26[58] + src26[59] + src26[60] + src26[61] + src26[62] + src26[63] + src26[64] + src26[65] + src26[66] + src26[67] + src26[68] + src26[69] + src26[70] + src26[71] + src26[72] + src26[73] + src26[74] + src26[75] + src26[76] + src26[77] + src26[78] + src26[79] + src26[80] + src26[81] + src26[82] + src26[83] + src26[84] + src26[85] + src26[86] + src26[87] + src26[88] + src26[89] + src26[90] + src26[91] + src26[92] + src26[93] + src26[94] + src26[95] + src26[96] + src26[97] + src26[98] + src26[99] + src26[100] + src26[101] + src26[102] + src26[103] + src26[104] + src26[105] + src26[106] + src26[107] + src26[108] + src26[109] + src26[110] + src26[111] + src26[112] + src26[113] + src26[114] + src26[115] + src26[116] + src26[117] + src26[118] + src26[119] + src26[120] + src26[121] + src26[122] + src26[123] + src26[124] + src26[125] + src26[126] + src26[127] + src26[128] + src26[129] + src26[130] + src26[131] + src26[132] + src26[133] + src26[134] + src26[135] + src26[136] + src26[137] + src26[138] + src26[139] + src26[140] + src26[141] + src26[142] + src26[143] + src26[144] + src26[145] + src26[146] + src26[147] + src26[148] + src26[149] + src26[150] + src26[151] + src26[152] + src26[153] + src26[154] + src26[155] + src26[156] + src26[157] + src26[158] + src26[159] + src26[160] + src26[161] + src26[162] + src26[163] + src26[164] + src26[165] + src26[166] + src26[167] + src26[168] + src26[169] + src26[170] + src26[171] + src26[172] + src26[173] + src26[174] + src26[175] + src26[176] + src26[177] + src26[178] + src26[179] + src26[180] + src26[181] + src26[182] + src26[183] + src26[184] + src26[185] + src26[186] + src26[187] + src26[188] + src26[189] + src26[190] + src26[191] + src26[192] + src26[193] + src26[194] + src26[195] + src26[196] + src26[197] + src26[198] + src26[199] + src26[200] + src26[201] + src26[202] + src26[203] + src26[204] + src26[205] + src26[206] + src26[207] + src26[208] + src26[209] + src26[210] + src26[211] + src26[212] + src26[213] + src26[214] + src26[215] + src26[216] + src26[217] + src26[218] + src26[219] + src26[220] + src26[221] + src26[222] + src26[223] + src26[224] + src26[225] + src26[226] + src26[227] + src26[228] + src26[229] + src26[230] + src26[231] + src26[232] + src26[233] + src26[234] + src26[235] + src26[236] + src26[237] + src26[238] + src26[239] + src26[240] + src26[241] + src26[242] + src26[243] + src26[244] + src26[245] + src26[246] + src26[247] + src26[248] + src26[249] + src26[250] + src26[251] + src26[252] + src26[253] + src26[254] + src26[255] + src26[256] + src26[257] + src26[258] + src26[259] + src26[260] + src26[261] + src26[262] + src26[263] + src26[264] + src26[265] + src26[266] + src26[267] + src26[268] + src26[269] + src26[270] + src26[271] + src26[272] + src26[273] + src26[274] + src26[275] + src26[276] + src26[277] + src26[278] + src26[279] + src26[280] + src26[281] + src26[282] + src26[283] + src26[284] + src26[285] + src26[286] + src26[287] + src26[288] + src26[289] + src26[290] + src26[291] + src26[292] + src26[293] + src26[294] + src26[295] + src26[296] + src26[297] + src26[298] + src26[299] + src26[300] + src26[301] + src26[302] + src26[303] + src26[304] + src26[305] + src26[306] + src26[307] + src26[308] + src26[309] + src26[310] + src26[311] + src26[312] + src26[313] + src26[314] + src26[315] + src26[316] + src26[317] + src26[318] + src26[319] + src26[320] + src26[321] + src26[322] + src26[323] + src26[324] + src26[325] + src26[326] + src26[327] + src26[328] + src26[329] + src26[330] + src26[331] + src26[332] + src26[333] + src26[334] + src26[335] + src26[336] + src26[337] + src26[338] + src26[339] + src26[340] + src26[341] + src26[342] + src26[343] + src26[344] + src26[345] + src26[346] + src26[347] + src26[348] + src26[349] + src26[350] + src26[351] + src26[352] + src26[353] + src26[354] + src26[355] + src26[356] + src26[357] + src26[358] + src26[359] + src26[360] + src26[361] + src26[362] + src26[363] + src26[364] + src26[365] + src26[366] + src26[367] + src26[368] + src26[369] + src26[370] + src26[371] + src26[372] + src26[373] + src26[374] + src26[375] + src26[376] + src26[377] + src26[378] + src26[379] + src26[380] + src26[381] + src26[382] + src26[383] + src26[384] + src26[385] + src26[386] + src26[387] + src26[388] + src26[389] + src26[390] + src26[391] + src26[392] + src26[393] + src26[394] + src26[395] + src26[396] + src26[397] + src26[398] + src26[399] + src26[400] + src26[401] + src26[402] + src26[403] + src26[404] + src26[405] + src26[406] + src26[407] + src26[408] + src26[409] + src26[410] + src26[411] + src26[412] + src26[413] + src26[414] + src26[415] + src26[416] + src26[417] + src26[418] + src26[419] + src26[420] + src26[421] + src26[422] + src26[423] + src26[424] + src26[425] + src26[426] + src26[427] + src26[428] + src26[429] + src26[430] + src26[431] + src26[432] + src26[433] + src26[434] + src26[435] + src26[436] + src26[437] + src26[438] + src26[439] + src26[440] + src26[441] + src26[442] + src26[443] + src26[444] + src26[445] + src26[446] + src26[447] + src26[448] + src26[449] + src26[450] + src26[451] + src26[452] + src26[453] + src26[454] + src26[455] + src26[456] + src26[457] + src26[458] + src26[459] + src26[460] + src26[461] + src26[462] + src26[463] + src26[464] + src26[465] + src26[466] + src26[467] + src26[468] + src26[469] + src26[470] + src26[471] + src26[472] + src26[473] + src26[474] + src26[475] + src26[476] + src26[477] + src26[478] + src26[479] + src26[480] + src26[481] + src26[482] + src26[483] + src26[484] + src26[485] + src26[486] + src26[487] + src26[488] + src26[489] + src26[490] + src26[491] + src26[492] + src26[493] + src26[494] + src26[495] + src26[496] + src26[497] + src26[498] + src26[499] + src26[500] + src26[501] + src26[502] + src26[503] + src26[504] + src26[505] + src26[506] + src26[507] + src26[508] + src26[509] + src26[510] + src26[511])<<26) + ((src27[0] + src27[1] + src27[2] + src27[3] + src27[4] + src27[5] + src27[6] + src27[7] + src27[8] + src27[9] + src27[10] + src27[11] + src27[12] + src27[13] + src27[14] + src27[15] + src27[16] + src27[17] + src27[18] + src27[19] + src27[20] + src27[21] + src27[22] + src27[23] + src27[24] + src27[25] + src27[26] + src27[27] + src27[28] + src27[29] + src27[30] + src27[31] + src27[32] + src27[33] + src27[34] + src27[35] + src27[36] + src27[37] + src27[38] + src27[39] + src27[40] + src27[41] + src27[42] + src27[43] + src27[44] + src27[45] + src27[46] + src27[47] + src27[48] + src27[49] + src27[50] + src27[51] + src27[52] + src27[53] + src27[54] + src27[55] + src27[56] + src27[57] + src27[58] + src27[59] + src27[60] + src27[61] + src27[62] + src27[63] + src27[64] + src27[65] + src27[66] + src27[67] + src27[68] + src27[69] + src27[70] + src27[71] + src27[72] + src27[73] + src27[74] + src27[75] + src27[76] + src27[77] + src27[78] + src27[79] + src27[80] + src27[81] + src27[82] + src27[83] + src27[84] + src27[85] + src27[86] + src27[87] + src27[88] + src27[89] + src27[90] + src27[91] + src27[92] + src27[93] + src27[94] + src27[95] + src27[96] + src27[97] + src27[98] + src27[99] + src27[100] + src27[101] + src27[102] + src27[103] + src27[104] + src27[105] + src27[106] + src27[107] + src27[108] + src27[109] + src27[110] + src27[111] + src27[112] + src27[113] + src27[114] + src27[115] + src27[116] + src27[117] + src27[118] + src27[119] + src27[120] + src27[121] + src27[122] + src27[123] + src27[124] + src27[125] + src27[126] + src27[127] + src27[128] + src27[129] + src27[130] + src27[131] + src27[132] + src27[133] + src27[134] + src27[135] + src27[136] + src27[137] + src27[138] + src27[139] + src27[140] + src27[141] + src27[142] + src27[143] + src27[144] + src27[145] + src27[146] + src27[147] + src27[148] + src27[149] + src27[150] + src27[151] + src27[152] + src27[153] + src27[154] + src27[155] + src27[156] + src27[157] + src27[158] + src27[159] + src27[160] + src27[161] + src27[162] + src27[163] + src27[164] + src27[165] + src27[166] + src27[167] + src27[168] + src27[169] + src27[170] + src27[171] + src27[172] + src27[173] + src27[174] + src27[175] + src27[176] + src27[177] + src27[178] + src27[179] + src27[180] + src27[181] + src27[182] + src27[183] + src27[184] + src27[185] + src27[186] + src27[187] + src27[188] + src27[189] + src27[190] + src27[191] + src27[192] + src27[193] + src27[194] + src27[195] + src27[196] + src27[197] + src27[198] + src27[199] + src27[200] + src27[201] + src27[202] + src27[203] + src27[204] + src27[205] + src27[206] + src27[207] + src27[208] + src27[209] + src27[210] + src27[211] + src27[212] + src27[213] + src27[214] + src27[215] + src27[216] + src27[217] + src27[218] + src27[219] + src27[220] + src27[221] + src27[222] + src27[223] + src27[224] + src27[225] + src27[226] + src27[227] + src27[228] + src27[229] + src27[230] + src27[231] + src27[232] + src27[233] + src27[234] + src27[235] + src27[236] + src27[237] + src27[238] + src27[239] + src27[240] + src27[241] + src27[242] + src27[243] + src27[244] + src27[245] + src27[246] + src27[247] + src27[248] + src27[249] + src27[250] + src27[251] + src27[252] + src27[253] + src27[254] + src27[255] + src27[256] + src27[257] + src27[258] + src27[259] + src27[260] + src27[261] + src27[262] + src27[263] + src27[264] + src27[265] + src27[266] + src27[267] + src27[268] + src27[269] + src27[270] + src27[271] + src27[272] + src27[273] + src27[274] + src27[275] + src27[276] + src27[277] + src27[278] + src27[279] + src27[280] + src27[281] + src27[282] + src27[283] + src27[284] + src27[285] + src27[286] + src27[287] + src27[288] + src27[289] + src27[290] + src27[291] + src27[292] + src27[293] + src27[294] + src27[295] + src27[296] + src27[297] + src27[298] + src27[299] + src27[300] + src27[301] + src27[302] + src27[303] + src27[304] + src27[305] + src27[306] + src27[307] + src27[308] + src27[309] + src27[310] + src27[311] + src27[312] + src27[313] + src27[314] + src27[315] + src27[316] + src27[317] + src27[318] + src27[319] + src27[320] + src27[321] + src27[322] + src27[323] + src27[324] + src27[325] + src27[326] + src27[327] + src27[328] + src27[329] + src27[330] + src27[331] + src27[332] + src27[333] + src27[334] + src27[335] + src27[336] + src27[337] + src27[338] + src27[339] + src27[340] + src27[341] + src27[342] + src27[343] + src27[344] + src27[345] + src27[346] + src27[347] + src27[348] + src27[349] + src27[350] + src27[351] + src27[352] + src27[353] + src27[354] + src27[355] + src27[356] + src27[357] + src27[358] + src27[359] + src27[360] + src27[361] + src27[362] + src27[363] + src27[364] + src27[365] + src27[366] + src27[367] + src27[368] + src27[369] + src27[370] + src27[371] + src27[372] + src27[373] + src27[374] + src27[375] + src27[376] + src27[377] + src27[378] + src27[379] + src27[380] + src27[381] + src27[382] + src27[383] + src27[384] + src27[385] + src27[386] + src27[387] + src27[388] + src27[389] + src27[390] + src27[391] + src27[392] + src27[393] + src27[394] + src27[395] + src27[396] + src27[397] + src27[398] + src27[399] + src27[400] + src27[401] + src27[402] + src27[403] + src27[404] + src27[405] + src27[406] + src27[407] + src27[408] + src27[409] + src27[410] + src27[411] + src27[412] + src27[413] + src27[414] + src27[415] + src27[416] + src27[417] + src27[418] + src27[419] + src27[420] + src27[421] + src27[422] + src27[423] + src27[424] + src27[425] + src27[426] + src27[427] + src27[428] + src27[429] + src27[430] + src27[431] + src27[432] + src27[433] + src27[434] + src27[435] + src27[436] + src27[437] + src27[438] + src27[439] + src27[440] + src27[441] + src27[442] + src27[443] + src27[444] + src27[445] + src27[446] + src27[447] + src27[448] + src27[449] + src27[450] + src27[451] + src27[452] + src27[453] + src27[454] + src27[455] + src27[456] + src27[457] + src27[458] + src27[459] + src27[460] + src27[461] + src27[462] + src27[463] + src27[464] + src27[465] + src27[466] + src27[467] + src27[468] + src27[469] + src27[470] + src27[471] + src27[472] + src27[473] + src27[474] + src27[475] + src27[476] + src27[477] + src27[478] + src27[479] + src27[480] + src27[481] + src27[482] + src27[483] + src27[484] + src27[485] + src27[486] + src27[487] + src27[488] + src27[489] + src27[490] + src27[491] + src27[492] + src27[493] + src27[494] + src27[495] + src27[496] + src27[497] + src27[498] + src27[499] + src27[500] + src27[501] + src27[502] + src27[503] + src27[504] + src27[505] + src27[506] + src27[507] + src27[508] + src27[509] + src27[510] + src27[511])<<27) + ((src28[0] + src28[1] + src28[2] + src28[3] + src28[4] + src28[5] + src28[6] + src28[7] + src28[8] + src28[9] + src28[10] + src28[11] + src28[12] + src28[13] + src28[14] + src28[15] + src28[16] + src28[17] + src28[18] + src28[19] + src28[20] + src28[21] + src28[22] + src28[23] + src28[24] + src28[25] + src28[26] + src28[27] + src28[28] + src28[29] + src28[30] + src28[31] + src28[32] + src28[33] + src28[34] + src28[35] + src28[36] + src28[37] + src28[38] + src28[39] + src28[40] + src28[41] + src28[42] + src28[43] + src28[44] + src28[45] + src28[46] + src28[47] + src28[48] + src28[49] + src28[50] + src28[51] + src28[52] + src28[53] + src28[54] + src28[55] + src28[56] + src28[57] + src28[58] + src28[59] + src28[60] + src28[61] + src28[62] + src28[63] + src28[64] + src28[65] + src28[66] + src28[67] + src28[68] + src28[69] + src28[70] + src28[71] + src28[72] + src28[73] + src28[74] + src28[75] + src28[76] + src28[77] + src28[78] + src28[79] + src28[80] + src28[81] + src28[82] + src28[83] + src28[84] + src28[85] + src28[86] + src28[87] + src28[88] + src28[89] + src28[90] + src28[91] + src28[92] + src28[93] + src28[94] + src28[95] + src28[96] + src28[97] + src28[98] + src28[99] + src28[100] + src28[101] + src28[102] + src28[103] + src28[104] + src28[105] + src28[106] + src28[107] + src28[108] + src28[109] + src28[110] + src28[111] + src28[112] + src28[113] + src28[114] + src28[115] + src28[116] + src28[117] + src28[118] + src28[119] + src28[120] + src28[121] + src28[122] + src28[123] + src28[124] + src28[125] + src28[126] + src28[127] + src28[128] + src28[129] + src28[130] + src28[131] + src28[132] + src28[133] + src28[134] + src28[135] + src28[136] + src28[137] + src28[138] + src28[139] + src28[140] + src28[141] + src28[142] + src28[143] + src28[144] + src28[145] + src28[146] + src28[147] + src28[148] + src28[149] + src28[150] + src28[151] + src28[152] + src28[153] + src28[154] + src28[155] + src28[156] + src28[157] + src28[158] + src28[159] + src28[160] + src28[161] + src28[162] + src28[163] + src28[164] + src28[165] + src28[166] + src28[167] + src28[168] + src28[169] + src28[170] + src28[171] + src28[172] + src28[173] + src28[174] + src28[175] + src28[176] + src28[177] + src28[178] + src28[179] + src28[180] + src28[181] + src28[182] + src28[183] + src28[184] + src28[185] + src28[186] + src28[187] + src28[188] + src28[189] + src28[190] + src28[191] + src28[192] + src28[193] + src28[194] + src28[195] + src28[196] + src28[197] + src28[198] + src28[199] + src28[200] + src28[201] + src28[202] + src28[203] + src28[204] + src28[205] + src28[206] + src28[207] + src28[208] + src28[209] + src28[210] + src28[211] + src28[212] + src28[213] + src28[214] + src28[215] + src28[216] + src28[217] + src28[218] + src28[219] + src28[220] + src28[221] + src28[222] + src28[223] + src28[224] + src28[225] + src28[226] + src28[227] + src28[228] + src28[229] + src28[230] + src28[231] + src28[232] + src28[233] + src28[234] + src28[235] + src28[236] + src28[237] + src28[238] + src28[239] + src28[240] + src28[241] + src28[242] + src28[243] + src28[244] + src28[245] + src28[246] + src28[247] + src28[248] + src28[249] + src28[250] + src28[251] + src28[252] + src28[253] + src28[254] + src28[255] + src28[256] + src28[257] + src28[258] + src28[259] + src28[260] + src28[261] + src28[262] + src28[263] + src28[264] + src28[265] + src28[266] + src28[267] + src28[268] + src28[269] + src28[270] + src28[271] + src28[272] + src28[273] + src28[274] + src28[275] + src28[276] + src28[277] + src28[278] + src28[279] + src28[280] + src28[281] + src28[282] + src28[283] + src28[284] + src28[285] + src28[286] + src28[287] + src28[288] + src28[289] + src28[290] + src28[291] + src28[292] + src28[293] + src28[294] + src28[295] + src28[296] + src28[297] + src28[298] + src28[299] + src28[300] + src28[301] + src28[302] + src28[303] + src28[304] + src28[305] + src28[306] + src28[307] + src28[308] + src28[309] + src28[310] + src28[311] + src28[312] + src28[313] + src28[314] + src28[315] + src28[316] + src28[317] + src28[318] + src28[319] + src28[320] + src28[321] + src28[322] + src28[323] + src28[324] + src28[325] + src28[326] + src28[327] + src28[328] + src28[329] + src28[330] + src28[331] + src28[332] + src28[333] + src28[334] + src28[335] + src28[336] + src28[337] + src28[338] + src28[339] + src28[340] + src28[341] + src28[342] + src28[343] + src28[344] + src28[345] + src28[346] + src28[347] + src28[348] + src28[349] + src28[350] + src28[351] + src28[352] + src28[353] + src28[354] + src28[355] + src28[356] + src28[357] + src28[358] + src28[359] + src28[360] + src28[361] + src28[362] + src28[363] + src28[364] + src28[365] + src28[366] + src28[367] + src28[368] + src28[369] + src28[370] + src28[371] + src28[372] + src28[373] + src28[374] + src28[375] + src28[376] + src28[377] + src28[378] + src28[379] + src28[380] + src28[381] + src28[382] + src28[383] + src28[384] + src28[385] + src28[386] + src28[387] + src28[388] + src28[389] + src28[390] + src28[391] + src28[392] + src28[393] + src28[394] + src28[395] + src28[396] + src28[397] + src28[398] + src28[399] + src28[400] + src28[401] + src28[402] + src28[403] + src28[404] + src28[405] + src28[406] + src28[407] + src28[408] + src28[409] + src28[410] + src28[411] + src28[412] + src28[413] + src28[414] + src28[415] + src28[416] + src28[417] + src28[418] + src28[419] + src28[420] + src28[421] + src28[422] + src28[423] + src28[424] + src28[425] + src28[426] + src28[427] + src28[428] + src28[429] + src28[430] + src28[431] + src28[432] + src28[433] + src28[434] + src28[435] + src28[436] + src28[437] + src28[438] + src28[439] + src28[440] + src28[441] + src28[442] + src28[443] + src28[444] + src28[445] + src28[446] + src28[447] + src28[448] + src28[449] + src28[450] + src28[451] + src28[452] + src28[453] + src28[454] + src28[455] + src28[456] + src28[457] + src28[458] + src28[459] + src28[460] + src28[461] + src28[462] + src28[463] + src28[464] + src28[465] + src28[466] + src28[467] + src28[468] + src28[469] + src28[470] + src28[471] + src28[472] + src28[473] + src28[474] + src28[475] + src28[476] + src28[477] + src28[478] + src28[479] + src28[480] + src28[481] + src28[482] + src28[483] + src28[484] + src28[485] + src28[486] + src28[487] + src28[488] + src28[489] + src28[490] + src28[491] + src28[492] + src28[493] + src28[494] + src28[495] + src28[496] + src28[497] + src28[498] + src28[499] + src28[500] + src28[501] + src28[502] + src28[503] + src28[504] + src28[505] + src28[506] + src28[507] + src28[508] + src28[509] + src28[510] + src28[511])<<28) + ((src29[0] + src29[1] + src29[2] + src29[3] + src29[4] + src29[5] + src29[6] + src29[7] + src29[8] + src29[9] + src29[10] + src29[11] + src29[12] + src29[13] + src29[14] + src29[15] + src29[16] + src29[17] + src29[18] + src29[19] + src29[20] + src29[21] + src29[22] + src29[23] + src29[24] + src29[25] + src29[26] + src29[27] + src29[28] + src29[29] + src29[30] + src29[31] + src29[32] + src29[33] + src29[34] + src29[35] + src29[36] + src29[37] + src29[38] + src29[39] + src29[40] + src29[41] + src29[42] + src29[43] + src29[44] + src29[45] + src29[46] + src29[47] + src29[48] + src29[49] + src29[50] + src29[51] + src29[52] + src29[53] + src29[54] + src29[55] + src29[56] + src29[57] + src29[58] + src29[59] + src29[60] + src29[61] + src29[62] + src29[63] + src29[64] + src29[65] + src29[66] + src29[67] + src29[68] + src29[69] + src29[70] + src29[71] + src29[72] + src29[73] + src29[74] + src29[75] + src29[76] + src29[77] + src29[78] + src29[79] + src29[80] + src29[81] + src29[82] + src29[83] + src29[84] + src29[85] + src29[86] + src29[87] + src29[88] + src29[89] + src29[90] + src29[91] + src29[92] + src29[93] + src29[94] + src29[95] + src29[96] + src29[97] + src29[98] + src29[99] + src29[100] + src29[101] + src29[102] + src29[103] + src29[104] + src29[105] + src29[106] + src29[107] + src29[108] + src29[109] + src29[110] + src29[111] + src29[112] + src29[113] + src29[114] + src29[115] + src29[116] + src29[117] + src29[118] + src29[119] + src29[120] + src29[121] + src29[122] + src29[123] + src29[124] + src29[125] + src29[126] + src29[127] + src29[128] + src29[129] + src29[130] + src29[131] + src29[132] + src29[133] + src29[134] + src29[135] + src29[136] + src29[137] + src29[138] + src29[139] + src29[140] + src29[141] + src29[142] + src29[143] + src29[144] + src29[145] + src29[146] + src29[147] + src29[148] + src29[149] + src29[150] + src29[151] + src29[152] + src29[153] + src29[154] + src29[155] + src29[156] + src29[157] + src29[158] + src29[159] + src29[160] + src29[161] + src29[162] + src29[163] + src29[164] + src29[165] + src29[166] + src29[167] + src29[168] + src29[169] + src29[170] + src29[171] + src29[172] + src29[173] + src29[174] + src29[175] + src29[176] + src29[177] + src29[178] + src29[179] + src29[180] + src29[181] + src29[182] + src29[183] + src29[184] + src29[185] + src29[186] + src29[187] + src29[188] + src29[189] + src29[190] + src29[191] + src29[192] + src29[193] + src29[194] + src29[195] + src29[196] + src29[197] + src29[198] + src29[199] + src29[200] + src29[201] + src29[202] + src29[203] + src29[204] + src29[205] + src29[206] + src29[207] + src29[208] + src29[209] + src29[210] + src29[211] + src29[212] + src29[213] + src29[214] + src29[215] + src29[216] + src29[217] + src29[218] + src29[219] + src29[220] + src29[221] + src29[222] + src29[223] + src29[224] + src29[225] + src29[226] + src29[227] + src29[228] + src29[229] + src29[230] + src29[231] + src29[232] + src29[233] + src29[234] + src29[235] + src29[236] + src29[237] + src29[238] + src29[239] + src29[240] + src29[241] + src29[242] + src29[243] + src29[244] + src29[245] + src29[246] + src29[247] + src29[248] + src29[249] + src29[250] + src29[251] + src29[252] + src29[253] + src29[254] + src29[255] + src29[256] + src29[257] + src29[258] + src29[259] + src29[260] + src29[261] + src29[262] + src29[263] + src29[264] + src29[265] + src29[266] + src29[267] + src29[268] + src29[269] + src29[270] + src29[271] + src29[272] + src29[273] + src29[274] + src29[275] + src29[276] + src29[277] + src29[278] + src29[279] + src29[280] + src29[281] + src29[282] + src29[283] + src29[284] + src29[285] + src29[286] + src29[287] + src29[288] + src29[289] + src29[290] + src29[291] + src29[292] + src29[293] + src29[294] + src29[295] + src29[296] + src29[297] + src29[298] + src29[299] + src29[300] + src29[301] + src29[302] + src29[303] + src29[304] + src29[305] + src29[306] + src29[307] + src29[308] + src29[309] + src29[310] + src29[311] + src29[312] + src29[313] + src29[314] + src29[315] + src29[316] + src29[317] + src29[318] + src29[319] + src29[320] + src29[321] + src29[322] + src29[323] + src29[324] + src29[325] + src29[326] + src29[327] + src29[328] + src29[329] + src29[330] + src29[331] + src29[332] + src29[333] + src29[334] + src29[335] + src29[336] + src29[337] + src29[338] + src29[339] + src29[340] + src29[341] + src29[342] + src29[343] + src29[344] + src29[345] + src29[346] + src29[347] + src29[348] + src29[349] + src29[350] + src29[351] + src29[352] + src29[353] + src29[354] + src29[355] + src29[356] + src29[357] + src29[358] + src29[359] + src29[360] + src29[361] + src29[362] + src29[363] + src29[364] + src29[365] + src29[366] + src29[367] + src29[368] + src29[369] + src29[370] + src29[371] + src29[372] + src29[373] + src29[374] + src29[375] + src29[376] + src29[377] + src29[378] + src29[379] + src29[380] + src29[381] + src29[382] + src29[383] + src29[384] + src29[385] + src29[386] + src29[387] + src29[388] + src29[389] + src29[390] + src29[391] + src29[392] + src29[393] + src29[394] + src29[395] + src29[396] + src29[397] + src29[398] + src29[399] + src29[400] + src29[401] + src29[402] + src29[403] + src29[404] + src29[405] + src29[406] + src29[407] + src29[408] + src29[409] + src29[410] + src29[411] + src29[412] + src29[413] + src29[414] + src29[415] + src29[416] + src29[417] + src29[418] + src29[419] + src29[420] + src29[421] + src29[422] + src29[423] + src29[424] + src29[425] + src29[426] + src29[427] + src29[428] + src29[429] + src29[430] + src29[431] + src29[432] + src29[433] + src29[434] + src29[435] + src29[436] + src29[437] + src29[438] + src29[439] + src29[440] + src29[441] + src29[442] + src29[443] + src29[444] + src29[445] + src29[446] + src29[447] + src29[448] + src29[449] + src29[450] + src29[451] + src29[452] + src29[453] + src29[454] + src29[455] + src29[456] + src29[457] + src29[458] + src29[459] + src29[460] + src29[461] + src29[462] + src29[463] + src29[464] + src29[465] + src29[466] + src29[467] + src29[468] + src29[469] + src29[470] + src29[471] + src29[472] + src29[473] + src29[474] + src29[475] + src29[476] + src29[477] + src29[478] + src29[479] + src29[480] + src29[481] + src29[482] + src29[483] + src29[484] + src29[485] + src29[486] + src29[487] + src29[488] + src29[489] + src29[490] + src29[491] + src29[492] + src29[493] + src29[494] + src29[495] + src29[496] + src29[497] + src29[498] + src29[499] + src29[500] + src29[501] + src29[502] + src29[503] + src29[504] + src29[505] + src29[506] + src29[507] + src29[508] + src29[509] + src29[510] + src29[511])<<29) + ((src30[0] + src30[1] + src30[2] + src30[3] + src30[4] + src30[5] + src30[6] + src30[7] + src30[8] + src30[9] + src30[10] + src30[11] + src30[12] + src30[13] + src30[14] + src30[15] + src30[16] + src30[17] + src30[18] + src30[19] + src30[20] + src30[21] + src30[22] + src30[23] + src30[24] + src30[25] + src30[26] + src30[27] + src30[28] + src30[29] + src30[30] + src30[31] + src30[32] + src30[33] + src30[34] + src30[35] + src30[36] + src30[37] + src30[38] + src30[39] + src30[40] + src30[41] + src30[42] + src30[43] + src30[44] + src30[45] + src30[46] + src30[47] + src30[48] + src30[49] + src30[50] + src30[51] + src30[52] + src30[53] + src30[54] + src30[55] + src30[56] + src30[57] + src30[58] + src30[59] + src30[60] + src30[61] + src30[62] + src30[63] + src30[64] + src30[65] + src30[66] + src30[67] + src30[68] + src30[69] + src30[70] + src30[71] + src30[72] + src30[73] + src30[74] + src30[75] + src30[76] + src30[77] + src30[78] + src30[79] + src30[80] + src30[81] + src30[82] + src30[83] + src30[84] + src30[85] + src30[86] + src30[87] + src30[88] + src30[89] + src30[90] + src30[91] + src30[92] + src30[93] + src30[94] + src30[95] + src30[96] + src30[97] + src30[98] + src30[99] + src30[100] + src30[101] + src30[102] + src30[103] + src30[104] + src30[105] + src30[106] + src30[107] + src30[108] + src30[109] + src30[110] + src30[111] + src30[112] + src30[113] + src30[114] + src30[115] + src30[116] + src30[117] + src30[118] + src30[119] + src30[120] + src30[121] + src30[122] + src30[123] + src30[124] + src30[125] + src30[126] + src30[127] + src30[128] + src30[129] + src30[130] + src30[131] + src30[132] + src30[133] + src30[134] + src30[135] + src30[136] + src30[137] + src30[138] + src30[139] + src30[140] + src30[141] + src30[142] + src30[143] + src30[144] + src30[145] + src30[146] + src30[147] + src30[148] + src30[149] + src30[150] + src30[151] + src30[152] + src30[153] + src30[154] + src30[155] + src30[156] + src30[157] + src30[158] + src30[159] + src30[160] + src30[161] + src30[162] + src30[163] + src30[164] + src30[165] + src30[166] + src30[167] + src30[168] + src30[169] + src30[170] + src30[171] + src30[172] + src30[173] + src30[174] + src30[175] + src30[176] + src30[177] + src30[178] + src30[179] + src30[180] + src30[181] + src30[182] + src30[183] + src30[184] + src30[185] + src30[186] + src30[187] + src30[188] + src30[189] + src30[190] + src30[191] + src30[192] + src30[193] + src30[194] + src30[195] + src30[196] + src30[197] + src30[198] + src30[199] + src30[200] + src30[201] + src30[202] + src30[203] + src30[204] + src30[205] + src30[206] + src30[207] + src30[208] + src30[209] + src30[210] + src30[211] + src30[212] + src30[213] + src30[214] + src30[215] + src30[216] + src30[217] + src30[218] + src30[219] + src30[220] + src30[221] + src30[222] + src30[223] + src30[224] + src30[225] + src30[226] + src30[227] + src30[228] + src30[229] + src30[230] + src30[231] + src30[232] + src30[233] + src30[234] + src30[235] + src30[236] + src30[237] + src30[238] + src30[239] + src30[240] + src30[241] + src30[242] + src30[243] + src30[244] + src30[245] + src30[246] + src30[247] + src30[248] + src30[249] + src30[250] + src30[251] + src30[252] + src30[253] + src30[254] + src30[255] + src30[256] + src30[257] + src30[258] + src30[259] + src30[260] + src30[261] + src30[262] + src30[263] + src30[264] + src30[265] + src30[266] + src30[267] + src30[268] + src30[269] + src30[270] + src30[271] + src30[272] + src30[273] + src30[274] + src30[275] + src30[276] + src30[277] + src30[278] + src30[279] + src30[280] + src30[281] + src30[282] + src30[283] + src30[284] + src30[285] + src30[286] + src30[287] + src30[288] + src30[289] + src30[290] + src30[291] + src30[292] + src30[293] + src30[294] + src30[295] + src30[296] + src30[297] + src30[298] + src30[299] + src30[300] + src30[301] + src30[302] + src30[303] + src30[304] + src30[305] + src30[306] + src30[307] + src30[308] + src30[309] + src30[310] + src30[311] + src30[312] + src30[313] + src30[314] + src30[315] + src30[316] + src30[317] + src30[318] + src30[319] + src30[320] + src30[321] + src30[322] + src30[323] + src30[324] + src30[325] + src30[326] + src30[327] + src30[328] + src30[329] + src30[330] + src30[331] + src30[332] + src30[333] + src30[334] + src30[335] + src30[336] + src30[337] + src30[338] + src30[339] + src30[340] + src30[341] + src30[342] + src30[343] + src30[344] + src30[345] + src30[346] + src30[347] + src30[348] + src30[349] + src30[350] + src30[351] + src30[352] + src30[353] + src30[354] + src30[355] + src30[356] + src30[357] + src30[358] + src30[359] + src30[360] + src30[361] + src30[362] + src30[363] + src30[364] + src30[365] + src30[366] + src30[367] + src30[368] + src30[369] + src30[370] + src30[371] + src30[372] + src30[373] + src30[374] + src30[375] + src30[376] + src30[377] + src30[378] + src30[379] + src30[380] + src30[381] + src30[382] + src30[383] + src30[384] + src30[385] + src30[386] + src30[387] + src30[388] + src30[389] + src30[390] + src30[391] + src30[392] + src30[393] + src30[394] + src30[395] + src30[396] + src30[397] + src30[398] + src30[399] + src30[400] + src30[401] + src30[402] + src30[403] + src30[404] + src30[405] + src30[406] + src30[407] + src30[408] + src30[409] + src30[410] + src30[411] + src30[412] + src30[413] + src30[414] + src30[415] + src30[416] + src30[417] + src30[418] + src30[419] + src30[420] + src30[421] + src30[422] + src30[423] + src30[424] + src30[425] + src30[426] + src30[427] + src30[428] + src30[429] + src30[430] + src30[431] + src30[432] + src30[433] + src30[434] + src30[435] + src30[436] + src30[437] + src30[438] + src30[439] + src30[440] + src30[441] + src30[442] + src30[443] + src30[444] + src30[445] + src30[446] + src30[447] + src30[448] + src30[449] + src30[450] + src30[451] + src30[452] + src30[453] + src30[454] + src30[455] + src30[456] + src30[457] + src30[458] + src30[459] + src30[460] + src30[461] + src30[462] + src30[463] + src30[464] + src30[465] + src30[466] + src30[467] + src30[468] + src30[469] + src30[470] + src30[471] + src30[472] + src30[473] + src30[474] + src30[475] + src30[476] + src30[477] + src30[478] + src30[479] + src30[480] + src30[481] + src30[482] + src30[483] + src30[484] + src30[485] + src30[486] + src30[487] + src30[488] + src30[489] + src30[490] + src30[491] + src30[492] + src30[493] + src30[494] + src30[495] + src30[496] + src30[497] + src30[498] + src30[499] + src30[500] + src30[501] + src30[502] + src30[503] + src30[504] + src30[505] + src30[506] + src30[507] + src30[508] + src30[509] + src30[510] + src30[511])<<30) + ((src31[0] + src31[1] + src31[2] + src31[3] + src31[4] + src31[5] + src31[6] + src31[7] + src31[8] + src31[9] + src31[10] + src31[11] + src31[12] + src31[13] + src31[14] + src31[15] + src31[16] + src31[17] + src31[18] + src31[19] + src31[20] + src31[21] + src31[22] + src31[23] + src31[24] + src31[25] + src31[26] + src31[27] + src31[28] + src31[29] + src31[30] + src31[31] + src31[32] + src31[33] + src31[34] + src31[35] + src31[36] + src31[37] + src31[38] + src31[39] + src31[40] + src31[41] + src31[42] + src31[43] + src31[44] + src31[45] + src31[46] + src31[47] + src31[48] + src31[49] + src31[50] + src31[51] + src31[52] + src31[53] + src31[54] + src31[55] + src31[56] + src31[57] + src31[58] + src31[59] + src31[60] + src31[61] + src31[62] + src31[63] + src31[64] + src31[65] + src31[66] + src31[67] + src31[68] + src31[69] + src31[70] + src31[71] + src31[72] + src31[73] + src31[74] + src31[75] + src31[76] + src31[77] + src31[78] + src31[79] + src31[80] + src31[81] + src31[82] + src31[83] + src31[84] + src31[85] + src31[86] + src31[87] + src31[88] + src31[89] + src31[90] + src31[91] + src31[92] + src31[93] + src31[94] + src31[95] + src31[96] + src31[97] + src31[98] + src31[99] + src31[100] + src31[101] + src31[102] + src31[103] + src31[104] + src31[105] + src31[106] + src31[107] + src31[108] + src31[109] + src31[110] + src31[111] + src31[112] + src31[113] + src31[114] + src31[115] + src31[116] + src31[117] + src31[118] + src31[119] + src31[120] + src31[121] + src31[122] + src31[123] + src31[124] + src31[125] + src31[126] + src31[127] + src31[128] + src31[129] + src31[130] + src31[131] + src31[132] + src31[133] + src31[134] + src31[135] + src31[136] + src31[137] + src31[138] + src31[139] + src31[140] + src31[141] + src31[142] + src31[143] + src31[144] + src31[145] + src31[146] + src31[147] + src31[148] + src31[149] + src31[150] + src31[151] + src31[152] + src31[153] + src31[154] + src31[155] + src31[156] + src31[157] + src31[158] + src31[159] + src31[160] + src31[161] + src31[162] + src31[163] + src31[164] + src31[165] + src31[166] + src31[167] + src31[168] + src31[169] + src31[170] + src31[171] + src31[172] + src31[173] + src31[174] + src31[175] + src31[176] + src31[177] + src31[178] + src31[179] + src31[180] + src31[181] + src31[182] + src31[183] + src31[184] + src31[185] + src31[186] + src31[187] + src31[188] + src31[189] + src31[190] + src31[191] + src31[192] + src31[193] + src31[194] + src31[195] + src31[196] + src31[197] + src31[198] + src31[199] + src31[200] + src31[201] + src31[202] + src31[203] + src31[204] + src31[205] + src31[206] + src31[207] + src31[208] + src31[209] + src31[210] + src31[211] + src31[212] + src31[213] + src31[214] + src31[215] + src31[216] + src31[217] + src31[218] + src31[219] + src31[220] + src31[221] + src31[222] + src31[223] + src31[224] + src31[225] + src31[226] + src31[227] + src31[228] + src31[229] + src31[230] + src31[231] + src31[232] + src31[233] + src31[234] + src31[235] + src31[236] + src31[237] + src31[238] + src31[239] + src31[240] + src31[241] + src31[242] + src31[243] + src31[244] + src31[245] + src31[246] + src31[247] + src31[248] + src31[249] + src31[250] + src31[251] + src31[252] + src31[253] + src31[254] + src31[255] + src31[256] + src31[257] + src31[258] + src31[259] + src31[260] + src31[261] + src31[262] + src31[263] + src31[264] + src31[265] + src31[266] + src31[267] + src31[268] + src31[269] + src31[270] + src31[271] + src31[272] + src31[273] + src31[274] + src31[275] + src31[276] + src31[277] + src31[278] + src31[279] + src31[280] + src31[281] + src31[282] + src31[283] + src31[284] + src31[285] + src31[286] + src31[287] + src31[288] + src31[289] + src31[290] + src31[291] + src31[292] + src31[293] + src31[294] + src31[295] + src31[296] + src31[297] + src31[298] + src31[299] + src31[300] + src31[301] + src31[302] + src31[303] + src31[304] + src31[305] + src31[306] + src31[307] + src31[308] + src31[309] + src31[310] + src31[311] + src31[312] + src31[313] + src31[314] + src31[315] + src31[316] + src31[317] + src31[318] + src31[319] + src31[320] + src31[321] + src31[322] + src31[323] + src31[324] + src31[325] + src31[326] + src31[327] + src31[328] + src31[329] + src31[330] + src31[331] + src31[332] + src31[333] + src31[334] + src31[335] + src31[336] + src31[337] + src31[338] + src31[339] + src31[340] + src31[341] + src31[342] + src31[343] + src31[344] + src31[345] + src31[346] + src31[347] + src31[348] + src31[349] + src31[350] + src31[351] + src31[352] + src31[353] + src31[354] + src31[355] + src31[356] + src31[357] + src31[358] + src31[359] + src31[360] + src31[361] + src31[362] + src31[363] + src31[364] + src31[365] + src31[366] + src31[367] + src31[368] + src31[369] + src31[370] + src31[371] + src31[372] + src31[373] + src31[374] + src31[375] + src31[376] + src31[377] + src31[378] + src31[379] + src31[380] + src31[381] + src31[382] + src31[383] + src31[384] + src31[385] + src31[386] + src31[387] + src31[388] + src31[389] + src31[390] + src31[391] + src31[392] + src31[393] + src31[394] + src31[395] + src31[396] + src31[397] + src31[398] + src31[399] + src31[400] + src31[401] + src31[402] + src31[403] + src31[404] + src31[405] + src31[406] + src31[407] + src31[408] + src31[409] + src31[410] + src31[411] + src31[412] + src31[413] + src31[414] + src31[415] + src31[416] + src31[417] + src31[418] + src31[419] + src31[420] + src31[421] + src31[422] + src31[423] + src31[424] + src31[425] + src31[426] + src31[427] + src31[428] + src31[429] + src31[430] + src31[431] + src31[432] + src31[433] + src31[434] + src31[435] + src31[436] + src31[437] + src31[438] + src31[439] + src31[440] + src31[441] + src31[442] + src31[443] + src31[444] + src31[445] + src31[446] + src31[447] + src31[448] + src31[449] + src31[450] + src31[451] + src31[452] + src31[453] + src31[454] + src31[455] + src31[456] + src31[457] + src31[458] + src31[459] + src31[460] + src31[461] + src31[462] + src31[463] + src31[464] + src31[465] + src31[466] + src31[467] + src31[468] + src31[469] + src31[470] + src31[471] + src31[472] + src31[473] + src31[474] + src31[475] + src31[476] + src31[477] + src31[478] + src31[479] + src31[480] + src31[481] + src31[482] + src31[483] + src31[484] + src31[485] + src31[486] + src31[487] + src31[488] + src31[489] + src31[490] + src31[491] + src31[492] + src31[493] + src31[494] + src31[495] + src31[496] + src31[497] + src31[498] + src31[499] + src31[500] + src31[501] + src31[502] + src31[503] + src31[504] + src31[505] + src31[506] + src31[507] + src31[508] + src31[509] + src31[510] + src31[511])<<31);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25) + ((dst26[0])<<26) + ((dst27[0])<<27) + ((dst28[0])<<28) + ((dst29[0])<<29) + ((dst30[0])<<30) + ((dst31[0])<<31) + ((dst32[0])<<32) + ((dst33[0])<<33) + ((dst34[0])<<34) + ((dst35[0])<<35) + ((dst36[0])<<36) + ((dst37[0])<<37) + ((dst38[0])<<38) + ((dst39[0])<<39) + ((dst40[0])<<40);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h68e92f7f29e2e4aa8f26a5c1d0221257a02f733d861c1828bfd481b36cf9fef1fc623412151ad42ebecd841d06c227d6b0bc8900e04ee5a13994dd51e3da0d16097487d1c40a6f2a46b2fb58f84fcc40ba8796c6ac782b81aecab53051252248ba89bcab43895dab608edbeb75633d925f85882a04d0c39d2ebe82a70f3543930e7c9bd8077ba6f8952f501d1abfa3f35426c8bc51c8caafb0511dc76cb19255cd4ba7d11ed4d7910360d9daba929fb7ed77ceee76fa81b9cd868ae3558532bf86646a4c786c2ad49281f993c03de33ebe7e239ce46dedfe43876f41512a8a38d69467f8601413eb1da7f864bf6caa2937e999ecad19a58f7e3caa4813cf5e1f55028c46a3c679f9249a3161c65dbadbfeb108fc101cd454f9656eafa78304179e76e6b02d90f851f67c630927ff4b477ebf24629ae600e3477ae67e7ec5dbfbb6bf569ab37da8cf0915c716780b49ab6301e064cdf127c8a9774a62e1731fa8491e5ce9a87e2d94858fec3a9ac7c607f5553e479cd472b4ec40025945cc8d4bd4136a8fdbccd4e88ed9d1639baf3cc9faa21e6692cf1f0be8a81c328c1804d1511afff65b4e1b5361ea268723f8f855324a6e619fd554a0dfc018c5dc88c39002ce624c7149f393328f1d1f5a63fedb48482e21e0784d368818d0d364788c419f5b3822d0fe2429b66e9d12f8f05d1f59b66cddb242a338131ae5a78ee462edf9cbf9b7f232c861fb7fd0c42fdd0883541707b7da201d93615e7e05fdca0bac107cb75ac83e34b4c35c431c6245f4f5daf5183a9f12f8b4834860deee50cd2d0ca145919f0dba58774e4d1b7abc1a3aa88e2cf2265fa5d3d44c20d952013459bccbe67f0d2504e00f1c460681d67de7c70a1ca593bf9be0cd05e390f4ab93f12cd43945a680b4d9f1ab96f018722ffdc976069f67fa4ef2a51459105d9d4bc8cef94bd9c60d95dfa738c4b6bd61ef01e63f8fa018b0345662ae0c9c6c1c5ff5d820071b665381a760e126036ee91f17debb323d5f207519c6a5789fb2abe86a3ef7bd2f855e645813e04c931068a4f78f47d987a995bdaa075b18d6f473f0ba27ab3e667ce5aa6e46afa2b93959ab658248d7246ad1147ac9196baa814b72fd127aaa9d135facc8dde78fc384ea2d12759ce33b0f03797eccd770a5d2dfe2ebb58c1a293517c32cc5f1a5cc78bc3fe9d0d4b17e4becf7290a6241e3bc4952ebcd848da603525d64116177936f000ef78807a8bd709e0e99d1629ac6bc677bf6d5aa86537690ac8cb62536f08826f28d57b9c2f0eb2fef4a85cd89046f70e2dda8c480a76d6fe5bd59600d9527736a07b0c0438ab1f7e6dc9060873991f465067042b7d36de34039ef8a4816664cc067676b73b2c8edc1c6637a33be3ae8a73ec75615284264671eb4452e3221db5b9f87e65c46d57392532bbad46c0e13f3e5f67a311b178c5711c2c205485f1f3ed10e050264fe695cd3788430823162aa5b8adaf140722e8d0cbf57b0f593258b8b1c74bab8041131ee201c8611375f701944bc064cfff97c72ef3027c4820f280d85076def76f30e3ae23f6d203f5850786351f4f72f5f98b94b27e230dfd449e9604d100bd54933746f8d009141633b2a3a71cb1007e5abde519e15387226638f6f280e12ac5f5bf7ccc389f756cae39f4683b1e513a48fb4b38bf5de107b8c63fbca80fef6b60998957743bf2b6ac75696b446755d083c3738875c54ac27fe733efe586ba961c1a363dca2fcce42d03862b3a58e26aa896a8e2ee26685e61425b72c6dc5c0a3e4225b5d42848ec29ecfd192f74d5796b203f241ebfce968c3fb413152d706062e038332f8dbc5e0658434e7f75f173dfa8637d72eeb24217999a05a7d16c0d85d8224225f868015e5e523ce5b60cb08a67365df73e2d747f1af44bd2e8363d8773f99ddb175e3d09194c5cc99eff170bc836a9170c45daa4cd0deb5179f3558859d1ed71df736d5354e1451c135c1f477f912168db0709d79285199979d2a2b168469471798abd9ab47dd30f0e75c3071829438a59d09fd4f28ebdd7d303c10a863a26afdb4cfc1beab134e43d442e0a5a82e6cc3bfd8771e1f61b004d4a7ddc60a9b05c3af4d5cb0520fed54cd8793089b1df005edee71d26baee7c4de79bd7e391a4a692047073f5e0a5ac7a934107a8ee32bc7d9da04fd086eb23812eeabb8c0e4256cc1fed7d57e4c6450fe27a8acb35cc364a36aebc9fc04763263a240d6c0510374759725e64527d669eb2c23a3db062899d88324ddfde155926ba4331622f5b62b2d852a9b477e7403f1374c42e12fb933579242d900e07e9445723ec18dbfdd1e5569baf81d6ac209014bdb437498cad1fbed1aa689730fe825d43def4c757d4639f1ff37b33357360c18ffd6337471070d04d0f76393dacbe084a3c04ae17c08fd5d34cf00675cdbde937c94ffda9d11e5083b0106f69984a0684f2934585e9d2e772dcdece87c11b51d3c3e73efb6388248a5b7b374d921b128e4b11d45c80545160ad57347c4c8db6e7e932096d5b7470320843669718beab97021585bb8c5cd2d03e0b44c3a23d53f445cecdfbd4a75d375ebace2fa5d5380a166384b6816088fdcac2252ac8302e5022c998f177f0f4dae280948d07bb237852d578e8e0eca0a2665692d2eebecbe8eb9ad086825b8dadd79f9406062513ea38fd2763428c6deeff58b3ddcc33eaf48604e2fdc309d09ca44a237bb844949da61b180dec165a61b93c208328099e84335c4448ba2c6120529f5aff64d71594dcb17151cce4a1aa0902e2ab107994e80cc008e8b6e16d19e1999d2b04fe2ea5c325d7f51656c8850614078331745272a67976af3af02e4a982c6a0d139392bbd4a717c5c7bfa29404c62;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h8acb42bf04281c438f59c38f1c238b8d0a9f65f48c0bb2b95eaca49bc50742884301c91dd4a1af9d3a63a64426f8b61aef9af42c7c96e261e6e0353c36d12075211a509c817661cc46215e57ef5904bca19d36b0290c70c4920da53487a1a23e16b66a0b9c3716b82886cd477f14b026ad981e4497edd276cc17fe0af7bd740fc69266174fa015813ed54739ee49f167b48d3028d3b67ae675fa60ad38a7f39dee5b9b5711c6e5dcc5041ebc3f7399325da4911418d81a644d275e8980a276a16febb06e6bfb956c0b36ea1e0204b12f1787c915f3268330e67c6ad39e009eae55e8044824e80993488d439e128e0590fd91afb20c62c823460217b7d3973fc739c6bcbd9dcdc323c2f2d126601114ca1d0fdd48e0463a5c375418f16fd51d3fc2a027e5967f5157705b27681ec3a9bede0ecf8fe3d2e98f60e18c9fa94e1accbbff6cd0598d016d8177a5a8ce6b5e1102429b1ed6c624a6b1723377dd3012a719ebeb6e26ca484ac5e8943a6bceef01b5a50377a7f11521224d677a3451ccd37f8e4e494c0b09286dada55c7a0bb665b79fc7cf10984e847be30cb0d296f48804a7eb648f1d17983d9478c7b8c7e7a952c8da8f5fbafecae85f18019476d040f2a79efcc539100021d66f4779cb3c11b6cfe08216dbe5e43d3e88ccd991ac02a8b36e54dea9d4bbb335d4d933e7a648129f8947cb0ebc696ed356e3dd7b147eba005fb0b674020a95ac6a3becee32ffe1d2a543ddd337cef5027d63a4e605427f49f63e41a7672105c3213aee8f419ff2b3f12acfc73ae9911a90e5a60cc096b6353051ff3c2cc09ae78888d3fcd5896368c827eda676fc4fa005a38dfffe3441026342df2bbf8535e823518bf79627c94b95f43789cd9c6a614624d4f03df9698f6cef93bc361ecd959ab24fe72cd252110171d8166cb92ebd1af072ec0b5479cc42b302c6e4eb1b442c236a9bcfca3f274ab46b94388192331909efc5e9652f9cbf9b6519ac2bd4f34626c4ef90b277b9e70f7a898c06781f7440d5eb5530835698db33ce6d3ef1eff69c60e333028a74ff089d479adf2c3dad4a1af530fc06eb49b5797f172fd79b11c8353f2a1a69e77675bd22a78794621e568c3ef6ddba76231d772498465c3525fc3a357bf9ad9dfda6ce4bf26d4647aa187277f78cdbe83ca5376218112918e5e8fae959abfe88ceb8b9f8963617a8830ad4f9dc815b633be6c7ed50570b139d0cf837ca5b4c7d1fd07754fa62a5511aec43d823d25922290c9fc3f0f9c5c902308b416a48652c9f923ed3cf08c4b760309e23b856d6be0ea95737132dd2a24db6ada9919f15f3841e3803e9922dc916984ee73e63c1b6f9868e31e2eb0da7cbd6613a550cdfb78d3e4229029fe89ef9bd42a9540956c0d504510b32680a31fa3eaee796dadc4ed002180687ace7b4df3420640f7e351cec78f89e41535774fd2ee86306a18368a9ab256e701512b5f489fad18d280034130eb108d48ad616d4f6cee772743ce6d1b820b102e27263afd397818b4a0611c06d3e12251a5ca04d3209d9114cdd4f819c67bafb8997d04ee66979eb4daba8fa3d8df19123db62ceed2959d651444cdbb86b3ce12e4133e779c171a12c8c99712af4f46cc7f1075a6f162030f9746143beacf7bd5819102eae248c63988026515c8019e436ad50f480397d1f269323820efbfb4a2b831620813accbcd4ef589d0ffb1f3d1a20d18e7ebb9f6fb3af7555fde29dcd5c2228cf09edfd80fc610b91c6bdaa260c1098a370fc77b396c7d6a6687908b26dce3fb3df8af666e8344cf998f3de0b210e6ba8c502ab74029c752b4e1271cd10f23555b181a1f587f0a0ce8351c0f0796f974402478d0245a74b725c97243560fe8fc8db6d6845d294c1a22e9344ad364aea80f300ea5dc87a965193514fc812b5b4f7ecc3d28870aab281aff6bb661f7d26d9cfa295846011be044aa2e7817dc25008a738b0d1a2e76764caa0230c035036d367b100e6d8e303f44e3043737d86520361b8bbd81bcc9ce33fed78d82ddcca3dd23475c77569bfd3a208991de08c5721cc727aa5306e2914c0624a756774a976ee52eeba41e6e18de44d17c11a5fe637ea3df3e1d8cf634a953a7865504a5152ee42d0c4a28a55bc66dcd364fc1701601525a8cf8dea3a93b824b386a90d3d5af45ab18df0a1014640d94a6cc7ab452e66598c5f9429c00c0f86a4fb3f42307481e78b6d6860bdaab3e6f00e07d574d3aa76aa9430a3df4bcc62e6212c45b7a0bc00c37d7f935cd66a0869549f70db2218afa51c67e6344960f377b0c1bd1e0657a09831141ba1074f835cb3702418f694718170117c4a40f563b0794fb4114884392276798cb03ae95d5cb2f76a95172e3b1e099412a831e9a6e14aa56bb8384e116265390135ba349f26e2d559aa2b663992337cf993800f4980fd978b1d6431e548557734dcc1387caafb589d1ceb51add857541a716709e308212aa237f69b1133a44d90608b7b1df035b53fe4908559ab6875e34c04acef0eb09595a0f02834e0dc7885b034c2f6b09a0c0ea2729d5eb9d65561a75bacc3dd0d85d27ac68e28109b195fcaf56481b02a98c184c68ab8756c49c3df32fe6526ea05777dc1105e452690755033254a605ad07e631a9f78f67a78f71942aa44616fc041d83692350cbd1d34c80bf21948155b9e46a0e57b61146e98fd2e13e444a9002ec066eab73ed353239fc6f9313505bf3b98c31c8976469a4487a2679e53f66e99c6d1309c4eeee20ec4cb57a6df314118142517c6e1fc0ebb4fc50e094fce3da4b0682aa9665423b52649ddc7fe1ff8bdd1f3340411b500d478f522615aafc7163f7f0e71424afd24552e5b28753b2f274ea9dee5d2be33;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h668ef69dd12883c980327040adb777039697435912c7da661ad38cf2a81550f0529d2a9d4dbd77ab907bb8b643bf30e5f835015f013bc2e48a905d6ccc393e86a0df4d5149654ffa037e7d419aeb95a7d0079a79cbab717f1a9e27eaeedd52802c0ce204328ea3456882985235e46169c9a4bca4d90c2a585ca62e7eea2143c8bea0d8a9aacecee1e2d2b9846130af7d51886b09c265004e682dad709537ce8ce50094606b589250e34e37fd4c788e216ce52cb4115e777cc86aa01d13635cc07130aae23e260867f54f021e84b907ccd423c0653632627ea1ee5f39d3e90125e6fbc9b067a2287ad0327a9ce39268ef7e9c6588d2af9b27f5e08211bca226be80846c65b005130bd7edc4efbe953ce879dd2b594e2a11f42136a1fe9777814360f71339f7265a725c2fe92676f1697bbc365f426b0fe418102c7a70f47f9d48eb8adb00834807e643d42b815f58da58f9e0ffef5bd3bf0ce7db10eddf462f95d1d37ae07a80e2c0fb14d9de94231836175414a4eaeae94ae65c8d8aea3fdd1d736a029008bcbf8df4e44c9e8fdd7d33db7e1e807b00fe45d38e28179874563fd8e63f46749ad7fba3459dbcd297b6c0d5822a41fc792bf69333b919d642b2ce37dc364328b0891bc3550818848e0e0ae2d30e90dfd89e1d6a91d17d2fd8c99e8351a8d2ba990804f32328634419484dd7ddf8b753ed80e7f6af114cdbe9100360ea6fbadc0f5eefd67c1c77629092e5727134f5ddf388e60af5697e43c60159b16daec4262dd5a8b9885af4e569f440c22a974817fa2fcc213bb4280990bdd8e2915e2e38d872889001e690638d336c2f7a4a14cc3e15b5f241aab5d6dc59e3c04e8f1f9d3af65cba3d7176f817075ccf88b2d9f78630e4dbe51197ad377388feeab27f0990cd2c66d0168198575729c11abc679a91fbb9ec98a015822c264ee85da8764b1fc673720050b259b725d0a8ee5ead7d32a9cc601059d80518b7454300ef63d8c86643b115ae1e22a43a7e8169f68836970d19fd7088224d8f0941994b53aab6031131c215b9029842ef3da22e946a64c2b6339263aa0d49b380afef2a1a8eaaba1a1590fad4e55e936dcc22c70495becb597fdaa7f383adc68352ab308d2ebc7ee2df694dda036f0a346a22046911c11feaa2b25f1f0d7aabcd8ad40b24d21dcffc683eedaf587080090ec8030d54df106f78fc97699d7b52cfe9dbdf3a02d5361e949ae57f95f1ee593a2ae35623d5194c63c310df0097a53be834b21e3c68be49ea56cd43fcfc98a6798b6f5fb3b71e2812dea986e001c48d7a5f8f22654b7d3374b3a13065d4ab51be610ab295aecd842c569418babe20645b07e9ba22094af22ea39b33b27023f7d6ad9b392249fc5560a3ae18b18949437dab32aab515ec40ab84d1b2a2e9245e5472121f445434ef0667f7d96ef890a829ad70e23d9b1306bf1e2145d2dc87a150a6098bc9ed380a057e4f5b38afecf776a813558262b68c3298ae49084349e62ee7d7db7117a08d6eb56aa6a9b2f8eb2c3ff5b9a3edfab5e69d7d1ce571924b4bf93bef71e9a707fce2f4353237020b6ed893ec7836428b085ebcfcc9d24c5cd8a0141803f1c20ad53b9e75a00199cdd867d333e30888b0eb9726cb3f602385363bbc9f63fdcf7437c5633d1164b6440e47e449d2b9859de9723b112101f93a2b922cbf690c4d4648ad87047e74d8f2d2bc03c59e4fe8c0df5dfb0598109a12fe2689ae16af8ba81802590d2503e7f900d71f868c3261e10da012f998f20166729263ec2734934f73a26b8eb85ee98d1fa6f0ec90fa93406d3ca69ed815237259245cc0152f827fc8a5559a82e171529da1097e0605f89bf424a54148f8d5eaf8156f50bd6209f449acd7efc94725a428185b9a0b15fba63d4d32b559e9ec18db5707a0f1666fa5b38e967be96dfabe548b53263e152ccafda79f22eea040f8f94f7ee9284a54134693fa3eb9d704a7df04c3e9b8355d97fa0050bd6e0c2a5c8f50ea10e63867dcb4fbcdbbaae7fe534fdc357dacd5ca92c775ec3d3ea61874d6d4d73336c2cd06eba7f4ab952384c00c367f14ad6abac0007eb43a99b951fde580d570d31b4dfa71075e8ec6109184b15296c50cc297ae3e1e3d209ab471f174ec49646bd0b015eccb4880525d4bf1363528bb6672401eb4cda7b6648e5bad6e0f01446053037b797203d9396911bb17e2b882da050972b1d20e2838ccc8323bdac4c921ad02243781214facceb1528a87dc2298a89c09df480fab5fb7a2adcef63c6aee7b589c06e30ed615a9fb9b989e3160093412cc9266a1616e2eb7306ba18136a0f9c22a3c585722edc888e1858ed2e3eaaa9fa3bd1c76cff338c282bf5b754b1d7ce7269550f2e14cb0b150a6c33ae74a7ecbd481d456bde7f49b2069363f5647e7fdd52c9737660a27c8910bce976d60e02244e07829901f2b156fdbda83a1038ced95c6f678f105b8cc9c65cc871c06f6b47a501fe59c8863e1970a47b82f73dbbbf81a50ca6d1434d34c741258d15137fd79c40e8a570a701339fe10159ba4b37007c162aea4ffab6e4635bbc6e19b7644774ed26bdb0a860046fbfac03aea885827789e35c75baea2b87fe0b8653391ba7a72ea65b439d71c8bd9f8a5552a1db7a5f3f64cf0b78166c5b4fd8994e556a15b984195a4ea7ea37dcdce50f26666d3cc2dc336458b49fcb5e2529408fd81414d7a370ae2e3aeb154104c32797daf13b87bf4da9e07a3d427fc31a1f8448f032c81e59095f7fd053da7cf77f42b73390882f8709467ca6e3c9310e5d538aa19be9e158f9a5a906bc96a9f80fabd4fe4e99122d719f2c88c28abcd0249328f66f218d4f03d870c4d6c8ba62b5ea43e11d297683baa7982b5fd2b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'hcb1e984092d96a0100d0a84daa520874edc8ca325b2b98453670644e6051dbbede2512b10cfff3fe69b58fc4905cbc822eb5930ffdcb4174f1cf33f8374c9ebb5f4fff8ed84d3aa1cf377f70a749c10d3b66af3f17d7b20c4a980cdfc836a4b78f5df24140c0ef4965cd61929b1c2ca4130424c57ff69c9fddf6ba21c71c87fe5339a58a4445a2489f0590bdf6f68d947f3a253ef56a5876b794cc484f43cb4e6c30c5b34b58cf5b7a6d04199e0fcb71d3e158530a954bc7e05775eea5363571e0b478456bd5b53dd17cfb074b853eaaef9b214e3dc05133a75f8ee24df77d91f88dc87e480c7f3170fe16352b04d543c410f0564f34cb86a3c71f078e39c96f81edc02593ec2f25b809a472404f114aac2faa8b325ee54f05d83866c9354a956f8958f43dc74c5d167cdeefab4414008c850313c9d8ff93b06b7e69911fbacddfebff4c397e7b1a3a480215ec720c8b5c49c63a207376163241e68e2e04eea4fd7c23ce901a2f8dd17564ea2b1b5c6ab2cf7ef46ad0b3175bc069818d0a02a5b5a78f0deb12e1e1333cae96a67f8d099ff346bc04ca7bb15037bdb8e9501b79612f4901313ed3431d7551e820c44aa36f479a38a0a090a2b2d147dc028b58e174c98884fdac2548343dc623c1ae0b4483705a889f2cfe13b08b7e2098b4ff09833cf347bfe49f302f9bbec4a2ab16078c32843f2312a332e223c3bc9f1f19d15613247e65ea4cf90f5e6cb89b63cd44a501cbb79b9d001d2488b6c43c1f4442b2bebcbaf39a68b1ccf8005d6777d43f2732232d0b269de48c6fd95f947ff847c1396d99e98c73a0a962411008f8ed8f422261a56197a993eec51d7aba077abdf5ea05309acb55fc054a7bf2761cb1a7f45ee62208aafd5fbe4befba22b7561779439cc695b98dbcd6e1ae08e4c7853797bd8fce3bdb5fff808e1db6e2433288da89ed7992d4d51a950c9aca9c44123c2282dcdfd78a5dc9b2bbbb528d903c6d2cdcb62e5e57b9837fcacddeb1f81d04bc9f3aa4e874ae72f49e118a0801aea3101bbcdb191397e1fc28629916c4002fa6a913fd743f515f58c74fde345db7c43059b987b6c15f41ddff0f94c67dca79885fe1e7a4711b083d21254fda5a1c85871ba4f7d557741a4aa181d3cf055d8eb2875e90f295348ff5e54a55d3bc6bfc05c848d606043b8a8de4c3f5ec9ca8c015ba82e9cdec8ad0ce4745e1eee9ddee337e1aebe90b9187fdb062955b5abff7a2dd1eb762d4ae2d6270a73678f3344fdac66d368e69fd0f1bf6e412250600b9fdf6d6e86f0254cb7ad117238b7d4385996f98edee00eed46abcc5604ee97450f3ad0423ffc33b0b98d039ff8e6a622679ac7d3571616b1a90fc091a0aefcc635d6d26bf1d179b664d145f2713bc8809a4d14ce8a7adee0186b1a7116425a512d0107e08845833369c1e040c7bbb94d3dee061b72682a02aed0e1bee7dd4ab54025549b70295b73ff27c7a813853e422ffb259947d3deebb0a9245a93fa7afbba4760880e2c08784eb8312fbb0bcdb79713cf6b524fcbcf13984a3d2a1adbc999b7680956180aeeff9a871d95ec418a4582e0b76506b1157e508249801e687c503c078eebb1e13702c3627f49de4a9ef810cc54bc221424d355851e1c224b758254361460ab42a93399c8b6d4a5b87f249bbc5d144555d03480bf003103cb69ac567b4c12bd83adbec6ba09a76af1950780e31c5663282de280b8cd26cb391bf304312024307af76a402fb45a3d97864c6b9a5fe84d69a2a58796d4f8d87780bbd41e1c762f5d9458c83891fa2a0da8c20fc53f62c12b8f8083e101008ee98fb280729fd13ded12ee8ae5f789a16a4880bad696567fa5eb1a2d30db8629f2f696db80462633e5fc5735f29b0039e608e28f0b65f2da7f9c58450d7eb7f613ccc05f4d5c1cbf92c062c0802a114a719bdefbb7b4258bfbe5c60029ced5e0de912929ce1a1477b8b4364ffca676844478ce6434c675054fd775d224e1a7f0716f0645178b9a537af20b0e564f1e2822250966ffa0b71a8fd7b788fc24dd99638c1c5864c9df56346afbcf71f4ac46ccad24fbeaf0426f31cb064866e8683f79591837798d498ac5bf070d1dfa712d2795cecd2eee8ee6d76a1f58516d60c0c3e4cc529e5589435ecfe57f6809df5266a5224f69374b0c1ed434f7c23a6d3156d2d4e17e40d29f4ea8a0ce66ca362447a87a62eb6d396ebce537c4e83d218948f7beca56f056208bcd88126369494bdbd82adf3e7897944f7c88f38293fdd1ae1601041fa2af4c03523232a86ce888a20d5eb5123b30da9c59be14e05a84e3800776eb55f9023a90d830a2b285d3ef3362769b281cb252dae85207026052c6a28d4330698c17b52b939171e1be8133716266afc9e1a2fb16e935eef70eeb1f89b4f88228409ebb1331a2be2ba4d754e2be55778c2cd596474af94339fdfebea2553b7b7c7f9c7b877449a6913112615f692d81267a804c55269e2aa2fa2806dae8cfe48f655e0357537e2a5c028dc382b7c6bbcff230e7a77e0288ca7bb77a8d6f017a4d91c3ec1294a9f2ff7538a0feb1b53fc39eaf51701ddfb6d7631f4c6fdb6f4228ab0e9b40e4d49c46c3bad5d02f6acd14f6d20e9e7aee14b1ec5af74254d73c868a009b0ac41967a038acbb94713defdb391b8931763edd35e5cc27d9a8c4478f9ed6056be38294ae759756004bf1694c02f65a3c93454ca06e8f14ded05f0f452382fd86a463c86073c5d82b6014e491862cbeb65d6672d005ecc8aea86b8d349cb130c03e477c7021e76a228ee2388449221d631a8fc201d9215a8534cc8993b644f08932770662ee6d500feb48c99b96f8cf6e0e30b1d604601a59c0ab8dd4046c7e41315ea6a1526a50cee01;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'hfada2b9f0011d284b60f512d183adc2ee5e7cafa7e6e838c12bac05a4c2227c2d6bff5e9b18691997dbe95cfce00650f94f40981d4e328bf8fc42eaebbbe0e955730f62e3aa1d50ff85b26f6d8ebe046eaae0637b48039ec2c7ca6c5611b68834b132aa58321f9e6d0483cac6b6a27dba82e10cebbd7225287f2ec380fdef1bb4c95ad743113270963ded4b708172f9167b01b1adf59aea429f2498c1a58cbb2e4f4e2131857804cc14149006f718d05bd0d4440f1e27aaadea6ab38d92aa3314cfb4854afd934bf611318bd87206dc58e29c11c117076c6bcc310ea76f1d5cd564a6d06abd7145e2ef91f9b22f9e571afaae93deaddff367da3af6111a912c5c6c8ec06b08fe6448fe26d4429b70e439995967b123b9318e15b7679b092e74b6c78507fc15b76380961d8eb7e872c7979eb823548456c0180d5b80c1cfd10e2981f13e762412945b545904d22bde3484d62b76bc2733f9071c41a5f294efd4ff43f10981968a96c7c7ae56ee36dfef1385924000c27b2c1f9f4f89e767d71faa0c166388d449555d14c33c2df93f1dd4980403729a90f978d7657e7296ae67bc45422e37d542a4917ea081e5d5a33f63e7738f43a230100e4b19cdeffad8ca062425639193fef06a752df7f57fcafdb77a562d8284761e20be16c3c282d2a9f720ebf8fe2f9779025e370c1f1ca011348a4e0894dad7dcbd227452431d1406c43b8e190b79f1aebaea5c15fcad1b42abdd6b894993d3859a6221115877cf9e2f40df67d820022ddf78d40072f80e5d301b1c16141fc253939259da22767dba45157337d08ba7d03ab79ad5e5c09fcdd53f45ab82f730875be8568a547c30502d1df59cdf530a665228103a987a0e849730def737d0baf857dee7009a5f1b5d70a918144e0ef5f218a0568c2a29153e150a85d44ee299f79c4c7fd344eb835a4b92b3cff1b8d6b084fabcea6839a188750955c1d314e463621e739f817320b6cedc201656d033524a410ae137d2786b03e21eca40c9f6fe6cf4885f47cc26df872493fed527fa74ea9d84e1eb4098aac4f951786e1fd14ee62aa4f40296d449db5c763649c2df85862c487215c464c6e910977a440bc26948c8ec687b86551bfc4044747121f8190aa4bbad0286f1932380b73317059fc04c577758f6c8b1ca2e22c2a79da9a5d63ffbefefaa3a7532936fefa27b9d2cc952cdb43dc0cd2c3f6a65d4d198a81cf8345e6f7fd7bba9b93f71fd7170d47ec67b8139ce0fdd768d424efd770e7113d472c087ede01a0f8f558965844ac36f0f860bee7deb45da74b756af51a121de859e8b2160a1e2a6e4db37061ff26bf5f82e965f1bb2dd1b5d9258a57ba5fbef0a05be01ef963019ef18176b4385a393f5a2479602a365daa35f9216f03fea97ecbc43e3b7e6e0c0591a3a52525b03d9cb2b6f5da1efc0264b4c8397591795e0bea6bf6ce674a1940f5549284c5d6a2d78ae834b6f1979342b66033bae64bfdd590e7d184e26961979a17c924b52b7e7f2a3d5aa4e1da9d9dbd3851c39f7ab157ae28d09db5a8f94c09396492cd5f67f3eb9ca28bccb8d0b833f9f893673f2fcd414a9c1212163df3d88c789cb913747c9cad5522c4e6b931b4d8e6806ec99800d966a613d31c97b926105da1b4dc2596305c73c1b9df563294851427a78afca691dcd18fac750b9c7ca4866497a97cec8b4287a2eb5a1e3588e55a2009d0de04e5c4eb4186cd87f3b67e29e7f6f9f2c8a1157e9ec9a477099b699144528a6fb94d1decb92467fc80abd7047e7723dc8916a50f3e0e48e2581afee6089641ac969932ea390348bd7bf892d4d9f8dc14a80f17cbfe0e977b26cfa4ae3ce5356a7be320d6f001da7c5718748a1b5de547e7e6e4c34c7b500e849f90abc23b1240ef2b86dbedb1c1b79cd80a07977838c2949883df70d91210c64b877232d34b8d4dadab664d0868097805fd84412b1b1c58ec7eff1d742a3e13415bb9b33b3ec3d2793d4308bca1ba8635470f6b11622e9652eaa6825f332c31b1fb5b26e52fadd2848d051dadb64a0d145385694f92c09ebaae818baf93e42beafa90f12f7ba17c4c89d424514b1791e1b3d0bb8747489c95739ac37c3dd25827cca142d15df5bc68844a5fe4922bbaf6a4e64a8bcccc1706e2a4a1bbf9525a6b61346c23fbefd14e2fb685dc31863f4ccfc47ac0f1dd3fc9d0b6640f4eb39592d934b10ee34b62ba253175c1d8169ae0786fc4738a238c3a5436de8ad867044c952841f1285802188ccdabc114e8e05a9f31be2a1eaeb2381e0e365831faccc916897ecbd23e3322ca408c8e8ce70243b764d8f36cd8d941907c203a4ba7128372ee6c20228df985239877769cf711a13d964e8be830c3fffc26a816630f69041bb4249685694f771db63f99763be6e3d59f3cb9c3337ea6ed6cc574cda652fb35dfcd19c8809479e1f5a301e892d00997f33e2b96f2990d3ca4855ecaab3cb4cba07820b2f25de1413e3b685d51e0faf9ac66472b5b38156386cffb6168f445f66eed83105b2d3d7a902a006a99279e0cc1da8e1795c381e56dc4d9b77cd048171cdff17441a5bf2300e4a9ec934a3c88f965aae051482df48bbc1c1cf01129bd3057201752ed358ceb559943d626c85ea39b69e0ab02596d51b154acae122e0524c04517ff401414e08da502ee10ddd456450c87107534d063eb8bfe8610930e4d9d7c3399b8bbb14c97dc819fc2036a722285617c5f39947669a18b28c138596fa28608aaa7dbc224e8bf9090f68e48a946f86c35b9f57d09789d6ff337e94c23099ac9b277524246d6fb509d1e558e71f09a5f8e284f98f5dc73cac68a59dbcf0635abbec886c7e01f0d3af225a1bfcf0cbb08b2cc7c2dda5095fadddf30;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h6922597d89764a50e615f615d0279e80e2df5be20bd7c28753a5dadb702409739a5d78b9c6ae7aa29fa3111aa5357b34d41a73b2c98d1c389596cf621a7fde148f8ea69f572a382ec89cc10d5bff5009be62198141ffe3bbdb81cb1af4916083a530b744a67bbc0fd3411dd924b0c6a0765a67971608221dd021d026bc6d76424847ac17d78710aa15436565296863dbe673d1154c4c9ba892d0edea4f64df1046462eb145226b7bd8909ee4b6017abba978aff689c6e43a470019565f279caf65fd0cf42d60a27fcf165bf202530e27a2bd79617343677e61920749cc4feaee6938097db4cb7cc8c3ceaba96eb39d39df76f60f7713002126c15f5e2047bdcfc8a1ec6fef9c829d6ee704ef033c4375bbf11cafd22135f9009b3025afee7d0e2b81523e638bd65f580a4a655d89dbfaf6a2ad1fd6ffb84f50309acead6e1fcc47c50f3292f5acb0a216057242854ae29f8189d8ecf59cd7a68e1b33dce423783901a98cd9740baead028142f845c253a78d482cd85f618ead229f12e75afa887521ccddf36aceba608d9c4e9a76e3b0e3fb73316fb737d2d4da61295020728caaee4066a7c0c6a0ca749a3c67f50cb6a44457c8828aa3a2575fcae804e67c6d978846d951719b52f519ed57a8f8ab40ee262a7db19e9798cb9395095903335695cebff0ad545d042f9e5564b903dec359d200ca844d9e5df5a15216907a36a895d7627b604ecd3ba1e67c6724a14bd952f6e15c9c16d16f918238c48263b00f2008c81adfd4b9bf1cd02c59588c7633f682d6d0009efb9dbe6fce16320a4335a9e817d651cb7fa1733c2fad329b5e8560a71fab6eddd0aace83c0b8d75619458b7a3e613cb7dd3c82e0db969bfd4cb526feb3267109cac8d765006e821d0f778c5035b31ff8120012e1ad4f0cdb1b998c509a6576f525d2cb2fe603cccd609633e0433305cbc97e25087c82838df998fdf0fe39041053961943acb43d67a09aea317e7c4a2472918c9fccbd774660cad1df002ab936b60499350404d65d02ca6da6ced9c9602c60122949eb54e24e4fd888d739bdb3c9fae8c90993672d8ba617c443b4f7ac6777e3a970a9846f9dbeb65d4a1363e7aff2ba33823429738f6719dbd075cd09d2e29e5f3c0e40ea8a51cd0cb8eab50a942cc377fbec7ab2fa9f9acc965a45b1c2f1bf2942658c03e78e8b281c2d8af416aa1e4e7d93c7f41f6ccf25f58a0caf3a3734053198f1b341bfd26a2c63c005bceb55ec952f34566cfde99a081132d6e41627b54a71fc7ea11b4dc6fb98c3b2902bd7652cdc887863cfbbac995801ac398f3f2eeecded2d39f6cf108c36ac19a20e1ee37628c8c2460c45f7572e0f45bbe6bfd21edb76f41d7f7b90b0767f7650b88a2fd6045d97325b3ac1ae2eca3db4f30a052d777b964659f097fa2c117e91e4861c13f10079b5da29249a9c22c8b91bd1c89c014254d3fbf7cefabc2ac0eab533c601806966b349a8976fb5a162934f07c2ea92cc5a76aae93949c44c0f8d0dd32ced7c60941ba69b717ab827f2923eeb96d5489712e4a3890503d983da38b4ede42f02cb58003bcb6f9b8fbf184be38d13743c62447bedd2fbeb697206bd31086806ca5e8d8bdc1a1bd94ed08f4f548aaa8221511f137e74b3d3dec5dae271715406ab392bc0751a6785103a8d2d79f3e9181d185c490559a69cad6aa6a9f41534dfc7dc8f6fc70618e2ea8d1e33a041e190da67d0e71ec29532da6d88671660a8c6e1590c7914ac58d6a99c6e83fa920024555d08881218be62231bbbefabffc3bcbc3f39ab0e9646c07c9c2d3bd5921cda709b11a7c48e1289703a3b31311855098d3ff010fe935686c5c8d84ea2476887cd0286db30e081114dce1d4ebc4ff3cc600dcaf9ed0a4e85351217dff9d9eb54d62dd939e37ca7933fcb18e1064bcb191ba7ffaf516454c04576deaf496a46fe9c408bf62b3f2b6c9624bd752bbac8348a42e23a7ee09851bc525a53f7445685d6372d51f222e54698df5a2a24edb3776eac4bc6bac0d51f04d8dd480da82a8ec4f1b8d6d1b092ea92d381e6341caa69da22b95f29368a5bf4ad3c0055f46a3754abd69ab881a952eaec1b53bedb862c28cfc6c9072fa7e87201d9a0e6523dcbbc8b7541cdaf24319949ecec3ec73496f590e3fb9f0fbd899b4ce891c7542feb0213cb1708f593616bd9b02092ef64d34556ded16eeaf5c3fdcb6d0e132ffd4397e044700505db02969b2e7d032a89284ad87e77fe08079f013c888d57e10d06b1a637b8334d4ec6eed83b332f93d87248cab470b6b02c1c8a839f724541d07b39349d8f4ddce2a4b8b88d540d1a169f9ca07838e81e152edbc1b7096d6db6014e9e87ce3b1fdd4bc59e6b1a80a3a9a36b14345c253e753fb90a84d19049cf70cd036e6c7e283ae80111d05f780c18fbfc67ac9a7366516f26c177a0b366eeea55bcdaa08910f9ee72a2081742e9470d9518297aa04e7e47e395ace74c334d367b3ec1a9312648bfa7614cb99649ec6ae7c2497bd13f9a1edb285dcaa29e2959bd4e7d9932b4672c2a279420838b92d965bdb9ebe78d5dcfd3d67a4572c2e57fba22bc5c945e2a486222ecaf6bba37a31b437ff5efc78bb561d3c0871e9505d9e58867613cbc5614ff5abcdbd89c9e2bd7e9cbd9d913315ffae8e8470e8adcc018e55a68857093791abc92cbcb1f69fceb9135ece0051eb003b5ae1e46dd7e82c84843ff1338f4ffe6b99f7d17287a366b60739258cf09f4db51c8bc57eba200a6204b5c02f16396693f234f59a916b13dca5b6564e7daa440ee3c2229d0f75782e1fe0ecf45b9b4bd7a1eb93cb6d46506d16a58c4ddeaa2c96291a5356a313900ea05898b1873e615038ed7fab3df40054106f51a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h68a360ffee500c71c71fa0e0bfc5012adfe8c8afa8310b0bf8b8bebd8bf2b75d1ec06db0100ff9449f5432097287bf7a327f565a26d3960cc39aa3d037b6fbc2dba001799244f06ab1c49cf7b4b6e03bceb43f59579cc524fc1867d06a6253290a769eb1b2649970777d9b10f71ea1ad5c5962eff7607c92a008a494706b9a1305856df204c2b7ca8319ea61c402ff8e8a6d36e0a14b219890c8872206788f6bb226863a7b8f3b4a9f2e6bf626613750c9b7011b27d8e1ce18f5f548330ef9ccb08054f8d5708a1d03aec83047b2ba67f016aafe351954354bd434a42c26e44a754d9896cebd579bf88bb9f083217f0ba178821e645e3ac769e60cebc612d198d494655fc924d8a3a8de046a09f69a881b3de1122bd8b5df12c629220605235183202e2636d998f0a391fa4bf5d192d41abe94655b0848162801b809423b317391e2daaceeb0c6b812ffdb37d47909c1b916f53803bcae3d0528add901f585629b7e2b8d8f6ef577e96497d34937645c15fd853e131984b2bd266e9049cebd5d9bac03360c4441a8c23763264bc465796864259472d548191c1f1513e062600cef5b5d0746df6a3432b5872a39ab617c79eb2cf36de0802853310a6b1d2a18e647a3d2761b42c3d260f5fc64816ea3a0f0b5e42af99e03f6060e0926885ca06d68b93e361ff1e2fbff584e85fffbd3bf3f90a075e5900967237e03cdc04d910ced4dc69d537911d8a16b21948d85ef11568ab133bef1794248bdc1229955080bc65234793596f166cd9d5b5f6d6224bafa18374704776925a1ef5c6a6a436e5e206f0ed5bd4e7c63e22f32e8ef43a0a5fd2a4ab167f3a8b3c0d90a3116fb67b68cfd730c2ab27790c60c9a1db9603edece5c48ceb0b7236be0dc266f562db39899849b5f7fe123b0e9c0dc9efec23b6c80c43ba34e975fa7ad19d90e0cc5b219dcfdcd033df320b34a9c775c2b0377a46598bb516b2f2c9d56aafddb353c35dbb514e6ac64ff3a61691c666d421b18cfbf547a62d5100815b5bdf142e535565d1ab4cbd48025683fb5cf11f7f6fc83696d45d6c4fc45813fc221eea4cc663cbe3f82a516f17852590785a78fbd214dcece7d300cbffb8d31a95b876505af2ab731ec2722b49cfed4873173a6a0cdcb1d433ee81c23540269e495ee24d0d9c9de31ac8fc502b0e0aa04f6e7969a9ee0b38eb77aa601e4c8c61ef1c1abe9f92ce851d37944c4d83bf6d468dc91576c7a818c72123afeca7d21ed019a22ebe6006c150e7a58fc9b1d6b165addb1dc741adc08b45e6289083b71a31680194ddff523b9b7c71cce8913825c6d57cc4c80f396d6431fdc51794c03a52185fb5fddb7faf08a5b1b6886afc800f378346fb0130b9e8cd783e161bf9058be2ce4a005de334df07e87de6c98b47499372297049ebf8d078e6a3245ee52c59efaa81abdcae9863254ce5468657dddeaa02e5ab41ef184a72881434978ea1d1928e150b34166505149466ffc8ee7aaaef1d9a8d33d0b2005caa9da7c793d5709330be0b43f4ce97c77c2440cbb7a3055e796cec0493ae2406c29fb7821dfe53be5bad82129c83597d181805df3f7bc90b0d966cd935be17d69b0d909c6b5877f9b1aad431eb9d8fe8592bf3f28bf7ae926266531700db75d401c2f756eb1b6f8814774bc69bf032a30e7a8b4a8d095247bfd3135768eefea4052085903280767ad652ea84790e029e3ecc7b642e02cb029533131f6412988d2499414e8efa8801eb157885a7ecf004a00e52f471a8ef61de71af9f1b0ea2b427be1615e13f92405c17974579017012508543d8c0bcf3f4c9f602661451366cdf0b3c6ea278809f904651c0c944b8250c27077ddf37c4578ceacee70ea6b03724bf6d8b099eae4596840586ddaca5096a476a21333e27ad9c74eef5046f7c1b006ee722e7782d7dfdf7fddd67757026653b777494c394ccd8a8b873e729d6e63bddbca50b80d1e8af4dbfea86d4523ad5537a025834af4e26fde9816a0021ae7d78c5cbd302ec7e353f4bae8e80cfb65216e2bbb4e76fab85b8b9cdc8df7901ef89ba0bb1fc251d1484b65f163ba1347e237936ff8fca798b322240afcdd6bcf886fb84ca7afb875463c27c742d23768bc91df0c170fba30a4d71fca45e0a7559d0f74bbc22eb9f62aaa477cf9253749d543bf02bb0b56bf082ad243d87ac363f96d634a84787ef2eb600be84f416090606d30c88110e2a9b1745bd1d7a5e9d3cadf84d3b01611b6fb188d53a8c48fbe824400435acb3ce3ca3914f3c4c2c6e010cc93d0ea1a9bce94a1c92d4021940fa18222275ca7394e9d13fe2c300a57807c22e360f1e551b7a62a4799fe5435c82ab26986d4a317dec5365aeaa5919cdf1231b082b4a44f5a26a8ddc17566ce29c03ad3ca319cebfa95377d8c6aac5dba8fad424a2555e5692e501bf9ff5861d2457253f8932eaf73a1097bc41ff5abea4587db39a28fff5e04bd71c1a5e844722e8c678d74769c0c6740584ba3e8627fd938f867f4d2b095f539bb51836580a7323f524340f5aed5a3b8ef0ea7a4a973e832a4feddd45f7d2179e8da63ef566ba5e13586533acc244ef0f008f999a7ec9e027978e1f73ab987afc152fa94037b504f215bd5eb0ff0853de0695d769b59e51cd92f73ae1578924df86cb6aff12e68b5514d86d8c1673290643a2a0a54e627167a010b3634056ef05427907a515181e38d68be81e7e51ccbc14ccae545a3359c7a8ee19ffbabe6a451341bc41b3058ef7a5870ac18e610dcafa214244f09b9d7a15b97e023db7f7d7d5eae8e454cf2760af72a7afe82f5a6ca7bb3bda62303873bc73edd2ec4b695f5ae80db61dca40939517d5113e832a7bd710cc93942cb2fd838abf8decff23b91e33f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'hd7ef7e416e444626897063180b7a2e5ac3879973105e5466869ba5cd4b6e65cc36386210e785cb8034bb7cfbcd53d3b86e861e7e63d14445265658186a88257bb22165925e41500762b0392eaa22d1df78380b27eb70ea5902e5d52700d0467e0b33932a6625e5062c7ed6d1887190922ff6ac9298200d8eec2ba38453c248711c3988e953511082f45a91a50e9b2643bd2ff1bd7252a3df2d91b568ab074b314318db9af6007916485ded78046d5a5107320b8bbf7fdc982f8a8084bbe78297f73fe3cf70fea0a88accb9fb64ad88e7a697fae1ef9cc5e9c6705fcc6d3bdac829174589fa97dd2b349f34b23d4b0146b13d03dcf78e13455dd783b05e82a5deb966e37963940dc08fa94ab6881d41ffc5b74a350e7885178f014e56a8d8d25ae1dd0ca2cc6ace689d6cb010046472f51e3fba5b71b0c521dd9d99df38461d1537f33e4b2f3c17955bd2b7c7bf741a1f501317220b91fb1fdcf1678184142fe91cb3c636bc6d19e2130623346a5e4cfac2e61be11b3fd37edd837ed037a3edcef76bf5d442b886b5a75b616d8a4ba0745d9032935ddc57d9c563ea413e0828781d235b85295e4b2e76a56d7d1570b4d559f0f0f79bd443ccb243ee76821e2d39768229b0bdd78c84dad122bad384645f683ad341e6b6f7365e01f1006022ae8212845326e623657eaa18c27814bc5ca7b14c07bb2fe2d5d4beef22dae19ee1d2b0e3b7472fae181abaa98fd98f96dccdfda6e9fa96d290c09e6476472dbda5210ee06ea17d87d2ef04e8143a55e624410676a05ff62fcde6709d7caef43c3c621630fc3c7c82479db8a6a41d982eef389533624eafd915e223aa845f587d0131035d774734b516cfc851830b23e7a4224ed250d9be0ca3e184444755050abb97df695a1dd57d55df60e0f5961eddc2a5d29c3f97f2a787f06d50548e25d58a958bd4e15c5f2e6c9a8598330d020df64a5634743977f15503037dcec01e7087bc429592a3c3fd0586531dd21d7acce0606cf4c590e4a9fd1501420b1e6f2feef729fc00f78469bc6d3640369d313d50149fbce31a084faea6c650337079951a463207f9fad0e68685c349c35978533789ea91d535a502a08244af058fefc1a51e636d5f0612a755481c439d2322d87eba7cbb9664edc209516161016c37dcb649a9b34ae70dc64ba30f0864393d1588c6a87ad781a735d704af9ea8af2da672024fe28a3d46964b2586efdf909a534343c852adb0902cee30dd947adcaa39a5e5e4ff43c54d595c830122fa60f12a4a5eaca1dbf521c59959779505e5a66826c25e92809c2505d11284856a2aa504436aeadfc79be1b0e975f4c969e1b080af6e4fd07dd883495d404a74f5cda5b4f0ef9b7975b8b5966e08fc8220d335291a81ad438cc27ef26aaf418b39d8a5b7e07b987db0694d05e175cae56c2e5b8364d845e9997927324fd8a99af720eb0011af7f5825ff5832d4c154d13dc46175d9ba5ac532cedb87ab34ab0edd45799f4d9151a4d4227bf4ac0111f57244a2a0661213ef2b8bc473b0241b979c2d41bcfca2ffafeb7519e3b85dbb04dd41dc82cb12e25f70742e48e5ccfddcc27812d9d931f7c183a14002a87d9ce48b56821becc15fde56e57fbd12033b2a960d3652873529048bcc7fd4f9790acfb72ad10832d7f7037d02ab0b227e11bc528e3e004e31ad587a3fda2cce06a9421493d288a9cb0adb21d5d646a3890cdaf9458cb02563223af5edfa36100b697b17374a2dbad48d74020c10a09093ae25fb8400767001ca62ca8f64fe34971bfdc3072e6e7b9133b90cb7406ac7aa970e949d483ef2920d2c2e848654f8cc58dcccea7ed95786d2fb54becc7eec5c24ddf730ccfd034641c47dba615bc104296cf9441f93e13375d34a94f439ba4f92736528780ae90f6815f953ce455342a7312b8c0d2303ad07b1a577ef1063327d042c5e73415db73af024702d43ec26a07670936c8b3eea664a0e9f04458e1f235b5315a4728f6472d1db212f43c3f9c3a6e481539e0233b49c57f9d901269ab7b5fde17c4dfcc98a6a96822c8dfdf8984826c1bbf29b82d181d360e7073c19da6eb97d2e0d24dee720cfd2e433d1235ffd41fa394f7767237730bd3d378eb1a3d53e19d45ff7264caaea97dfbc24609738f54b3dbe4b07c54158cb0d1724df3931951015209acf8827291b3877db540ddbd1a3d596ee478bfb1169e56d03d5064ceaee7a7b2a916d82de33a1970d2ef0e415f7fb3b600979c3d55006ff484e93ed7f6071da5c5b1a1e4c2dd5836e423bf2cba8f13022909d05ad778c0cca1a9c6d3dd6be58c6d73ab523ce3ffeb505f44aa2a0146de4400fbaa1d9badbe580a674a8dd39b7da6529ba859c76b2e91f448a604f33bff81dcebd7e066eca4241bb43d762a5af8e3eec114604166451a12340485717e8766144e597f9c2247ea768d65fd993b4982f555307e14dffa65e3731c6f4519987ee76cdad8de771634f4f430406b1642131d8308e12b7fc8ac0f5facfdce4d250fe5c38c7b8a3d0798bb2b7c22629e4be9fa4524c3f3899411583267a9fa5b1d77754979b7bf5934643e281c03c178b618b52311442f3d2a7694c028d374882a1595a95bbbcc1aa9b84ba2e830aa23c93ad98a3f3baa819f9b43d9459b4d81f6bf8e5c36a284f6f263d9901882e1e21fb94fecf2807fa007bc95484de81cec2ca77cfbd6e10863177fe9b8f33f967b18f04f858edddad4831bcaec84034dedcedd1713fcdb16a10e87f254fe26b05a51056e418ea8b1255169cff45ef2730f1de2e0f2e452cde3bbc1aa7892f3df6952efdf6b45b42f11336d7e4179760fd6fd12ea6468cdfacc5e2652dce29a3e0a6d3f9ddfa5bd44de77b25ca492573b8f0782;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h1b799d4c96a138892e46cfdfc93af2cfadaa4bbf5423b03b120887b4645ead2c1a2847b8a8c4b42ae1f5f0cfdf1d029279c00ba199dcc681044270a0460e413e21d7ce74ef90174e6920e9c4b71be2607f72f3b879b35e0a0f258a8fd754ddfd3575e9d22048122e7781d9c43196dc34f8ddd12e47238278fe1e786b47c18ce113795c2f7b44c1455a74c5e06cdaeb2a1c3d78cd58607e632899e0d2248e4a678e776db762f71c170faf05837515c1c382090951c23d906f385f604eac1902232e69da8c8e3fe5ad685e7a31dbcb57b97a1917780a940090d844b50b1fe43b0383a1bda66496ddd81dbd08588361d393cf279062f00bc1a7af1d427d4e412d1ec4fb02cf5dcedc6159c17ed93909ee05918619211bcc323248efc2bff732f2a8b97659c4180fa0edc88ab9c1e26150801edb1949b7d79072c2b0b2b48e81cfcffac1bfffcc1653f7e18f92cc3b7e852b32318dbdf0624ec305890f1186c6692d03643d4b3fe66942f208064ecdd73f6cbac60484adfcc149b60f920298d764b41fac8baeb8b7c436284b13efc203be2ffd69158c68b13436bfb40820c7a005b268b835dd4b17a9c6c81834e5a3931b19cb3ee0c78cb92ea843f870988abc42066d22914e804baf31222491e83f0dcae197d2ce24e8476aa3ce32e5525cd614f7f8a1021223c0ae4be10278f459007f5f44167fda192d0477428a37af462805df33a2c1b969bb8788a75484fb9a50a29976b94317ee2f0c8ceb78969d9abed47af5147dc14164f3ffb9a91386cb132f236a66adfb297b53d17594b1846e1626801eb69bf563b34e5e11952eb5bc18d9b012a64f7ba1e8cccb01b0c50860084aee88e068fa3572cfd14c93aec5ce0c9178b3c560bc80654a8a9dad6697e0da40c09a7a22b0df3b8cf57c86f37698dee8ccaf5f474b64a530b174324e43cf12afbeca282c4f05e51a2064c00232be268f1fe3e3fb2dbc129b977df0d835ddec54ff97c9eb53d2e893027b3195f64b940bdfc6f1255f3e28ee932a9a54f2001eae54c7f41ef3e3b03b2d6e35b4fe51042917cb97018637fb26f8994139fb09b91014fce0071178511adf47ceb90632fa6b944090df955ea39422056e22810c0643b8ac6654e21e647c6e85c552c3ebc6d2f36731827b16e9f2fcd4b70ebcf8a8c7ba427bdc197046e6a7b874c4bed49751af9cb4d8a444aeda528c90300fb8dbb3b0d7e83733829766d4caea84005f8570ea75fa61f44c5ad193b79b772324d79c02b0a9402babb0af873a2a0a6f073f40835c7837db1beab1547f0c9ad4e07c886af8f5cd4b074bbae73fd117fb494f9d1c37d00b12b5e84a3dc8c7404397d9eaa0a4fd5f05ba871dce3689256e91e5a793ddc0bdd7c54297c718160fb55ecd5255b43e6159b0dd24cc7ab702ee970b868345a4d1274ccd177652cb19c6f254d9240bdd054779baeb8c661671decc5859aa8112065bd7b6f4d4d4c15a60089d8e3d0fe8d641c82b9b8fb5fae38a88aa2ca5d25d4f4d8706671c80c8e2a2adc82020d393ae22306ef9d9ca3d890053cd289e8a1cf233e7adfcea834f65d5a97ddb05f346e88c328469220ecc41d3f671eaa5a5728577da224c6ba99a2afe66602720d0b7307749f53d4377886fa25578d69f89f76deed85837e699f95c5206a032d7e996ff5b0cf5d885d772511030d699bf859a90e136474026cf1899bc58557f327acf0296d039bcb89493b0ee19b002b45382ccb398cd1fbe23a61f01c3926d00ef8cc6346064421f9d4681cab5b33cdbe0e935f694bc549dbf02859f9e4649b5e2579a5a277f5b14be66e940a14bea1e64574213208e98da675eaa7ec3f9b79e674795f77e73b7fdc8ad07ce00fbded73f0a29c3f2da4f9bfe87cc88ad54216572e96a1b53594f847778c6af4c2dfae970c57ae90f4df7ec27f5c4a88bbc6527b3e982f1c0ce942bff118b468f3dc535ffe11b3085aa8da7c1132ed93b83b72ea9f0e2d8800f4d2ecb26071d2635f53a59a755dca9cff5e52e468030ec65ffda073b3b4c41d3f065e3d8b0f16302d032266af9825942dd89d6ed1efd7ab33f0abfe0dc7f6621e353f3ab81f7dc51d3f8f03505ee21bf8bb6abb1642aeaf5c2854c520e37ec8f9c5f1b40d52a78b80b22bf319b878a06938311e5d32c1e34bd356a5338113a24bf3efd5b5abed7aa35fc61c6b1ffd2596d33972945f823a8b9a00a2be774866f78309327d7c2a37192cc286b5462b899eae31357f2710c9c9e530f9a1d99d865a7e25418f5c8d15a215d4876838e38e3514a7da4d1bc5826e465a877b898ed539a4564fa1059748429c3f30253754986a8146489adb8f77e7cc2e0c2fcb219d9499f6277c66afc9163fba007cee8a160977f42dde424e8bd798d56d8d047543d47f714e803beabf2aeeca0ac31dea423d6f02b998e81e6471fefb7fdd4309cd99c6ee6dece83dcd6fb14638fdfd54bc7c659b2f7b9032a29f1c9f845382c7ce18934ecde4d3b20aa683cdd23afb84840a6e3d26bc46bda4910a12bdc4031caba7205c2d02a092744660865c8e72650c3d1eafd39a738e735b9c5cf934abbe6d6f5b1c792589e784f6877cc7c5ce4bbe144da1454475d3ba1949fb2aa8d2fa2abfc8efe7b077a7a54b66b77c464b0d99d06137ceb92a895c50608422dc5a67496aee96752b5ba3f67e3e535f75b395708a51748451fdf021eef00fe9faef57222261c0819f54139b1add310b213a5b8965146ce65544b460e6c63d44c4f59176009789544128abba54fe20328570fa00230b7191b5e4f651a91ab37595a9323fe002bb783842ee78825a0a27028fdb731974f3b347495cb703df2b52545fd0027ba5e4d231fb85084aae3164cbc491d2dfef741dad49b5f1fdb77;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'hf4d62ab1cd87164853c7a4f8438e37a0e7b0b2b50fc89689060d4e0b645a31fadfb73b57b3b5ddf598c6230e1cfdf3578a688fba5aa4c14fc92b9078be136c58122be08f132823b3da7cbd435f293e1eae871a97525bfd4bd665e096dac2662e3968af24c2d25006648dd8c79c361cbd5412c2e8080c317eaf80edcbd4432445910c02de8b14bfdb908c445ab6ca40aca45586330f744dd673754eab3f20558aa9fd6fd16f9c5a2366b62b0c595d46fd68035675c2a09d1bb106269468c445566de035a90ed198a91b381bb0c4f9ccc8081c7c896deb878399277a4f2f173c02502d8cc02639bfb4ce1869d0bdda3b1552f778ecb99eac6e48ec0d97e8433b4129bef5fed00e916f5cde60a877409ca16e760caf89b46d0d37768761b53a30ffbb5f4eebc089d0a20d8b28b52bbc827cfacdf727359e3a59f67f123f9ba38ef6273aacb9046b586a88e5ad01792cfa591780e2e84c69b7b37f2a959c511322ac3d32d4bfb68d09b30892724ef9594be74c2141dbf7ed52d43c48f5969e32c00c00f652d5022fd7d941b105b46f520facc6e8156a6ac7296ef0e76de6c8fba7f01f9dfe01a026cef644a40a8fb56e13dc6ec0dc615a1def312dbff0f6cb99f5397585e52b2b170b4b824d6e9674c556420313894627c0470211b7ee7e00550c2693205da9e89036d3a9b7d816e834d2f1eb27189c1bce077f39aa8b497f045ba4826247661e2de5e732551be9d7f6a1d322d10f53dd9bdc0f16073d2b6d99db264d13d2aa56b391b4500b8c6ccb65a1eac2e450592284401fe5f6dca6b3e52cd908a26672a8cf3c3490414b6cd603c4ac5016aedb848a3e742f2b4edd0929e6099927aefafc53627a539b6ad8e7c47ca04983cb4ad407b549d3552688b7a6878c6e26dead72ccde90906d98d6746f7b061ccffb031d2531c7d0bb870b3e816faacb539408686f4c05c1c21763fe95513c746d99dfad69350673a423b77fedaf948a234c757c909c58ace00e022c87c97433feb9f4460601f51f0659496c6a443c7029cf4063d7722fb9366b9d6388825a51a5f8985fe839d11161d282e2fafc99b19d3f917ccd2fb090f81b5e65ccb7ad0d91a4989aa110a8b70dfb8e432d8d01eb8eab180bdffbaa0d8d48f9ed6ff53532bb1f9e204d6b5b13eef13df3f3243bbeea94f8a7f0e9249931c3949dd7d0c022c485c3a9cc6635eee1fdf4bc216277118a31d8fed20423a64f1cafeb1c5e0f1663c1fd7d08b73d74ab53e62eb4ab2d145e6992281152051d7eaa352b06d24a93545ab3134010b53606586475c7626ae9e0372f3fa48c3028c83266bc314c6df252b04c9d394a2a2a341e76d47b85bdf5e881f33b8f5fdebd82e3c98ceb63d8ccedab528a174741cc22b696afeb0686333d1c5c607ff78082bee233bd959760d55458b6aea04234eef9be6022303620012e0c3a56ac2315de00d0c178d55064918872c10bfc979a9a2ee398c0c3767b099ad57a3ce2f154c5b55ff6335ee40e6a85c06ea22ce2a92bb1eb16976272c84005efa4075c7a366fbfda73a46262fa104b2dcbbe0509071c27d3fe66ca479d5eb1a86d6767ec94b22dd350224dbae49b268a5ee9b8b522627701c306f34c7e0bb56ab5376b1f7d7472f4ac5d8b8300042cae719e28e9e4a590a902fc5bd1fbf3bfc7c2c6adef9c25089cb515b0426783f78cb6bb4e62eb63a0b526adc0146f8c0323f228d2ccaa91cb32e6921f9e1c014195e715fc959e79d0d799a7b2216135b0da2e17839ec3a01571c2811205c673a97d3c3284cc952cb46e6e5be4622ea240973c34f31533eb936ea6c4f38cfabee46ed52ba1230d2676ff42161aa4683bb7829fd9cc8867d821deb55369ffb845b1cba83bbbe906783dd69ccf2abff007dafc662c1a10fb35efd3fcd0c24b03a161688b06bfb5590455e65f1847a22fcb6347363b7cf391b0ba6a3178acda4af9050d7cf80c60f2fb6555f4a89c0979095c27788197936de4bff4fe541ce08531d29c5354b71067034d0fb9eb218b6af6f8bf5d637121c32baa75694d965fb2f1a01c4c929675f352851a42830ef62a23a3060da6085eee442f78ac72eac5c438859889a6bb72e1e523d19c6e8ea6e015e18ab6628eca00ec20a1a78f0a8f83f344070034ff5453bd0db2c28754b14d49aea2266bbc70b7e4300284d8e19709dff2a99be7bf1f42be27a317ddf9458e939d40a64b6e214bb11b0a96219108365b1dbfa317535cba981f28669f9e24e4f4edeeab1016ee1f20e29b55fdaab909081303f0df40c9ad41b218c9f1fea8e1928a77357e5f2ed3129b7c767be79d0a81bcb4a490cc570273048141823eb9facac66e4c618197b61f01a46c5e5791431c8ef081008e060e8761877b49ff6b91c6d2799413523227a686c68c3d9fd581d4b52c2af61c78ef3dde177d1e0dfb8eaa13614e312622d89be3785e70409c9a0e8b754e7745d72a55d04fb4379df0a799044f2c804b5e4453fdd5a75884ffc385ce9152c8ad6f0567c7594375f1db9fbf3211a42d5940916c871c7635bffd945813106c2483f9211a9115e6b7f977fbfb6297edaf2efeace5203c7828f7f091de06ec59ed8fd795918daf651b610e625913bfb33fa815bfcef8faa7d39e1508b9d691801bb4686fb31a9c33e8a951eb0a5f587abb032388e36758ccb99c10a5f9a4b51c4e2c62eff4d4eb8ba777f80e39f94ff6afdf813e3bf912e3c918956c59d5c2275422364960a4cfa79ed4eed317a4b184b21b35799f2d5e482e8d623437a913e3ce0d6a8a8bd5f718c8775a539a890dd7a3a457e87fa1ff37f9502342441565c0290618088f008a038687a82b648ba3b1183b6e656858d7601f1df3074091390562eb3ba272843dead4aebddc;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h227a4c10038a881fc638f2cb64b41528de861c7d6adf3c6ceff5418a7b919d3b3e48e80d04e4ea1bcf43f6a5ec9ce19f93a9e9b5ea6c591f51ca88db40ff41f62ca651e1c75db7ec4d6d7eb7b8cf30e3b6dfc49255705a729a9fffeecd47ce7bcd066d9454d944496131e30ce80b55a3bc78b4ad6f6bba915bd65cdca41511423a749f5f604d1c0a8d36e6d080574fe97736ec1f5d11e7840b0c2c9bae2d45bfc9f25db8e0d4030a07000a8bb34d63ec0f78de82ea6e48f7f4d1b75f379f46fc7b891942488ec93c08eb5fd1ab2c64340de2b41ca526bdae160551ea4626f50fcf7607643bcc24914ab8126e4f99275f74c8ba659db14e50e0215821a679b52100a8aef3064a9f1b57d1ecd78af11a0bf106d13ae652e5d307d0a0168d5ef746a2bcece6162649c051d7a6fc522ffe8fbfeadefa343ec94fa0da0f69196aeece8838a6552df7f83ee510be032fe9215447e5c9e41ec47f2bf8ff6e0633b96c1244eeff99dbac5073c944e3ca45da860febaa1c0da0edba701936718d55175beb8fe8a0d367ea85b52cc73c979f7a6123986bcdc6a60ab0d9e13a09348937146d418c3014e8048a4eed6acb5826390f04727eb70bb0066a8b9b562ea9d563f05470c2e28c8efbf9936588fd1a74ae92942b12bfc285de1bcc904b4fc9b9df9dc759cd21f237ca52c2ee149de98ee5d068a76d4e66de6b0df60d39588e08bf73949201453754d94fd7deea3d3856ee67aa63fd54e31a1ef09b019e9920fe6c54925151d28129337b18d9e53d0f3a37210f2b29a30f743329a97104ff024523674a822df6698375e2dad2fe233a6f870864232c4edba8e5c37c52fc7fac8792f6faeafc82e6489a520fa8e4c775c1faabe4c3184d940ae411b28e3cbbbe934850200f1c36ecddd039c5779aa0f88f3214b8a96f700e1fbd45196f7441b30130acd747049339fdd52c499d45a54e6fc5948d5dae6844e19b27b4530155834fc3220988cccc0f6740febcd243bf8f92d98c01b61e201a4d733b1d0d79015ec490bae1629c1d21a0f360bbf23d662b0ba7c5da6fa4543c96126fa536a7b31c882daf733808ecc8c67cfa571243a3d790dadc1ea25499f9c2958d14a900f89bd60db116e460bb9f365294228ce6ee33f2692d155add260e53f4a04ecb80686364a60b7ae062444bad304c6cd099a6ad61d514bb1d905be99a79209161b42cae6926e68bf84211ab445c5d6786c708d4ce91b6b1536b061fc563d15ae20a60a9a086c9a13a13569ee4db86e2008ae6d565a43122cb1b0c145117eeec7f5927dde334401a86640b729ba6f8df8b806f8fa8751c4b2a079e3373d99d737f2c0b81ab01f72b5b793c241d5beadceba10ae7ea149f5599496e523db92cfda3e0de1eab6fc009d0f5edcddb01e0f3132874149bffccff3825af56d6ee82c544feb8922001934df9a53a7bad8c693af0300d9484c4439710285d4adabbd59e41e9d5451b091daecfa172be36d04b03f938df18503569cbc8bf1eb821c21eeb25bfb16780f59ab7b68009249a75ddaa953cbe704a36a943d1ee83164c416569572a12e440d76877579c174e54dcb344a852a11c37055ce3f9dca4902c8ced8d47ec5e842afddaa1135a0bafd50ea608aaca2c2326a238172fc5748fece0bd6c5d94336ca0a54e065523c82ca6d7b21265d0d85f6e9dd0aa83c80aa810b30f808ab59c0d724a6e3391ec8167b281348e905b261e19cc5dc5586bae8abe3c89faa2784ff8bc9bb08bd7e2fac431b527e334e1f6c47dd6fef8c760e925c44ff4b51905cd9f8802c5aa1fa16b1460e7aa619db65d2ef7d6b5bfd5f0349006503b13538e06728d609b21a9ebd0f28836094e938a25610552064c8e5b48a626c45aa7b0bf72aee34391933d3f9ee8dacee5bd6d98b795803448d7fe2e40afb114ff3f37ac0e141047bf226d1898311dba4a062c6e8bd96f7f5fecde7866aa1b2c06856f3bfdb3600676964ce435ec4011ece18daf682bdd7740574ab34d956c144f83053363cac539c60fc4835fcd864d99e9205175b67a022a534c41a9fa131f8338f3d7a17854642ddba0c2e1d7edd4b6073c5428d9580c778e0e56f7c4dcff1ac2263bf99dc293a01de4169661d8407e923d5debbba898417f213bdb825b94d5275f38ea62d42b2e9c46dd62900ab2b373e8bbf604011f6c58cc6a876ac11cee823aa65c6dc4aa3bf848f1d8f287ffbb3d7dd4d464c6c244f332eccc193f80d7167ad71a2f99712717a1c8d35bbacae933eba3c8fe4438261d634cfc97be18d1fcf11ac12b8f3ee3c36d56e1a51696d9d1e9601a63be3573b84e4db5223449c360fc963acd416548b7d31de8ea5c399a171614a2e1b983ebcd525c70597621d37f137eba38680405272acbbbc771729cd5296c0bb7669ba6974bbf5b162c4efd38d85282ca1e331f5fd51226ff2cae418a6cd9647fb9e7c502ab20b70ad33545d9d3e040b8f289da8ea54c5576ea48a2aeb54ac96b013b94134017a04bad650dccbc50f00b0df33dee0da54e5a0bd186bde24c87aef8cc53e9bf370fcd027629ebf19991da413fc01ee82f46b28b0a7b294f2959afdea96b2df5ffe99fdfd0b9ec14b01c5d5d085076683014b0572c2016a1ae13f1b7570eb0ad5082f1975e6e8f40772c49391f21a60460ed83abf0bdc9adfc1388ec113dc1e856893e1e8bfb846c8fdd253a9d05b0c445608db2279c369497c343701252ee669328c900d57ad660d91826a45b580c4f39c1c13324ffebb097eb2efebfbf93a565418f650c9b3b22aa14fdd47b8857e5fd4984fc33ceacb519627aa29b57eb5dc3800b4bcd35e310614bb3d9ccfcda5805dca09fbf837b2fa1e9bc1b58e7b06a04398a4c03cf21790e32a94b72fa1a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h1116bee5e03266e8542c95fc5a59c8b97682e3846398e963794fc8c7816a8c557d56b44d3537749685e1aa0c3b4a7b36a47dc4f867b28d0b2fd98cef07ee652c10d073167c370b1471440b72848891412ecd9c727078b5965a75ce93eeab9e488f73ce7d5d618f75017f12f6184e9680cd87d4a0003c485a9eaa1e9355a66975a90c166bfc9b0b1a9f6745d8b917c4d8f0056bb4556699b1b55c8c54ea3ffe08b24bc24662876f4bf931237cf3fe7544d913a362af7216ebca02b8c2058c75de1a9392528198e1f3d46fab5f16b59af508475e36f5ecc311500c1df7c73308226b4b48b2e2988f425c4b4c3ae093bc4f06ae52f8ca9c51ea50af29c829a059b1f85c4f0fb245ca015ff05426681ef245d8010b03cf26c5c836404bed25589e835c2edcff683c180d0cc3ddc53f86d432c162d77feaee30baf050a7bd459cb30c4f8cd72b1781c606606406e66b7e64fa282282fee3e1223e24b2bce3233866826a32893d446e982673e1de6e6038828455eb7c5f493b0df1c1fc4e1f301f50def4566911ae23a1ef2444e031edf9b44c397d2df5c0a5b571721e6f9cb03df719d02d6a2a9ffb781bc376008fb624bc6b532ed34da1d96bd584b09ddd37dc599943354c997510d4c5ae93f5be8e2d68d1deda2e989e2ddea0bcd4d25d531b27a5b35a65a872b8eb5bf10876ed5104e69db94b5d5e5a1ea10785826533b3cfa4c44332b9a7db1d5c7914c73690d528f42fb2a9abca21bb79d5036b2a34905bedff25162ec4b999c9952375628a1520a3d793903a15be03225cefd983c4b9112cd6958bada61cac00ea69288403e7805dc6373ba16bffab2f66e8cfe1b34fcd3b089402eeccae82127b4f96c25d4e8b9c72d5725278b6a91c0d422f78d885152d5c301a5af65fb1fec7ac60054257fc1a51a230b7521b5023751231002cbf88bfe01403534f1de343befb8b8e8df823a587685fd98d81cb76939771a5b0245961c9fbf6a7d3d61d58075668708036c3fc39d1fecf5c7d1786fadc5c91e27c30e88fcefb79d0acddb5f18641f48b580ad9045f43477a0bfb45c765d2f6afc84fab5cea8599f297b0ca32907b5a13af9cf47451418892ff9f746367a4114b112e7cfbe664068f23de3de2ff5466c09625beae741b648f6f7637f3db2756fd64a633f85ce814d54ec35ee8c26527944a2b4ca50ff41983052ca7bb95c95fd310a3d81f73c38c05f6c2b7f07ea379bb6a0c02df4e88ec6943c1e32cd597fb74ad4058786a07047c3230068878c5c88e1cf4295499273bbbbf0e486b9e95a8d8426ec987481bbda7b7f6977c22a436ed14373064f09b50a632bc1e162e9a9dbf6ada3623528ca7b9639c8c76a602c8613f789c8ca55468fbcbc117028258e4a4c274931bbb60ceb6e7afe0120a39443a96dcb0ac3094c33a83fdbdc1ad22ea1bcdd628ceaa3b97adf4788cbbf54598e747b06aa0b66819928733f1d1390bcf96609cae5bfe163af6e0e97b7f51967a6f22eaa961e4cc20f83e219991b17bda4316bef642eac4630db2ed52a95803890f4d8e80bf3b1055b2aac00354daff72978c49c9adf6a5ff759e846f27508c8fbfc37b38961f7293f5efcb283c5af58aa6a7aa764447e41b4545e92425e32d7e8b26beeb177d2295119de12826dee4aa949193e15237992638ca8051221978721d064677fec73964b58eb4ce5a673b8777a9cce43abbac3c44bd5c55561ee84ecf6311c8b07a9cfbabc57c9fdcef6bda465e63e8aa1f3e2652a21533f434da7b279843d60b493e156575a1fca1dd963356bf2f65949d39194a8698bac72d436097a38db4cf917948d072bd05df1d036fe0b1e44a308caccde40f5bde7388593416637676525517636519034b59e2845b21e689c34c2f144aad98db9d9c92a228ee9cf80d5ceb013189be73133e397f73a52fd0f64a0277c590299c6e4bcd3073aa91d5bc2adf167545c2d1fb1ca6aa1caf3fdeb4e1d83348ca68a7412b769c33820ef022ad94049e4af3e9d56d7b51370335c1d657f218560c184dca2e2f3e8b02b7253d5e34f6fde031038f05ad37740fb65de3becff59338492b860ac992243424a0745b1d2409c8f14a430b41f405a2ad9e9c9eb45c3fd991147f9d69e97ff1c6dc99a40a3aa206f62bc4e7af595899d1109704fc01ba64c5191d3f5d22a2dfa539ee649ddc8336b7f70f3405fab17d23b8ead2ab7235f836e49097f6b705977142b0a13d1578bbfee00b49cb1f773b22b4f16022278a6f9a2585ba7a0c56837022920a7aab26f14f575dcf2c48db7906fb5f58d6fd992369728981ffc7afbb69b02f5d215cb49febca8b46c84fec1a13aed5baeeaca1d5b6d1157a28e2b4bd444bf70db2f7fe4290e9df80d1378e8614c8c9f9c018413a9b216ca036bfe7abdadf69d3e0055bfdb0083531c3bd570cc5db6bfa827164aca9772ffb3543c60148294085eee962cf6790139aefce0e18de9849887c70812a1ab0c3fc5a184ab51f7732756f496a2474552c7d53441a3109f22e02ddc3828f1231d2d3d1dc793099c7aad2fc07e50e65ccc2922e8e90388f23042ef626f1100eff91f23e38a78b17733b2d16a22f8a1e5f21f996f931e0d9ba1a86937834bcea2977a6da0bd321463db776661107beed71950e1fdec1fe204e7ef5a20759d1a8a938997842b331282455b12fa13a5721692f599a16e3e2c80b5f8be4eb8940f7e22dc819a67b57723abaf7cd8a27eb8f997f9aa184bed0b9bd282239b3da639259c96354c230a4e9501427e4f3581cecf9c614ed0db0eb2c5ddd84fd8d81bb4c6af5423e4996204c63b4ce13bda2836a1a43140e970ae84ce53d7631cbf465695249639dee2f1e60ce2bd831cc49e71ee249a3d60efc3fba76ff27;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h295b17cfe320b7550a9a78e7f5fc1a3a65e2bc981473fd14f699c07c12ff138b61bbd9d31160473464550149f11ddbc1195fb0559ccae146500057391a86153ba412edb49385397df18b0187aa8ff85e57b4812d15b27cecc060df8091ddbf21df88c484456c27589399ec25a63742587b6069a195aa16510c9d33f58ab4eedd8699c4b11c46997f1ac8efa65138db0dc8261d52e5eeb42bf3e4e51f55990f151ae72486f88703218171d65f28aac86fcb6c4b0973fd13267c91b6a83d06d8fe320bd6a9bbbb4e87d25ad59baa9d62093e5cbb99a0573dd2c93a030e7a956dfc5bb19c43b67835d65943ff2041762a282352b1ff51d4c77b166ca616a6159c62d367a133ea9fbcd5ce16085543f9c5cb2db5727f02cbb6fea5c9df344f508c6213adc2982405b8f5cc1b48f7db51d171c3039f4ecb37cca9722de59c0c1adeed93c3d6fb26cce7916dca187f1bd5c8cde9edad4dcfb6c7e8951de8d9c9f264e18c812fd925e00152d92fe6eeadce712620f3c0dab4a0004b5de68d2667c62a825622cf29a0ae19e832d8edc89b583e1d30bc5cf5e17734c6a4c393ea9b514b5889c89cfd6dfe503feb74bcc77b991a4b6e2f8d63c9f68a673b02604b6b199879a36b1e5e691935455d29a742a02767e53accbf31e5a244391d094e6a0d0469cab3270d1c860840ad46af8b931321e0083ef26db9e54207d1679649937c10e2e3dad8406d8b5fcdb19360613cf135ef65fc7bd605decb62631c839757e061ddee5311208c053f413c56fe48f683ef54d9c0c35b84d10bcacab07b73b9c1bd2a7226e9030da824788dd9e9545233fd519136dd5da61b733abd70c32ed808ef6d973997fac3314b43c6433619944c55ba2af9a3e0d6e9feafefc918db917416efc6caabdbd9db3d1072cc0bdae80ef22c2207e2b813cb631ecbe3d27fca76776e22a0c55094b038805bd004f53465d70728d96901915d2454a97bd333a78da5d406f24945ba7ef0733eea1b88ab9d30da8864d4fe45185eaa88c8927535cede2b199fbc4c0adfd7ed925279a94312d3ed0e1e498cc89957262f9913e1b6b0edbec049e5b4e9369b264d65e12095c1b0cb8b349f7998016bc7f948b5643e11926f4c3eb82cba731a34da386631b4a9bf6a75cf4aadfa7bf58d6aababb54fd798068a2631c1ef543fe01c21e11258071b065aa30bc8ed0d7578a8a831952fdffbb66d39439f3c474ec81b9fcdbfe289b5875415d4ee56bb3932b6793db2038fc46783b6283027a8c3a2d2bb1555a546929b4ccc005a634d80074214f9d3b218c29d1454a4c9456b3fa202a68baac3dee3d0b1a0a25f7cd32f55a86c5cda2b1f374811ceda6ce5dbab581c348ef030028007b0a60a088cb2e03d28886e68390ee893a33d90ba5ff514496d2cfc6474a451a3ccf1d3b6c3bcb2b46f5ca7d3c5920a0659c47754a9e0ecce98ab0a155c68132f8ae825d4e70b9e1e91e046a4f230885c1d4c7fa5dc0f6dd0664162762420957293180fb3bea3f3ca19f192634570bcb468ed2e877a462617de5c3311a007da5b347e2fddae38642d257b2fca30fe2a8829904d8aca20750332e782c560fe06ca3729dc5abe7614bb5bd36e9d4d67f9946ba191a2249287026102dfd329796987cf28cc2dee460e2f4402dd0342d14aee049ca5fca8dd4b010cbc83e4c084197c06f045b6e423bdcfa97bfbd2f1e54f1890ea5637bb0c647adbaa6b38ad97fcf4d9c187b66d416b6377f64af1c597ccf9ca00b10a698878c4285096867a2d292b62e5d1210612528e3ac7bc1470c5c16515dbc1bfc035cebee10fb62f09a2244f32fec4da134f5a7fd656afffcce39f82fbd6a9bfe6b8768478f04cebae981e2d98b640a50ba68fafca195a57db3525d92149606625c683a5477ffc11ae9b06d30da83ea1d1c91ac53902a39e0fee6cb9cf865da6fb6f6ca08a40bcf439515a8f7d40805881e5b7e98c0250b954533cada1315e056b5471d32af562c5a3b0b6e0f3f395c089504a4cfbd7f7a8ddc9e2f3d3c18cadd2f848e732e1fd33f0eadeb52f4d5c6367b6a8cc1d6731081bbd6d1ffcec19ebc39b567b3d712c85497003d7976d2108d12706ddb8595f8fe2252ae600b427a887cc68cebf204c7fb8b30098c5052808e02f7ea9b6d2284d57762521fb67d05d00d6148077d4a5fdef5db3205172f31ab774d1604959d28263c91025e86daededf3b92eca8feb3f4a8b3b52b1568434eda5fc4d7e36af6012342380f8b261bde42e1da777117b90ae630d24a980bc62824724953a8c891208f0e5257c4bf120b4e3cb53950be61e519bf62b6a227e37c8439ca53c0256464ebd2bdb514debd35223d54cb93ed7f57d61461b5dd53c0bd362a5e33ed6983298eaa7bd2922ed6392c8fc26665f96602f0b0809afaf3d5a7f0cf5459f652aba5489ba3a788fe3870d4affcff4fc858a1def7b10e1fd66750659ce97651ef6d09b7c059341a250760eb4079edb3b434a96fb86823269fb4fd41605f33e8bd832dcb3b67bbb393790e214a260dd5f5cbbbccd0d5ad1199c46a64168706751ebaed5a360da60a56b60c3e8d6300307496e599c76afa82780760dac3193061923cf890f2c4875ffc2572ccf8e82b0f76ca0af30f89f23a3aa378559b7c552f3e9e30ff115f1b0b0f8466b9a1164f020a4b2380675f6dc7f40018329f9a5d6855cf81bc78c5c5a0f6452b59ecde47bc5cad505b16a94a76447ffda17766362c002eefa5c468c0dcae8075af80616eb2d434fb97ba7712386926ce48933d7a54053122166d1c89b6a6746ef81588ff4ef90a13f3dbcb42a40e8604564c128e1aa348d86cec7be630df88bfcba2f19e275fe6f4374e40c5886e946c9487b89bfc1017f6a4a7d63ce8;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h68421d2f75f9c90fe111fa2901f8a0f74248c91c893bc8fb66ab7a6003dd171bcc79a0f630b87fcb8d353179602d83f07e1d613e1f59ec0ca9267a2c0c611845ff12eba0152eb3aa47c68b2eb3cc477b997109234a342d09abbf54c4680a86f3655257862b2b700ebc7d9a5a6f7b4d4ca1d556c0ed77c1205bba648eb0d573c45a4b93337f763f3c4d20b896623743371e91858bc2e5d01b02261d9f8ac4d021a6811ae0be5c7fdc09bfa788c08c6b59472f87199e2e72c44d06c5be5f4d9b62615c05706c4a87cd38d3ab672bf31a1a211504e62e28586fc166d90d2e192b07cc2e10ee172e0abe363ed5101bb1e2fad699d368756ab53a46b846451fdc6105496a4e78a9f492544e01fa767a7a1c814e399ee038ee9810adfedd69e0513a15d2401352842177afeaab80f63376fb20cb2a33e82ef8f45f82d7ef78403b4d3ccc83537347c04898089d7252bc9c3417f75e8e5f1722094fa90b0b0e10c2c5545de8dc027540934bca6e10c57c4247cbfaa93eca7fd92757834e303493d3f4897bd58626b6158d31505f17acae158d44d8495e7792f6b446d3e3ac6c8680649d94b82a305c4db56e88a2faf6986871cacb34a79a4902114d634ecf19de824c64d376bc9284231567f17458498ee756adeb1633d7ac4af76c4aaf246264f83fc4410f15f65a6ae0db24e02f0c4e86e0c01e1064dcd6bed674419b5ac767cb5f332426204802005fc8233b40fd237be268f836d048a90188dc90b548214f99b60c140741de65138d5f019555dba715b7c3ae414b59d3da1d302a8fa588695c0b64be66eb261cb630a6b51776ec9e5f8320918e1ebc4594f1994cea8efb1667054ae084196fc72c38cfab3e904602b234d34f6aa7aac92186c00058da7bf5700a0f825cca83e35a683e30d76903653f1a5912b8eeb703051bacbf76917c9b7155b7da1e72e421ed75867ab2e57a4c449e1aa777d45e32eb8fb07518d0094952df834e4cff903248d0425f2a2093c0937446edcf7548c0c91a0276dfa4da93583fb7f09b1ad8413605f4551808d2b22b42455cf9ca9bf1f111e223c8a42cba49874801ede17cf74bc3c82f7bc26e23751005042eab4a6c5f53890dc458d2f6edf9e1a57defe50438f9a33476f73fa34b1077755e45d55a6cfdcd7990a36f4e631450e1d39047ede20dfcd21a42f2612ff4e37b1498b9e1e6e50069a19947675212e9e07f765fa6d3db188effc7c234bd357ae1f16e05d985ecdf45e0fe832879aad6e1eb8a14c5a9a1eaa356823607a6e41a17301d22fc15472ada26614161fc19f5728328e3969d7e2c048a5c264878b82b85dfb25e6303cf5ee4ff2edae2735270ec5ec7e43ade4e9071621805130ce51cf4e279a3874141eb9690e01f2ae87e3742968eb5c3fb0bd1034cb7c39b7148bc6b5eef6892f51bdc0cb71c0fd9b7c37599c7bbd4b8e351cb90daa483f5855ed3dcbfbf80593335090f9b8557c5e2df0a74480a879a4cb7cdec70bab55f5085e0b91775916222bbf5d311783d4d22f576bbec17a2f31828e60826a0701e10eec19191d11a2a6827b09840a8e8a3daa820f931caafe65dd4f66ae95dbb228d90106877343efe6f5216029287d8f12102156489de6575f354fba4f1c37739ca657021d0e763993f3b2de6f7f82a0a1aaaf7557d8c96c0373cea21b959e07a1aabc5de2291b13fd90c512ee9fdfd00198a8aa5c89b87759543852acb1e7412592ef5ad6572c5a773aee16dac1827258d7f5d283ef7f27bb1883f9a3099b01a618760398c28a5b937589973d780694f394538bbd2b2d832495b6131fb8541e714f2cdfed8dfb4982df9414579fc9fddbbda1b5e59b4eae510ad4e320da90469d2a23bede3c845173599ec38d29049a873824a5b7b7e46fd512086318f30d2565c8fb77002c39fe6dccf7cafcb775efc1106efd599946c1be57c41867805f55a72d96f23a8fa39e91ebe0c5405fe0f9f72283d10677406e1571c5e810b7bbb0aaad33c263c8429550fd3500d49631f989fd22bca45d78568792715b6dde49590ea4d74b55bd5014abea405458fbd71a5e2db9d717b11bd13a9635a9cf70b6fe023f288005732336a819ed38bee2094fef47f2d70fbd2cc7bbb4dd8e5f0ff5d986d51e4f4bae4bc3656a9f48f86664950d95b3157043192f4da70c5cc873909cb1f9f03197f33544afe05d1b766cd6d518f8165e395eb20ab57896f81d1dac86b5da809e03056e0f39a041c15bab17b5f3cb40c9cb26634835900f41e9279d575bb156fe4bb6674f8570925e6ff0bf45a6dd4ef1b72a566f80b14881e23c7032047271c2264658bc3c755acb1d4195cad3a6b1bfc782949d7ed411f50e60fc08064d3909c9bcc54299b8cc1adb2aa9c85ce2fe9ba4f9257a9aeb3cef9d12af86d205b50b06743a1bd3d610f179d9690af7fdafb45f8623c543e38bd7f0ea1957e68e0a6c70b94344adcec5b9014f5e46e7cb291988084446d83821ecb650fe41fc38543a224d762111fe15584a2a046175da0795ef25844d88e99554d119db12668073b030b627680eb8da778262849ce4fcd5c2d88ade2b3e64b5e0a03d03c9c8e00ba4211ca6c051213bf776f4b4ffcfcdb9d07c326723d1ae1fa1d389d92b0fb29648eb4b3f41e4a4a51c3d6eaf8188d220510d537e1c0fec7fb987766a4d9c72ef1aa45ece22d136b85c0677ae9f8c30f88b89be7c2dd9ac915a8b6e22ed6327502d3a30fc12ec77226fb1bdec93ed45e52b87a78194c275834b65240d37868881540bc731df825c9ae0277a53ba9ded7ff4f0c1eb5a5f709d14a2d9dc10a58872874db5ee6e3e385fbbcd1354133802c7d55bb1bd374e130054522872941258b614d7b49a001249ddbeaf5c2285c0248e8;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h2a1df6762a21f2088834320fd3477882c43788849c47c519ef016e975f3391195f4bc1d306e0397c68e3248c212eaf2f7f86be1684380cbcd07b68d68f90e98f06d96a0e94435f7550cdaa2a78e1caa3a53699a3a89481ff40067108c2e7ee56b5e4eae6fd0ea4334a943ae64a33b4394b46ef66919ea93696a0c18c9247ee16cc73ab7ea6736493f67936211b4ca3e6f888868a19ce907530cb6402a0115859c1d3afdf125f301939c76425ca2deb0745321074d615358e7028577f748a32c454babccddbc43acda3a799f142fffe7f40e5e9e304461c7981d96062c77a4f86e340ebe55e31655367e8c8c33bb8e4198054dcf2f229a7e8304713b82b87e3afeaa78aa321125bdd2d413b74c2d8021bbf16e45494032460730ff0df651ac3ba8be50c59efce2baa0e6140fc9649c5630ffb193b42458b745e241bb0150032d2d9c73c216b8f40500728e0b59725ece63183e1a6cab4037c5658d0e09fa937f203244f7eedfec1bd11abb04ab7d9069d97a412f04b024d3e3474ebf4efeb259604bea5910b5073c40a4fef0db1065f71cf3ed68151b85f6d7d760f1e2c84127415a9694d109549dad45a1657256336551cebe2928d22364673f82033a3d06a3d88b18586535a1295a58c130c71c24b8fe8b5eb67eba2c76e3aa631ef439bc5f690dbada128252cb06c3955d8f0cb8d2839d81929678fd34c691be35c4bf337d58fade8656478ce591d8e64bf3f1f88f3d7da221e9ba72095a56bb6f0a8995b33951afe58d6156d524b8fa899f574a3e951e427f0403d837bdcac3a9145670d9ab407702779d5c574e8c5a8497724c05c2eabe4e93ba4202965c5fd0ed0ca0b3ab90c1124643cf07b1c08267bed0316ec0cf9cc44bdaf06d049cba7d4c12c2feb559d53bf9c64837e3486dae66df5c39b52e165f88d619b57a138cdafe4afad3ecb53b17b2ec80faad96dfff3be28b9ca679bc400e38eb02d58325e74ad8dba6bb2a524e50f2048a8c2855c1147ea93aea286e4bc135cabe6d69c8ba900b773debfcf11f41a1e89a18b52619fc91916f7e6fa74303a1612ed9cd2ff02fa04759ad606c6effa5f5d13121622e73b3d295ef6dabd67820751479eb663a97ac4488d52b84dfd9bf204891e4ac1be90c10ac51baab14a08a5456880da0a8b15d4cbf886c9bd4b8a44aa553f7e7990acb53f7254740362dd406fbcb2177d0823036725c9299cbd357c5701d9368328c7df144d685a44ddb88a2016fa301c82e546130730ab75a54e6231afd6791236a772ce48a6cb9dd0c6eb8116ae1011690d0f58894836dac646dbd1a185e1d412eab46788b7e83ac3bfc1dede8cb3cf288f6c497f2c4cf2182c6f327f801bcf401d3114adc7892deea244f268fd64412fa36d10ec9c798156a8be0d44b3edd3131e3aa25e1505e10dca62ad7487d9bcc7937ecb7ebae8b821ae2fbac2a2ce521e74ce3a04e78910b40700b0a96bf7e4cdfd2eb73ee3b3a438d17c8189bc49c778ca2cb380ac1f5e69edc410023127450eb7b0a4992e06f93c79aec66f719d1c8c602a30d61120671deab6fbbf2cf2f5880bc4d179171cdca414a31470abeba05470719839b6c19e1a6db805ef1e710ed518caf2be9bee4e959d2e86e3bb8d93e1ae408cfdba644e2bfe9a8c0a7a65a3158d885256aa9a9177bcb99da65a705578f9a66076e7e789191b4e3e01807686705248659de334d0c6074baa79b9103fd0b6eb914c2c6a248dacb75b11267e3b3dab279a9eecaf67df92fd84a902fe442131b426cb606bc13c91595fabc141bb64456d53d39104eead60ae274aa6aa17edd20cae78c1d9b2825dc7d77f09464b23b6a6eedd6ca58e7e8cd96d4bc94eecb3389f1f1e693cea27eaffaedeef8bd4b95d393d985563a93cc80c99b24c5d91015a179a120076e63a780f3192f9995490ffd4a30e4dadc0d4694510e0e0da78f1a9ff2d453ea349542d3f3a31e068b14c7499b0b266137e38dd446f9fa5205767ece4f74c797590253f7f0ebae3b9b60970f63cbbb27c0fcc367161f22675e455fb06cbc2a0c79ea914f52106d4c58a9b95f9dc364e972fe16b49f53e86900fde2c01447e69ba7fe304ad14c158a32884dadc41a7929d0277a4c6d590665513366845ea6e43339201fa9e841d60dffdfda3563a727ebda74779ef7337eb17dcd2cabc1b022708d33a64f9735c5279ce6868d1d341b74a903fde8d757dcdd1f974b5f200e6f3f84d0d25a5227017bbc81774e7031f9819bb18c84c10f3ad094dccde49216037afece5703f379548e8756d4e03cf31e463e32817847ced9c7d5794c5fe7f3a1ca5e077c8eeedd48d7e4d14a9d07bf41974e51dc4e0431b3b165884411b29cb2c488cd03e60b8898dd59394af4610e3a0e6214787b4796e58c0eed2ca673b6cd569a1b01555358eb55ddc0b060a71f5a881d19d75fac069367598330022a2f69f2aecbc36343cd437723bf380e14a51e16f907ab994da202cf80eb75c871f76ac0efaa77ba8f278763772b2ce1dfe4f6407af9ba36c9e0beee6f7bf48eacc824dbcf0f359f574d0ca33fb385c35e43e3be7fb45cc59f6bd94a6c00ff3efa62fb626fce28445447e86ff388fa58414ad2f2ec1dc5b3397610f84cee905aa992fc87c54cbc4ed43b2314aad76d1250cb0bf4b2d295e2146ad629132135ddc30593840d27dc365adf228c384ecae1163d9a0ccd2f82404889292666da46e568ace16d02186b7918978ada106cebf348432f693498d8c8a98c83a8dad663a95aa863d22bed66565ff83432475d91ccf390d6b1802c3ecb47a237b23fdcd31f2615c8c16e80ba3dcdbbc65b14b894a7e2997fda25998189502d4eae56e4f9122a071998dbc38b1301e4049062b3992b99213;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h9e8bef3cc5f98088d8f9d1ed9c730868d191687d9f026d7f5acb82436736cd40d9559b6642733d35cc4446c711a36000ff7fd3b83c9aacf5d39c063a40be832b72968ec038f73161f65b3911dd7db2a2a39e34ff4d3d9f712efda0d096d11e3137cee2140f406fb14fe9b2e36875e00ec8eb2067914ac02788067ceced43d310667348ddeca2b92e4167526b22b0cb3be08e26996eadb5ba45bd1ab366063c393572de528e0086d9e7e340533f5c9d141ebf4ea5c748dc249c2eba446f3795f87a07ef60e00d8d8c3658a417419bb02816454f0a6904d442a0e05c7018ab67d53454aff3c290d3d89db83e6e23c259f0eec2a7a73af2dd67eb241d5ed9fd2dcfd5a2263af9b1ee5bafb864ea72268d1ffa2aa67448584f0eca0b3725105e38dc8bf3e91fff4a8f226f7732d22a9d6bc86b7445b61b634e3df1abe2bfc163752d9e7ae486d796ceee1a50564d06c2d4a8c7a5af3957f258e34c94987406ef7e836da1e7c4e5d6e3ea3220ddb750e289c0058a9af24e89ffc04fd6858ed92415bb69881a4327d2b0fb28a9a0cd0d8e0f7ab8bf8a3c7b6090f379f838f66ddcef6491773b1628e463ee051edac3b861f0aed18cba8c992f47320e9d988454acce265a02b7e0fa48b1c9c21d01b9692d4ac6d9c40e7e7bdb51eaec63ddbddc93dc14fac323ce87466f42215b978a6b2a18d98eb29b77135ea0514d22c30b94a7bb9be47cddb1250ed567f67773b650bdb3f92260c9e72c2bf15e5a9a4b898a8a81056ae51dc390f52a11eb43c4d7651b8af7816f84c25cde7b3b81fce4d5cb89ba6f7e935bb04a2bfb205acd1a1f5504e8c1ea07fcf64cb5ed2fe730ad5bf90edfcca9e98b5bd3987966ab8a6ad62cfd9e054e2f2fbaf7df4c61e32ae8b095d1c8ce554246e6f7de67172fc5ced4f7f9d43578ca43024ba589456642bd06215df1b69834c6a97ba296b8d7f657a9222f4095c1c0ac5ed20b689b6f2ed26b9b04d017b469e78b43aca412f413cdd123667a112ea9ccd619b4fe1dd217c63ff059017118145d610e1cb0f6d1ab95d2fee52fa59a1544c34f4338e5249af6f10ceb8511ee374a1c722210d187694281a9ff46931278c3d31387f6e854236c0f80131bf869754e54c625e50a67208ce8750993c714cf221d2ec431e442fa88e13ae0e236e6c6bdea961bc7422a3b7fcde1b37526c2999df5b22fdcdd39cac9caf31d029d6a30deafe32c7a889a448b4fd0019f7075e90184d122950fd8ca5cffa3bff4f50cc55fa1ea2df0850a3494bbcca9983471855f9886d676e55b60e732397947cfc5f781ff88598484780210904c90d01142f89ca90ee71c8fdc27af07ce50ad73afa1984c5dfae3a326b4cdd7dd193da80df00aa26e6747000d84dd797aaf917a80ae86a92409f85259a0f6634c9a0ead8d466abf8c6650ebe018ace980a7382dd93b7dd287965348c453caa1c748c4e0b4513eb5f4af3b341d93cb8b8c753ff67ab034d898574f60735f6bfb7cc3d5881971f8d0a2c15112afc35aeb49781b9baff3a3238ac882d93f6667289e03f32dfa59bc07f2ddc60cfbcd716d628a5a5d255e1d45915197cb8c016bf89e59612c9f71ad686831ac5e1d0b6ef2cb014408d8476936c7ea8409d2c9682fde5944d78748a692f477636afd4febf942f1c3c712368dbf9622f25950c6f083adf0b0e1a0be400d8dd322d8ba2b6035050a1440aff6ef2344551679dfd45492d47b5a796a91db98d2c772bd23cb4a44ed57b3b3fdbfe5fae34104b0e356be6809b5debda7a35f4dd1ab235e513509883009643696c58985793c8a5e7edb51c3c6b4f0d7a1580b72b5e4eed61287c419f0e608ab5eaca5e504d07af83cbd10929a00fb0167ebcb1a6c2251549557ba166e48332cb69a5ed25967b6852161af22d6a34abef98a08e48db0dfa771851fb794253621ffae0ef100044125be84677df40defe85c4995d25ffaf8e8a9b7e0e8a51401363ded85523e4adf8adc8381f82952f318f15e2297ea81380e8f681369bce0730836fdd211ee55cebd8d158bbd4eb7da794c198ffd56871856b143969bf8e4b323cad740aed5ab9495878dfa8385c06e999f674a949bc817e3b3f94f3d81b351298caf3b77b2b3abd95e18da885421ba4a0fe69cc32c0972eadb72849af5536740d58e699ea5a21ba9c496274fba8fa8dd07086205b4ffb4435477bbf4d9caf3e021a7bff404357ca8f7448b970bc2023f0f51337bb382e59d62895454677a9e371e30b835634e77f0316388df21c5712935516c0b489c80c93b8c7c020986b2730d224284a1199299697a23e674e461173715cf79b131a45bda50969bd46ceeea56cd01781042a245fbd46c7ea5977bffff07813162d615bd8c9db5268337b10ab9afa1a79b57950b691b97e3b467eba6ec27449f26924e991e239bdbaa227fe214a08171becebd6b809828760661e00142eae0cbce8e7e05b64b9bdb4845797448914770017ddb94ca6a30f56d1bf249c7a688b61dfed369f7fe4f5eb3230c66d7b453ba8d2e5e930e0bb1de6f1170a1c539c97ae3d9bfea2247169dc5aecebdde278c9012baf6064e591f61a19a687479c6826a734326f183f72f7b4de3c6b3b660987850a932f95641d001420681772f82df839872627192c7f03aee2d2378f6b998cc1f1e8277c5cc88ed40b84700978abaf1b112c65049ba34273647146ea76cc0168822ced20a2c77e986fe429d4b153d7f4458c8c6f3dbd5a4db6108c144e679ca8414195aea4ad84aba952a6b070dc0dd321922d3cc38f2b14a860066ccea2254cf811457ad624767caf0e576cb92d4b1c26dd061038ded59692da8958a149975e185ad1be45f4c03e81ccda878a7fe32493b3a86a49d8bd091c4a000;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'hbc89069e343a71ba257e7bb01359e0a84e640150a2d67521149007145e8c59fe971d5cbbe22a3d38416dc42abf2dd6701e1873f2b13e7be74361d25f46bdfe4aaf23e86f42222e3c211e6f230192339f4cf0ea13f944f7a17cead80ec81b2931fc330bff4745a23cdbef05361db5c3e6a97c574fa2fac3d48111fde1227f3808fa0638bddee859237f7b8ddd1d243c84e564299ee3c0522641e8bc241a6c1a5c97b6402566e4f6a0536c36dbc9f1453a2d2aee6b2b009fe79ed451b926f65ba2d953fdff98baa8835049b5aa0b80ed4f0fca7d1ee31beea97824c84168be37876e54648af82c106f3b0857668857fb40a8ddcdc8689b3e672513d958a08518fdc7c9436d14402e81c51e837c71bf497bf0931bb1c6f4490a8678394fa5a91fbe646540fa5427feb102d03a705559a3661d5786c81a11992b89ed0172a6c3966459dc6b04b48f0e7c8806bd9acf20ebdc2e939634bfb95d0b516f97f8509700b8a0f718b4501c6f024f5ff71e5c82f52df70f4742202c72f3a1b7470fb92451bfc7d507e4fa9bccb2628d5a4c0780692f98505d287a20847923307bab7d19eb0957284500219bc6a51ce3bf37b5732d576d9a0406b754d477d3ef15e03d93f392100cbc52aaa3135fd10c7316177f10607588e4f7a96a7cd6ec328c9097707f834868d06c1656f6f92afe09d314a36a54652b5ee02bf55aa8a93ab50197c5bdd37b11c2c8acd01d66ca77da2aa58ca603a78f7cb7922eb02611cf083da6de1e2c847af3d97162e12d57fd2da896738f8763285485037781e754db653a96cfa0a1662e3458c204177073166e2649c041e1450fbf02df0f516a5400f277ec5bb6e30f9c54dd881e189c0c58bee17e31199e7625422f9e6976ba956623c10bb5739479320cf98707c403a8d10775b7a4e8b344b9e9004a6356f968032f948266de07e2bbb2c4a7c9f0452d0fc077da3281e01e44872e0572ce85dc5a051ed88a651202b0530728e566465f88ccc2911180478937727d6c1e58c11f05f6adc369cc0bb2db021868f6c7136c44550707af0968f622b070db515cb394bcd859797a4b7b872ee8a41ff625426d83daf0f222a56f6974cdaef38736d1e3632ae079c3a9fe803808e3905836bca1b2d6bb48dd46b37c3250851b9d32884ca4b9cd3c66d71a8efc77f95e3c246fe15544c296b4bd39c2627f5897f117c1be56022270e0c4c907af77a3d4c210b6e6b6f2c391e9115efcb734db5c9d52094ff0b268a11a48e328cdfce4bbbdf219faf793ab3bbfa419bd4114d9f83ca52be818114a2d0ccf2fc02e76b3b2112be437df8d031415e9d9407f8d10a84298e2bfc067efaf8b74f0816311f0c8662dfba736baf8b8af124783015271f123b36cc45ac878b01f113de400c54d9fe7dd8a218811e73a4562e5cd35db8be21711c5b245720c96e651289332001923e9a60cfbfa41b97e10c18a9172d739aa880af03e11e023e8d060753da9cdd40b51e2cec22c4ee65d823a537209c9c9fc74d826a301e846b587446b92e9e3288a3c5cd305be0fb4880314211892f6613ed1e56c4f81104968a76b433b863d2a24b9c6abcbca9b881129ca9af15003a533c15f32a02085cb39a026f6c7886e6d79656ac7485cd51363a5a26a472522e735d41cad536924231e9c4a2c873422fc44a780bd3646a8795b0eaf9219a542138281bf87c16e983d2ee01666d68bb8254c6e8245ca3ad7d4b86409fea8d6fa274c7efafef71b8a2034d48814e94297dea73102003500902fa92f165c89e24d01c215078df7f09aeb8461b031118ff66f82b59108f08125695a801e7c1aefad1e8832dff93b5c2d7c0617110a46021d14cbb461b0801c23768519ba6834cc46f996c37c5cc89cf43765a8d7cc91224c024de91a4ac154336155a720664969faf8d828c1927e7612c99c6aef897c3ba881c5f1a1148d8cb2a37dc6161ae11070e747edf19f13ed498dbc62fedfd8f9c0217eabe51f1552bae7a332a637c052a5b78dd06e3e338f9fccf271ae35279cdbd76df58e2123b9919d648adee50834e5c3375e2fc6dda3cbdf5b3d8f3d604d119584909aebcbaaaf339c8b2e39a55117cec6a62b70dd1baedbb94abc3f8e2a14b9ce60430062f66ab06e94f5e40e44bdcf0bb6f631c9379b0083675ecb995be0040e9248cf6b09318ae7e00acc12456dfd3e55131e8bd4414f5013cfabdca7160a33406b4c235f91a5358b5fd66a808ab1f1bf3587450ef5eafe069b92ab957ef8914629930da9f1632030a1edbf051ee41d3de8dd9e3ae233320e8fa702b2ece7cb1ea05491544db351c6dab9c23a91eb61801ce838c507f831223ddfbabe24dcd8052470c607ede26d5a09237f22e7625af5729016ac5c6a0ca959041ec41414bc5575fc4217225a55e54800da87b94febb5fdb942e49b3aa00e55abb2b4e789088ec2d4a2090b1d5e2eb21aa09e0c3fd0f17c83e6bb4e967f393a52cdd8e78116e04bb731296b6b442aa55de6a1dae366623fb4275efe4ee3aaf75ba6d1c748e0bb817b65b1c201e29a6ed9f2a33e96f2f9ee08457ad895753ea30b30849285cb3240ce54fa38f02d7cc8c28fe95d59180d52a8f8d7b86e481beb126929d416f8b6b0e8fe97a24978687e2d6e96a624624aeda4250b78e38e4ffa29cea8648b70b140a64ac8f8ccae1d352c355cc70d5f820260cfdabb0489972f227f04ba0c5d7c50e24ab6189cfa7b6266a00f8d65b57df93db9324c666c487e226d0375682c404b146f3fd38f7ef503b1e8115a4b1f7873d894598f1981010385f63b2c96fe130f8c9c806125e4ed370dce0b91eec022aa40c7d19ec79d695b965bcf6c3f8a0a2c1a9a3534edb9b4b80fa275f78e73891585355a36861ae6156c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'hf82adef8dacb24b3796304bc50e028048076e24d31d982ad3010a2c087deb496bb9bc22b8ceb465e428f2d8308b1483e599cd752f5bc862fc4afe5a27a1e79c88ed929dd387ae459a464bb5e61459ef92df29326c95b80cd384564905423bba7ef90b92b962fcb0f1c780b0224629df0543900479b4ace5198a2a6f1b79c5361744170b697f649cad4ff158b67407c9414ee56e8e030299bc222dde0ad5d3fb6b543cceb647225e670fb6dd969593a83cf9922beba3ca7c7c62797ee2c541049bc20641b637b928f2dd9a9f367c7cef5b572552a52397d612a8a10671a1bb3e09a000636a1a6df4df5089384d64a968c2b8cc3da0c936aafe4288c18e8bc217ecdd73dc086955b017666f3c1c2f5c525524892f8f46399078d01bc7e5a1a6b236f5ab464f4eb108be807348c32f2f360b9d0e0723a1a7c3b8cb78040cc3918883539a43cd38c9d2c0ab959431a5b67452810ee47da2e3e556483cea3e8879d092522db5957ac321919485d9f984278b0deb946c4a488a28d96188c4b648168072914346cf55a8e22750f6ccb19d17619f99253c9a5fea3649da0d5a23ae25b639b5e7875f4caf2714f008e3b08d79d848c83c7af57076782c5778d5ea285b2549b4470a1d6831a88f1208334528264eb145a4aff9bf37ca1c8515bd008c2cb258f4c2222246ad65392a74805a6f683762f6d69f9b60809dc79015235db3ad86e49d96237cf4b1a6eaf7703022736979d69f28c716d04c4d5e0ff27ae13a14943605c010be49dcd4b1b5638a2a570ac7882c120620386d4b4c930ea60db6a26e47667f571c10dc4656a344f78b948532f45268cca0335af3fdb53bd7c59780654731256f5c61f76ef674d165b285708c90418933e91aeb6852db36a6d5987947e0718d7b8c0a7d368b884b6ffc4ce817ab462c38d211e00772e50c6d714d97a9f6e943cb5428e00747d8582e0663b41378e77619578a0272da86c39245e7eb6a2194ac4ebbad73982e166e8f970619d5c44d343aaf3182d4b0feeae8872f632b4abbac074d74089eda9baf10e5e4e1957c1ea6d4bd2a9ed0b787e70f9c8aa31f943ea8b0530590082c39d4ae8c77f2b2bdb7e0a76b461409e35f8396308c5f4f6596ab917c5199e0ecacd7bf71584c92f9e146886f65dae227fd8fd5a2c167860681d1255324abb5b8840e9de03dcd8308aeefc32e7c000f42905c421bf058fa682116a4ee5f9aace2a045c043f749d1a0f9cb3ec8f4f623bbd699bad118025f95389b464fbb9e1932a034ed70e6ae7bddfcd7b80dcaa8c7c5e9782eaa2ace97439064ff1b96124c9920c77a28d16806ba47ef35c944ca29e6d561eb69e6519da8b6fdf454e495285194a947ab6417d101a49a4ef8ff3d493dcebb4d9283db8a6348e5da967c017456e473da8dc901ec80389ec263b2b1fe0e197558ff1aaf79bd1f9767ebb402260b4af81e05eb03261f18d234c9e3591b9c128db8e86a948ad113b1d22ebeb91db11027ff05c776c3065e5e1fc26f3273e78f84ddcffbd0413e5ee6328caae40002ddb6286de8ff116684b91f08502eeec22ec104662d17e903fa9fed76a0190a27db80fb0c293072221b867f58b6a2f6b8045e005f4dd815628e972e51ceb21157e130835eddafe10e28145baef7aea76dadbc7aac0cb45826d97b84df3a46210eb3d2d0a5a99830cbf88ca56d6c35e67653576cf2376c9307dfcfb82ab133c0a79d48bd54710813158af8b7a164d5c416dd9a058c86c45975d1f3c71bd31e4cdca5f4889f09283b37fbc914dd0384afa9060ce2750d59c2aeb6e5d30237b84b5f9942acef1d2771badd4770383f9eb02ba49ca0b235c9ccdd43bd8f00a2ed3cfcecdcdf137c9ba0e30baf87f4ecac5fb4275ea26832cf795f7a7249d76d1db7fcde9bf068b3fcc99e2ecf37ac6b9c35a21ff9f4d9a0378a9b518dfb25d5c995ce0c57e427f844229c4823935ab14d88d5acf0dd57433d8690c4e885c633ae9553fb0ee8125ad2d649655710bea50b058acfa208282e8ccc886c8c5a34670c125882354655a6fbfae8094501ebc641d6ff5860a3a58a8a9188af27821263153ca32c9cc1c2a9a6180515ae61e2576fa77dd759ec7afefd921a84dde286c6cf7278389635ce6fe07907d4c868a91acfd4bdd27cefae5e3a9dd4108e387e0b96df266563803a48fbb6881f15659b5c6429a53ec385b94577b824211024c386ec2e81981fc4d459faff01e3f7d4d01808a14385c6eb02ac5ea0b439b04a0956e884e70bbda5a20af5ab8f554f774bdc4251878c92c240ae1cf8a3f69ead337d5a7ad8030738e1252d43a01446970f3f334fcb98e3eeceff49d92163ebb76758026539fbac73a02e68bf8c61ff023a538f775b960647d360cdff4454fb6cf7925498a061212543eff88403950b0b138d04712250d66a80e9cda7de86d40e378abd3b3715196dcdabe74b575c843451a053ac71e74307c7b897925c42e3a6f289f134ad7469d771aca08a47f883a46fb2e13989c00e1626943fef529f14bc6c72e995ea65003ff9920acfd1222233278debc4132bcf926214db495d8ed67a0ec5b2cee4774ac1d15848e61e3f0a5f540a148574a220f287ef2ac3c34495108223412f6b201dc7663fcca14754fd839a887ccb238b0beb8be00ee2cea477a26f6f3a1be9f7ecede23ee2dafd16399ddfbe86d37f0e0af02e0f41897f4c596f1e7a0e8f692e33d50d1833c06853842d3d63977fa1ee98979859b23c43202b744b9219780b4a2d93baf639a4ccccaa9029696fb4f5e64eff627e9d4a95f8b7f77c17b047e5bc29fae513d823274f1e46528bb40d032ee5432b03190cd904eac92dcc35731ee4a6bcd294999d1054e68d2b6a73dbedf00b6fbe33219ea;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h43f52bcdd21b0af0f8afb586f002c40545aacad986ae54a4acc81f6d55a10d7ae7974400d3fd01da9fa8c45e5bc3d9be67dd5ec8f8c1e3a23f92fdf500c32295a6c046aa0ebd136307f9b8f216a1cc3c44f0133608ad5dc59c25d2627a38edf2faa4b0d3db4f5dc639300b0fbcda124c1c3e9bb75122ae503aa3eb48a3eb020f1aa514fd040359913991a63a250e15e4c25b023a7d7a284905f81530172d70b3f643e7c7a04490697a711b3ef80f2739bfed62d6a8331d48e04d037ce1e5f64d89e2c4201d5d3a446e91738f8d042297c026a3a9acbd6b9f7e5ef5e851fdf572f82e9f2a948e722594b2d1b3368c4691fbe7d85ecb36dac9650aaf10b9fb7ca963596b09697a9b7dd50b55547bad032900f030a1b006101da20ac91ccbd77e6607fdd172e0e01c97703c8afe436d56e85602b70298fa19ecc6e1b46a0ee2475f8e36d320ce457adaef32884b52f8188eb4c53af7efafabdd5109030973263f2ef88970f253aacfd9fe3377e3565b47962f96dc3727173e5f42cfc4c481936b2594b661784bd59583224058709ece08c8840f5f1bd2ef5441e0d4f5fe8fbcead7ecd488fa49a5977d136443617fe8b6f183e99bca5b8223add1a46c3bda1b3e09a31ce9060d7b59ec8403f283a27affc9b62edc175d0b88fa53ebc45d2fe72c33a31dd97c9bc5d604aceb32235b418c7d6e1287b4fdeb4781ccb867545b7318ee5a03b3e519eac265c180b9873298f72e72f5da6f964138ca490e5439030b49f2112dea878c16b4d5d040d0ed19aaf24767145823473437578dd09835a8b67c736011f8b3bd3f3878643b39d86fa7c02d850c235648bf4d4c01051d5a7049bdf07bc0c1a00cc88b3dc46241e6541441fef039dfb72a45535be0024c864f17f5fd272cb6200d33d75b121b72468d68cb7003988e70eb84ba40b90124750026fd65974a79ec0bce8cfa3075244715f8afa5d9531ff76f5ba6756d9229da1a51dd81e26269b97d4e2667cb0d8878fdb461539e4f8c5f12e4a53170121ba973d720fa88165ad6dbdd7e109a3789c432426746b6e075b7f3045741bb26e548a27cc69838d7753e327fd4eb49eeb69241029df65c0207c37438e042abdffecc45cd075267a88061e6c50632f15660e7f288fb5f3c50aa755da14c6a2d02db9776f5b8ebbf024f932b2e1ceda02223a4f5862bbeb6fc88a23bac7d12bd9f54c0119062bb63ab22432ea3095b7521a1126b618a735e1b59e92ad7b782ee8a2cb46e11500c79681232119a61f2d522ea89e23e685f159098bd6338b94cf3c602ceb752a8b1f8fa07569f3f18aa2f69e509c3a5a70ea4bc6f45a388d27360e68fbd5fe8d9819253cf1e44792c6e9359cbfc24c7785304d9f1277f65da518806d807db630abd34e6441c6b422480483e92ddb026fde401ebf9fefcd8d357ba44635acfe3503d543c8de26db87e305126fc5b9fd2b6db52a77b87f3cf887f2e735ed592ad9f0a0fd479a5d51b3953d964d4442d980ac6ec10a2354297cc936960b965129afe4b76131c5d180b1381ab91498d368aee543e3bdeaed4d4ea8e1ff3e367a331f74a6442b120b383c2d9b456efe356b5fafc86a615c3445fa41f5bebb75364cbb400ad7d030686645c048f971d033509fc13d33bc2014633b6e77a262c4b07f22c7252182776fb023e1cf92ecd1715df301d58818ccacc964438dba587119a37537082b730997f0ad8f030cc9dd928b09822c7963c8340667ccbd9c6615390a481b275ee4a2ac029799fa67df50319b99083d71e7d21d3518b1d16613b28941656bb61f671e149440288919b40c812a7155c1daaf4d379d16f2b75924cb6db93151783884b6fac7fac900556802ac8c19c234054ee93da81f44f485242bfd16c312dde2e2bc44271d684b9ffe9a171352c620b505ad5509643b43cf55e96c8daa7da46b6d0da898f6b86d30ea1e81e23d39d9ce44d7ae7c2f7c81b96f76585e1840db09625c423ee1aa150a4afdc975a84a1ebc96435e04ce255da98994dc48c70cf8684c1e0cf399415dde432ada86182d7dbcd18092ebec4f9dca9c5461a7d4a26e7c9670664f073a05fa8542eb0ba941acf0f789968feb23b703992a699a33cd31b55cbe844400fdd48487071ab017061285a299050def608f6749c2ee75a4d2b3b8ad29edb041f7b7a7d62b415f1cba4a97b757876222f1672ad1081cd559f5525bf56539e81fe5574be661babc25816e007e94ee286f165c3cf21e4767b373e5668cb89da588b9df82d0a108bdc74d6deea48fef3a970ceda58d5d1130cdf36afd9aa5222071ad3c44c7c212f66a929ab2d50c029d8f28720626642ea5817216faf545de23cd70e3fb7d6a67e7c59ed0b345c5a48ca5e725c190c16d33cdf92631a74eb42d4915fcc2483ab09c8b49ae70a71e4ec996cd7900bbdd2ab981f84f316d3dfbb5f2375460a87657cdbdae652d61e4891d612bd64b38c6e1d3958208751a0cd013bec1bb3e5ded9010489bcbd6d1aa075784242695ed607cc8fec94eed34015ce4d3ebb1a81140346490f3eccaefbeac0569b0707728d2a6517f6494360ae8c1dddf43482481cad8f8ea213668da42d8e3542b64caea5160a8a54ffa5fea1151004ed510f9c9919b3a2f1feead206a99fbaf9c98ee0f5bfceb019476b35b87dc663b8118258841f2671c417ddc2683c89095057ff448f5d5cadd58cc128da7c4c6803ea282d9975398735f492409e9784ae15ec08a57e057a0883598b2e50efc5fa47e1c9ee8ab35750b90b7b53af254e74aeb6f477f4e8d0ab63df78dd742d077b57cc0cc8d3a00f69049223e53a33a99f215c30e45460dde0ce660c0cea99b935e26441fbcd8e26cf9489739ab4010b629058438889df3d786ab3;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h49b4df25e68e97bd54cb7ac69e7af600df1848f58f53b59eb745735cbc88edd89fa4328f34ad72f12cd7aeddc984c575bdc7be5595a855e0e22a0d59ad5e333e13281dc09a3854a4636b2e0b69e1fb21fdcae0f892c459ec8a928e1827bf1cbe21b6479e0e5f22d2767cf5145b8f3d1e1b1afe374a1f982560e3217b25a26ee995f996700f3ad960d7abafb369059cd1e5cbd6184d1ca608ae31c9644216591a102e8e0cc221f71859947a9f00cde8111d75e25e84c1e3cfeb51fa211edcb76cc74a1bc78f0dc0dbed7003a058717cee0e27f5af7796cae8ffeb2c64b0cb5a94c1abffe896c4eee85de17a6fa6c90acc8775233eff581d140864d01d21d959c36aa64c4196a602f2c828de0e31eafa62888ba0cc628aef05fef5f76cc119fc045f9b42842a89456255ff7069c85f508ad5895e9514669bfe1b394ee1190dd27c16a27f9f9ff9024e408cfde06d9eea713b6e55535d290b373c3da90245b92114823def4a5fad592b1a7f1bce5fe1fe3bd938c84c4f0af16c02bbf4a3e85109ec03026fc07c94c4f8a0457c8190679ebfa501d1be2e3eee577897be3dac2cad9d7da580e24f55c48d3a8a63d7a69ea1b508f02ea123cb650e89b07f29d16226d3187d7c8f2000b4fe7bc848aceb35c9860f823131d5910e749e79a535a35ec9d5c698235fc87a18c5f5819229f2efb114389b3f5a8b3ca836e11e568e32a5509d0436c3503df1f814ec412b045c95e415b0a5ac4c464cf3c150142d5db092b0e769550704f4eaa8133658ad4ad4ef9ae5ef2cb3ad4c1992a3dfcb8c76c49df29e72ef769156f63fb1247e4a360af7858bdffe1a3b6e5756f9ae8db332e1f241ce867fd5eba0d0ea72cb9eb5dc576f1a0fb8511a6db0c8802b76d2d3ec6452193eaefad31ae3e696e694070018d4ac28fb6e219dcccc9c26bc649ba27c8362a28ebbc57a0132248e481c311daab17bdee978c75f68af5e18b992d80621fc891ea5713ee3d7f3773c5b669551839e26257df36e8ad12a09d6a3743fc253d5a4c36aff6b0baa8c6101b8a0f7ad3248b76fb353f9e1045707e7dde794a0fc8fd772adb28b3ac4829650cd06f579aca6a80d20e6b4028f71cb5c5e7a44ea76435e31d765a6c7a022d2afad28014f394228a693acb5fddb9d548ed47411254dceed080169e602e585a503b047ab0a6e1bf6e615dee7dc4160736d0c41a6246d735cd0a75eca7bc86203ea61aae98745198d11dac9c2aa29e1fbd6c3af0f631473bf1b35feb3486d40967d7fb0a71b60d675194bf81bcd6fbc465eeafcf3dca704ca5ceb37230a93874b7cbc4920928e093f51f56020aeaa2152377d65f15587b71b384be5e627f3add398b05c341df2fd2aed92b6e1c9f4ea4ccd311f36f424286988c3febcccb16dcfc33b62c84d939658be10140b6a03d5b221a670650a9fcf887aed8a1d70b334ff381e5010acd9988fb80ee7f24e9998c24b52193c6acc54cb3aa23590496c1dec6bc0579f67889e2b5a8fa05037074191a54b6f0c92dbe77c0192b41967d83b748f43d1cd48d9d45af787b7debbd19645008c6dce765c4871ba9a115df5db0e5ad8cc6d5a05627a398770236d4a72b89eab6b64a53ecb2f0bc9842c13f07ec943cae600b25fd1039657e90796df62f8d6433e7af892703a8c101facf0cb5e03d86529014ef1913bcc232d2fac09fea79ce9a474c607df8087e4fe55f5231963994f8b2f0fe6ed6ff2c159c3e359a1f2af71a0589464cbd7debed46f8713a52636d279d0af187e20efa35652a564cd3765b03865385558f0089310a67c9988fac47a751a83e23580416839575d625c301d419d4cb591cea14b23bc73f0a80341473f13143fe0a4442387efa160ee2ea1df492a33a62c90dc8ddd3f8e03537de267a0cb74977a8fcdba5091af9b00b7b6db247b19683cd93859f406a77e2a21a5a77d387a96aff843fc01fe706adf61935ae21d1658d15b8fccd68a639ec1c51cf25ec237bf7fc5c6dfd6058e214c8e99609003f38d4cb7d8a100b71e5fd80692d6af0230fbb14c8d80875fa13795decfcd464b309748f4a214348587140486f118e61c414cec6a534de70d5a2f10f7406370c7e9b2037421bfc81753cf2d33be9a583878d7d0cdeaf56070609ea2e3d8ec81ed3b814221451907a11b223d4c9da28594f34f14c0f37430e35b323d385c21b13ed0005166c3f4d69f860a4206d42d3eb5a9c8348ed78da4328f1f8188a9ad1cafc747b5c8e0ea2be7f07755e74f47ee694c64d3f57370a12fac12207adb91cddf5f9f24ae0d821eae333b01c9c00ea8044e10eb6b1df247b66feb707c4812dc7e3dd0875213d715970880325e5f8edd85d6d2a2042a0422ca6e2de5358bd997abf11f0a447b6b6900cbaef789a4304785ea52efcd2e3cad00243df2d23231c3d4198ec1e1cbc0be29e2bba261e42341d3b1d44e0b29715c470c9ee1004c2336afa1399f6f1aa3a41d678d6ade73fb7186990ea5889c0a58c24e9c75594deb6e5d754b64f5495f94b25d240b24675c060017a78076adf6a2746344477e2390251c2b64c5fa673d1ba92eeec00678a34104e9d675c7c86de0e121dfe7537e7d7c8bd64671560480ad2fa0f228cf0d82c3325069aa5e221844124f84016a242dbc8db473ad9c4c6f309685190603dbb1b70e3b1b3fcb810f155719a0ee8d110ef063c04b106b2b4dabe3528d4d9387c2fb42c9831c3cc7d60ff67fb4900d6e4ee652d076b25d51353998b31dea843c666cf2dcfecf174619a5d1a26e1db1b31ad5cf05d0266bc57cb6877794893c03f4c2e0ffeb8b899ec2b7196eabeab9f1a3ad8b6ebe6f9f5aa1f7a47c1cd5b42b4666976ea20dea6e26abe839b34601d76bf4e42105a98e1b450807;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h23465b96e1ab266d947df87eded4bec42b478ad2275d883b8a9e58e9b715442df36214293f9b74f1c1cfd33dcbd06cdecf5b9db47cfbd6f6eac6270d26cf67443ebcb51eaad706e4425be6091b097cb0f81c2b715847f9f7b27ebf6a28278389d6aeefc800764c6c0127b643e7f4b9d7cfe9d05e8a38aa35e7cd5f6b200c31098d437fb25c05fb0ca36e37b174402b92efa95cd900f1ba98472c1a0c65b9a1e2ab76e6fefcff009e040fc2a6f350ffd502d3f6fa628c2b85946b9bacfd0e5d8a543422423a9688443c6162e478eec71c815df9b2e9445a79f885990cc11c52c26cf221fa012e44e5d08c9b29f64f9455869d54411f2bafa0addaa7e3b3abdb93567f0582cb5be42ef567e656a7bf103c7c85897cb52e5d3d6a7e1c20c5af815c8e6b513470c317952fe9500769a9bb3af8d241ad6754b9d8bbe54ca58df905450993fe0fd6879720a4638a1f8e3c9e97c965f1f30f07624eb05948de40deaea87c4ec1065cd6b5532f2394a370bae50b89188598d284d2f5a563fe56d06ac61e7d7e7b90fc86002b18313c59a1e9aacbc8bfc26e42d452a2757b75d30a1bcdd3b4f01e7d6e86b049dcc0e2b6ad673bca0b9f68da54c41f420d08cbeec3c40bbfcfb8da2afd4989e730fc60b4ec7025ed776e82d3837ce172a92cc53b75d5867cb6375cd48e2d15335371b2b0bf8c30ae3c44ad231e891d582d062c063c2de68810313dbfa9cee7069aac132f9e49d397b6b3c19084d02c471e88569f45ed5e76127ad6f5b21d4842b32c1b7198a318409fa2329827d5b1400c046c06931fa5328cda0118356bb97752046a69e6123b619e80dba71e877acfecb386fe0af294272125b5535e32b1143c6f2445c7eae33b1a2a942daf6ed6c6412c230135e9cdb601de74244ba4ac278a31a1a8b56cde9f86572560906fcf370466af573f0068435308d48327d56f9bedf9050a33f4d236f1fdfacd9a484094a966c2edbb3a48b3726d43ba57c1f4fb4f2c0399ea8479fc8d28d2cc58c459df50fb899e9bf1b8d5023fb1bd6e93af07e0ae85a1ef822bf55896f211eb76a1434da4537f1875994e00e0b6c2af543d483282a31961deb775c36adb6914bd24f369d0b035b51edcfd7b18a32ec856f7ab1b945742d9dd4d82118973fd2089f3d8848016b11dab6b05c66216552ca3049b4cf694c7b1b912f31ec2320d9acd36b86f73ac72f5b173df9b8b2f67d612a9a1ae9c2bce19c1e9f372be5112de2fac54b0c505ef2cc358afc5b460b609e110e6990bef8418950a80b46defd078f28f5c988bccac6769723f5a30cb4c99fb51184e4c76ba878915cfff53a18b3baff8996b0b454515a10cee64475fced306ecc346c8f330f31e741bdf0d6dc1e4724ea45e5e1b18e4a6741c4d394930db8a892c70e22558213d4fc9fd6af8c3330c9568ae39897095d8a3bcff07c05c26a7e7cbf2018c18f1a20901585f578697c3870fc2b8122a591638a28ef8c248f0f7855139094978d4a9e448897798ecf812cfd291d6429e3b770287db1322411b571e1f87cbe43ea1e36c1b21e853470a00ef67ec7545bc5f55edb53924148947b464e2153629c502c6661324edcc77d24a0de0365df57159fec74aa5dca0cf3f3557b4ac5a4911e9e9eba54f761426a676e95e5bfd8eefe70bd745d91faf0271be941c83815687f55c201e3be68bd47e4f171f25a9116a5c50cbcaaee850f8a35dccf67acfc4869b6ff27c03678bbdf7ef0c4fdfe7aad5bc86a18afdb4b96ed1ded0e78735e30d2eaa6345fc6e18b4ecfd0e399e67e970d68b89e902334cdd02ebd406b2c2ca34456cd9f088193918d7eaf3a8b51f2ada1ed11b3759a71c0ad111007ce821de9c5faa3fa9191ed797357bf26598fed79cb8a4cf2bec26f6e64bc0777969aedb3bea57b7b3c2f5a42ca915ad6e057aa8cbb73a8c6b90a693269c1e9cca239d229ac90d235eb2f660a919ab8222d6f2ddc67e12191c446d1bf53fd98e29ea8171bebab7ada3c7ea3709553ada46ea396669fb591f1c8b5ea7813e5e68c50b8b5ebe3d71fc8355b271ccf60f363663fedab3ccce6493b33d6d703d8bb7a51ca16971b799a50b24e4f853021fda75c7fdc1ca981046649573be64ffcbc0d26541e1fa19565887a37ea8c6f7b734b71662edc41db3c075d9f014a35acd9bf9c6cf976129e9abec939e6206585a05ddce8be529cf4c74ba94417e7db6ff142b8e3fb3c232bb46f170295aee1956a1e71e2fe06d52d7d01d9f0bf0bbd277a07409dc77ac0dd8626fdab52705114c60752f7d4c10d95960276b9e3f8faf740db736cf18964f8f007fa2eabe470a3102fea1848a12e9f9d62bed7016e4a1f8996b2a44106acdef643f65c2f842b3e6d43b5184bcdc5781940db6d7687b90309be87b83291f2dac633d29dc37d15e4b065e6049731df941eaa5bbd2acb1f8cba8916213f25b1b3ed7c0435ed92444b5eb1c51f239835d16d5f26670508a8232b96e08d18ecae291e89054d3a02feebea93049a83ac81479f2b620ff4153169f878b58a9805b266ca175000f37da1dbf6b973140d85c5e59db4139d2f32bead031d296a79bea5feed7ba8ae1acd6f70e24953249739ed83a50f6af49b560fcda7dcc3d43a03a0ce5eb89f0cce2cdbf623c023d17c3af9a0acd1538d1e6d51a8a29677d623d8027e2feaceabf1bee8953b0bc8c916cb9d4f1709cc22e03b67cf3f282ca1a6290e8f07389cf3006e76a4c1d236dcf82fe0f48c556cc281d9ae52285f2944d7b12ac38473d7e9c5af78acb5c215a964cc11205b005d2537964f10236c930542e2471766bb167ba939775e9a4744030ed58fa0e003ea2f5cec5305b1a4d39202ab36375692e9ba9ed1d420db980dfa7b91486a103d3;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h69500b693ec7310641a6beac692bbaa3c335bd4737a67ae197135fba5ff98085818673fd6047c4b9799e47cb48f4b522a1f7834fc312f618ebc9eb531879684963a2e99f265f9877cde10c32039c25351e47b2fae5a667b4bc3ff9821b670c98fdf1ae731c7607b72198384c79e9da1026ef1eb1c703eb3cf985b1a401cc57f3c1623f2ea62d7b2808b0f2b6baa0ead617f6ca76dd62ff2ed1c591fb22ef84319c07d4732009af0971124e390f6cd3b89629d61d1b9c3e268895588f20fb2c97d6a665b09f249d073ad2298faec8b9114ab3cc9afdd5f3e5f43345b73efc701d225293f35a7a2e36395445755a756ae332700d7ff29730e805f0a0a9bdb909c89293288e4ae5c0e4c2cdf99ee2d250c4898b422167c78fd9baeeba491fc47b4f6e855f13ad450f12abaf69eb792dfcfdf847638360ef6c50bface87f6a1431e83d963482caab28ae8a70404df410d416e96fa408af585cadf1de7447eb12b170c17031c45704942fae73cea0d7b4bdee0bef09f6dc7b6cab4efaebac26ed231948a65f1f6198f753f410b835edce24d5574db87558c892ec627bc06325ce3165c97f5c2b4bef767b69e4601aec3e25032d9bc6f83143f045556b5a4973e8ab4ff4fb96804b99802aed16adc44befd1934c836c3970639977c3e96de858d018117f90c62cd63ac3dbb633d3591900ebc882e2bb803434667fb544ed79bd8760ee33ddeefd6a7b8a97d88ffa57ed36f2261f387c20292637324c324a8e53903041c23254ff6341e6823822e87f91e14ab83733be6c3d89d13e411330d148bee419a07487310df600f41f215cebd06b2c98cb502efb4950567b59442ce7d5ed6b431a6892f0f89b5fe3a631ef8e5cd113315c7ddfc52c274c4ab3da105284d2d371279055d36840eef2b1d86a4c629e41942cc0bed744012e0b4aa20704291e1d5a9702036dd2478aa83e877c712cc9772756331c0c52a85e220983e3d6fe69edeb7e1379e16a3f394a72b1bfa82935ecff9a667de8ca14d5e80e626285020ff7b9a990f7b64c72c2fc7901c55d058419316ed4c16b669bc63c3b286048b981d511f750c128d6f01ba66625a3bad0578df5464ace77d76a5d8af3bc7ac487c3d43acb957901dc7f9f478772949474fe80265b36d576fdcbd924d7f1b23b13a2d9f7d373f6ca00310af21cdfdb6f7df8c329e742e27cd24dd066ca0704288b20ff88f38424639b6e005568c1c23eaa74aa3bc325a99265c6a3644b89ca5c6cb6f068c79b922fa6f3524e23490d8016c8d690bce44ce9c6c72db7e575eaaa98bb20c0d0cf02be26050cfd585859ea217aa48f6a83747a5045e8664073400491d5177da22587f355c5a4091f2869f2616f9ca6ed6562f6f34ca8bf1407da8a3c5f7bcbf1a49901b91f1e1080aefde67c84f131a6b1acbeaaf4421c32d86a97d077c882d702b7d05ddfce8799ea29300b857977d66f1de39a2d72ebc5896a521a1cfc13a976d34bedfd04886ca176bcf600e46434c6b4dc3e1a61e98c3c90b8fedb0b6bd228294caf48f54efecd9cebf94e925cd85ad5032fe2a235b974489ede78b33989887eaa5804a443d2c111ec899d23063d6d7996047100b2fb7d6ad0e24001f66e8043c04b41171dfed4d9101d62758513d067ffd06a105b68d8ce8bc08c2913baaf451c9ed262c2597caba069978051adf175dcbd4ae3057b24be5764fca14f4c7ce0c60d830ecbd1ee531a3d69668d7470efc116f54a0568042cd2c32bf12ab0b3d5666066efb731c4b8f8190d32550407bf9039d9f00fea2821cfb03665aef689a25ceb2baa3617914557ab4fa8ff14c965bddea4556193f74294f7fd5a52f4b4e97d32f814fedb03117a8dbe23294d8b737eeb5af0ee9f526a6eceadf40a19a4ab56369002e293faadab9d87f5c1f426c3f7892207f618e14bc0204e7b8da65615ade1087f4a5ec5e0598932050a2c55f4e6ba35e45ee686db24eb3da656d01b8d5ecdc97d5dbee371317db7a6849923759580c1522b1baafd9779e928d412dd9091ff9baaedeeb9ac008eacaeba0cea57e8b5ac730fc3b930a121381843cb7921195bde9031ce8ae796df4d91f921ef668f64e26bbf54e3ec49f0d73021fb943211ed2f0646fd45c55f3e9a25ef05ec2d10e26c10f0c258bcbdd30d7c46136f923f446ba4ec184428e9a3d4f6af34b0c424d75b175c2505dd65de90c9211ccee0825bf8cb6a9489d1c1deed2c281301acb4fbe1129d9c4626b07c2a91bd5940a9c183d87303dd36fa4478c5d883b1628e1fd9701c7d84b358e7ac69ddc5347edad03dc2cd4d706de7a80327b85f1f6b2b5d2492f1049594c4258b2f3a3b4cbd23d95024e57d0938bd41525db3c49d8d46828e4f101f22a232d2713ce11c53e4b3d1cef17e6199cf70e7d1505fe07495822da6290ca1715a3c16c2043f4fbbedc41825e0e56594a492e468ad6d1c649649aa0e2d815e9204bdc4be54d55c74c052d18d2b1524a0aef0a6c2ce2413567d678928652d21513d88e78ac9e68682cf674931d1f7b86ed3545bc494b2028b253ad6983c5add72ec8cf5ee83d5c0949d2a46f5c0cd5e3305494dfab8334de4f76196d3f6505d115b4dc709a453ed710cec7edb838510ad814f2053d7e83adf999fbacad41675287508228b23336973785913638b8fb2af93686ee530517b005b479cedbeb56bbfe00c6478e4d41b4f835a7a8b8edfb72419b0a681aa40c19ea296007159951ec7ceffbc94ac7eac0ed63f1700463ee1c1883b60efb754ee8992474ed58ab0e6c363a9ba4bff4f8c4f34f0d7b7d4be1465abfcdb5ca2d3527067d1553334f591ca65f554a068aa8430e39034fa1753589f488053b48d769aa53c39b713060a9af08d974a4afc2882;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'hc15a704e264f2dcdbdfad1e1c54e41fa5247bed9171038ddf109eb3559294b99b8fdb0d32ffd289980bcc174a51fc490987383f359ea2810a80a7307805746ca2ecf4c53dd7e04b61a8a00e681a7e054a124a67474678442d2da7fa8c9cc8ba218bd1594088714a976c310448c421654bc754f126f9d4553cb7f31b13fbc57e6e79297b113d0cce2e4025f9a6c556d0a6f900d97e2912de7eec51dea58cc55f21642191571e14fb36b679fe540de9dbf81672a86f808615b051621e4977047cde74e9d5b5f2d80a77f4273987480562b37ac41e4beb84bd29389df7adc1ae79e66b8b2dd102f368afe6f3ae3d4e1467c14d82df7383e3c787d634d6a0282373194c558c053aa67d1029bafc4e9610906d44b60a5c2cd8f26283afd61bb216d4e81f43374df68ee5104d92dffabf8d6ad309ec46418515f1e402574d7cef4bca85e088495e6484da94348c663ee78384387a41d00d7be870a74cb3d117f71bfbeec7de83e8d0efebd50b454aa8a45d6c7255e29eb661a88f433623e87219533061dab88b22fa4257ebc5aaede0e29d12ee5fe3f8c7137ef559eaa656211bc37f308cdc0e70253a8ac108064afa341913d13d86d029862a759739684640720f3d225d7c87d0a8793d8da88fdfe6951d5e0576b2897dcd399bb8357abf830bf71eccf3ac1219af90a1986b44f52c32804b7a0b3d12170329403751c2f13b4cbd8359fd69b40953aad6b2dec50b64f364e7c4c743969d7853c527a249f0a3aac0cc22945b9ea21043efa2f62d62cbb93bfe0a06d95d0948ad672fc61495f2c22bb7f0e008b2c8cfa636fab28baaa71e0f1fd0e68058583e13a0a42ec959b4035447db8ed3cef1f0c5e67f3e92a92919118b3e9405dced71030d2336b42882f1db39988254f9da189904f3261bee8e65cded5bbdb4eb5eb54054ae09f1abab81f2372cbb1f46d024ecb33bfcce31af0c7f3dc6d533e4085422fdddf1ed00b71424c54b5e50699aa008edbc0da91d5ef8c522b8b07bfa81071d8d2cd6baa464fd75395effe500e4a0eaa6ae564f46633757607758c3f54656de6609ab5cc66f40f095afcdca6a97c9816517237e08b694fea76d58dc70d33d2cbeaebdb268ac6b58f988b81b853023b4be094c8e6f0c7606fda9119f637d6ae250edcd40fa971db7c58bbf9b0831e61e10a9d5ba0f8ed7f7054214f8a853d76b8dccb4209988aa11daed80ba9fc717762d3cdc395e5f5285a30065a9b81eab7e7e81187f331d1a550e94661864179428a05f6abcd05a901349269a29ce7722f9821a9a46d6425c3ce76bbcf2c16a7a1f91c1f23410fb861e73cd3764382d20252a683f814912109f443d288112b818f9a805beb35ac8211bc7e3304441059d7daf79d20e72008794abf44adf127f56ecc23b5e89af609ea154bf3825361502c8e519496e1d03f32fbff72d6334742f162d097860180a8caf670c7672caef346200f226575603771785fe838db095d568e21ff3ceeef4a3fc12327f045cdc42dcb84957c896e7e3664166eabdf981acb413c7ef689f0e8f410317176680368a09651e91154a892b204c3553e6f9df6ab3861635a6ee54cfc856f9ae28f919be7fd68b51165bb1eb286c460e41c6141f937264201941fed238b79527f715f21d18b28e6cec0d94739a603ed8a8757a9dbcf89124457ee30ad9fb78d540af801e08f82234673afb3e173f7537a6327380128ca555800eb6c6feffa345f2fc58b76119c26d17b8ef9f674bd19ef07ce946d47424ecdaa93efed7d8f7b41274d1e3f286f1759ae7480e18893562371894d957e9371efdcee54d190edf6233048aebb36d9bafd1526888d7b152877c81fae7903bfa2b8e0e703b3f1b09eb1b56a55229b9b36ec06cce10515aa4a86f553a12869425c6564c72d18c9b3fbf7fb35415d11d75d99c0aeeb8fa76d48c1a52b2068bc4829052f4bdacbb0e51411a7621e7b785479b88101bb3296b587ce3f064766d9985178b8eaf490871fd462f80e9f034fbeac8eca563ea06da99eef067d0da34a905162a7da5623b5f93c46843901ab7b1c0612b5c82c4c29348797c6b9ee376b4315f7545840e2774551b1f4f92480871f8731c3401d7f9188e61a9630d361ab68c06d6b9df92ffb93edaef0daf49d2394d144633baeb2f003d1cad8483d10572517ec1a0fc2b3672426d678b28e575f57a301a0668b36fb496cde4bfdb2f0689d938dff5e42b39726bfee45aabd6b78dc0125d7532c867739d1cf3a03ea707ba9073f471da5d10c647c1eecb94e374ab9bf71f86846be7740f298b79c53ddf4f35a3035fdeb54e51af4831ce7a277ba83ba49afa557f6decbb572e98625c7a7fd4a580ea2090c98e62749bf53a04da6f374b349dcf8be389eebaa11e786f828382bd55da77f1d0e1a7bdef6d6a0f04b24ca5c00a2ae51a12db853f6282bdc5f55958949ea56de795e9b699ef487e7acf4b3edc75e6c218dd9c002d9f2ad832307f1ddb5b5f452f4741c602aae18092eb5e48d0b750f9f2061cb831d24460bcd30c14fe3f09416b443cc990e7fd8eb1a9f56be42fa84884bcd23d11d276de60bb25ff1e97828a12b49aa8abb56b65562be24e1bc733bd99b92426020eb18b210d0ab96d2af3c02e3d5ef640f92bae71d234a147d1799cfaab95600d2b19d2dc0c0f74069809f20e7aca187e25664bf938f3d355be6e8e6b81fe6e7c0275b6f1b2742395aeb068a582e4a7744676ddbab6d07ed5064e5deeacd6b2b1ccdb7f8725a08918313499bfe7f4ea50d84345e0308c0c23dc4ff9ec4fcfc58d2b54ab2d2c123e72bd4b0b1ea4a94d0160eb80f3f9a684b7a6608bc8d1509263af3dfbf9e2dd92097b8ff0753ead37c9f22d12b60fcee0e806ecd5b53f2;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h5c299211db364ebc4ce733bc21a349f379663a152abf01689ead3cdbfa1978a77cb1d1038bd41aefca65209f098aa313d619165d91dfa48fa984ea0332dd86b4e7f10adbc184dddd57e03bb63e0f1e44406ee11315a2ce2dacea23e7d71b556305eb8a16ca60a0f25c037ad65d561665d59c852ac0ff7589e74070b2851867562c3d7fa883aac342f3eeecccc1bd9a5a9595cb643f6c597192cd1d1efaf724fa34a661f341ee29503f112bd7b380d31767a603a13f556f5fcd54ff43330202202c7b594f420485ac9600e48d12f0788b8002f536d64c0b79c60d42594023231d585c3706992cb9e854a2e75cb017ce9d4c721b695af194a750b5ddeabf649eb2ac63059e2afa28687114ee44245aaae38bddd2def428f6d3f07b7dd1ca86ce420744597b8987a9261719e96d86c370693ebe7aa58eab86c714b182f932e2c1e237ceaa8525c987632c194c25e275c21fedd473ba3d67693d18f3a2f82069a826de1ff749afbb10fe998caadf92ef38f618fe7c79f4cf92154681faf63e7dfd2e553cee4dc57a1739359df833c9e1fa1d4d690635159e7fff0c1506386e1a8d7429f6db10db55682566e7254b69b5f8ec4e46b94a8d91b7f2dfe6ebbaa34e9cbd0bab59c895e36d6586c7374054e3d0d52dc79fcdbacad8f457dd53e9e46ecee6a2c837e4ba63269e0e3a9aeeb7c9acfd0aff45c5e3673ecbe68b9dbea5448029aa83e15cde2b4208c73f316868b624bc630a44db7903d29d0e9967d111d79de2dba3b01698b3712a1afe78e219544ea9fdc9d16bf653ed2f662844aa16586335845c5d4a7b800232ee24655cdf3ec2e61659a4157c44d4f804641b422509bf461d521559073bcb1aedbd7b1ed2c2a79d8da8030f4961e792314a5e8c6031fb8da6996a2c6ad4f6dfd880e13806ce0392fe9418213f78f53898a5ad6dbfbef914c416e2bac2fe73a1fc99a80029fe7513f67fb52dfbe1ac8ea4bfadb80ee765bbae8b5cc06c8a53b79bc4d943a56792e6f692924b457c84610b9a96c76b3bc5a35358cc011c24b26a66e270c148bca0a8ad4895f2753c98cb525838d3eff86dc01f4c57b6d739277aead64ccb07eba30c581852d62b1cfda1a76946ee7202560995c481e90452848629d5bba6698c3a87297c3e7d79b5157c93d54d2fd6c16ced29fff99a5776d68f5f9b20db30e518ab432140c2ff48d2d6ccaf8474510477da72b31c0a246c702d716122f4e7e81b119e585cf937ecfd3d527b6ccdfa45921bc6586ee5cc1869f9820718089bd05fa79b6ff0a4fd767a1ea0a8c8dcb8bd4b056d6b12a7f80c8a71f120f93944a1c31009029904f6891eae11148ecda18c8998e01a5f4f84956d855f05198146ba1aa5d64428839eeac31e88566b737274c6652370475ae6774292db4238c2cab3d446c86d745c30fb517cae3b72a9fc0631d51199388c096286e5ba409c7e7482c660626370bcb9b282a6f61f0d5b11e5f3fbae31f87e7d5ac97e346c8c6ccdd30d3b80c8f4989797449c0fd5fa895f337256b62d5c1b3e7c7f09afa0217a3677e9b034b70cdfa2c1d96f53e17762dcfa491a3ce7b539f966766aa9adf6caafa4b197d3dc4fbe5d2fe5141209c95db3af5f8d4efa58acf445124fe51bf0ccc311bd3f85ca3f94fc350026391aa92da9582dcbd9ff94ad8214a139dc49e8fdac3fb872d202825e4c6707c4a508a268178b841ea3c09fd5411fa4fbb1c778b873d159b6c5dae91c862deb1b606d8b5347fd5eb9dfbc2e2019c55677e2ad9590000223cdc181dbe606aed4c18485099b340cc2c9cf6b9b23c91a8bc4bfaab419a2eb4112fbc9a4521bdc109e7b64088b9879d7e67349c11400afe965b0aec2299a7f429197147370b3bd4c38fff0a30d7229a1b58fb451aed75679ecd9c8a840d0c255e8d14f466268ddb308a45561a6adae55ad123cf2072e279d78f50cffd161f986eaef3b80d23222642c2f4d1e6fe37f0fbf83d3cd9a32aecdae4b8ebc98fab23010030b010ae6b29610d6349fe8836f25f4dd9cbe6379f4785c1bed4aa7cdcb5730ad68d2aaa30d172144d45175b1ce08bcf149d906a4c3b474278af9bb10a226452582266673c6c53cfa33a607f3285d5bdf3dfa924cfc404306697fb41cc1d54fce1b3f03b03a4815990b24c7645084cc7c27b6b538c7b282ba3823084f7ef09bc2212a112611ffc79bde9d1aa732027301e2151eaccada1a0dd5fa463f20370948edd665c9d1291d3d699db9dc6f42b7a3d9da27be3276192ff37418827ae4e9f02ca6d044b1779ee67eb4d60309eb95831a1d59dab6e8eeaf40df34b56aa6f025652fe9da5aac6f75d41442085dccaaf07b9ccaa9024e96a5096f00fa2c680649f9bc1d1457166d07de8bdb89ad6b9a5a687c9fb30ae6f47580b66591f9f29ff1fd7ebcc629e332a6c85431a14586574c7cc2d1eeb507709807f44fb6494998a10a9ef0a53452592c397594319c8bd2c89b302b8ed0bc6d7fac4283fe984a401b7e3e4b8cd368cfe2251b32d6eeb34e3036705764d181e3088e09b98ce95d8479a811838fe8268bf9ced0602d0f910a87596bce0c11815bf61f70b0737ca5640fb6259679685dcfaa40c43c94d4b2a8db95fbad3d15451113a02807b0a68008d8eb7280d4820d6a921adc1f7102e87529dbe803dcf98c903c71f65602cc2ac3d6f1ed50f6b2ec7edb45e20401142ea2155f8cd283eca68a1ac9dab551a07464605e28df2a088b7e07d0e13eb955e7c619d3a55e9cd8a8cbb529451a74da0ce37c1ee03f221d7099470037cae3df0a46b88183240da13b3b84bc8cabfdb4eef3ea20179f2ef7ea5245fa1daed485102209b570a8b36a17cf845bd2652efcb0fff3336ba59e454a4ed4f40596a284973c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'hdd16cdd9f90f5f085687104ae3fc5012c6379a34906909725d99025f51ed31c129c5d0c1d460411f21fe901f16b8c9e6824cc09a83c120bf3970e1be369ec9dfa636a6167619c62e232d2ccc37edaaa058e052529fbfeac2f0ea3f8d73e5d8ac2310fba8c2200053129b3bc3e2be6523d6e00fdeb11a2511124d4f7e303dda2f64769c94c5d2b6f3c124410f443d36b81bfa3a51ed64af7f23b8cb0ed72f4a98532819946e4d2dc2d3c6bf41fdb2dead2b0abf2f1debc2d2c52c49fe3cd39174dadbd2572cf6d6830655249f48872d77850eb415f10b74ede722384dff84e862aaf555ef9802379a85e3bce251a5c8b7c12eeec35a2b90ab398068001d54ef22484b7d7dfcecbe74a31e7df7162d51d7246fc720910d489cbf0e080df8e8f1ffae9ebaa22b122805957dce4e7d413f8e8ce52b89cd29aca3c744d7ab551c6c3263875e5b5ec7913a91e4602c6afb54fd24f25a1860fb64810e4d3dfb8288e9f24848926c3a7b703599b70eea3fcc338c357bc0323143cf3cfb4a6f0756151dffbbf9df9f436244329d27ac1b311a9ed225e04ab1a27483997778e64c233cd5010ade9ea8f7f4a3a643820851785ae15cef294daad756e2316b7408472fe79ca2ec0032e3e7d2918785a9a99a2d926c8d7f1915b7f095417f0ef1708b90bd65860cdddf5048c05b2f1327491a20f7b24aada7a32c26a354df0da55da152370a1fc23d7351f47c481b7f333321f8f841023b69216727253db1e03a7ebe68733b86232999835290b0c29687b8b8bf321122b67ec8d96ee819c3aa4eaf0a5913e19080ed4b988344c0c92515d0c4cb233788a7608584c239d4b3c686f73c3bcfe238ee32f8a4cac92bc60e28bd8b5cf6c5d9d3559c46ce45e3934b5d373fc3e0703818ae5b90e0a96100c4002944efd2502f63642b50aac523fd5b721af40a93af9ecbaa6d645fb7038a8da86f808a900b6e54e0fb9efcf53f69ab48824086ca1d506ca90f44a9f0ab28063a44eabc88dd0fedc9b2c2184f65339e08a55d1d592ccf6f2badf3eae00a29e76b420e76372e86ad406affcb0404264331b5d2cecf5a7fb96cd415e4504549d26a5978119b98e0ff78ba2e1d7391e54fb47973ba632beac781f3407e49b1335f22072fe9e22c8f0f705af44da55b869c22ff1424ed1517257772d0d1f84d2bf4ee7284ed2ac83d2f5d2e9bccc4cae9dd3ee956f42b8836650bf175794507d823fb5a493f490a99afd2c1486a20ec62d3d5d2efd0f770e7828cf6e7e9ec471c2c84af394c6793716c78a78d64110c9626899d028c51287dcb57bc30000344b293ec80ab410c1bfbfe102746ca6b56bdd09b046ab821c26582c1e97a6023a7f1fe1ab57f62391bb91fadf82be63705f542b1e838848c3f8f71aa5494f047d20eddcce9b383431ad4835d699d684ca9d6d9996d48b904b2da13d43e08d3aca413171cc250c41b7ccb15e3970052e16f5015f5edd84a90642ca44419097da50468633359c71a35def8e19a6ec1e8c2cfd67060a2e2f7b40db1b279dc739dbb90b6b2c354c62552c5ccd3c5bf4ef3d924925c3a6c65e04ba6f78e716d859e945643def5613c9ef8f7b9e6e945e6289220dbb7d70ebf30a65146b1394ba89a976179228b0a31ec3cc9aae7b9508460c90163a11229ba20551594c6f03f573fc4206ea5f5ce70caf28c553414d71fcfe6572b36ebb4f239ec5222de7811cb5fa4ca5136dd174e8f3840c0e2050a1bf5fa0820a81da07fc890b2e5b20b90ae156ca5b96866c5118344fc7f472903d2ac0f9b38284358d719ea0775290fa6d641f74c49b3d2a87fceeecdf3155a94a904b1a76fe32c423f790b81b3f92be466454f05f7b5d9ff52cf5cc1f1936f051ee81a72cffae357d26b831d059a176cad82e15dbcc08bb9c75c728c3e94c55faac55ef8a66afbe938a8f70c1e6a81c4a17bfb767b55ed4967aeebd8d809e733351236dfd434a669d2d4b77ff8937fae2d85bf53c78a3a3e84f0c33eb9348ca3e416f3d5b302671c0330d597afcb06ad80ea89d0071d81a65090f9f2e35626bf18b8c64ad159fcad8b9f6eca13d2f6b8f17784d21bc198097ef6df84fe29ecd442d49c30867623e9044c6d4fd14666fcbb098441d938add7fe2700ca8804f61001e2da5f1d26fb3a0baeeac360428b2308c6b2238ab46afc669f19f5d4e5fa76ac96383cc8af3c2854608cff9caead62ae676f08c05511e9d8eb6901d53b940b9a736c9367364eb7efa359573fb3d650d729d79b2bc267e47cbdfab5ae116dcd2009febd2cb6b8f2acefd6151322ad710971568a2fb5542be85dff45aafdb39638fd1321cccf5c01982dbd594ea706c1a3f30f1c5533072c8be433edf488d1a029c0b1d4a9380d6e604248529a8cbc60a5c6978eccd190c9ce0469ee5063b32f8b79b9ee69e6c37c2edebf07a4988cdeb7c9d13cb8b1dcb82f29279d6a947be8d5a1713d782d603ebd96cef785da370f3a09dd7c6b89c83c0208459d83f9a35595ac06069076c5990c8c7cda89c375e76dd33fe8a9c2fd0c887e18826b76a4078f93b98afe3b10240e2a3d42bc560083f24c328b27b7fe9c17ed52194734014ddfe7484fb1482a6b4cd551d0238567d9e03e149b87a886cb77325bf68c9b68b5e99c8e019c1b21e02f8f7e31b41df840db46339d89f7e43b8540a18e2dd87a79945e38c57071373f2c41885990b036947896c9422dd731d3e657e6d9a9d7416af0ad81df1ee09ab957a3af783cd8af5104522f3289452063dd3f4a631f4362abca5b8b05851904c45feaf9a6dda013366789d5fe54f0ecf087e70c474c1bc8497370e6562e9e70f757af35b7e9be6ab7cf5be4bc64aae1ae27b9c0b8fa75d95c5756212f6917f4f77eda13d7e4;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h7c7fa05080f6e7146cf6f45cdd8169dd47d7af8dd5d30c3130a2047189479ba5d64467462118899b26081716e0f2ad20506ee595a160f860d53a17e067c943136e38bfd1bc7fefdb2ab1c63ccaebaf049dc1b3c478e2b06153357e3d067bc244a92cf73bff982a2ac03f9289cd36fd42b132b49c753f5c976582b1be345a57c2e394fe091491c6806e075e2ae1c1ef5669c22efd9ccd99c0f99fd57688199c61fdbb8d5fe92e262e4b245598b3a823707de464bb2961374209e302cfdf7a3bd5167c0c92f3caba2f01dc2fae1603b254d9c9dce45912072a98c2f919ea1e293f39cced6623953460829aeb67b0691218959ea908b52d322308f845a95dfc6a5a00e04888e81d828eb72fe0eb3fdf2f5bddb0aab91b9df22a32552c5a1cfbc64654cddfa8ab912a796b1a42b4b8bf9092da5d2a57f17d01918acee9d33482f1275982bf6028f8aa824c033e450e96b3ce63c42618d0d495d1e71e2b79b60a6ca8e016e191103493ffaeb5e57ea2ff11977675a49f8aa7efb1be2a6df6b46d4c4abcd85d3d37e6ce0adae18f50b45507f3dd97cf5198667904702ddbd8cdc851aaf7e807ea02c1013297204f27d554bc7f2b7d23c263098613cb8ed0e3d6f8a09ecbb33acc21ed1236ba34451fb836887247b2de12b0ab5f9dcc9d4dea6d0e177f452d95aa45fd20495ef548ae7ff6bd7158f698597fa55fb941670e009f8c6422697956a2073dcf4e3ca1290277fba4a35ee3e1282ce74f48cc85a2612a99735f5d80ec5bf91af566430cb798f14e8a3fc1aec124665884c9af02032211f9f63efb35ce0e2a16322b004237cf1474dc067434cfed1de963a305dc1ae6ca75229f27068da01967f3125592dfdb78b2801912e216f30bd1248c724eff547c2c1f857c9498ff1920d8b00fa60a0207a009a364f2f3545c499234a59120debad074d457aaaca3bb367107526f824a164dd43a8ae565035059da523f1d4e1e0e8eeaa0658890be068efc845f614355441607782180b6f1d69ff1b2272bd35da585fa0a6491fd97eb417af5945ab9fec3ba49635694f649bf7e842a0783bc097210dff71b4f63f39e0359418340bd4d7253f05734815e36d20f7ede8b06cb70f288de61354afa8bfe40475c71558fb10b9b1b9328526663babf4c46971c920ccfe8f32df7b399c1173a001204ff0ed1419d68be5367eba02bb07a2ecd406264aa0e48d6873b84e3a0ef893e03333d66edae76ee5b4f988c67fbe7db2b6dee6a0c52b10c1540f3f9d975c3bc247b265ae6b67e7c4596f2351684f73ff9a0c573918208b31ce7dd8817174eff4b11ffae52e9887b2e4a7436c478a6f55dd008ae8c95eafea3a6da6f3a558316d8cd8a292930c2ea29c5bc68fcda3eaf9162f625dcaca8bdb1ab35415536a7e04704537251f1c1470bc55320806401bee8eefe0f6cae912ec2e7949d1c23a4b0c46829368109ddaebb08c94b39b4a654042d2424a5cccb89dadafbb889418841284c974c0f7339e48f08d57a07251249e46be257f64033f55720c0b37d43abae16ef06139efb5247872484da80753c001c0a9cdb603298a7a3363192c3872a4fc6af781a4a09708ace5de9c6ea653a4c08c6c581f00ffbdfa5c7dab6f3e35b2b329ae63257f202a2ca5cb47637b4bdecfd301e068cb998ac45b1f71ed484053e0b7bfed4be8c61caa74145ae4f6ab926cc293ff182feb6f379b515f165ee088be13804465ed873576bc50a04b72bff2b784b00e96ebc0f99264df6e1220edcca642a222d87ef671a6b3ec3f71582a2b306229f02610980193f1f0fd2778d2f89256a8fd59983ebde9124741c53270643778a68ff7d3035c83bb6d5e54ee7a65138cfa24c44cfeca36aea58347eb75b31431cdb642e0c4f65bf384a9b9e8520c4d3d0a7e1cdca6a6588fc4a43493f71ac2771bd743794d2fb36277cf8016d74333a270dcfc3c26adc4ae9e3f2e4b0a190f9aa92ad01f2bbaf7dde94e425bb0b92cc5e16226f9aa12450f3c0dc39d2364285240f1c9ab37f668a90fab89c0d218d6fd8be739f97297e29f473005f3e7a6301597f8fdfd698ff180ff1701c09a5904c0df0654f61c180704ebeb6c937155b7d591da6cf8ef6e31d761b032856c79c395d67433b78c8067139e3b1407739992a86733a30e6d62d2cee1316962067c84b12118c2e11fc262fe58d01a76f4af6279e7d3c5f7c41840396d8ec49ca687666e34c1a0d728da7043ddd173b7425dea817655ad759cd4799116dd1defd065e3b3d3e08e5774ebb67f5332a8e990cf08b8483919d22836d1be93e4413bad2759df498209d8fe3d22f6a2dca01496cdedceba30fe1ee0fc38484eb6ad8bf82a863424682528e994cbb2f5e311c2eba7df0031c95c01d42c534ddec8e63703768e2226f8d581f86de06d7d79cb81d369675ef95860fbb2d37d156f593bcbca45a05e2114e3627fb926014c394a026d346b781c1f382ff0594399026c3f9aa99cb14833223b58d94837d61b80b04170a4b668420c1fc9a4b9350d04d8cce1f166e135714e9af355399e4e804070db00495489437accddf1f8ecfe8adeb7a95ff8bec77f30068f06af1f3d5a234a5844c2b53acb333de30eb5d7f81a9df974afc44e3f802f33c1970fe389c7c7706046a18edea06150f47ae8d70ebcab140dee6aadca07d9af0f18c61d068d004740e321719fca922614b10158c4cb281d21679a696e499ceed3e901646c00f0c6a30ff617dd09dfffed3d09acbf2c9d3c46b33073c1eb8aef4616e920b89613778913d2e72e6d66c97d0e24ffb66cd0599e9979d2c72b6a601919f447769878902b5f0dbd555cb05cf061fd90e657913b66211267827d286b68984e681febe1024c1045f5e604dfbc64a9baa;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h5a259dc33c847edca56f2be0cf75060b9cf3f6a7989226f4a793f624b4f0d132b49e78ac799dd342a64eec81132976182306c44931900d4b4df8617b7188237da2e8d7d75c4678f0778443d7ede2263bcf560c1e8cf85c20bb20a6ef243b417c6456e5143407b4bba8d470298b0bf7d2bd34c5347f1cdcc643cd18e583f831e7fc4876c4f2da78939d70dbc82bdd746f3af84614da4faa6ab87a03d73f64575d36f876c3bdd8fe2b9f735c1c219131edd10fae45600189492abbe029fa5a20a6ebec4967a2fa4cb6682942b7566cb7f266946dfeae6a53ccda4f512d1f04cab189ba1642d117330b364ba58ba5b9f601c3ad5dab809b68f55c257ee135e070e114a8dd3a41f885c5c4c67b58de75f2b27b9af616d0e7c522ad1c9e016f079cda05bc8318c055a920908e6e432c37e441e6471867a780aae5617c2f827fd1d61f80a0060fd4b1ac45f6c81bcf78e4e8940e58cba64a60c3b5b8d25098db5757bec0a533b367914f10557f6942f3cbe16571953272f32d51a4a7547624214f8489176288f4d20aafa33f86951ddf8fdbb49fc51ccdd6eddd463e85acdb29f764cd171e939ee9f8c5e2671ddfa3f17e23f99ffe561902f00c576a3cbde7fbd142ec3a80fe2bd86931217e2bd60cea0d08f83dd7aaeec617df68005f9181e253837cb2a0939a62439ce0dccf5761f3c29734a3ea892a340ceca6315f0001a071502325618fb332a6a00d865cae9962ff790d0e3a7d5bc2709703406dd2442839b9c7f604ff76fdf9d78c27c8fccef44666c1a211226244c14d8fdd3ece6f577a8b2442484574b468ed54e56e57c6f6cc7ba5320ab5d00905dfa8c5f185c7541c154729df4d3f9e0f3b96f2a3b3bb3c20bda8f320c018243a51d0806172bf1a94cef62c4549d9ecf9f0c278deed0250c1e57f7b21132539e2bc4a11b7a902e6082614c64c85312b089299a84c96b71e1808cf483f1fad1cc51d1fd22ac7c8914ecb60e0b0cc7c583f8d61d050cf756179c0c190b1ddf9ce1ff7959ccb97d90199aeb5705f9502c85039e13c3c24911ea515a3520065e28e8ebc51483c8a5685c9e4aea9881e9f45b46915c932453d3dc01eb3a5fc8696371afc7d13d959db9d2ebaf0b7737ac9285814186d71e9bf9b7935f082579b7cec6a04b981c363593b82b4f244c9d6a31d7ddebfccbef1b18fae2bcc5512494083ef30b6a990a272db27a42a998894808a8ef47bc374b64efdf84f71932efcc74e3bbf4852c435378857e9c02936989a3bab490be70d3c482052f25edb4790f539a3558af80762f82b878a33fee384deec85fe9ec4503901697434b932021ff21dd0185636057f0192adf623c2fa41d7fb2812fd954eae646152891cb8b0306da38838e356f13ab61e4ea3cdff253c7048d5455a7fccc9f96d3c7fee3fea83b5b87a655ffca312e1065119c92b8d5e9de96cee63b434d232bc334a2b0489796e67ba0ddbe725728661abcba64b8c531e75ffb48f1e3b2c6f16303779b535a1d8b9dffa8e4bc2a11c458e36b3dfe7c4ea7c12cc661429414fdf85b117b00abc8416a8bf33d4fac42be43ac42921e044cb6e8c1129ffdeacddeb0ce6b2416d22253d248bb457c895f89f8940c3c33a0dc06d33bdf952f79f06a71a057a785d9fed4e156802a7d1fb88398c98dc86e63395da450d96af72bec42f61b46d1468d8136a92ae5d5f9671fb1c6f85d0d0711fd6d6a0dfca86e1e0e9c97c4785ef4a6a8bec6832be0ec08f74abf7e943e69b0e2a12c796166bd7ebf01327ea829885117486d9a74e20570dada42eb7ee1b779a48c825b34a3ca02ac66ca49d20533c2f0cf57189bf17384b3e8ede33b54b8a877a4a07e74e00d0b32c6d343dc7d7ed1b44f3a69412deb899ca66959e162c0bb522a0fba8f07d1860458ebdf875b97ba120530c7b18c93077ce986945231ef89efb952091765bc3249ef61e9bf8c7fb626e0022814273088b524a87c80d147a3a9be34eb71ed39a8aa55d683f95e525f089a2d12a301b9fe154f9329a1415a3ef2488bb1f3d0d6f2157b110bacde5f0fbc5d9cf271ac2543b5304e726468b5df835df7fe71e42be020f4f1dfc728484852d212b688cffde1174863d9dcb2b8250ffb36dabe441f06860fd0f5615daa56741f9359659d921a0e926ee1b4d3905c783347eddad54a1e1f2c8443976f65d1d5096b515acedb52ddd54e6f10039bc8fa883c66e9e4dba72ffc8504a5388d9f2f81000c1cbae208016f7410da3a6d1829e81b5df0e15c6aa21955fdedf7222c4410bf584f614e3efc7047ba88122b447d90e7a3d0c6be419232b87c3d1f7568b61ce90f7830625fb059b4fa9348ccaa3b49fc31416da744e76af6d50d2a2fddfa806df9608a2834d9be3fd5c5bb6d12376d78928bc882b4e8187b0e5449e4b3e075e214652ac49b711df99f85cc8b263f63b75b8210787bcdad50a9d16678f38eea83b9893762894187ef9d4742be991e8c29870931adbe8d9275731b06d2df9d117827bbe7a1bcc7da229ce30ac4dc854b4500c550f369a1f16756f121f5b8e8db203bba83e96da54c29aba48c216f7657b666b1eeae0535be44b7020bca715d056580c32514d4dca82d8e3e7f8a2051c08d60d5836e2be6ed77bd65d1a1f23994b6798e792addcd4610279db81975d856600e4fa1960b39dbba00f3b2b6681d394244f44cfdc20d818904ca09ec83a37f5c9840c44655692dd1788973b65cde43740a0df50f4519a97f6f58237a931ba2814cc11eaf53f7a7b14e240a188a312c947021f73890893458c6c7cbd67acccad9eeffdb3992bbd5dcd492460dea35feb5a8e8c088db5f5b80bef20d777c95c8b142cac1b042330b0d34e2a4b7607baedb7e403c672d1efc2f4c092;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'ha800f8274ae33401444d7f100e5be76b3e4c444e0bd909659a0e1784c0cbb070c38f573d40835ded7072775f4f59c2ddaa59690d4194a0b9f7d2fe68268578da6da53ef3e0e4f57e4d699c97c283acb5a4fa894069840f20651cf386c0a177b57fef5f3767dd42302073ec73f93af81bc87b2defeffe58f3c7fd9c6f6b0b74be1bcf78a3fa463dac78d9ac2602ca2fb9beeb0d2f802a27ea05bdfe1b3c3d2b51be1b38df410d263efab697fab6cf9bf8ff542b4f4b059371d5d036ab65a40a953b0eaf437f0bd8454e05e06f21ed93bc408c757c55c624db23b9e0ce2e6eb87bce1f7d9421efd3fc2a17e5731f63ac4e794724ac787e7a7acaec99c4c15fd3f7d7249bf4878ccefc628e1abf7d4202a987d0cf3a8c71e2d4af8a3ba2de0bdcf3d28458ba0a54a222121a469a75eb9d900dcdb0548dbddce2613097f5abab8cb59ea2b4205e733da7b06f4eea47c7d1da783c363838e8978b29ef8fda8143f591eee319a6aa3c4f236583cd84ee2a399ca5dcf7b8bfa142d0e14e74230861e1b08b2cbcc49fac0c35a22575c9ca1c40caa0c458abf9f7a9af1fb273b19e9332041f25312955d8f152715f69e9805130e1b8172eb5d0f8fc3bb739af4739d9cf490f69abdca3f859866475c9ad690bc3c33f10a47bfd574811682d0d4a7566bbf8e069270b8923665ad452e055f1dc636f08f933f3c862cee5d1d2d65e272b0338b9e9a2d993c5f2d7c2bf4ec9dbfb7628a9fb87de917da16718171c55d225a636c7f51da63bc01d3ae10bc463b733dbc2dc813795e3a46a7a0a82386d0e9221174a12b50e4e71b75d8f0846a36893a322d86ccb3e24f5b6caf05ba71a2448e3eed7cd0112f83513cccfc7783960ed972bd3cfb8b901e9a2292958c0a5de91d48f17bea91490517f15250fc30cbd7eeebc486bfb6d5075c8c7bcbe80ac06d3f9d590e6a42d971a4ab780dc69025271d524311398513247c4f5a0b23eae3b714dcd92e3efdda51beab8545ed748f1459e61acd7810d57542594b6366696468b91d398f98e06cbbfd6e66b02aeba539ead29a9bea7656660cb8e4fd0d50bf436523684e11327fb448224d4d65ad51e6e8062931ad1ec5a3d8e567b930daa05631b8342fa0e08632fea6e43460056a46e1e332502dd66d6a9fcd8d7b2d248fc5875af6bb2663f815dd7a815b7ad6082e4a9f7628bfe17800ceff355f61526e3b99261649f2982abe021462e293e3c7a51e4f8f22585fc97c76319053c466b88b1f4825a516a3382e9065fb72434aa3da6b98a71a551edc8950c6305409ba6d8f081d0219f03beefa59e2acefef0104c3fa2b0579c6d2661307e32ac33dbec594fe0a0dcb89667325824562926276a3ff279a94b5f183f4f0197d451826286f9fc62b4230ef03f6444f4701648abb72ce19c3fd86598600f4a0ff26b78c90b38d538fb2d36fa9ac9d0c19bb6aaa6f911656c5db1668c01c178a8cb857c5d42a796ddd08504a9d71c21ed721e92d42bab2f6724e2176f09d30dd42fd2b84deb1013c4d577dcdccc7129a0db266c9c3dad946324b83d6f7ce2422150e93ce940b244a591c230dcae4d2ede220fff7fe764c9f4f84b5b88b7ab493ecafd03356a55ab545f19fc444ed79e706064c8dc267af98e8a1b9b7021100ffabd419be18f4140fa168cd66102ea00663499a189d09588bac674fb742c2b0c82531b3a21729acfc67272e4b2371ba8eefc134e490000cd00566242fb485860e522d1aa5ae5bad275e74b05c02c877bd226fc297c2b2995e9b1bbdee7f685ca43b390964f0474de657695fb9152dd4373caaf869c309f0944266f961ab2c5e78c3e8a0caa5901fcbd6f5bcbce4db3739a99428cead1449d811cca3bb5ed70f11bb974582d64be9871b0fdddbf041979094c8ab83793f1ac0f99bf650f398b8697a271ab782fc3ada5fbd1179046b6823046a640933f442b61d11d22b6143033bf84c59dc0861c9f7809b61dac78307dd2404e3ab32e4abff8e6ae1934887403ffc0fd496ea8626625e53bfbc551758ddc317c490ef4a2af4de5a66bb9f3e04e49cec14fcf16ad1788769a82c8b7e8b62e01d30afc72fd983d15914b07fd36d3acce296684b45117c07efcdc040387894f36954fdb5de37c6beb9dfb7383c2a16def7b6da46229f53f582aaeefa11bf8d4f551c83525c6c1bb140d132282fcaab3ecebffb94a16a005be353dc9acf288d110242c86fc1d42305c6c85c4aa212d9856da31bfa54acdf10adcc04c919c7e40913d26bc0f575afc7d911a47b1ecc129ca8ba4717e729e169c6cf74ff706f52dda2b944c079d90f30d3ded91644282ba1109eed0d3e44cbcdb7a69debe9e07cdf77a7f0672780ecbeea0c1887b7baddf1d84dc0e762acfe056be1156c7dea269c227c41ff28bd9109d1eb6a94596c81dfddeafd2f57abcd70dde3afd73f8c6d87fe0b69366fe69c27836e7b4e07e607303c346eea7907a3b0c687655b6a1d0847b11b292f23725a02b5c93268269609b469a054f0dddc3bd0a963bada4dd2ed6129e2f910471e902e32f43c88c2516dd42bcc8611f1e7e65ddd7fc04d107e97dd6eafde46bd1c11db0023471334376c44aa6e6cdfbfa09df996ba3de8fb941082b3d2711a59bc6c5fb364ffe1458c643312d083f9fdfaf6a62d52ff602870e184a16f5ae9d57169d52624483cf62d649d90eeb0457242a8dc4fc015af28b86168f5299a2f6b2718cb6cc6587f9dcf9b57e8c24e1feed9b2d28af77b2541a14f4149e703309bb1c6e7ac88307f14ed3a1695d77e43bb97f3771de7b90484edde5c307571b67a99b881e349390454cfd6567f6459360dd150d90d9374dc46d17d826665d70623c00168c8da270c51aac025b1cf0958d7430d6b4;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h8480429db140f52f611a41e51e7f1a697d77fea87a1ed67bfb52460cea6bf59ec3501203973cf2dfed258c498d92ed6d13b146932a5ed5f3953d562014345a314a431a6367a6bf092156327b9c3c97529422ec9a2692615906894aa894ae0ceae265ff6b00946172fd75b19b34a104730a6fc00fdf60c7f991b879c3421ff5d8f2a12641965d87ee3ad967d8bce54e687c7032414256979cb40c1d453499571bf64171cdedf49cc6bd9b91e26b57b6ef28f8721aa469f3dc5179f18ab70bd21b66bd5c3da18794e70deb0b39bd068291255a95a89339583d0d785e79ee60da41f52d30ab681c4922d5b9cece7b8cfd707e299da757535bdf4915a46eba86edde0331a79018c8fade8ff9d6126a2858591b5daa08cfcc3ceafe0d1e493e70fe8246f79a968089043719a82830df532ac590d1239f470af23c931f597aeeba1e4908c58174905500bfcd12fba08152c347298f832f75bc815cceb32bde28bed4da74e244ef49100db823a230f33d00ee76033b2797b55bbeb419ae46a28f4bc14079e061edb80edd0e846ca99da42d3081632be97cadf3e5b7f6e43ee1169565d24d2e0498674ba045258a25fd5c312f8013b7313e533fd6d18cc7c0b124a7eede46ed9b268be907c364ef9644b7565d5aedda0a0a81f45725f5e2a5c40ef9e6f782f9567f9263a23265e4cf950456ad1f644cb190144025fb52deb12377b2d327298b716eab46be17f27cc60fee64cbe1c571507308c74169d393e7fe82c010301fb0a61631ec20f778786dfdfc786f00119e21b8002dc746330754718ae81fad88dc51d25c9cf7498acad78462ef2dab125454396a6507c425ae00bf765606d4cc91ed1362350cadc7079ebc3b38629d2f4f116d910326044855bac03c3cc5c1f96cd71866e5ed5cd078e0df31db8327bb4a93c040bbbac85dae53cd61ad99bfd9646f6a5f20787b11170364773ccbab8764019ce82f29c6b39ddc832c2f3ae72fadf16f6645999ddc7057342cddf248bf34a64d03f555771deeae10bb1aacb2c88aef3a549918f7223298d682941c3a47fa1299cede5453b25e0d1ba48f0d4cd72d61fc7686c1c53ccc9d9865350313a6f2ec1fee3ce72cbc5989e9baac0ad0055ca11ae4ea9d093b6293c078e47075478802bf75acb37a08c27fbfb3986190a4b3f348aa13f7f8904d313bd7eb1ac4ee137eb5c08f95be326a9035bceabdf219fcf0d4f387cb099dc4d2d65c210b67e45cb846f0d53a2a3089d9ec595fe3eac1461491026eaead2291e1a90814a0bc0ac9569239cd82531000a803584933bf119eb552220abd0cc9cec29ca4c9254c1c905e6dd498bca7dbd75e7557304d53b5ae9983caf75d3da29214a613c5a0de6fcd04eab8e0da87ee38bc095d31ad24d782c8f6c57111cfd4a3473cdc77bc8e3bcbab3a774ee4b1823150b265400d94db083c642bddda40b2b9e4789fd4e4738df89c9e1c978847214a7e6af5638fbce76bf6990c8ef1fe00acd82dbac7ee6ad3400e5c2bcae30f1df8b8ad8c265b8064394040e7740aace38b22d2294f36788b38d2542b659d6e68bbaf772c3e43168ec1b23bf0353d18a18bc61f2b27c5619440670c34f066dfc78f998862df06098f67e10e2bb686c52d163508bf0f7617a77410f993b498baadff209a3d9ff75754d5127d71c0e4a6c6c2e8ce6a22d0ee13ef09df4bfae4b8deb32db066b458bb9f1ee95e5ebdb95e676085fd0cef2b8893885b15523760a67affbe96cfd120016e904d6238c624566031cb9ca6e2a848c74fb782b9bfe1e6830e31e71feefc6827731ce39bd605afe1f6b79f862f91859014fe148ad455d32a41606c204b0ce295e2fe94893cdf0db89555aab9090d7cb24b94cb4c64ae949321a152424107516a2c3ca393ea6680b1e450fa756afd5534673fbe94bc1dc38c9c0cd31e124289caef0652a91b7538d2678a3ab199ff159f0a839e3612df8d46c43f9a4d7d46820e92b65047bd4d121277e4e901856e5468a2bc1e05870e5c8ae523e8ff3820b017b348de0111bb63636def514d0f6503d0682633e878088396e7ae1e3d1e8183242c640530946aa05cc7243639e2947e428f5a2ab984f67c49c1d21e60f779f8eacc92ec11269cf895ed77303fbf1fdfd4cca30053dada40dbc96655c3d7024c57f03dc6e1608f02af24fd38e13b9cefe07038d149facae268de9a270b259c884e73ad1ac0637d8e85a90917e704bdfcb62046bbd5ea99832801c2900b059888d29e7446731dcc9ad4185faf2d71a904c482a9bfd78a589260eb824657fa6ebdd03371d554d216fc3ada5e1d4fdf6e5bf14a5520219c94e630b333e9b7349576f3097df425f5d8f825174d625f92e844d2e6ddb472722db98f099d5e17a3b262334b6903fafc9dac0777c5f219e545fa2ada22a516f968904ed5f805f703320438f4f18fcd109f42995a9f4952729328ae612fcdbf863c96aaae83580c54498c15b5bd4b10e338b5d275dc7fc5acb72d4d5ffe3764f60d055329e2c7eff30e5d6c702c9743fbab08fb99dc9055b9e05e30e25dcc030b1536f1e65dc9101fe2b08af01eac888a265104eddbbe415df74964f0223a1222d3efc27b4b9307f30c2271793972b4eb48140a26369bf470294481fc6ca187d980cbfe0b940beadf88b7ca1d035ca3e8b433192fa80a904a0d7987c542dc3985d0629fc5184beb9e6e5c50c80e778eb4a3e79d458b72a19b796b2a35b22ae01fa21a6f0edb53e3fbcf46d6905276ba9155c26571f2cc38539f61cc76d254c2cdb82f7c245db8101cc00c85fe79517027c1ad1635a267d481bd72ce97f306482c3a3ea5d35c9a13819111b18182cca454a8668db01c96e624f1d1fd283bd4324d185f3925dbb846869ccf;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h6284a485c0b25d038029c6b792e060835db15c9910521224ea5960895ada40b9e56035bfd8ec637c102a51090482a992badef09c383e9dc27d37da0f7644b4a4cc09ed1b0228046a970696ea7f171e02a1aac42a092532fda413de7b28e715ed95c690ed4dbfdc5d9e928cd4cd423480b918a57c822474720d17f863d8ca8fd96a01c04203adcb4200c264c8d5591d3999c4f1d946edd953ed3cfde21f7bd6925d892d361c36959a266075a622d2f87b57a2fc61c9b28f05f5dcf474dac3072e4b02220a325ac46c04b540dba3901cb8636c9d7d9078a3d801209eb47aeefb20893c8e6482d13e4ece1265859aafb21f08bfaff592b3cf75866ce06b553e142ce9d51b9cfdca9b484eb5108e96dd8fe92a478f2dc869011296ba574f278e7775ec1d6cbbf21fe60e5a83b4c6f8c5591a010061445281fba3795353aec9355c368a78476e51557f7b56a97929054da45523858cb821ac31056101804fd23a7623b89cf0b9717f7191119db41628048bb1dc6d60f9664b1a4b48912c30d23bac8b6db861aa20cd7a01cc40668cee4da653a7cc38a735afb480075997718814cd7539450c06c373b5d4f28d37050774bc42b6c3a439258ab9d9d3daaa176ca2af55661e5e68086cd150599b6347c829308b82d8c4e60ce8f95e41bd7a3eae937d916627caf364ea4dccd32f7461184113411b0e89ebf4fb5ae2c9fb0a6f47a6622009296204a3a2eb6dd50bb80486b76ea9dc446512352b980af36c1306fe0156d09ba199314d1f99e7407b6287f36d26882c395c6f9fe44800ce1454ef7b325a9ae0cb413b986d2e93cf92dd4d7900779f6ab33cf5d59d9c3eea08bed12ab6f5ac807160d1d4afd1118f1f3687ffa12cb7485a6dd6066a85e059d0717d857ddcc0d8d97406060f95aabdfc6286a913b0fe4796c579776091ac1fba205e190c9e94d11fb185fff0bf4d6cab04f4b20364189c9473042170be4f72c357060d517146d93f38786dafbe147efb999d4438c6e52162d03a744ed31c71ae49f9e9fbfcfed1a1db17585db43d3c2b5704b87f41f478178bb8a849c15f5b7c2dfb457bdeaf6bb727f63112787fbef93fddbc897be3d2ff32ded5ac71b860574f1059bf92a2c0b49e528fc086901a8e3fe9265c00ebff8454b6d2d658b42d8bae9b0e035e964712e6239d397b4d8aedd6e40c01ef5febc485aacac3eaf3ef6a69326fb83185209d7df18cc846a86b7d30c57880e7ee1495f6434db06223ffc50ce3800b23215c602b73b165c415e56ff6a59d6f0abf7334dfd9a2580e25ec0081e76ea63f6a6f97e11b53a6de0100a3ecc26399a016fcb8e88dbbf105968e6b60fdd42db95627f7ccb5455b8095859b55af88f3cbef0fb4a5e101c79a956165627db8054e4042b4916c2dea2552788721108dfb3bef86e7d6cbde8965e66410fcdb49c32d3285d28d49f53581441c6af95e312c56d10719646d0d02d2432f6e4a034ac3274a3689ce8bf43ffaf469c1e59b73e15746e31802f81347ba3452c0666f5596561285609ed8dd138bd19ac3870cad27daa9a707b5dce4fea9e1ff643dfe29df20b84bbcf388a363ac2d4b601bb09c9d5596b18d523a3a71cd8d66d62351dd3ba40d761c846cd4c7d5a31d80dea5e32af81167fb897b1168db3b4f41adc1f1f8549fc5ff56413932586d5414a1d6ed8f95e3653f9ffcf6ef6018953845841df53ad434332cc9e67f0c169ffb03773de61b4f795c0bc756ed2baa98222175c13c20ca24e67db17e3778da19e9f70f5b62d3b090eab240810af155048dfe4a717a41301f2a2235badfb90460d3f379972a200938c1d27079356aaa7b64e5eea77d2f56249d6ad33e4b82a450de6cc962bb5d6e509ee84bdab49bd764a8f2087fe7702a03c107bcdcc89d3b069d1315e98c33a262c1a92c38805961d3f96ce4afb35a7a54eeb243f856231d665781b0e75d9c6c9f787df70cc2a309ce0ac8dd93af1f3dbcd0d357b9b94a9ba4778b1d82ff01f832d233f723db328da5f164f1fc58a6dda2b0463b4d03021847b3da6a5efcaa65dd32ad91e8daa6ed252e52d85afdfdd41711eb343461c896226768feba86e237a0fc1bd5b36deea1872c78c63ea0f81aaf3e82d5f5794bb4f488885b67d7bb6dee8f3febe9df6d1fbb7b51af66e8deb0bb428b4ec0d4be33220fdca2756b544375316028cd2c56dc6db5e42f8d42a39dc682de486ffdb5cb156ccede3c61f17f7c619fe532144e1793935cff5afe88e097691c1d4561aba9245b1635bf02cd02e7a0eb015c0ab0c328d64683f07aca1ac16e27be1e1f07876456b47eeff5083060b39f5710d65ad6ab4fd99ab58189e2f8347cba2608fd34dae046a33afe6ee335151c75ce7795bb3b4e44638aeb96c01d35db07327bece952fbd7efe57b6f753c92abb71d38f1aed67bc558510f2795a93b7ab7979877778bd10d2fa51c9f32ac184e0cee8128a0cdb14f570b7a57bd013d018bb34e3773711c81569b0d0e229651fe76a790c24132f30e1a593bcc66fe7992ce0ac90c85cd322fe9dc3b786140faf69bd879e2f465d9dc66b5b4d0f8970c52b7454dee6eb7cb2c475bee86ffd7b1698b19e3bdef755482d31941066221ce632980432459661b09d6a5580682e34f83f70ed085ced88db98739ad9014190206fe99d902c95b599c49bcd25a1d04aea8757c171f642400a5c2cb115ef3a996d3011f3cc3444845e4146c6a3b343521c723cfb86fe4205f608f52a3894046188c06f30c0d5687265d7d638ff7344f62e0c8b34f679e1363da37e5a69ab24d1429b8edd22e72952bf9af446ada400cc3fff06d75a27c926c0f1fbb89c5c788eb68f4fce2f970a1329e8450e0641ee8cb41a7d91514a7b1dc48c4314edb74;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'hd90c2ef86750043257d0ea634547cc35f3f4b820bebdc1801406021068111c4229b32832306868194a4a741bd510812d67900d8d0988815ccfe14360235666ab2c24f318c953adf96a0150e2c4c841260386614f589d37b078336ff0d20fd2e86712670ed35afe797dc3eadde79c297d854747587e1bc7c83fe13ad4cb1a3d8396c11df5509e1dd9c46a268b0e48fbc3f92e78e7fee19f18563bb48cdf8fff09215f1215f6ebde572f581005651f9b46b82a6b7454471a4120626787eea7b608fbd04579b06030729edb69d7ea1563b96ac7b180e71f793733f90a3a7d72e09e46778cd06379157e04582bb2296b11de433643b90d54295c733e61bc34acea1a678564396e3a996dc5c3fc28223fc2494302835fb1defc9551184e62cdec65b0139dd16d315c14503c51a8747db91d9b4555085fe6570ddfc0efdf421d1532898ffcc76f91cb6ab02fc3ec519962f48ad99930bb21e8e301485e52d0c3fd47e5b2150f30f5efcc270c22372134584f1aa26fef6eea213f05e8f5d8b4a20d99f9d52870f314648eaaedb505e48d269fbbc9592f93f873d739bacaaa2ec7f82661a7a9c3a43a72b54eadb2fe76a20eeb782d4ac2d5e9117e2b158c6b3cd3a40c57ffe36ed4d5b8e6ec019ba428ea5d87ac0aec03c02a5ca4328fa847e905cf0b4e597f924d70c3efa0ce634ac83c7594cfe86b4ae7b5bfc3516dd175157441508c555bb5f51927de2f64bd3bcf5ce7d3015e499a39d0a19190c9ef6da752c48216166b503da5fe4abd7ffd1cc8b87d3ab0558b9340511ec6ef44f4040591a537abb04b5e2050d6ca3e8018f859d91311d15afe47a2a157c8f7c5607ad34002a5d9830e4cd5733f31da8aba5550fd25b11d75aac043f07bb5a198f2817f4af4f8aa3b443686fc62b8f5b6f8ee2c04d1f7961781a1b9ea3cebcb9b60bae21d9dfc492fd8ea09d6264afef462d645ac5cf5bd01065f4df8571fc8497b938070d4fa5199cc00f33a229835fa603747a6a1aa4f2c1e8b9d439061af513437668c1cb39787ef99792d43e756c80fd06e99d3d80e0d9a81fc2ebd6577a5f797a5cd309e22c1e871b4f4fb2d74761818ddad1e1c0d96746f4cb3b5652bac8e4fce78572a29b4703c7311516eddc05ab6de6d1ec63077b6a93e542e0f52a63a66553eccb670b90579fc9519da02272991d1274bd77c82853c8c93b5c193b714dd626db12fd49389829d683396be811c7e78712457764aa135d388ab4af264ce2b6adc8bbe91da6ab05ba3dbc2d86e753bb5ffe1f9da934a3ca4220cdf576846a7a3e9ac4e9e4eb84e63669b336b5237b4ffd92d262b5b299e1164de592d23dab1de4f9efca5fe6bc5da515facad0e40d58659a483f7e39d0fd104540238adbdc9212d2cdcc0688bed16c87a5fc7c6b004c9650625ab5ecd5c41c9b59ee353ae28169fdf7639afdd84785bfe08f4ca2664791924c453910febfd7c5687e6b6609f3688e76da7c97e50e182f1f5ae99a41c9fd360bc725ecd2ecb8e42b0dcf7edb6a34855f216ea35ef41e200154bb50dd2bcde9d0e777517246727f9197c3e596494e687bdfaf545ce36247a52bd07b464e58e427b1c31592b128edcb751a4bf585e80bce51caf194b8d561d35dee47c939a6c05ce8617f698dafc854c90dcc2f8582d517aca238addc9c645650b5e0edefdfffa78e2267e80d18afee40050cb161a7ef757b1f9d916750d54aae1d14cdf8c6c62fd99a8dc611e842f1fc04ad96a955edd235107b8424c22dc47a226a008e562c0d9e702a070b9b929da3807207928500e012a2d938703f5fb62221f5adf2ed22bf58070cb7cffb61d10662896bddb62341ec501d4ea63d2b4286194a65cedc4e14951bb9747286c3069386444e362166258a880cf0007b8916eb459ff73bc236332eacd72ee5122230b19df5b96899598aa1c61605cae340547898e5159c3b765cb6da13b62611236c123bc6cf61e7e46497e46427cbab52a2bd63eba510fef3a0611aee95011b2c74aff93bc53fd335a8ed3f00f0f042085c152139038feda670a89468a524e48c23eac7850bdf34cb7ffa47c7f7a65d19b0a0532666d6a51b2e5a672d841cb2c1a4b21bf52fefedb0aff7cc68df179ef1fdb728fce5b4f04892788b463932c18e831fbfc3c8b59290157af62e855c1063359cfc670ce73dad79c0d4594dc363704886f3de070c61fcd9cfdb6fed773cd5f3265fd9eacd4145be048940a21dafdde2ae4be882efa83016bcdef595a5084feed1b285260d5f130a16cc6c8301818faf99072452ff81e78f1ef43c99f74b4eb9bd2f2c3c4b371da1b94ad95a099f2868a0de1bb19a8e808b539cbc8848c50802847ac7b3dd4455b7687c12c18a08de87fcf915ce4b31add6d8243be5cf30253fd200adfd8dbb2d691110d2431b45a4f06e231220764d954676d28f61ce4c929ae3fb94fd24687310094c96087d4d1489e040b9370e53bdac61129acb0acba6669b7b45f9550797efd01f2d82d063cb13ea2b1b54ec42c85d7021181164079bbd85b170ca1c3aa7528a5c8db75813fc0b20a10f23517e9a7b551be59916890e8e352298f1a60aa087fbe0926ef43642d5b994c8756f3449671076cf849cab2ed11c2f3c75527f5b34de85dac48806a14cd8ef7a9657ae929ae3d0f0acc10e429e929abc6f4a06a7e45bc27a6a40779f3d50a38a50d29b2f91a4ccdf3185872cd1bb42fde4dae29a318ace48781e17f1dd4860bd91f8b975af8b9b29dc1619477529c48aa73040b9d192c33b54737fa54a3d9a495be64742ad0638be77f1528e3930e64ecf74b5c0e7fc41419810ae8f729de45337daa448c62d05a555d87272c0da714d48e492e89fcb39a47de73fb8ca7bd80814c032744b60f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h322bd756d7ec0050ddd643bedb940ee3281a13736b5c3c2a2cc5b6b07eab0e5aeccbf47be661d0398894ca806638668951021e8ec94247e61b903fa6c4e40f2aca0d82f1ae4eedad4b77d305d535410dfab5b2c27c7ba53515f7ca8d82b5b4baa0d9425b53f23dfc6073afab5abc09d3b840604d21ad8585499cbdc130396a91e6db42725f9474c831454d47edc2db41f683d4de34689393460e6642b773ce9e2b641309fea6f47b600861af5d8129a53f351e79f7a36aa3f49968e9f4023caa5ef63f8760b0cc3e58042e960cb97390cdc9160b0ac82a6add8fa73d51ebe1edaf53a1925dc5a9bf8e40f12f0205b02d6472229dc714273f964a0385bb7b9a6f994e8793606828b62dd81f52e6f8f732cbe194c6b5afcae2ad7e2c64370ac2a9f75ee437b782436480a4efd7fc98be06abde1fba9e06206f3f0c7300bd855ea0804669a972a6021b9eec413604f6515f83720d0ae20020347e94594e5536a31e94df7001dda252e396f18d5a78831e53b37fd007ee131d51332c14baac5ccb7296df14d0ea23bd63e71e7f6996d531c012df4d0f2d326985f464d9e7cc6206a6bfb96101f16205c1048d368dc2457bfdceca524c17b74f99ad9a3c3a23b28692d1aff3c89ee45ed072b22ea1a029fed5a57b93c1228608f8dc32cd5ddde13dbc78e51e50f206c961a671479278a30509ed5575224953e72992babba3692cc29d04814dc5c9959a7f0faf4068d2d7769cbb95a1f73d507ed9a8b3d02c5db2e452cd186430145cf9e4b82700f96ea60349d07cf27df830cb9d03d07ccc8d35719102d16c51892bdca863a46ff950eec136a835e9fa05131255cee2ba7f5a732aa186a7274ea20e302a84ae6e6997d7746de2e0a703fbc03b6c185c9bb326bcd06ae54410988693ae7473c0804e2a0512ea693071bf3fb79eac102f4f5c3422d9b0bd31745b527fcbc92d99a720ec3aaa42e416408ff60144d6cdec5a760614c3b6e14791e355908967c84f9e24b8760b5340dbaf96ca716bd5934331bb34aeae5d20685738058052dc7ffcb16d70f690426a69dff12ed485a62e7c2d19af6397e9ac99cabed29374b748b0e20cbd225b9a55babe019ceaf94df292115d7ef05ece324948f14347698e91f42c85652d840d26bd4d8049cf39cc22fe9f34859ba72fdf3ecf433b3cc29eca1d6ecebb45f8e83aea0b19794d1ea7ce927bf1a41403f4c98e37bc667b06f8867b2006eb436412641b121667ca3a073935d5f516b0b90a4e3ca7e2736d798f8360b91dcdfcee0f6b3a9e4afdaef1270c950fa06697edaf9fdad906cdacd007cd5c38f33a5a532a9f6b34c2b0d72c62692173a633ae8305c08eabe166761b3265449866a2b2fa8ef571683244032cb0cc5555ab9fe87d2c17185b051bf427a9841d1607ebddebfd135991ccba44d195e25962cdeec6accb917bd89c8dc13c77e6f46a4884fc57fff50cfde31bb6599c63440e860924f5e508c7f25463256847bd70461e4b80620f542faa47cbd02250dbb1bf2c8c9ce57e432fd54ad1ac0253c297a8d10d6ab6bd8461190058dcb6e952d9d7b306188492fd5fc39d1d9cc657ab94737bc6768c96b476377d3d129cd75af47df358834587af87bbd0d57a7df9702a28bad5b2969e4b1e4a688526b66ff2cab05fcc11584ede93d67161d9b4707eb19bd82b505aca9fb924f98b6a0f1cd1384feadbbaf11bef4b67eb302720e726142c7a60b737f5d2cd87da4626c0e44865498c899d221c0e32fb99bff2d601842ad04561ef0e2019c3a721fa5cf7cf52e973591120893c0c54c51468af5002cf8b69edd59c225bcb341527ae5925e45ddce3f1e127559c6bf810b2c756cef19e590a7e57ba8bf4215c2f37ee6f4abb7998146db81c13940d4e902b94431db5a4474c02de800bcc7ff51b4e38b502efc1751f99ae37423283655b6c0d995eeda3b6411f51d3053a32466510bcd286c3e0eb8fef13f07eb868a484f62185539affe4fe8f1e341a98d140ba2604e357dde3ca824d95fb5038005ad4c09ff65f1662c6c1878c461a6f8194505f2c5915f0f7138842e9452525ed3596924ea8f012cc4c399120710e97b5da0cc64fca6d5899e8ada59bae7b6a253945998b0a819f10bf103d8a728aaaaef18487a414a47542586d36d7d40ee43ea4404a47b28dfaf4d7a37a868ae231f3e33d0419c4967bc9ad43384ccf551585b8a1a025a67002e0c0cdbab2d11aae8f3343aec9e84a3387d39fd10fff514efab24950e74527ac4dce85beb1999d9b32a7fa79f0f1a9563cfd9b69643dbca92378fc492802777af769b1a30679db794695f4d7e175a831194942accb66698a9e25dc76c59cef69e5176e33688f9745a76659130be808b7aefd0289404ed6506da4df2c5e5cae6bfa6b6064c0833f11568b002ec0857b7632152a4e2a10170cd6c691694c1820806e75cbf2b34423e9537167ce57819f0e0dc9c5c0bedb7c312f045658fdf240e92ecd63a8334078cd21821725f143b7ec169dc83cc408715864ba635cbbb7e6c6a376bbd8d66bfb1d0d98b24949cad8043a72901356a32c7c5d2cac366e9f8c40f1a08b2057939ddb9c14496aa89690b9fb8160fd7cea0ec3488218449b9e53b4adb16d15afb38f2d5879c540b68757aa409a5ba6d3ca2e67796d70c9f1502920a3d3cf421a31cb7d345b3ace725d214a21ef78922804a2ea0dfd4d5b07d3bf0317603448dedaf74781240d3b5f372a21cf0917576701d0ce79df899a48a6e76b113fd2bbfdbefda082a1cf787e2e5a06d8208a7e6c73a19ba3de29b89fc9d3346ef711a6736b73786babc398ef3c56e220cb6d56d4f78b517c79065f3a17d35246ebcf1dd5805847826e03b7f3c2505afb27356a189e2980;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h2dbdf50d92c0ac300342dfd340ab4448a5501b3acb3e26845f2a8280451f2eeda7cfa4450f8586a11e81fef46c9c03376453df9e80011e767647a5f6b064325e2f57c7d59ffa4b8836a8ed203672e10163d36c693ca690856ec5e1d801f3cb8cdb4331a746292e9b08a75e3ee202f74db7c9a57ff3e9643e397e833710eef2daf4b4af318b1f4b0cd27146f1ca005f8394a71067098667d74ab8e22d5bc9a4d28df4db4dd601d9aa831372616e6844c92db87da72eea6d253304cc16e65563903269dd7c48911a7284d72be997f1ab7ce558d45a6d714b93fd6880ef315c9e4445fbec359abf81c41f992c9370b7b8f163bf370098ebfdb01780541d85f9e8f67974937ad5af896d76b660b7d2066b2564ff196610019b377ec7b13179f53085daa19294caf1ffab973b5f5d435fb2721388ab0b7e79c59b544a944c9c48304eeaa69392407f1e27d032af3afd5db6114fd90ee429f081901535c942525a5f1e644149ce4ba648773c71e9f3efa5487dc327785d666ccff643d73a14e6688dc1362500d7a7cdb83aefa226ea7bec4035ca01381e2540a641959ba42a64aeb105704343b93898f1e3791c9004838f0b6a7d90f0987cb0f3f2beacfa9361dcb74a31e4f4ebeeeba25d269e605cd4021915d3f3305fceb531fb54f1071e003eaa9c2b899d7c7ab5498f1f5ee062bbe66c175fd4b40f8704c17060a93bff9c2eedba270e32e33e8d147a9d1c7bd77bc4b0d7cb2916f58bf100773ea03d84c59590c18ab073a06e68b6f2ea8458b7991e479db93b47a1f0703cee1f9595e9305df9779a428c92b3d51142a218d0c7bff6d9c57481bbbacb7ec4634ea292815188d07788d4f5c96f2a5aa6dd6f14c834d9ed5d2d6980b0ff497b5938737fa96aa4dbe520661e72fad0cc9227cd9f749718cf6dd47fe5506f8badc83b26727502d76a715badc5a631ece34f771d4464b19f82db3d496e8321afe773f6c25d69ce927c113edc792ff4f082ee9e166ad8360ed7692a6e8cfffff67fb0ba7cc220620746a729aff28f6e42b29298b6c172f576bf0edccbf4e3e858d9cf4050879699a8dba0a44bb9e1e26c7d792f8518cbf620685a6d0386088d33fbf337f86c94d2f956d6a43bda8082a7ab24367438967117ae1774ce8eb1ac3e581efb7b01c93aac798062d0b2bf0f0beb5ad07c011b41792423b4548eb7d50b72f76e0685f2191ac6c4587063d7b9818b8bc0e1cf50908d228543a6595db2737936e0ba1226f106551326d90421051f3a530496c63fb9a34ce36b0c7fb7d553d9b68d8b616728ed5749916e928dad4786307faf824839cb506be42031093e77bd086ce5a532e6686f7f53eafc4552ab7d7899d1f444d4656a8eb7b8054f401ddde2c1f5cc5577efacba9f5e5ad7b5d9bc929851d1f3dc21e79ccf1cfc5515f37143cbc17369a87f6cfe14d7cb6a8e950c83195f6ae866d7f644282cb9aafec35b01886306f0c390f226b86762091fe0873ca4ec75146538deecd0b339a9b169c23070b66d199fcfc0ab24a965bcb101e8f8673d36b661c831116e318b152610287487e2c6de67fea6a91174ca13923fa7244a3506c91cef255b65b611937cc706670003bbf707c0cb1f1878d7e64bbf0706904f2c3eb605dcf5a7c2d52fbb7ff917befe458055c5b56a87f68c4b775a62d72cf09dc6003c6e00b967b08c3c67b271b004ac671d74eb2af221dad0a512aa96da2f050e97c9008ef33894fc8c73f662887e39b0aab942ff5a7cc800fb7d1f91f2625f04c2104da2d82109768815058088256989e6b1e9e7149e670c15064cd9d98b50a42bdf57d236086a17af0b7a661b1ad7b1b34a4351c619a64ccfdb491f44f7cb22f9eaf8c31870759925855c532608fdd325bd2257635edc9603114b180003178f15cba100a90b7150a2a93441ea31fec8dee871aa6299b406ec67c0782260590d096bf697bd2f85602853a6600a51ffb1a359eb3e7a28e49d30af18eafe619f0caa7274296fb35722fb18d1dec00541d8d858555b63e6d37c0a273607008bd1f9da09b58db4017f9a75c78f99914d1792a4f94abd462fa33de18787e3e6821b7f489e5dbcc19bed1ba1db74d43e197d4b55691d113ba3a0fd7afe8b706a2589d5bb52fdabeec96a81461128281bc30e64b076e38c19fa0072567b82fffc9d2d6f3a1eb818dc59567d035e9f64eb34aa8d7648a1266baa5c18297d5a0c7b18e9ffc8f4e47a5a4e1a039e8c0ac0441b37ae1bb2ed8c294125275790217bf1934192ece80d54be71478d36ac4a57be7231d49d9b81aa79ad0e43ee8822a3e8c8eafab15a6606813acb622dc47984ad97c4f8c84b758cb2824bd1d1d0c044706f2c81a68806b414e911b8b311393da1f1999e4e0dc34e852df50fb55555537d192b58a7cd1e70290dcc1952edeaaf991d371b02b83fde5435aef05d25d85660338d0dc2571db2afaa4b5169bbc2f3ef0a5585ab8c8a4847a60f5db75ab8770db1f748115c581dcf91b194bc989674a1216ee9989b04ea4e238082beeae81e59eac95a22b8cf1c87875a3e95b2c416e217dcc7efe52340d80e09a7cf5e889c9b62b7206b400f2abf855cfaa94b20a45c6db421958108578636c13ca9411b0bc5159097fd166da14c1b662528abdae64e3c17e428e964798ea18d10022bceecef8ba98f18dcd7bd4063dd552f1734bda3aef46a54ed320f384b88aab142edcc636088680502dc7c4a7792354be2def6ba04403fade1fd721a3b2ef8adb93a57bdf6aaae39c9e3882f03223328e8e5aa694648ad138b3d34b68af8b2c1334910393691f4c5a48578a27df2184c6c94059c94d7bdf6a6249fec2653a556b2737e4354d9d07602d688cb05338d2946bab637d468f14b5f5e8b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'hf7d82c4fe1288ce7073f1554271c963bf09215b240d2b14ca24353b4949f1cf395e14de231bc7958913e68b811d07fb845e6bfdd17058f0f942a351b69077faa78bcb60afe12f1c40f15be01d9148fcb2180beec68dee9ee027627e40b531c13de4fe612fd9b21048002aa1cd639b09cc68995c44d4650174d52a699222377684d25b601f988efa0dcc71c6572c7d2dd29420bb46b4eb84d2ba340e46321eecaf0b86bfb33994b4f8488f306e725e213f78966e94bd2e7652fea24bff383f4783400658e103d3ecfc08c7466f2aa16105762943a5f48d67eefe2030074798182a86a12aa90557eb2e8de3d32b3d458ee10f1f894a528587de0de3a153997c5f62540dffeff67c4580dfaea096faa6823b3e7cc20101f1ff3128f31fd6e19280e810a9f7dc7dbdf29aea7603510417732f840e3739217ceb129807660752efd1da4fcd2ef748e19c28020eed592138be89ff995536dd438010c880c60e06803837f38e23f6109bd9b5d502c4cd13726c97ccc0da7b73d4128022bc2bae29a30698bfe68836c17342bdabc088d2663260eb0dcd1338ec28db2e2d16ffdc2cf89e567056eec6573733d2dd2b4a9643e5adf239663e3d222f4b876cf9cb3fddf5cc0965d5d02c97cabecdbb70053ef8ae93403f29c7bf8054966861ccbb4df42d7b2567e099aa8e717c8b5506f9eb552a9bacc2a20d0a6e60b6a0a6e7d6b88c48d0056432497f2656a225c2b8da9b8d8b220031a74a064d4ec7f369ba97be2733f9f625f77010a2ade3fe564dd4b161ec72d27febf74f65b681f6457a67d635beeda79b5b36284cf2cbb19b9a82568f8aa6a2851300d417b3c59cea38f629b0457bb9d8d998becfe0636273a7f9f1ffb505676863e408827090691b82358e878ef8ba8b3e35e4709f1d52c5d0d373806cb841bce2b557de3d9db0665b8f1fc01e9c2e48c03ee8208f017b074b8d92ea07d9d175476276212c47020c1c8ccbd3cd8c69b9634326d8239abda4de7dca0051f6b4390a19b87bbcb3b5943fa21dd633fda01fc156b1e7f8e1f739961d80899e7c690c00dcdb96ddebc44bc9b91a30ed3d485e39c518fd4f308b2203d81817c6df5cfa0849a54764dcb10890af082d477fda31e777a1cfb14d60f0136807a4e25a087c06e8cf2ce7e600a77356b8bdb288675c5b90465c2c3e8082985aee44514f526db3ad0770a4921a5bf1f1969d5a37b047a6da517e29364e04bfc105c83fc81598d4afabebe29c198110ed0747246b6790e153beced0d6fe4629369299bfbced0e87955fce3e93bbfb8e1dcd9e74f8207e3c34148e1e10f134fb174851c4a3478313bcd76bac975f969080dc1282772c11dbb1fb3339ef4b835add684a67fb6c6055a8b067fc7fa210bd7a4311edd5b058f718b2f70118a5c3b150e3718e8277e130ca9d7dd5e9d54deac36d1c437d290630820f2584a44346c3668bad7aaae7e06a0b9c2b33e4bd868174a976874cc7b3d4f318cdd01a83707f41661c51f231fb71ac830379a618ce40bb11a4ecec5a9408e7ca27b54a511ad1845d29bd19e76b09d690c1cd58ca29619641968e4f04d49f2cee8323247b9f69c1d4a6b97f0e2edd8c90a76de11a17e5c6ca30628284cc9de12cbc07817be5c369549ad151986af184585a49dfbd5524745feea8d6d863343df7c8fb7108abd1794f8f84961f3ab13daae1364cb73dbf5f01dab45508e99982a6ffeac2da7490c35bbfa16c07b9c4c21fdc81d648739fbeafc97bfd165b53689f2b9494504f76ca64fe48a5dc12926fd1be5f38035be135770e7c8d054d144fcf97d8959ba9e2a822250bc28675f627a94b7fc371d06bc8a16ab139b4e1fb453c5daba7531e18c323501ffeee2e15791298edf49d8f8b8df3767529d6fabbf470a5b27dcc74426d91882a361bc56c76a2fe1a499874b02592344da45d2e4e12834124a6335a0980d3c6a45f4d0c465b164a992999c3601d1007016f8e6b2b0f1e0728e19f4247f34484562e0133cceefc914845f76da232391d27aa19fea6caf7945269231990bee1d75fecbdb2f13a7e23e8b71ef974ab194d4dbf3deba906556cbea867a07edade54c5d6b471fa6c0fa8c6bf961b084e4be340a636c7fce85e8717d3a510fa4d83ebb0ed6a9bdc1b3aea1c9bee6d0c04625c47f80e731b83fb88c99006bf99916f4a1863aa7de06bc0b8f861e5c0c6907519c14ac5e9ce4e2375b486fcea796aceaa55896f204e53a9dfc01c34465c0134bf74780e6ed4519a14f45bc4fa6d6375eadba404d3f16a73932f45552035822fdae1420b661a1752873cc836ed644c468141fb65f98fb227e8d1443b622ed52c91a61961dd338d70b54fd99ddb65b29c1dc9377ec885a49eaf04c20827f0535c8e4e948298c42abbf71cfb7c9cd7d5e670e1a9d2b631124320ef2fbf2895b2094a8d51369eb9ade37aac2555fdc2386f237905162113fe6671893a8fc80c7eeaa6881cd0a2c27b02fa706a7592d4b57df90b79ac57cec9e35c12b06e148e8aad2b7de77d44687c0197c0b9c4cb8e7d108f4103f75f26d5245e2d426dd6c8260aef9fa6c1138f90e25bfb90c7196c7829a71cd42cd1ee73872ee27d3c5331ed6ed63a5d64a06caac1f14c0dfa6f72ad831bf42c72b72fc74d8a373cc4de683bf39e6e274d8b1530a39c0c726410995ee25c5cb2264e2da98655eb53d62bceaa0427a7ef5a9cdc398a9be75a6ee6af3c99c9d21d71314adf36a156788bd2c4d6ef5adce5d4ffb8075c417d91179d0e6916dfabc022a50987579dc3251b3cf1d0942c913b7c3d25c57ac0a3f0310aaed12e35a0604b65e92370d64101891c0685ed29c2b287a4fe74780896be48e130e8b668bc3de3226360efe97f1e04061ccba73bdbc92;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'hdf8b96913102be1faea37796cdc02a3bae570e38812a681cfbe41d1a3fc42724b99a19449f56a332abe2758434958b3c00fa1d22dbd6f71c2957f0ddb3723c15de23542c3eb11b18964261c6daec188d3d35f6154784a98ce3550d768965644ffa9e6148af6f10a34bb910fb07287f0e5a1d4d7d1dd8e8376ac7be073d2ab1f2fa669c661ab15589eba9436e558a7e21b329f607533f9255e2c9b8134561fb2f304fa1ab8d069ef200a8d00a918a9c52bf21200bfde301f29910af7c077bc06dc809a6457268a690efde6c6ed98110b2befbe5ceb3cb3ece0819a6055d9ca92ee83c609d142f9f70f216a1249002ade7b6c8dc23ca28984ed0a43952199f3f136ce38809e744bb57a43a570d9670631eb4c4982d8f9f22f430f7e2a2ec007ff1bdee8942e284df892505b87003499e1c4662047efb8c5d3a05e579e833f3599b3b46bb71a9c9e72b6ad6a326c4bcdde55151a9f5668ef2f663465e4b552669e904a4397367cd194c77c681e9a9795b55aa26879ece12bac874df28f0832a289cca1d89340f32f680267af388ff003f21387bbfd2d20d91fb22c233329721e7661c477655417d9cdacded9cc1e0c000506c454debd6684d7acd50a74615cc064762ab2e4db8a7e172b44ae1b3fe39b883fad63a457bce6a36e0445a5d2f59c75678a5e476d15c3732548db3c3afa8eba96963e23725555a16e96fb0bcf3cee7d1470083d27bf594cd845bd92f1b063fb6dde24231fabef3161b49d7b3a4dfd535dece7adfa8b8053f525874146ef2f117ff56f4816c1c72e4a9746a1270f1ef91826c408b39d118ce9b3aed7acb020c8a3ff7c1d2afc73b3f38a66e63044b043093b1fda93cae106b7231cf82d8ddb9f40d714f83d296ec9a5e5e3f119a75373ed71f85c16f7dd0e87f1dd66e4b4bc0f2eddb7a29f59013b221dd81cb94f7791d1be65a0a4ce93ca87313cfca17f980449950fdfcb61047de2663da8991c74b727b750b76ceba18ef2567aa9ca83a67780630afb238c0b02a9c6cbbc2404bae5e304f72ba1fc0c3a3265090b5733125beceadf874ade1ca945a32477ad25a4748ce023fcd80c250714cb075adb2e1ef4349b4228f97e0438d2220664d5e76b89ec4b8d729fe3e7f636104657ee7ab186eca15f181bc885c2232c09d6a5d3fb943f53e26606da29723959352a12d039ecb330d8d4cc7860beabb2388955e01cfcd1379097f5540626fa199dac1ffbaebd449c215a66608d227c0a0aacf108bec835238537f6424ae2d78e57f0d69dbeeccca8fa9aefbbadbdacd382a1c67ee5fc082bde15bfdd6531588181de960f276c74c902a3b2ad1afc306484533073a0d370aa6b8b70a2150245972d675912dd15e3c72f53907babcfb0b3d5e2d3e7de61f0c87f0c7f0092a12a3e89180b456b5d46e86c398fcee3a2cf93df6d81d44ff6ba88859ff4f6739a34920933dfde71a32dc324b66fe08f1418ac87a7c3d8f324b0ff11d055068f8be049889dbc1cc732e36d8d438d974010924f01a81c4afe4c905befc31d1f3f4f46ebb2e5ae690e3f8cede737eb8e614d058f7306d8342b4f94a51232ad39a3aff8f22a3595e24c9af5ef8836dabe46e379313c029a5e3a38bbde246af6c62531a271163cae58e772c11c2bd7270147ead71595b71b183001b7fddddd1c8d52c9c94dd54a52e7eb297f350aa74e86911e8d47bda593d663ce9e1570435a9aa1b45068b603fca47efee06a9d4b8ae02f18e63d4544811ce045f69cd6a3a66f2581f996d9659d596bed6f62893d8fd6914954cbc93d0cfae545c317c21039f2068b15926feffecd366fc1559692209a51705e3f0a418f6e9f3ed7c8b80e139f120842254f88a8f5dd428cefc223dd526a06eaeac7d85a0074933ed2c2b72dc37dc5a425a0915b994b9e88ce37c7fddd4772121ddd419e3ce80327a142fdd1ae4eecb17c002b18a90662b0a51e1ccb877b0a861bd4c77b592935151950e5f655f51100347a55e69e92683fa6df337776ca1070d33ef27bfb4cf89c385029e3b8effceae490de26188c37dc282323f28a03f97200dfa0353cb5ea6578056b38d7b568efa4d200bae2ea21288c4a8d3cb8d634ba44a18b1af0851dd6450ef171294a23ac4667fc1311e44e3abd88df4d955e56de849f4174cb22391e3afe2b43516c2110ac7c12422c859b9aea59135ca037576282f9fbf1cd914b7636188924284c83f16a1320d39051a12191d7000a8b26cecab329b93ee947474905201322efee15e3de0fa7426060af381991313e23935dbd6a1446de95cd868f75a5cf568c0639edac7f234926a477b5cef4a8a8912ebc58388e1491d30ef87f2d0933732fe5398b9988bdf1c14be4b59c3cbac77efc7bc22cae42040ee3ea352da635cec10986b42407e516a88cdfe6377700225e59ab4b98fedd2b3901ded05f682e6423907cf72e9344a10f8c944b3de87c184db8e17d643ef5195445ac519b34b3937375f061b3ba3c710a7d1e4601e1d29099c83639032003ef6c53f8b0b5eccec6545892b32bcc61bb74e3512110c4dc512b9be8c25a1eabe65ba1cae69d408e8686b9ffeb9b312ee5467d0a1bd710f762ee9cf943ea5ee68c0eeef9f9690496d19020a21bcbf7f866897531c42207056c494c0e27fa590be2cf2280e8e3befea2c0eefb8d29b82ab7c45f6fd2157246fff0503188e9637c53bede04fb48c6436b42b2e2b2219018a2ede95c0e9d18ba4d1bdb63fbb3db91e1d88cb9ef82d1b9d7e29284e7a9d5da2a9335af1079c537d406316a8293a7649c09b3525eda5d081d529a619cd8a120b7b0736afeeb20955a56f8096ef3107885632ecb1114772f8065595e9d8007d17c6d3eb41e53c27f32bda57cc48a2f7dbee85c9f9;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'he0eb329f0788ebde418e8eb934089a84a1881d759b0b6a697467be654f15ccd5c2c3c93ee23212b494d7856913a618b168e0faeaa73ebc2a8131776b4fca6370526a6e2fbc5a3298f1a6d6c7d90ee71757e59dadfa362f8cc9bec93400e3716109f33a7dc6f6bc2732c0033386980afab1ab9245bad7000a59120488ee9762b9c4016ada41011cb4f7b23c7b7d3a6a34dbfd31bbf4579d5ad25a371e8a0271a136c46bed73769901d924ab691795358a65237dd5156f58a80a5361d3bc30d73d8fd6ab0e9a00575926b5926e454d6abef174a18fa1795942469b0db20db86e2b4c9f145de03d397c05ebffe1fb9b56d4ee8226ca40cbde64ac45f0c5fb1e740b7d14b4240609e9baf5060e51ad00dfa076f7df5823502b219c5a35f6c9679c8af399e77547c298391fd7dbef7de081d163d9851e977ad45513c15cdf57f6cdc6ae9ef35b8f87c4c2ebd7fcd740dbf991797d6ae67195c6ccd0a28007a1f90682843a1815c98184b9beab8ef77539c28a6526a03c8dfb16804d81dc4483ba35d349aa837d32a1e252c907cd7db20bf7f65fd13ab054c05148f548d61783c40683e0c073a45e93995111aebcee859ad24f8b65b1d0a82cd73788a2afd78116d5bdb947f89e6b6a396e084c611fafce997efc8eda160610fb65ddb9c502141abd89df43c9eb50e264d745af5f353373b79a9418335263eea9faa57a635627cd43553479898f6165557705e5fc3cb6db9accf22127b9d2ae6c126d8a8afeb603e95bbfd9813cae3ccad483c98eee209ab6671b15af6b8bccb027ec3e20ced3a5492b552da7273f531a1f636c29eeea04955db8ef00e2b570e95d4151a2679a408ca68d3ac090d311092d148c2241f59600030264f279c0c0a2c4d8bc0523b74770157579d9fba7d86bab8ba2682218625bfc40ffdc37e2e776b9cb50b168f7231a2a3370f75f7465fcbc085841e95e82918b92607ea82af0feb544cab7edde5d5aa79916559cc6e99fb5cc819252cb6960bdc066000922d680b44f59cd43062807ff6b3953da40b2fec85ff29ddaebd24113ef9dd38caafd3aea0e31e15ab37c95aa81eb773a3e8ec7e075029cf679d70e2ab429902bec2daddc620a6ddc87203577d36922ed6a911af57d421a28c02d9f39318c27fe6e3ed7ab8e214ac86759d92c27d51535a1a99caced11d42c3e47ca3734daef8ab4fc5345a902d8373a62f724370c6c08e284ac7ed39a91e801076c133a6dc2d91aa92aa00c768f3b1bc748a8b05c568d5f365334d7bb938491ebcada2d901caf07bb09269f9b4b9ec9474e19f797a9cff80e832ccaf87bfe162d6b0d205c7968f16e5331d6b46ad4b9e9982a46add27e2ebba30621260a6059c2e79548dc2f5114a1a66b58b3d1a1ec906d046af64dc029bec76df4eae0195f4bf13bae25903594cbef0619820e1c5401a6ab9209319831509b258383f5887913a50b91c358fd875426f978f6fa72c43eb1bf64e35c74aa93c3cb277390a7343620b397646523704036d0846ad360567857dc4315b8d9556e36a8d0d70db3e20c25f51c973df07eef8b6bd93a5ec331a8bf1ea1bcf508881a3c129fb039dc42df0c9e2f09597cb0cc6aaae59bafa0dbf84d89f401ba4da6b221cfe003d53ae1c5969f60ffca151d24470cf6138d6240be849520855bd43de5e1c6b741b574efd153ba7c8ef181014919637edf7b28315cc03d5e088c52e20d959046524c63b59b4da0462922e867da27d82c247eb79309b876adfb6d1122a6a76305a7641dc6b108b183c6f0a41bbc90f6dbc3104cb0405204db2a7d102e2026aa924d940fd77fcf575d9e6e4d1c5272a9c0c701725dbe412973893f0b275ca6d9c2d1fa422a5eb1e21b3b0a0ebc745e8efa7efcad2b4a62f1e76b3273d0e0d8a930dc7dce314406be8afa91b34a6a9fe5c528e089b73a3a5067145b8c9c90e97c8c41e3c4a42cb2cb1a935558e42c0049a2054ed4e8bf5b5b64fdc973d291d4682d4be62af7b5bff9e65406277424e7a95970f8133171af8f78edee4d86c3bcaee3df9aba22e1921524b0c1aa925d28822ced6f1ea276af06678346f9ac70c99b06405337564109a38824d84e7c0c193b27ffd4602560f91430fe302cf59cbb4f108b6fc57f98bc929caed14cc0a76e3697feaee7fc46c1199f0d43e7894d4675910302b943e6f51c66fca6cebe72720bdc9ff14efae3f7396541347eab93d0d8d8752542618d4a0739d69b0bb39ab5c85a61ee6acccfe2f64808ae862812a02d862b7818e3bcec27f2741926f81e09b26c7503543f819ab45f454717d544af4460c4492e498c47fa75a17a0f8866892cf9ea64e6978ba00f4004c81e41b4b635e04dcb4c4ad968ca5349ea96c89861e6d1a95f59e74fab523d1bb9608a3911a03b2c74bb5347967af439f8f6f6dc31530451f77e199571869e8661b3dd551b0f9a12d155e743f43d045368a7fc672914edb603d6519fb780d2a80d180bbfca916bdbd8f956132943c1468f5e228ae92ce50a7bbd96049bec650f2983c85536bff55c76dcd8970ec912da82415d6ff5998310614bd359888c6d73f92dac5c304baaf04861cbc474cbfc55a46faa470351c5ac9c5ceadc848023689d47192fa75c55f392938707f9a75b2e2ffd71bcb21d82c1cefb29719e6cd59c5c366b6ad124c8883fbe61ff41695420f1c9830acdedaddd961d35caeff00e9243c308d94729eeda2566f1c093881d28431fa341b0de67859df4da7ff4e7329aa190006751cc4c502490baab14ea53bc7d539c853b4b85d811d87c2d22adcfe48a00c86567f7e9d1c75b9697a393a9ac5f79c2472188f4ec360ae619825495e318729d5a4914b9a9016afc9e5f7558432844c20417c392a7e9149663c11a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h7fd3da96ba432de589ce3c7ca0a6a47e624235db4ed42811cf950fa5708e8e9d8015461642702483fd4ceab850ae53cc77a055b090ce6ad289cc0677439607510d7cf39666931fdc60dcfda2807b35a66b82650a3e240e0001d56e11bd1b39790e4fce801a4a76126236cbb4cf8aa835ca9c8c00c338693e12f6ee77c9b9f4d5a3fdab4fc9320c10688112d5037990642c36462e11b46e718227e0cdf7c74d49d1f5a5051c87ff006b7bba18f21dd0186a7e7450d9e7e81c84b487997f96f8669ace82fbfa9c17f019b680dd4afb65f7c3357dfa5931cc6896976cab2ed8f7916e481013a53df8751fddf93583c684f947f782e9174930245f47cda4c2c720a01c87a53851ac85c6606325892a925bf021bcf8f4289553a7a763636be36df0e3538fd60f6688e8f9372c270643be3b12c25b8c18a1717bc64dee956cece347c9a3026f4fccebb0bdb36ad354a4c9abf0c0c6c910456c7a6ebf06ae040894b0329652b413faf8df9cc282d3bbea4d4bddb1714166fa92479f8ffe3073da51ac02412e0340d327c41464779ea33301ac2fa5f97c19e664ea3e0b7be6dc2e293cf38d2bc3fda57e4e48c7b3f31247162d9fdc3f91dfb70ffd5f9c30cc365555b66297f3b1a673bd23dbcd9737d2568fa717f77f36f8caf2a7396df1e2c605f865088a26cb0473ae987cdf1c454aafa426e20369adeb38d290bc4ee505b427bc7ef8e8f92a3593b26313e6cb0331879182716b79f1fa02ad3ae657c6df3aeda692412f5795eee1e220891a286144dc2c7e9f15e12e144ef96dd4e8fb328613b054f5aa6dfb0a85a6ea72add83532caa0fe687633d466aab115953e77472aa227c071b27072664e841f56008d6b98e8f17f82dceeff09e77e8c6b21b838b41ca8dafb31c52b8a08af4f981d50ebfa7c86b2ccb72b67f9c487b347e1b33f4f0fbdb08b39e234aa7d1294c80430c72e79fc9dd99961909cd67d5b59904115caee1da7bc927dc20fb24d8737ed8585bc95e58f23a37b7835ac86bc6ab58e237dad12d3e506afe67320d34bb7ead436955a4ab346eab2918e00c596724daca6320898e2755b19030f714ccb73935192ce87c4cf0c6549a6eb892859d396eedf6a0a3e4c86e52d60aa8b862df897374c62556b18821b99dd1be271b563cbc98ce10628568ca8ed7b5450a8851cda1421b4884be21bbb922ca72c13f444266d3bab233cdaa60603394437aacc75d197de2e588d622dfcf5a08894e9a654c990f36215fd61e0a6177edd8b58fac8c6bcc49879d2156066dbc976b12b1dab3baefe6676e2953c6f2dad20f0e8cae9480b30c57df8995bea29865be69cead8d7b986f7323723333a9ccc658dcd195d4bd93d829d53f2999b8979000473f7c8979adf49f1c419306a3a4973dbdbb94a2b65e9b3b58818f6ce97b588851fc0d2d66f7f68175f697e96c71321642f4e9683429a0193d72fac8682d19dc036f8ce0daf9cbd649521dc93a16c1adffe7497295738adef215f694cc8b388f2bc4d4f1128fb28c17815a0fd787341508ef3e791e3b7815e99eb68250b2abe8d849b8a50127723ce066b5316345d12f55a925cdf396ce92afd2de092cbcbb0bd3fec8cb87ae6cd02393aec416f9b31d161cf35989f6c7245b02093109c6f12cc5463282d0a7998279875444768d8aba443aae2182b7f3ba734012b51160e2dcd302d42e0645d963e49ff8f61632ff1ef4a7130e288f93958c0401d5ffd60cb6598c801e16cee78340d0c302152de8e4a28259f65c775cdd082ca882e0ded3e7f635a18ef8e2b8c08cbe4fd8a7d15f4d488a369076a211749b3308e3fcf23d3c338dc598d1bbd03dfd4186fce866b550a93baf8f501298475d86c73bc5f8c977a45bc4aee1158719a1393535bc5b18d8b743f46e8d4dace072bda034b4f6bc23040c423b1a8a0e2594ad6c0651286d88451838b589fc635ade2bd8014972f96643fa9177c58254acd07ead0b9af2620fe8e6cd13ad11696fca57cdee7f56463a880a409885e7dd643ed07c2a442e7a641eb9d827919c346e29f041a07b23a0d05de30470496bbf9f6e1c5cc4a535283c4fe89591e62bf9b50b409cbd2ee6eb5c798e1af6c3ce037ce4a48ccb4c3be6ee825cdb8e91b4d610ee21ea54190a58221f245284f5bdb1f4b3ebfc9409adecdf26610be9b250b31089b95291754ac8ec962dab10b42374d0b2c60f2a7512dc041c04a30fb5e73dba55bf3cb81ebaf4c2e85daf044e94ddf6b207a5dde172a5e3c376f4198d8484886f6e88744692f8c4023c97acd66a5f251132bfb65a8b59fb99e14a5c4160d8f53e0c79aaacfdaa411abfcf019e759324a96899c77762e397f21f540c7b5e42f821c5788a49080b1034b8f20debc6b1b3d9fc3e52b9325d753b22f0c6310405a27cdd2045715f9864c0be05af5e217c5a8df1e70ad3e5f7e438ff39af755d0d68cb9cc1f459fba5bdf6771850a8e49f2b8a9d127a4b9de6349ef811728377ab3d1b0e4c9c4acca175d7b34a1f4405f193a459c968bee54265fbf60898c2ceed46643f61829a81becd1ab0cc9ceb44ab1f0165d3022e225ee876ae99193b7425f21e186b2221f45521d16e1af531934863204653acc98ddb98fca915cdaf4806b06049060ce0fe4170b0901d94b85d303ab92dfba78842cff305150ab87dc51e6f87efe4c5bb0c9302cf9d8a6c60e8f1869c97c39906c019805740e6d34f9179489b08fae2d4f8e8a040d701ee72997592b4c0f3402d7bfe6dbd6e5c0d89f01c2f389df1ff4e8c23d9561f82055c73ac49be9bf3aef55468f3209645a34e4a20883296d59611f8087437c3834adf9b96a3826a2c925794f4ee9c5afe7e4c00ae9de446133f9b935e497daa1c61f1c05cf46a402c4;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h405a682b1e176686b81ca3eb3951d9e3fc49dc3f1875f0b1f80e5b3ac94fa1e08f2aec5896dc1b144b65c91cc17fdcfdce5b93116a9dce772ab43bb60974a99c9d4088cee088594993c5e5dc86f9d523603a82502598084f4fa2e95bffb906c427264104c4e237b1b31e0752474b2f70a6dd15658e0520c210e69d7cc47063b3845bfd4219841aa05cec407b57c5937dfc5108d1935763d2ee24beece002a51bebb0eb6260c2679a49ac9a16c89bb13c0b8cedc9a886161826195a988eb50b353c6641108e3820aed1465015e1e857ab4a93b14b08f544e8689f959eeda65d4d6281885d4619876872a01be686db4a097ad23ff12d268a2791a277570dfa72fb290a7cadf7dec9d546317c67dc635712fe52719c3c3c8d958885076c2ec833b5396cba9d95b99ef665cdb81ac9f02b3687e0f15db0cae46162aae4962e92ef5df7cb129a1d6fb7b7aa6f690e389ef12ea4fd3d4b5fb2adb10925ccc3e6bed094c6b26484f18cd822003357757e48390f067cba31e24b0fdc598348ce04cd143e7c4d033a983dcf40f4820737ee33e23837b7243a9537142739e498882cb840a70d8bd8a955f4776203e52b0a413074dcb47ad8da1a892ad11cd51a252762f2f6d1862d75ab55e77bb07b6d1837a9d3eecc3161fcb4693f951732f1378b74325231cfc12f259a2988c124c1418f171ddf9194abd7a522feabf8f4dd5c448c8748dede76672fa0d5ef31fe505f743f10f7ee2c306e0c9e0a3d052cd2e8064f8ad190a775f208fefa8081907cc2d330163aa0c65a062b5ad11fcc080d3af61df664c219a992cf827cad3bc125cec24c0c7fb8438e9d9a25e7f78e665cbaec2589fb8cdce4bdcfebb7b10436afdc115e70abe1bedf729f9bc0d20440b48bd7e41f0a7a3fbf3c546170f47030cab3106fcf675c403c4716f211e6943846835d1f522a0ee7f1741a066db79fe57bd9d91a505c0cb4631ba132cb9045c4b17b05e30b8f7acf778df65c3982a3bcaa4168e05d00e36886257d49533cede4375f4a6dc435721912a4d54bf9dbf7e0973968ce7824001dd3c9cb3c360d56416162ca301aa700fbac270386ad6a7d38ec6cecb550040027eddfd355ecc477697ef0862602339cd37386110cc2ef66d75140022fef7e4253634f9d9ff4e89a14f974c9691597e7563b3f2aebce995c75599be492af4f1867d96a66e9ef5e2101b22a45aceb024fa8ab5b8c9d8217c7632eaabbb061ce2bad9e7dfdfc782a28d9d678f7e43776dd9f01063443e9b43f6aaf218cabb743c9c0ef289496a32d561fc5e30b6f6e6d1038d3b18dfd7f5c34284072390b84c428e2ce69597a2d54ed659070e9eca2fa5c1da592aaa97420ad103a8828230fd0b284c6c8b2e14550a6dda3155ebd1070585583b6532d52eafff4aab15517282da704e695c9dc2f76fc14119ff637967100344284ec1d6ef4e15ecd4dc80793407bc7db3544593f97e6f0be7db7b6040abb0d3fa4fff726eddb445816607c600a3057bbc3f46d73d289216fa0de2bf4f4ed93c8028e981821d49f2a65c55986fb91e5c8b8d7574be57dde4ff6a4e700483ba292c264cc1f53c0048e96ce179d6062e60ee51530fea2ccc97c4baeba617af489941fdb038f9d0a3820a140568a97c1ae2694120bbe2113c10d61630049af65a05a5f7c575fa4acecfd101cfb643eb03d36ce3881fdec97fe08fda080f695f97ad1e7828614c5b188337a89bef6a2f7d81cbafec3a681599f1fb70aae1c1b8d47f332978f78f57683585edb530ad42319ebc3a6085f029c1562545c8b84d25ad7065e82c71be8ddbab95cfc400db96f7098904eb5f8cd660ac52d8736ba8b56bae480966257c1b3941d853d2694d360d5fe17935fa246bb306f53495322756e968c5144a88ea06ae8acea053f39580349afba1fecb951347aba95ac95bbc7bb077cc47cdf33ac2141d86fa0899c7825e7999ca4f21b81dba8b210a37027cd8be79f482471f51cb1387b13e0a9117f0f4c278b1967ded1a99ab30978c7df6e0339673b678a1d3090f36114ef2ecbcec50cab1c1d302f5422d555d4ed9b352db5345c07136505fe99075828f3d01c591d9ff63ef91eaa3112eed6d9fc64d6bc56cff068e815c531fe732c8630dc71d61418d438c488070aeca6e32877a15f89e23b65aa6970d31ab30d93897f4e4c1813a00e7bf05c3c2e2536159a41aa7bc8bdfdf4c20b9f58ddf408e993e2b8477971eb6fa56f17bb239d55564a146ba17f401915b5e3532fdff4a486ffff24265ece9d674a3ae111231aec103cb3a8027fe8fc336e5ba54215ae4af86259e7c0ff89edf82381ed470b963bfae0b58e2e758edd0a8609d7b6fa107cf7faf62737de578f6526deb6c2527c6dbc8a943fecd4fa34e4ca4b1d523eb014cb856b050da2d2c9cb0e6bb20df473b1589a1780382cf954ba8e030f212c0a70f7b1a0d7ce6147c8e23f2b1ba735fd39078962e413a52e5781c9a26c0ce117f05957c49e77f4369e0a932e8705a984c97277b58bd7df6f190551dd6e5ad5f61d27ec8eaaf971498779ee1832fd00ec7fe57b13696076450effa6e3a9e50fe8becb099afe9744319c148db6364a3b0ef988fed7591d0e04174d73c15fd7ae115f40daf03e86b4922b07c13e1daaae6ab06a4d7ea6715161c68da29ad7b21188c74aba24c8e33102c7a14cc28d3a7de1eb6aa7942d91961fa35cbe30f8b25df3cb16df53e03e1fd05280dd46b2617dbc93cbd6d19b582a54784cec4e54b8d3b7c5893b4ab2e71e3e057ebe06572634bf7ae0530484b1ed3d1cff09272fb2192545b985d0ac33697b73e711429fa5195c264a3eed413d6d887423237b9dbb4256cc50f6ed312da101c1ce05ff3ed31be5e5aabc7cda6eec;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'he678e57aad56254e624250e3f4e5bec750646063c82e61504400709ef1872cfba6d733f6b41c69c06a1502536b3da0016e7ef0fbbbe4a7e21396948d82c68d3e199d821f40668d060240d312470f47eb8d5e2798ab72ecaa8bda93b482a5a213187cf540385423eca8e26471afee2f699a4aabeaa3a868f7aefbbee05c32aa39ee99b1f35798fddf641b4cfcb99bdf72a53e7cb22a7a539cda993dd2791837d4ad72f013f1be2aa545886a4c00a0297fc9c155f464c218e6a1a5f0931e23dfff8951ad35ddcf16e5c08cea7ef35a4b0ab24dc073a6dfe5257d7c7d2924a4616acee6de6e25d6bf475f362d3cfe86d3a84f3ae8676baa7dc47cda1e68e7a2c57b1e119fa13d15daacae9ddd49c86669f754da5d06521eaa5d0ae86be44e53a905574c8ca7b66acbae709727ffeebf8b1947070f7b2516bfddab23d770e3ac688c28618306e5500ac9ac2185cccfce11508d8033c757eba37ab8c9f69fd2b7499d0dc490529a03d1587eb0ede259bf12b3260de3f4607e8f174474c013da362aabbbb2462dbb37af91b018bb8bd247d221b8d05d64d9e2405316ac800f2675f4ebbf1ed8f6086732e6a54bb3326dc6877a3e118dd0af3e2d3175396d4a4714bb027b2925b6a25a165d89729ea5518e7e826ccafde77956c8149e90ede168b2c316b9c83cd53bc3224ef797bb0b109d15a52122d88df13120c4d7b376ab0e667e66278f991198f8393cc48551f8fc08302d4b366a67459fb39bfd65601b35950f1dd59326fd68088494fef60c942abb23285e12d968ce2e0a847fa7d80d8607a31ecb5709fdd840397bc80ff68fc8fe0e4336ad2e86db050fa13ae3c9a806b7a83354ede0bf119e2056f987cc46e8e0ee8f33f8cdcbd902e6d23909c5b21844f1451ac440463abbc90aa99692fe4219efa10aeb08db2c0b2475be6503775fa7c9638f8e694bc0c043736b7fe01b7327c497569714a3180811946d49425c0840f02ee91a49046c74037634ac5ff4225d1fcea82c5457688cf238a87259d0afc1150c2a355f66f2c7642102efe8be0e70412ee4ef418c3f59480f6fe498230313e51d559af7105629ee46f7806ffdf1e4884cdd80166fe6e45ebd23b310c7734968e2a67555bc4c6c163bc476fa9a270b63f62223ce294158f590b158c59dbe70ae85675676d2f8a1fedd64c9a24f82563f67789e4aede4fbb6f53dfa4f4fef0e307bbc933b3b854e89f2b424d70e3a4c848a8e67206281b2dca5f43273bbb8e7242e0947e4697510aff24c8e0fec1c1c116b121c3e8b9491f194e89be3c6d41f7537b8564605d6a31407d44578456e9a675849588a5fdf4d9cab969663d530dcdfd7cb36f512ab0291f1bc87b19f46c79c3916cf3e105083934ac7b4290693330613aad3163e3e783727dfb3201279b2cc220191b8bc4c4da177f246499c9be9ac5160daa199f55dbcd275059dd0fe0c73833e538fd598a72f10a2d18f46c491bcc672f0b78135ae0250487f86b2b81c77506a6f3ce1f1a64402fca5e49b63cbe917b8c02898d3482faf6f537d3998a2620d765b35b9825f66d3ae4397ba8d00a93fc15f447b5a9cc1f3088ea1846bcb87a3094fbade30430b8ef1cd7d2800d25d8d1af3561fa7dd15326a2137bc9a0c3b6a320341d2782d11fa625d6433ebcacf5c39e50a76fb1b15277ca41a0f37fd9b18411534a6f24e5d91d2806212bdfd74e558bcb47cb9f39eea67ddae38152d0aac4a1a1dce0a758b5c8950c3bbc96c13ed5ebb7cfa1a155d4385ac415a65bfa6101b7b5912663d6d18ebafa128cdd9603bbd69c7a1ee3ed2e5b428992b223186bc0635973e8d438d2847da3d97781e3edd58ccc6a4caeef12f83081fc6116be39779936befe50e267240ac10b8a26679f43b23b26e492558cf50efe8162736cd16dcc30d7c5eb2dd6c912e95f8ce2c4caaca2cc3f7564ee57a225992a8497ef1ca9e0c45af9ed687442abe48b53fbf70dffe67c7d2896637769e19077c9090dc4be80469037186a0b2e93ebaa51c10d301d4adb472730d0ef5605003d1bc38040fff337775890b4633e8ba4db1655e19547bb0341e28852a26ec6c020d2a2b026f56c4b224cc2dd683578cdfa69269ecf3e42175c17e814b52efb10572b1021f2d4239acc575c7cb6ca79d35d8ca29d51c99ac3afa84f744a6b9406e20b076b41eee53400fafae334386a157c5f2f93cb7df395f66268dc36dbe9a42349a4e9172dcb279de48d37b2c62d60e92d04dbad7d71f392afa28ace3e693cfeddbe74b0eb68625a0a0d7c334eb6b846d5efe847d70ea4ca95440706303913ec0c0f3a55f4499cd887ee56eae1b783d3d30f1375e652b7a5a914fefe042cda8c5a4af9d5cbbe16267b1ab45ebb52e9a4c9ddd98bd2ea2178a95c1a9b4850920e376049148dd8d111b4b3d09b9e08c6c558e18ef11b77b5618246aa55a5bcb59e228c76697d0ef947ffbd5c0740c3c2058af32e1d66d6c50cdc9fcb7a1c0f9437f33daaa37d6a954616488d23234f98a4b76ad5ee02affdf3bb1bf4c00ce5b2bc077aa9eddcd2131aefac7c1cdce1a0aafcfdb939b98d94b4d991d70132a24e8257534bb11632e1cdce4d0296b5d13f9379a957b730c6566cc37734fd7d39f265043297ca17333117c13f208da9bcd557b8fc993f6c1c856f26e89d02cb69d1675d4e53cc46cf6b6eb3812f740681c2be994e7a23c1ce439561fbf0a0d21e84794a32592df8d4a153219cfeec7c0ef9568275a0ee310f1c15aa42dd75c75fbc7278ae02d7db5871fc86d53fc9d0cbe3dabda0508bf1bfa182547d4ef58ce87d15058395ce6cc076445d74a61e40569705cb4285f497f97f5cd8e6a4b70e33a9eedf5b487a397a3afede76f3ae2814dc9d6f15fead2;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h741e43043a454274ca63db47a82e3d65a6b0c623555664ed96c1f33ba20d4cc49e8aa2ba987e86db26ce16c8cba05b1c4f849e9e98131d58f49276fbc9d1f791ac8c4a018f37658a755cc7bc28f59c79a14d9357ccc9772f05f7e21bb042b0f0012cec326567c424c96eebe76dbed378a8f8f65cd58c3cac11b95e09395853fe3cb38bdc0b8cccb6beb2ba30485284122dc92f7b6694408a9d45c0884bc34f823e1007b1e562311b120c1e7856836428e84f470111371bff96e626247bf83500854dcc9d733b835d2f9dcf7fbcd1656b616a5df8439f304591b45fc9e4c32b716fd11d0d842ddf9532560352beb89ad023d333d3afb0b38ddd451a9079654d81798ecae1f77fe53b95167dbd420dee8fd743e23794f9d5de8ff135d35cdaefd07b6552095d4ed2c55d4275bc1e76f8e56dcffe4fc57cc8ecd593a63076541c50504eb2daae624cbd213f05f13494928718cfad23412484d4142ea38918df3adc9d045c8bd57305af8e7a516c576142288fe6ee5687551c6bffd5ae7ab0781ad698b0ef7c6087dd64d11c2c02060b9c094396439032c0a760d4accb7f7558d2e67d5b0048eab3ccf57ee0ae9feda405c299c2e4c007285b67d4645b8bb645d50013248d420e2a812a2222bf8dad1020166d70c5e4306a6669de931d17348f8dc0b3992533c1a3764711042f0a0f5f93170647f5e274e0750fa112c73dd6e7ad79448668422b9d939eae2cba64c5c46c94568d01389dd98ed6bd83355d81f69f19af7e313cf466286b84bc1c1a780c2bc40312fa4a5092db53528b4e45624a520cf70fa030650a822a4321f76426479a1b4c1ab06cc0338ac19717a67931645dec003eeb75cca77d69882b0a4678c4cce89026f5865112ecd7e6f9124e97802e828b3e20c145b435f5b731cc4034b0838565e22b1779df6a4dc9e789d5c9795247c491a909b03f05e8dac5aca1edabc0ffd24634ad90cc6c840c906ef6b9318712804c78f52bbe1f99afe9d9df9cecc6d33e53b7325cd3b796844f61bcbf6cfc63012769c80e46cf5412bc4f04df79d3091d21f79dc66cfde532361b94f52f060226e52e01fc9dc8ae4e8dcbb48c940b970ef0dc4f3e68884ac898f11b6dbb93be2cebf9609f9dda07ef2c7aac39fd7c1743ea46594b954ed5391e5f9ee51f6b3b3a72a36c21ea196c3a3bb542ac05b27a8984852edce63b3abf6d2c97c5555176114946038b33e6de3dc7a621e2e6d2bf98c4e51ea60855ea4d0f72de684ad434b2dac89cf7192a92183ffdd971789e9ffa0678ca21172be5fb8fdb624d49b5162349e11c6c34ef7e7b987068e298d7a692d59eb7b10dbd8bc9daffee60c4081d93392a4aa8ab85234658264e4f08db6d0b3f44ffe4ce1f427c0cda1d46f41b5cade186160813b8de3b151e2cdaa8426caf007953b00e31a7c1fbf89f2f2313c0563e63d07a6820dd67a9c02c9eca634da9ab878eb055ddd2290e52c6925e3e655f8cd70d5312bc3c54fe427a73ef95347c7735760fca118d4e8a0707bf7230ce504f62e52264d73a683435e8ab688b14f2c89525dfbf6ac5954e58ffacab4bea54f7bdc4ec4a1fd6986df94b6a67f07786b8e101307c07bafb4d3515e627ba182cba53cc368184e3679f189b889c1bf377f78346cd92a441dd1d9eaac4366a60b9153c0ee71c7e75ac679c54aae9105897593e72b8cbc3fa708f00db1d19f7b7b341852373a3b311483225488612e0c9e767225de0e6f3fbd01a581966f16eabb0a57ffe33db09fb0de18cf417e46067926f28a93fd77f412016550ca7e6a580cd79cd800346b93330eada167b89314709867ad17b631e45a5758e103f025bd056a231ee192cf3f74a72323fa15ad98b3632faf7e3986e1ad336c6420f61b755d553c06111cfc071c58bff677920df5cbc65494a6660dbedb4c99c24ca2acf2befe502e289f48cbb730dab25e2e06832a3209194971b6995ae09a2bb1ca42d0088a18846ad925d16033bb092324b4bd44d355647a228f3fcbd431a976f3f084240594c0e6cce8a1e872e98ddb50e7c2e1c2fc0d7f9522222b566ba99a5b4e5a7d74a8288b3b812d3cfa9c0433ddc48df1eb0c30c5de5164a2d22444526399c6162ff0d4c15ed1deb50bad4d2ad62aef20f18fd7ee2b6e0309265986f04c6e5d7e8369c2f342c2269d3b80b13b28cb004ec3bf7b7d944cd50e8a6b7e35763dd2e55ddba4dc66ccc6ed7ae2de6aa4db34c52357b12d273abc1faec3530e076cb1c0335c51503b8fdf29616ad7c400ece2b49aa28deaf2c11f775d1ecff303cdfa229e408e8378e3e55c4b553055176421df63d37a42ebf412bfe75d35d0620d10f24d0fe7be4372b4d4d640f263fdd4058053b96a4490a8dcc8529717daabe7c3fa226612e5ad2a4fcf15fec8319ba685cd9d614c4c1ca043d616f2da514f48187953d90ad56494e65dedc3baec6cb66b6cefcf185f220536d334343c029881e86b95ae544fc04a07a1b4a97750e703a164d49066cb0dae160dc08d70d1559cbf3c58f0f5ed63c4d5697f14955d07b3696c776ecabafbfbee383bd67d60f87bebb8702963f644c0175dceff8de12af415afc933558a3c7c82d59208637d78b78eee6bdd0ac43507e658ed636ce212c3a5c46531e5709e99ba0e5bfe58b356062c1a3bd219836f6ef01b837a7de7df962c6e76cbe124e5322bb1e59b06e658c64c47d638e535c5e41de155d8df3198802a3ec21bd74db208bba776ff41dfb8b53831e80ce5f30896ce7b9d0b07f78707d96dd3ab293eb313b13ebe0d2fddc182b628dac126c39b81c9e4af45ca499b0f930293c62741c052dc3cd431bad1b92064d933801f30f473a7a1bc503f9ab44156889389b9509910ea127994b99b1eeccd9;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'hc459b28c0035663ac85ea665ef2dc6a53accd2f7aae9e6d6cc0dd838387ca4f8ee124626d36a45b041595cf61a48a1683132356c2fe21bdfac39c67e6306a61c6136ff96c1169cb746473ef81a67bed3662e046f4079937ac5ca3362662f923b15e950d40ff1fe23aa4a76be8e48af7f3e3bb14deebbb4751f8090954ad2edabed00f9259916b8ec7d7e1dd02676300071fded6ff8d0a37fb775fc89281d0c84455c0c20758bd57dc33f4b62d2f22e582df00ac13caf61bcbdc824d263f12b46933209928bb48a0eea80effad57e07d6143930366af11a955fca8280b1b724ce3f323020b9ccf4aebfc4e88fde87569e6818f04cf7aafcf3708ccadaada8aedbb504f0577ebb10364ff5055ddffad58765adacaae39742265dc27e884674b47268fffcaf2362ffcf46db1bf30d70b8890c787947e58dc243e7392b233c0dc5df36426a281d80ef546199954d50a825ebc0180af7ff148e323dfc2e5092a777797c2c533e9dd85013bbdaa56a4aa7d8f80ef06a348e89253ccfee3df8e3d31c94c6fce40737b8a90cf498a02efd2a17e96c50044a914f6d5d78cd7eaed12a9bd91f6b2efaeaff75a9288d1db9fb5e27c62eec27ab99e712ec096dae4135bb09ef5f1a3f8f75a0b64b21441488f314d7ad998bdb1177308cf7b95e02e1463b000f958a1a30c5bbb57642feedf1ae3e21ca83b62ba03c8515a672c40df3c0761e1602931cd968b2ae21a7219eee8f410fe58d6be4047856135528fb29d233b53fd24cf991dc6081d3242a8a83c527b08025b1302a0a5cad63c3454201217b3a7a4974439bd08f80e434497ee732f0c1626e3b8d74031796cdcb7a682868038a5d51b3834837309ec3946c30f03f76b7ab2fed8471e981642d308ee504f58cb6e8adb95366a7a6304ad442eab61653eb3428486dda582a0313fea3ee0f4fa74e72a866fa15993d7b2328233c6bfe6bf56d704b5669b6c85bd51b2a2a309ead11d765031851bf47140afe205dfc3bda9a1cdfcfecfb0792269405e9fbd1abdec3cafbf2c9a9dbfe2f32a54a24055d069d4e3a7b020b737ff0bfff0186a565772ace8153a73098b0710556a02db0b5eed373eca8ba290f08128d7f187fe23712342c7d7e41799c5245f7791ea85aa734f70cf657986f23f25eb5c3a55e0b319fc5bd6e476aa1f0439a118d28588fcf99d98afaff810989ebec70eb548bea83476671c4c633c921db91cba003d2548280d3ba85fc480d7740f9ab7857c56d2b8171d214f5c4da30844b22d081a4a6c78a9267be8701bfff8a1167ba463750fabff31c336db85362922459a759106013622229fa14edace0df257f8a13cffc975ce24b7d65d5f1322cfe20b62ea679e60119ec611e608243d4c65e29e29f30110b710e0f1ea8f37cfce8b3a7ff46ddf809b7f79dbfa9d487b3176558752812d75472d805e7dcfd0fd0caff80db74d3b9b1298fd5c24b7bbd00a045d740cee95305fbbff18d2b17447098c447a01037e844d575d5249b71ea8a49a54b52a46c24d1f165aea64eef619302066778398074f9e72f9691a104f32ddedeaa9707f44ddc3746ba1c349d793ceababf3b1b65b1ccc56d42947c6b8e5db7354508ec7b7e91540717107fa8c537b5034333b9a0c410229b777edb44486b2fccd1a7e09cba7c707a8f99e9544d75af5409a6c5748f84b6bb63c8d0c0ff546d3e9756c8d9455acbd4b7a0f3e1fe2dbcf4a8904c95703552d069c28535715adf644082f6aaf8f131cf76a520a06645d20362e5875d5951d281d632938ba9d0c4874963635479bab0cb1e6af8685d8274d8466e98489770c7b5251daa17b6f2a85e132585b98081d693cde83bc37da2e1bf0b5514495ec44b1dddc71de6006c2599fb683be596c6a99d126467590fe36e9c96ca3ac5725528c88dc07ef5af0f4eb0d626953c67f75b48ceff132a96e602d39a579f28ff43d59d270ba99199db8e9b83b5d7b4803019118c8c6cdb55e1c4f4b21e77443ba86fe1e372467cc379860f05b5a6b69889738aeea5169cdbbef8a34a564e09d4028aa54fc9d1e4400e1905d6f76f5dff709a8a544b0fb88192b61955d1863734cd2449b9640487988a330c47e6319c78211aefc5b9910cbcdb26afc9566e344219209ad4cfd818f5b1204bc50fa8dd146a720af617589d989d9b78961686fade88b769cc084f2a42fb281e9d72831b63f0c36f8818e63e20b3c51a4e81d44852696994e213197d9988c1893d9f697335a95eea9cd434cbbe2c27588a5504a5f2ae525bc7438b8e51f9e2dea52ca0953012a611eb2457d07351ce3c3ba6242359d7dbf860e1b761b5a66152e0ace0feb5df8888b71369d461d38ea07ce35ab83036569b98bee9e2c858cb06b5991330e96e2a5209482559dd73e0c15b2412e1dc8e8356638d781efdef8f9ac55e8bf5afcfec3ab107c9dfe97ea7b7561b8b092724e3f7d67348b28ca634b3f2063f5c3b9adaa780d59474aedee6d84003ed30a1a0b872655484c66d284a5dc71ad75e932d06f4fc9d5e64f605a7ab87870710be16869a67f665301405a0101c3b1a7c14766745e440bc709b9f41e14ec4ee5e8e772e1d85a234b67a6d23401b9814a4dd60adc6ca3d354fcbd8ef12b88ea9ed06d0ef74a029be1cb2120a6f33010ccbdddc507fe159a55a1b705df6a49985cfc05c77fda17bd65aee19744e780961d67ee8460d3e6986d7436d2d5771f71ce365d6ffcaa74b528f83bdaa106a24ea98fb0a87f81aaa6e24b0b7014bb95e5d45412b3978069cc56c67821c3c1bf2822541b9dcde8cbf2082441d2e2c9adfaada7f93bcd4af42a079fc03cac519bd24a4def2c58bdd18444116591bf89f2020b13611b5a87c7003a537ea93cace5bec6b327a307d5b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'hf2dfd5935813749f4d76ad37739cd5f71628a3dfa3e0adef4c709d350caf0a46cd5f24fb7d81f2a5f4f1ebaa9bd83eee30a09a2a19c278ba678e9a330fa50c50f4510c41ffeb83938cd8f55b7bc299b1509859efbcb9084e91588db995184d1339651ec4feaadf6d749ecf00e43d662b285408c0d90dfd762e11f060ece8d6ca1187340541fc9022fa75a0b3283223347c67ebb0fd8adcd17bcf659a83ed7ce464b14796533ab91afeda188ec00cb695f76b8523302f721e0fdf85a777df0b1ee97ad442ec08ba2f35a98034222112ec24a77da6ce7555071f29906f414602b6281fcbae97d797d54c55710e2c0e4a6940c13ad7c3fd1f79f1a233a3910c8d412a931d5bcac409835e32eb5c3bd9efaa867d67e9f7369c5323868f2cfbfb79ee5b45428cef6385b641038003065079ab8f1ea726cf0c4603c284abde096b67116296d2be74fd0c5e3c187f16341f293e0e4fee59f3a6098935f2348dc3c53cb667597c8394a065f28066819736a59d9ce6e5d6fbe10ada589bb8f00fa7932d5427516cd6d4e61661a0208115bf53fc0095ca9fb75facfb7eae7c0f7b68933c1826203130c98c7d049e3dea616e048fac2049ab9ce53f2bfd523b0c27ad4506704861907d3b94b7b65d2d3fb6ef806f021f0857ec5ff0c567042f3056381c39079c0f524fce223e20ba8717e596450d6a2e169bcd4338af5fb367d3827d6ac66b11b3ac1f05ea33aff29c285b01f2b6e16787174f1d8d76c22f2b127fe2f80d0c061adc6e2fd7b67f5037daae0595cdc6a2d947c8f6d379e5cf62e5563072ddf1ef81879a6e68e239a400e2f87abcd21207714b72819b836518d2358a5a1d10203b882294184b2e4c8ab5dfbc581d4faa82951040b6ccafe72518c4b416ccb0713760234cac9690593574303622bc92314e19bba503179a2f9bcfa4ebcc995615234b1885d9f75ef733c4ecc236449c0416814dce4b86a42fa0ea84d7a53babd3983d74c7e754afd8b68a148057b739ee17595770b23064760e819bc90a77bd0d32c433216dcdd5a81e154d44ff16d24c48f428c86f2c101afd2c92c5f9c03c2184b6c0b7287db103c560c984f4add7e05a02f0b9c1f0d9fa417cbe3273db5c77ee535eb1844dcffb9f33c7c2b1703cb6c9bab12792954de16cd691c22fb4904d1fa3a65806972f66e638ca9995a9e4c6a7138c69341c1f8440c96147b037cdd4477d78177e1e9a388914a5f65f97b2ecdb0f93bfa5eafae95782718133e2bf30a0622826e5d13feb0d3a1ec394282fd3d60d5679c448340320518923995b10ae2ab348163133dd883ab1afe4b0a06540ff575e44b1c38ea2f35fec5497c449bb80f8c93133b973571ad4c0b14d7b04428e044909536b2a0b63a4919491b994114d6238eea19705144ee8d7fc8fd700b6663c406a8157ce1c52e8f2fead2463ad46521479c5005981b66faad7b2280500a9068c9e29fce1dd86d41ded906185c22794ffa0ac31a72ab90e55b94a353a7431666bf862ece67e28c59830fb9db12086bb3a92576c6e493d8058dc09276ac22b85de21c24dc6b5b04d54959fc9f926f9ac032e9db9f1bf79b33d0fe01f60c3979fb91d7e72b8f79673ae7acfbdd81b87fca7aee60e99ba6bcfc64f2d6c88e11a664e72aea196a5a5e0017546f9d5ede078f66581fb9733c3a455590ccc5ac57631169c03de8ca8da8b8a87741ed86d33b4e2076f4e388d0c2172a260ebfe8c538c201f10a059beca9a217a7a01e94eb8133df02332be93bb2c5ae0d0ff8ba5bd7018d3b8b2272c5948b10cd72b05b78033d8ab72c1710f58850426911f2d8d8a48633fb91c65e147143d36248a3c3f1d4105a19dd984d43439896dfef3dad55ed28e7c6babfa63a69f4975a9983215c1e394533d459b8fa581aa71133f4d9197b4912d477a49335fbce9f824953a67bd702dab0b1bda2f3042c83423ed63e7efe901c4acbdc170b5e4067135364211c58665443fb73f20db9534e5d89a961abd6b60c46e9c25ca035a8a7d4ec403e436f240a3a053af28f5a390c71a60f1b0789d153c3b514cd5545ee5934c13dfaeb14fa89f6bcc00ead2daf2ec44142dd3d4c9b1184ba3ca93449435eaeacbe3105081a68eba719f00f8ffe122bbfe42a2019f51c3af4541d920c5221373ff4c46382cbeee7625cfd4ebd2d8431088e8aea946e2327f844b3f63e69052d60ee29899bd53f3a9481e89833559277d8b2749f7cd9c17225be02a5c0690813a94360a543ab9bdfca45ca7209e58889ce60c3e8c7e2b8998175b680dc40444f386b67537f4fe139b06d4cdb013e8dd61b6d35cd09b483735e2fef9b6b795f7a8d2702d1ff304f40055c4167848adc679d3ccd34b1519ad69ae8dc8e612777a9ae9567df2b6798688395a3cba64be1ccbc0735dd4348670421a95969df55d211716eb68527f1deebe6c837cb62bfb8b57871659e32d0a9b8c197d8ed626ff6feb618017feae89a1be2c1711ed24346092b033e8f80d9f484fe04f63d16cdd891093ac2696527742164a1989186e23de9ac664cd7ced25333a37ebb054924fc2485c443f31a4f362716e93dfedda22e5972616313c7b3c5c365578ed5399c1c62ad7da8f1ee29a61e3601023b32ff8fc10e0f73e49a08e410fa71b40d0f2e0f20bba0c5ad47bb7f7f4f909e67a7677dc9fb39c8c1f63916fadbe5b9daa36d910ed6773814c1b7a50aaea934bd7aaa81834d0b8ff3b1bf5dc6b5936c96876bd2b23e1c66edfb717941d1e87fd1418efa442f38d3c435695644390f0ca8e2a39ffecbd10c47e71cc4a0a801026d914b1e5d0f47029eb6224a39c459f33b7175f1324893eea3ae547cff2e524b5994984a548fe600a2f7b0c6dc5890b044707a16cfce4a392;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h45ebd0d57ed196dbff6383cdc6aea2ea92637801bef47cc2cf1e601404066d740eedcee5b70b107d7cb979b9c6e02c2eea4a1c579816b8e3a054e4fd053aa4ff6907858d63f66e792f6a909e7da81aea654d0165b42bed3193a6a2d6af95a992ce237ef7486a5f53c548df4388bb071b967abe62f64d6521d90da1ff0b30312d26d174af00f0f6148e5603c49246c2de2623176fbe14a47253b526b6e72f3aea491d40e59c639c81300d42afec5511f65be452faa192665d705452677d308c0a0a79a8500be549263d1415f054c72892f3fb07ee8c3fb072f4755da4c177a65dfd270d6b4d3622b25487aeeaa7ced3724570b1e054a82c0ab7dc325234fb017a6bc1dd8903cfcbe0f2619721a7de6e0ba2d224df145efd6e297acb1020edcfd149aaa9a8a687b5e48f507eb690ba12eb50a46b2a25586a9c5b79cce0dfb8d8230a29fa06aee4666b95a113aa037346774fa92229cc5c7f268ebc351e6b7f60d9068b7f732d0cf53ec30b3a433cfa628b0c8c7edd43ccfa40590daab68f46ade3280313baa9ffdcb0ee00ef6128ed85922ede8e6d2a00fd107f5379f399c1877e14341b32a2f2893ab9659cda9b01a48a043d04b5c38e25c78fb26797421778f3fd1024df19c59f11d37b1946b8cdb5a284a2407372201ec44b87d3d559179cbbc49ddaff5e40b52bed0d173949966d94aaeb42b3d7353a1e5665bdc8b2050648613e286258408576fbcdea55e8e6f28c7a7e5595549b0a1767c90e66919418085c8167c24130988735122bb92cb3061ea6440772952bbbd38edeb339e43be4fcfdd1f6c4d6daa20a3eadc513c3ce8ffc3910231250d89b52a8d6c76e861807ff822c21334499ee6996707b9175f9de04e88f114c29692d91f4568a856603cd97f4f63435c82dd05813b15727acdd07b3683ac91370e3d763c5e3b51dc21bcdb834ce2b5f5e4e5b8ef61ddbfdb421cf5f818122f15f36781da2c669aefd196a65068dba71d9b0baeafdf0399681aebf6f893383baea5698d44cc03045fee0f9dbcf80242e24702eaef35d45adb6d57dc9a48fddabf34ad53e32dde0180de5deade5f3ad046f730b8b38d58a5642d615200d9f4396cf027f59a42bb5469ff4760289aebae5ca3e64eee80e09a41a4942f9e76eea056ab8e96f8b4b8b0cf2919d6234c235185b09679dd8bb49a4b1ee30a673cb9439a5b2d9dae0ea0ce8ae12000637507126843bc8ada484ca7bf7638119398843a0231cc025378043860e340c128ccd96ceb495e342bb4005beca149bb2eb91363af50b6c670aba882a052a0b77912754f54d1807c74f7e6b5442a3fd7f61fbe20069f4ee5db6c9b94bbbc299bfeb0f1954af1ae83554f3d968798ecfec112d37545b2ce6dcfef2eded9b16fc5ca9aa5cb4d8ccf3ce18cfdfc6df4b933c3b3b1ab9d7040142b5c64fd97491174af7b56c4d335766be2bd59e79fabbd08a0c5ea981662ba045bf05f6599ec2136c280f16aaeba59dbe27c5ba1fdd3b39bb68a14ec23a64d1bc39b3ca6af8f832a61b83380aa683b24b3abdf57ce11cfd0156381ea238dcdee111d0b9f653f7f63d2115db5ef8e5998dc9591cc4f8f4e55a14a203a0bf7575efafdb762c141c81e0a7857c2ebe0bd0ae1be32aff63f0c74cbea25da4fb66f2b00ad3aff2bda999a51b3e6e76065e9f3d5ac24537db6589ac816510e19d465be3419a3b46b943fdacbb27da6a2ec94731d49ef60c1087a1b3c0778ee1691b3f98ed5ce83acc66d125e92b8f1c87bd55c677caa863821b9be1cf2bf15ec188dd2adbe6a158730e6ba55e34f4ccb62a2872fc2b06705d5a135fab270422c1b06fbe2f4efe9dc6e2af737dee0b3248671ec19439207ae8fe4f7380217986817c8b56c4b39314ea6031f899682b9f71a166eb6072473042879e7471c73e95746fb918f62833b4207aa8dd24362cb5333898a4a97107982e6b5ae4af6b2fa80b18953640abdf722421ba11ff92dfcae07205082f30e257f8d036dc746057e241fe7c935797830276a2c02fc579991f6b379a5abf87347de48ff7179891b47fa04d85996bb6efc629cc8ce0353ba211e1a311c9ed1d60dbb00af4238672ae536f9bee21f63467f8c4f84efb26f9ae1ec3f8d4f3ac6c3b4d19338f739584d8872ac2f7edeedebc3dff5cb1c107c7fb82312fd257e30ac66af94c3b16accca8a16872ff01a761a90cf20f404f94c4409f0773dfa33af9624cf83f954aaac7d67636ebf8563c5fc1bf37123a66ff436a95005d1a37412c7aa128e0bbca0a732a70610155b3074888a5806459c5f1b71aebcebd21b9ed152215905032a8915a1e7918a539a4bea8e1d45e3e9035379a426801ed47af92278e517293843c9c2466c35625c9aeff8ea4c6a7583109202779049cf2c75d5405201d5adc0d33da3af2ccfad6df42c1dba6f1ed0d02decccee3d119378ee6320a6ca5d0b88e93008b8744d4f8bab97aaf99d2bae02eb3582d06b52f7a0092b104ff0903f63c0c766774249a4d0303a944578c9586b7d62b6434f784b4e7f53665ac535308ac2fa1067b28d80186953108281d49b80d9e124f91d3efaea31d3c7259a2a14c6986e75ff4eb7a05514291f4788add35a82ca08e7cfb9c385173a129da2e0af3619e6241015593201a97ff41aa1db35cf11432726d03aa7ace37d61875c2346f3b170205b0e7d56561883f74788dbbed6e66fc6ad26007a5edf7eed080ddadbf708791e7d80279d6b60947c4a73d5c6f30c71fc4d0f10a17d3c3a3d08973dcc2e71e1c299625e4cf4c309dc0083fafa24420d35dfb13b460b09f1619204cc02d34740b8bd376f05dd0fe7fc1d36dc52dc3805ce7c78c4113bebf66f8c486dc21c4732ac8be2a7450157867d5c207dcf3701;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'hb9e22cef1c864ebd901fd1f9df15eae4fb4f514d92e0b18461804fbb4d14317b3a04add3590399504efa10aa8d545ee7f332cf9a766505c6b2aa91ce25f3fa819500053dd3fcf241fd203deed3a26c3470648c447831a05694b1cb02b8f00bc2ce110030a79e9c628040d2ace66b05c7f8777077db73e96afd5f04aa32db7ca488d741818269bdb0a2aeaf8c613558979a1f9b44e173c2eb3857d388e401f18eca56a452f4a077e543568a5cb789fb682c1c4af8344b964d57af5b112960c9ef99ece4cc5c73d2cba5a4af89802cff56f1b41dbbd579f02e723314e38fc9ce8a545f3fc575a291fd072956e21277c2973cfd60b52d4fe9861ee608c635920fd3ce6e68d0931f2a9bd3943427718630ecc6b4344593737d7bdf8d96d0be5d996055c110901048a209e78c5b5d88677b64e9771f274ded4a31be4332804842ef737158dda6feba52546209ea0b27cf6af8314e8bd07ee96e1644796141e4309087081ec03306743f6d9efa9d709240371ef60078f8dd3f33d1a4ee848b2e27b3458ddd6b07122416cee826d0db621f790ff15a3c9f8478708ded24e00849884af04c036ebc24b0840e3b440232b2f3f8538883d54827aad627d072447b791aa0849ba0c154465aa28dffaecddcb4620ebe1f4a9d4ad06d4138d66c3b181a8bd01f09a32ba4ea3e1590a48b0716cc87cfb6970d20455ebeb27d95845b2418152ed373d15e299215892498e64719c50c3303395e554dfa533df8a6b838e491282413be3dc5ca456ceed131f6f816e94824b0d7d5fd4bf4657a6e6944bd2098cd231dad25050cc681a08dfac67fce47453bac08f63ade9f8871266f1959676563f8189b38d0da89a215694fff5d8ff98bce2b47a51fcc69b17c5f52506990ca22e63f099f2d22a8e172ee98da5edf8cb5d7240d662a513ba9f45052033b0027db0b408df7c780480b28487b494d5517ab63154fe7c6cc5c79ada74058257b572132e9af374e85d51da27d3655aa013314ac8bb8ffb4837f68c2964184515d3c960942f0e2433f7f1d86cda502d59ea32fc1a2d8d6d7cc51908d3e8a81c4f9d3dad87e8eea575a08c09f1d64f5119506e4e25d12f74a1f4069361c0e8de92c84cc88c112763d1b30a56606d46ded43d84d7635e31a899ee9fe6cdd84c68bc9c1f11dce4fc7dc7e6bce43df2b4921d5ac3df534672d2fcfb9cff9130efbb83cc010f3429013d3e42d2545de0fdea0f19b16c9e92fc6bff178e61b315ead5bd881d6f1b4c83635d642436a0f4dfe794e71c564b98b2728877fa2a2bb56a1f82699d811623ece5e0a292058ad36d817ce1aac20a9b7baf82d0f8c6a6cab5fb68a8fc06dff2040b92bfde474ae0e4bac37d364af3f71500f70b91600b6fdf112be9709b6d9937daf08457e886ec540789ae750d2a60e0f11bc3ccb0ed2ce30a9c14829a267ec4694b4606d48120f96a3f4c205cf3bb2dc4c9a303ea08da562320f3b2aedd808a113a895d58cec05df7caf496dd5cd2a72dc4bc3e20c43a52d5d4a9f3d46dd2b1e721d21dfa2e5fa96418dc42365999406e7d757ff8af68289978c14e7458956a2a3df32d82aad00ad2c81a1e6b4d27aedf7134a53669a73fc4d32af721bff18428857ec83600166763a7477cff942e992882ee6f73bf24ce669f5121e088bb28af3caadee74ad2d7f6fc9eb95ce4931ebe45e52e01caada841a5cd6f9a434ec7ec5b686a3268f5d22ee392a6fc4893297b6177d3469f13d3789e6c4c91e6ec984f045773cb7788f9599d7b67eb1f82dd0b9048cd982d8da81e6140d44ab32aac4e0f54b5ceefd9830035d0ebcc3eb3d9739aa151f150ec99072e77aeafc2edf60afe1369d998ab109456fd4db1f284a8a1417f5659b58ec65f32765f99448b631fd4d003afc410c816abf4a7a33b519da09508cdca922f3c8a3c139d181bdc66adbf3f714aa4f90b0fbce3b07df5e8bca119788652a9ac1316ed43e296d68649cf7d742bcde3f5b8d8dca69646e99a42da3172bd9fc4c726e87d7841ebdbab6e7cb96594c17016b6f1c0639beb84f4d863fd5c6822320c8ffcc49be4dd1fe3a3df3ad6880c27bc55f9a2916d533e633b8b071fa2a899ab13eb9ba7ba6031a7f49425f2d11906380e9946623ae89b6d9a7a38c7fdbbdff3eebb6813523ff118823439f6611d6daf623ec7988c89267949b2077b98eefd5611e3f529e04261ef61fb4e8af92ad106059262ed33efecb956eb04dd032ba3f45e225e4f177d60ce70ae548473952c68b5a5555fed2e2adef1f4eb34c584183f7f8eaf80af6bfbbc6817728b2953df2703784ae386455aa8d6382bdc71b077c518327642f3f0cea8b04d2ad983021377c9dcc6e3f26983c252b1c1b0dca7f41843f920ca3dc0d0f7d30621f0a9a45ec225f802b0cc6b3245c7c4f25ad66c2939dc96fd2adfb2ee4a0293390b1815de8030cd1088d1d49383d8e4fff90553cfa71703f8c49afa7740d2246cfa8229f1761239f4e7524cb4966761dcc88078dd2f05ac148a18ee80d56869d87f1762f65d0685a7a66c71fe62905b8bd31818e099d1a470ee76b76286e9e68b0da69d1508cd3530c1744e861319d208477635246e2e5353a92b0a36ff8c21d3c8fba9dd655badfafbd7bc00acd3289bccf89ed85dd09bca14b1eb3e6955f08ba4261d6e49285bfeaea3163ed1d29fd192655b4736696e4bc5949ab9d6e057346db66542526dc5d8967d456d8810d0dc834113376090365f272a2c0d704fda72af64b5f67dc7aefb93c4fb138a153cfb78a8740f89824cc175d4ef1b0f9dae28c997d5d02b06c806216212017971f4ad742b3e3a396539d4ab6d3ee912bfb4a02379fee0b6440db17160d560c2492854958548674cf5af300e7082fb7;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h262cbf5827e0671597bc384b1349d00e60080a7023c201e2bca807d5a1acc1aa2dc75c1f93a0cba9a0415c972eff005dde088579c9483888fcf41e38d3c096105f6a7800cdafa225bfc8b26e3febba2485f1693eeb6257192bb4161accacd856e550aedba33cd81c9ed7eb491d86f96a8216525a9c7b274f837ba8bac61ab4f944f0048f3aec64d341316f60056653c997efc976add318c3cd9404495d9a4d92c36a0d13c5e02f391bf25fe2e08d38a3dc927c73884435d9720666b09607e75826e06b4b352d9ca70e92a67d390d2af609261eefdd82e567095bbea97b83fd4055a3ddcd55523e8238efe60e85d616a04f4485906d5f1607252ef1895e46a38dd07af5f5580aba5e8beab4fcb279d2604e3dd4fa3e6c81dd131466fd4eea3996c70f0272f8a649fb1d6438671de29747587d357fdb3f46320feab38b6f1b78983767bee5ac2aecec7805ca1ad0802dddcd469f20a2c7f67087ef95523d9424c78c18274f07f108115521feb12f19f2eae54a2458c0c1b47a66f1ad30c12080fa590666b076fdaf226067d7316426188cd67aec640566f24bdb966dcd742065cf512eeee68696d2c1eef68b477195197f0beadf90ae7c4abfd6b2cecc9bb62886babb457c3fd3ebd153e38663252f268046e4276c85b8484405a162ad9911559205471bc5d4b4810bff9e0b618d1fbc0e54d871b90b4447a53588ea6d511eca3bddcd76caab824a3e7ce8e63f85a0f3e38ff52ed3be17c643d4f9e1e58de7cf827d6badb7de613934106ab8c2675cc20e6bd7e5bfa4b2e01c43263ce46f3030f80db0b7842fe4ddfb1361bb7bb763ff81d5b000d23d4262023ce5f280611beeb25f95b2c04a32b085547c6701abaeef8b83e324b8aedcdc38ad6202801780ae9e6ee42d59b002383a3d3ac3e20e65ab9961bc34518a134ffc08ddc7ec0451649426b8e570d24408a808c8ec8bacf6828f187f377cea10fc089f23760e1926b55e48d828bb02d7c017f44629cebde53d151ba00d85dda195d1a6df71e17bc5167ff999dfe602075b021b5f9039d4188322611e6b251d7978e65fc09785cfeba5ec97bf104be76627ed38789321f566b2bad9daf8cd7614b9ee301f68cfb66e635c23321596168f8650ea9b90b907e1346a97ab8fdc94c994bf4e95d72e2308e89739779c3e48ca45cbde3837e92eeb618473a3edcd2ec20934e1c88f2119f7ece267950be6156bcb3767db9ce184ea98cee10663f7088f18b020b114e9e54a3be8697f841c61207477d457ce0e0ece670a347a4d34dca54b5eb3508ab03763c8dde7cf6fd36732729df95cda03e05a3ffa0124b5e33c6078f3504522a419253c7f276de72a66d619367d791aeb1201a5a3c82179730b3f20052b488a82e7e1480c14159da7c36a61f254a826e523d6b26e1da99f55c17139257c9c0a5e065d103dc1ad90c499186ae8d780c091ec2129291bdcc1ab67635ad833ff6764cb0116ec1b78c32a94e355d78380348ff0cd338a4fa3cbb8c24ec78f108aa242cf820a1a0e1f25b835928b8cac2d2458fb00d57a7f3f1327c95d1c58c49630fc002531ce17bd2e8325daf1e9203326d054dc302a5fe36c216b7ffe813b2ee881fda9e319b9937e1047dca4b08822a2d90e8c2806efae1e71b2ef6306db1fb78ea2baa38b0ca49195f0e76837030e3f1510937694163bb4f9a52dff41ef888c867a0e9e91cdaabba9bb5480b5d28c5eb6d19e905a82dcb0b71af1a1edc8bf86ecf35b09a60d8a7a7146e9c06a28696c11b70965ef62977ef1fd06aae51428a43f86a6c6e3d681e72102587d0773c92259b9c9df419a8e2e750197a2405025473cc854c64be579533363408dadf882c78b870d3405d402b539762b152fdfe6e22b9a3fa6c42f54d8affda956e68a95e453437fd9d8318abe9893ad7a0ebec506204b4adf9f6959e2d74f6f0dac6dce2fa5e58a9e99da9dc2f6af25d597e9a5ee071ac8c062f20150dd0a8a56c4d5db6f5806b36ded1d5c420ab699e38ae68f3834870a7514307a1e15e094327b2e3731cd0f5d0135c46efac9c1e0e32b3fff72cdc01c67f05cdc899e7f7d3510739f5096117a79734b94a4b6083a7a8e8b0fe2afda1c691224eff21c7b0e94000cd402a667828e23c0328638aee410d2b6a87dfb7cb85f99cc8c27ea01e30247a57716da3fb940c1b6bde398bbf07fa45e3789e254760b9d6fdf1836f37dce292f893dcbf8a003caf16e145538e1a433185a7d500fabbbdee46059533ed7122e4ae01ddda5e7e89ac70f7c0c9058e37908b763d79281f2652f2f7bafc9c4d04a95ad0c788c06852e1db8c64f84557ad67d7d825b17989a496939ab27370a08d4df8cb06c4ca134c494c421f87ecbbdba91203884a045dfb02e8704c84540c63a631046030d1809f7cb7182202adc6d9385d2d5e5a52910da1cacf2dacb61e512068061cce52fdaa1be4a247c4f3674d58bed56c4cf814b702a20534df37fc82b14473db8aae4e2e0d87c6a1f25e6bf6ea6e656c999f7bec099074e39bb1824f69cd1653f9bfa73fac5cd7b2b91ef7b160ea70635280520d499c17f5bab3518d610b148c415decd313069850946a8cda2de68a934d056232affd5544ef64f223738bca00f42deef27f9ea425f70b3da46a66abde5f5aade138d6ab2cd3de637f9a95d13c1e3cd5664e5feb1b1f93d82def279a97559ba153f962c2a23b0f53b9d92e71c13a70e56dfbe9c7738c0ac70357e7e94e35d8bf57355cfea2ce179c43a564b45fe33472dddaefa6b4108148f772719844656912da392bd201ebe3032e2c709d9b4edba0f6914eaed30db9a00492a47438517a43df152b2a3f7316f0c773c7225da813eb345de717ef47e32bd7b80a7daa435b30d3d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h26efeb9f4e49e9c8c4177aa2cf4edd2b003fae7b1a922aca584d23751bf69bf466aa879d3e49efce948be046088d932c6ca9717548f5b8727e5393676361ce12cce5ad5e9c0a4c5dc5c65a9724e3a16919ce5b751008848960a75f7470eab89c77d76e917b0a0fdb0def86f071a85aa6c07632eb7192b100e24d5802dbf48ac9a639dcd6b597b5b2674cc98bbb66e62cbadbd520d83e2dc4ff38cc1003e05af1f5d00889bf8580591aaf13a10a83ab22906fcf8bd6e56d9a34451fd55178938a1376b882d5aeafd4bfc4e8f98077edd421fe786a27a2ba969d6e78d0af2b69e1de139fa09878ed313080f2ab0b4f15afdd36e2b1814073fb4fdcf167fe97fef062dd94282fcb4fc9424281a9992950bd6b40c2dfcf09abc4e22926131b4087d26d99dc2af9babb7915111ff5ebb25c24fccb7aed1087fa824abd4a20ecdb71b6dd9c1699f4feda43f7ff3eda21e5f5a116987deea345bd232c27e47bfd26f6508c901acfe017ebcc3ce82387f5984c0705ae9c98b21703670bf8e2ff1efb2971023a085eb38b9427b8c91ae4e0b9418c78e27b2b937b531521dd04b3f3142aa4a0ebbcc6ebcf6595349b6154b4242a43b2f04926342901bd9518add669386f4fed190fcd0a6d13ce62ee5a52b7d9b842870d6682e2c9995b61c1356806a14919c0bd0cab613a65cd134cc90f393529efb55fec58014847b4197321f19e2ff28528fe126a8b381cc2535a6e1845415901811019b1bb50333aa9b5f7edffd7af14135b43e4ef9881714ee9ffdc7059533ebf65ef49f938022d90b862a2ce5b31a637195e34fd48bae983011a5266753f4009ebe4948d5febc7995c9a9f7eafee585a59c9e284afcdc8e9a458c162b78892762677bd536c9b96cc859d83e0a3588f0ced5ae8337205910828986d180bfe9d4d1309fc3f87a273f390e1a09013be83b6573ba3e4a3116a592c98aa3ed616cc31fdd3e5cb906ed36c2cef139d699906de92980941faeb1b03c6cfcf9c3e6b49774234df7cd76c955c84fb3fb4a837ad17a107785ab00ca30ff61f3aac2d2014ae529a3e4f53b2a65805af4e75fbeccc3ae881ef7fc34d9e5e763f529c0303ba97598bc1a0365e4c9de7f4bc3500dfdffc886f3e16416e75e75ec4bd5aaa2f226d5b798535096bc7cbbe1d8b3d392af59c010f615d910e83223f8ec32714d7d4084a76abe5f473415f6d22394277a8d0617a23359a74b8358211028e4a9274dca942b40b881fe0e1af82c4ffa82a9342ea03b0e4f115b082bc68b6067f6a864f86daa1a523a3cc116a3ae5c5bf96eab002890867e33d86dfabe1238bdbd46abe6b8ed16c5fc7734b9b094d3e4eba8ecb89da47317c57c89664ee6c8fe33fd436a21202d1c2e550d124e4ee38066ccb5e5d26483ad4a541674af0a5ff3eacbcbdd6f7d7aaec37b78ce6a293e0ca01bebd875cee54bf4afa4a99c892fae2396157b08c47fc456c721890bd2e6abb77873276bd7c81c8b5bf93e39e74c1737794c52e16d3468ab5c3ddbc197a36c42d1bd1cee7d4efd4331ea158895dcca4613414a11b45aba864653f79e7ccead1db6e4eef003df4b9e35c3e7a6651e4002e3bfa521618834ff45816411d3e8fc1cebbcea09c41f1fdb66485e5021a98ce61bd249224ceaea7d47cfc86e42147b89cbd79ba335be980fc141cf6763858c7a6fdfab56f507105bf3e1c51f47af17eb47d801d6ed16a5c9cc80a73593689ea5203ad4150d87264b7a7476536130715b19aa20dec58ad8258dc716366450e69647bc772bd7d19bbcac80f0b558a6ef4efce1430895621bcd7b33657db6856d6a89e6676fe9a8f4136b1fe68f80759352b7f2d2034cccc7ea932902ab957903eaef61d9870d6592318de8676d5c086fbc40c0385fa82d1b2bdbf8156a873b0187fc9fbd6f108d89b3a5943f47f0b45c950495e2ab7714ab15491560adb7641403ebc380237897505bfbe85b70e883dc3cf96a39d3d3c142d9e91b661368130a9ad0031016848c4a52def10bb79f5295eeeebed6ac235ed4cd37985592fb36bc9c00d0183203cf75077a46edfbb3bbb0a41c746db19f314d0db1d1e161058d347696ea8917430f0100a26ac16b54cfc6f7631a0b64729068a369c2ea3f2e937bd48a47e2af1f481e838785f345f3a07ec8490036ffaeea18dd404876dfe7cd2d9de590c8a0a74473498dc3d4e54944f9c71b77e6e0f17b2ac189312ff5c37685a621dbfb075663e491f0046bf19cc883bf82c50f989e5568eff7dde12cb2a5594885b6c19ddb72b5c817454e9b11fada404d9cc769dea48751c34b29eac73304523695856206dd529b0ecb2c1ede6cdfffdd7f1f879d52f819975c6d6f9ca7a6f8fa81e3c6407c9280e7b0afede884d41dbfd5e1cd15490794c7eeefa61b6e623bd1d4bb63719a7f928de6d2669c8fb59590f99c12dd9d1fe4f15f9a2ee3d5e23a51ce7a0cf1fcd9d77726740588f2bc6378d6eafbf813ac4c58f5e756296715ea6fb7987b85ae0d42be0209dae683e5143439c2de48d460de232354f6df46db1179c98f1eb2eee0c774171c391c62d10f4e007293c8954f3c111a6ff7779b42312fc85a7733bb896e86d103e074f11380f736287fed7e617ce70d44cdd76043cc1a8c2203230478dccf5429b61db78fcdf471f4fddf831262ef7b39fbb963d00914f02f7d1b649318b5a48cec0846312df06f8a14fc0618d06fbf065d9a8e1f84a9cd89b94cba7ea42be6b04bd5158e537af4964bc80a48860af8738d089e070a2d5c824828a2fc3b021e053bcdc68bffe8a632f115241a237dc4db1cd349e9c142d90db14af97d64067c31a870147f7ecd62effa0117864fe8cc1dea042bfdf652bb0276657a642ccfe3fb1b5933aa52cb223;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h2d93b35b5f39428b93608de79509aebf1929f4a5845befae6b83b304b577970a04460558298dcc126d345b616e9fe1aa40167e142618a4d285082f90074979d4962afb45551efe5964bf1849643486c052980c2cc7aeee9cf4545b639bd2fb649fb9afefdb52101f77cf4d92a52aec7549307224dc19da6115aacb956a7bb5f5326e1729d5c6a9a3f10c09fcbc2fc6a61ebe2da0a67fd41540ddcb45d2c278240b378dea51fe0b73930780b39cae769064db9e4e80a2c0a8bd99019a63c60ee90d91e66f0375e20b91181bb7dc37911148ac3df89d81d50050d9f85835cd6c9056dc2b9df410c9e9f106b7358b0cc9971bc20ada76885397cae4ba9285d4f909c5da212d085873ed502bb932df3f20a4c40817fb7e28faa4e173607b36751425f561ad2206d17a000582caeadcf98cf03c18e85c433c5dbd6a9777265d915f83870a1bb7c276b832a974ede6d1e3c7c383cab9c13b36c7af11bbdbb4c73b2dc3a66b01425cc7c2906ad5bd140df188037fa82d92c9bf0603276f6ce9e3bee1360d100ec19e898c9a9d615aa62c76d8e572c3527af38f9536e4cb601d1e45d17c17a58c054ac6c0c78455549520d9af3a0403a82ff941848ea5bf90e4942036783fe4c72e0fbd1bd2e318beb83a0d0807c65e9e49ca6a2ebf264fd1f2cf06e8058a10bd616016a34227d117e3d655f230587ba689384d0587df2f768215141cdbc484328a27edfec947587cce083e97eeb5a2b8fdd3aa52b78cd9d1800a0c6b0bdfeb7ccc2e89ab2675023fe3be702d5ba8e345b07e77dad352cd8d4754c786a910abb4e4eb2676a7372f8236e79efda823992a9f7cd15ede47041fc4f9db3ba812259c0687f57a21ca27f9a1da1860072ad9012f47ce55e37495faa142a8e1ca15678b23817818416fbfabaf31b55c2ec88cacdb988daaedb1643146a47f11defd3b3c4650e9b7b452820c86eb4db404e0b425c01065786ae3a5bf6a5b11471e45be7c99b8808c4e859459449699e54cad7f2f6072e4593b1bee3feeca9d8ad45f02e9b5c346f23ed3be656841eee5f96d7302ecb59d0f07568fafef5c2a94d5fde4f12c0ba6de75653d329d3ca2221516fa08a2f23f89a27553fed986ffcce46db3f2a0184abc0a808dd260c797716b8c117a5024b20b1b7a22e119243fb2ad1c775475cd71dac826eef36f0d5a5c9660e8ca56bbd92abefd6b8610c7e81f9504e12a13c71f739ff4b41b2ded6efd7b503ca4b6e7169d941d32920057f90dd276d1550799f25de3fbcd63e37201c4f76d3ac182788c2d99eb2a4cddca792c0c7ba2778aed9294299f8cc0498aa0f46d517caf7f1159fb38896f731e4a28ba3c7b6d9d97bd46a0c47b8c3c968fa5f2f92af84aa794c0c8751734514f1549c47614979f73fd64cddc949e5a896d691d9b57ae3659662173b9773e5532ab3fa514442f13f8dd143df295b5acf7c38cfc5e1ef0c33ffc7b0a91db58042f8248b354e9ff949295e934fffa7c670a78142a0f4f7da8ea131c120f64b4736ee0b67348c99be270a482ea8f4fd4e642f18126ba39d55530ad18ec9e8782275387c37ad021c4d6d7e4ee740990d0f79e6ab0ce6d114de974037fd87982089a3e11c98221e8e2d1b89fcbf1dd3353d7732df8652950cbafe7bf7e493826fecf6fa41425e3547312d8dc9ecf0eb5b6e5057ecb290e3371aea226f9b235b7fabaf73508f5bbb47d8022146e58cdf44b2c850c7b940c004f1ce5b7a80df2d94ca016691286d0d65c97617dffe7273e37cda969965f56c31a89e8838caa4c31ea6bb7abfd3eb2d8587ebe3fa91a38f70b5619f6dbabc87f796afb9073f5920542d2d2297d96b3b42bcf9707cdbb89a9a8d4991b636d4506d1ebedf8adfb97926e318ac84b0ab849948787137713f26379061416c2df28019dc1b7e325b7cca4532d7a2e45adc15250013b71dea0df174b202a0fe79379baef575f83217eb4177acc3a4a428f37e072f824f3a48ceea61baec5ab27e19c2f03cb00a5740726bf5ac47f3a78ccd1db3c6fe71e4fd54f57f9010b60b940d873a4c84f2557788f867b88febbeb6a130e44dad4f25b71a98cc9a3e39dc707d24a11b5b446d3b9484fb7d96ea66571a41d646b5604a2ba4bf8257ab6946009f5798dc888c92800758f1dde19b55adc156dd39f6893d36a98b2ce716bbb77463fb210b57695a6e64bdb906f7848ab50a5b8be6d67fbc5191192167257aa831168b89a2cb4e1072e7d0ffaf0c30a9f90fd5a4bfe1034fa587787910d0bf60af710bbe8840a35b5342705e09466d2d5802f2b5c7042089f67e1fb77cc6a140dc6897165c29900b147109ec8e0e1c17eaf0400a0608123e244a17e237f2e36aa00f0906a35996a26760325cf2298819e58dd071f117f9680abbe4fd9ec512c75223d2cc90f4dc6834ec115e82247815d0228aa6d7de3968ed220d4d835e39893bdd19de75eba2be07dedff545b9d0a38d37ba69e09098f2740521eb735dbb159a54771dc0b9529b65e4d46ebd8ce4fa09507548ea0299323f8e61a4d659f954a3af1636c46bd2e669bd749364a2d5b3afb8f32af74aa7559acf315c0b02da9ce19f5e768eb9290bbf2fe92ef1976fa73f74ebfb9ab5bf5e2d4c13f2d0008eca84250b792b0105a4ccd8bbd7b722f31dc7d903fcfb65279709e586524dac97074367094e4bc172df7c374d6be8a765691ac864b48ce52f4f1561e10f06f1e266db802667984426eead100576b05f3ecbfa4c7fa91e8126954fef3292374101cab792fc95adee418250d5e5f52a1069dcb792bfd93253a457c7c0b763196c852a7ce7e06350a7a1bc4fc29561f60244d04e7db58ae4fc78a361e1c1474873928b2e3e748215ac2614161a24d0c4bc16984fed9;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'hec7a25a9e8d6bbe54263e12f059400487736a4c14d8f5ebeb393973ec973ad0facf3e719e318aa010c2ce4cd6fc0b28aca3e6ee6ecc00a5d534aaccb9594351c7057edfcb68578a7f4d0ad86bdc0e3ce1ce547f9e4c086d28839352d5dc7a205fc892fefc5c3d93dee224b6257d6f2970f848b080f4a4793bb985b6c325aa7da2c4bc7de0383ef3822f43df1861e6a1fc2c21ae8a2280da7225c6280c80a8845ee16fe67a0885e3625ca0b2ff05acd84921ee9076e878feec0b558e19ece4731f1793a995a98ada250f58e548f065b35156db2ea8e1c74ce98f296b8512ff5d4092b4c2a570b7e90f6c712139c90dfdcbf222c4984d14e7e694ccefce1ba9cb9f33c2b927acce48d0b84b204fb12ce0bb04ae75fdca5a0ff8fc388ef439d04bd76d60a4878c9d1cba9b6441d8fe05ae0ac75479e1e880becaa7a6ee60236a923b6352cb0a8e314fb5c94caf2c9a76c6e254bd8357604fb0b53f182904da5648b52060bef911b0b8e5011e219a9dcd736a8bc6da5d95829b96b5473643518fc2e2ef823f4f4ce937343a73d73d41e1282d764e93cd3baed58f07dfd61e98916e9279a904e783f4ff636764618e51c1a11f564ee9fd04a0c0054bcbd9804a387df9b4cfdcbf0867096f29cb2cc993756dbdcada5a0d1ff8f896f2daa19a0ba1850c97df33329e4d33c485e0b5053b38e3c290fbf85f7b6255175cb5aa9630657159571210c0453228033e8e5d96913bb4e0885a92a7ac07e035d891c9ad8a9974ba75f2f669398e137b01c903d272f9be24a14dd70cd316c7b47e20b0ba3edb39924abd12e2457edba3d65c72881a5bbc4fe67d6e14eb6aa0fa583a22317792a7af44b82d8b08a0f16811ca9ea9ca6b9f737c53f28c4563987379cf5a9517bf95f933eeb5106bf4599376e1b5fa7d7857c4e9dbfa6641c277b38fe2b1c42e02ec4494e6855a448e852600a6984433f26e4cfc43fa9febccf30a206ef0aed0a0c91b7286cea178dc3c606052396c8a2f12ff44b3d353fe81cb17c4f4666ac749ffd801c1e2073d8522b216858946fc13001fe00e1203a1ee46f0c9b5588206cdb6eb979407d561612297b0580e4eafcca8a64eaceffa4081164bc7e48cdca9f32f02b058016135d4fece21490aa208897ef4a4a8a15ad4ae544c4ea546a7e56f7280d225be13278b51f78476bb70836c8983a2c2c317d5a5fe4ede3670d2c4451c250f5cb9bf37342bbbcb7e046ff74c45ba04be27cc9162313db7fcadb28e9f8bfc0f56c9d64abf07f023729b9f9f86985ccc2e75803ce80ef4355b0a68dd7c4c67927249f0bfc4e03014a6d1a4be9dfe62e1885a30ab0269179389b57f6161e6e8a646c2f8b2d9210931a013cdbd7c2b10d783f17a4faf0997dddb19957572799db579b87666501309f00419326a8cdbc6befa67226009171a014eb6cebedab83e28cb9086ddc6c709f0feae1d3a59c968974604981e7299b16c1a4d65c4d72bc3199afe54a1b00a4c90250720d87e0c171989d1dc5042bd27018e0333e28bad743bbafa135ffa43f8622b24b58a55765cdf4a8c943a8513eab72beae671266553311162565aada92463a07f69e59d7f0c59ed6156bdaf4d05bb55e52a93ff9147d38a2afdeaa61fad559c631b3aeb8b704bff235cfb4c8736433a174ae8af4bfa036b2674ba116280f8755fa3b21b5b699f9097ed590196eca0de665245b0c9643bf06e081ea51935df037e2e64621c3bb3b0422d2de6e438df3363563a328e6c4caac66680bcfe0a09c395aafa1514989155aa90643726b7b5fba9a47054ae384e56a582adc4fe5d90b3eb800e8c6b1580b0d135b931f83b3364fcbe80b7bc4162a5695f5a7596855fa7e98e9c52ffc3107a606f0c35fa99a0fb0f94636d14b1dda813d24a6f5820a0337567e74df23cd79faff5c8231d2ed3133d5875559d6b79847eb153be8fa1e1797ef58b21cc2b5318a89f8ca9e0d85c19d46b41656df7cff7da1635f4a9c49d9fb95b847f3a33a1054cbcee09f74953786cd8cc9710a882eee30c9f13dc8497d61951132dd75879298ee0c27b2d17c132066abb8b34c8f323a92a95698b609fb00442e143ff67699bf6dc49e64ef81d7660ac7eb78cf12f8034b443c2d847a323f66e25c57289df73c2a70685b8188e4a02c38cc556072140e92928ab97ffa5a3dbab526e7364c6f0bdf455eea589247a00f28bd447c04aa86bb748831aa07f7fd249a635307823b045e9e34c591579e49d5f2ec31b685fcabc03c54828480e90773ea330bf2871d100b7161fec6c4ae30fb5831b238d2c4f05873adcd345cad5c310ae76bf67fa16ec6e3e09ad49a2c592e81f657a048c64e87bed960eedb5a78a6573c5028f61b8f5fe49bc994a4bb573986b5ee2a6e4679b78a3123ec5847024a5a9ae613f6431de18e67e74dd9c1419182e0502d52d241b2b51b88489444547258f9f978bb9f2c00bad6820ed709d477dfc0212ea5456a15385e81b013b4d779a094fec2164959caaf3f10aa69fc20448f565f4b3a10ef5ca0a6c00888258a1b3e5e3dff30e384f1253ac742c49284884f93ad20e6be25b69000c5d2587e576e4a5866bef56d63c6779ce6f1c6035f81820140594adbdecb287b9fbc9706615dc6c5b7bc8bcf953b9c08bbad13e35c360a1258e50fc64abc9c4b8cd52a2cc673f860aede70385440fb1be948b70235b876a9e350db3b3fc4a6187c7549aa4f7f9013291f17061dbb489117ad72d8aadf39834d15be7b6ba41bed3805412449d1ec0fa848e4b17f19306caca7ee24fd580df72d998d1736e086862e2169764e96e3720cfc8bb283cd9df9a6fa1fdff88d91a23079b26634f50924a6429e39710e3af65d92460672fee4fd5ee3808b3bb4bfee0229;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'ha26946156364916b10d2e608860f61761fe9e25cbd512f8221ae9364d7601bcae9af621655655a67b120aec02591f868fd848dfe965b49dfdf7e82748cb642735a2f3661c75c32def17509c30282c60a207422e80e1385d3f9b9d02be312614dd49c149acb2b2b357f54aab883a8644be87532c59c7cee6a3f5f848bb7d9e5d6b4af0c793c8ba0787647b5f26d5871f048224956ed3d028ba6c116d5ab51fe951ac6eee4039d0f85e53cf88e14460b53a72c5bf8538a35eb84e87ab9917fedb7066de9085e16d97c980460c9fd9e1a41c2318a4a1f114402f09e1b16954f86030c7d02b91d57e78c175afbcf3fa51e86c695cb291e659a66a8e0677872c28e28895f23461e10cdf4d833a6b30b2479e26a49b2946c16b4d4d5f0f917f103febb3dffb5ec1fbd654ecb34dedaffbc7ddb374ccf97f66f99e7581089007f182db6b9d33a244204c303410d4aa387bee4a49cec6d21310ab56d5b15f17bc8f9f764721dbc0c0dc96ccc83d885f3d788826a496bd188a5701925484e711a230d39f2ef87d0c92edd7d623c923ed1ad5239036c1fb901345672066f034a839de0bd93b3e264c0af1fed5ba863723e1c5fe498f210531a4caa91d63de57605197f16a52ab7283ec881de1447579ab81e84ba0ea0fc749d3cf5fccd3fb0120253ca9e09e7782b6d821dd051e806b8b690f259e1652b40b73e7c040e6e58c4546008e97abef0804968297bdf4d603424db1eb6894d7fa6d5d3da97c0d36c7c533f2874b537e2609a1f984738e289d180f3fbaa44a0d2a0fba08bf7f4cd7e999a215567fdf39963724b9fc9ff940450bde5cd11cae8e54e4f5b36bb050ff96634ac20fbb50570e0949b1dc609c1f44112f222b3ca2da341293b50a2427b9a4ca9441ba35a2f4c0a0f59ef2cf96a9f89f90de0c44e1c1446eb5d8ea8fbade78a4eb2e0dd84ae6b00b86919f584f70df1923cedea9466b36267b7fd946ff827d9b1885b727b5c1bf8d6e9c230109de244536bfbc5a317639319cbc02d9cb24857042ed27533d0a072ddf8212a57f0e0de8cd6808de6bec3602ada32a855b33dd75971217bccb5447de6f4114c676235d49fb4631af80f815a0bef22797adbf157ee7c45a86ca8c52fc727e8fb85a68ae41443da25dd5b05ddb656fec85d088344cf66b624fddc8b54c1589420a1f3407bc3a6408c1b27ce1c3c9c3f0309accec583c858f209223b8b753414c5c830af75d15ddaa9a4f6e5a3b9edb68858e04fe4834b7a4e5d9e8dbfe22ae5bccd5c3b535e88c02dd4c167c9b48f461f20a31650be426e0fc924b36dad092497e830a1e7de262c50c5f8a84d510aa178e0bbd70f3a2983e046d32c6d7918b07f6b02a40b226e1e7f3c833e187908a9017c6bc4b844748d4291568b06af3f2a36468bc67a6293843fbe74d60d957fa572e4f08ba1f6416d28b13fe8f0e57e53343e70c503c5acae56069452fc637cf818da72cad9b4a6d185fe63972044a224d9e6e3d52236e8791cd34f659ac16d0ce85332006d939c5eb70fc9fdda12d874ce54731176f9ad46f9878d5d41b5f28745ff63af2fde5d88423efc1d80c9a67a6bebea8105b66e947de17e513deda7ef405520b988be9f038a60944a79602662a663d7dcba825bdab7295f0eb5ab6abcd9e607e4f43c479e7a69cf0289082e80db4b8d0705cda7322ac1a16daa2f9b1ac90e7694e04a105bed84ce7e70f53029b2222e6d21305a0f0debfe1d82eeb7fac82d3f085136b69dc41a08eedacc0ec9cbe86d853d4f4a67cccdcc6e128f1a7bc7923cad2326af73cc5218235c6424c70067f6e2ebe4256986ed0ed03db0a5f98fa83d12cec7dd62f896cca1cb41f35afb92c383297db6827a06fee968fbf6953e629555f262eff571f51c538664424aab1b95a723b2a2bfab7fdd26707d5330d9879c6125cfc4aa583c0ea657fa7db7a1cb842e3d0463a671dc4777b58ad9bc8976b2729fd222eb3ff49de05f2581728795a80efda61284fb087fd949c0b3f78d96d592e9d51c672ca7b5c1e670d4d6aa1cc335c5965ef8a81aecf993ed95ea4ed26e21c486e90930f2a5b047751ca9a01d83d0429172a7b72ca2b0b479692073c62251f76ec36c1396b3c2d78c1b8458ddd27c2491fb018983e8374abce4f12bb50f550f1ac47aa85444c9a3045ac2d1362e7cfe44b123d227d437d5c28be0933601a6291f3b036c5db1a41cef237f692bd1100c4ab39bdf9487c52cb5925e34b1a4225b21fb16d6e1cf98a16ac6c555d77d66655e1f4d6e01a673ac93054dd88bbe90c1a841f03ab46c9ad6a097e4fff040050ff91f8999d282dc42a5880dda440af1cc838f0c059a587d5e67cdf7eecc64b61e0b22da65fe53416896e11895a002742dd8e08deb2846b7b1f1402643d68ebac230d748d3ddd61d66562a7c9a79af4d89a591b931406b51950e79481187ea17a83764d1678da970ac0187b8aa674a796771b1cf227c7566bf8372092bc8fb4ebcb74a29cb990db788ede34dcf0a8381d1858992f091382c6510bb485b25f98cc7b8c46e6fefd744d1de0965643712d919a29c923d8a02b508d9933bd7175c063f6bd5740dfe6d5ec7b86f46f9f917b5736e3df2b9a1fad9d602eec03edd8af4dc97d804c5da5d5bede6c78ae0fb19755057e94dbcd80d7b8e42fb6be4e37cccebc65565fc188765df06a0bd031a38a7bb424abba851233ecdfd793d8d9931e3edf441599e297c7a5512ff3104e98eaeecfbd760f133879db7d3d150760168366019fc209b2d00a656e0c0c79806a8a51f5418cf8484c7b217d936610175ebc9b5487dfb6fb637e08cf7eba3d10cd2d2b0f4f932fb9c1749be378885a6dd4459c523cc2b9a9c67f70f5587af13e8370be724bfb752ec;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h377b4cec9a97456c3fe8d945fe28c12a972c22915e1cc48d97022ba8483fa011255e9de1e132b695a9d67151dd3e68750be2b992ed902bb90221fcefd7a16bc7458e544bae78832de8ba08666bf8539718dce204104a45e271bc14dfa50f45a2c5f437e9bac23ffd3ac6a57f4516c2bb1a85d5e2e8f6958f557337f7b5726c0bd1ce5e92c4a38404ca8d9cb0722ac2170b73da70722adeb29c7d51e721afe7c2058040c6b7dd73eeac499bd62bf873accc4db72d6732660504d9057988f07d3ffd7ad232f279848a3ef892d8d7fdb16f1f80dae6871958104843fdc9f1c3ee2e7b8f1e7a2bd003a1b92cd8259ead9c46b47cbd1894b6712323092f1df48b53b95a17041072230b3e82c2b5cf2f0a1eebf29392f49dec8921037482ef31379a9d67927dbfdc32aa50ddc4076d61b4a366676a72424520c50897058c439fde0bd2560664d5ef856563005311ae7ffba976d4b04785f8584d952372ce91d3a97ca1384a765b18489d4025f1d50df4408f2a033656e733240bb2e744fe18f867b0c92c67e2e7a42ce47021b19394189ef81f1867166e50f06e3d0d58e510507e041a9125958f2a5b89ac22bef0e1c9c23c989b74ac5d56c7cf566c0a7e76502dde4ddfc35bae351ff0438c00092c485547879b5490e1920b014e8e97d275453d3f2da02fc10fbb1e391ec7e067b0ff701e9a446495b87fcc99674fa14e39d59c4ef674fd9affa0207804f84e7f3cb6204dd95933557c8408775ff1cbffe87f59f13089029a645d3afe76c6e11a9b2138eba0007e20453a4bd84ef9b713d089e5e31a96073faf27431627323eabf78c1d6362cf3283d63770469bcfa900b56f6e793b12ea141c214411cd1df3c4e97a56e92d482263eb4d8873c5f2ddcb0a27d18e40f957d5e0410de60fe09494bfeecf1b8b551b63c73bf1d4a7d34deefb4e5c752755738c744ae7e19972dbe5b1639188242476266c3f4ea841a066e4f5d8d29b72d83c4c0726f20a6319da1e9aea1558fc851f5ebd5e6da339188a119a6e2910aa9253bc56da5b18a4661a24db85ca758766060c0640520e6c4ff09bb143e9cdee3d1f43dc518a4cfec758ef2a050d86a49a76e096581ef0273da21858a81409d42a1da21e26cc887fc6fdd618fb4d92fde6f7e0d8f4504c1cdd54973c7ac5defc4e4f09a8c2e67aafc61ff0443bf6f4cae05aa999b32d35f1d106048ae7b5013ad14bcb577f016b7f72ac4ced58904a288f76af2fdb5cda9484c84103682d57f2e467de70ba8bcc9bbea07961303e9101ed55959b24a25fb39db9cf6bac29cb2eb6be6dcdbf367822faeca62596f70eaf7ab54051453c8b3235440f33bedb8379fc29d0db17abe31539b94738e3ef50cec5b71f62dbb81ce150a81ff00652af80300529a41adabfe89a38e267df11155617919082ef6635f62ecdb4bc374496301eef5e0e39f201192f498090616ea0608841a7b86052f89672f06b8e6e845aa406e6ebf756b7b6f9e3bd97e1d6f38c0d4550c7cbe61eb5b4e6b7e8a252fe32493c19cebedf4060f333b0322cba725bbf310b5f2fc11cc79e4caedf748167a05590200a04758f1b3883a763adddce27e491f48621197d857c92398a5d961ccb7432d14ea35c2190d660067f6cf8c9f430539653d7eeef8971ea57900d035e0de7b1910f968f95f7da33e57cd37697a7e31ce7f22ba593242121331ed6bfed4ae592011d8f9b77c110c38ee24f71fabcc85cd1d6ff79027fc452e90b3be7938951169fc074d0952e5df4fa6478c7c8618af6907fbe09b613cde53af95a6b377c863c3468a2dc5368904399b08c2da2d5d6df982a0eec361806c310f5e75909bef957775ab1a9db32ea9c4eeba1b0b8481c37f5f4de3b532957625a4904eaaa1b5f001344363201618bacf1602ff47288dc547bb4d41fa1392febceaa33249388dfbf96ca26f2a74d879855db2d7ea7508ecda1b7c6d57627b7edecdfef9b5c69bf7e7f404a912554d8d39041ef912195ea6958d938bce86987901770322dac174b8f97b93622725f87ae5fd9fa6b4359fcae2958a29da28ceabb6fbf9f8c08c1586630170ca73ce036107882ba760d4d7bc3f40f88062d6cfa47710183a0aba32a412827fe46ed7118bde0aa429670ad3c0ffbf93fbd51d1d15dcffa72df0f5dab83b60acb5f40fa333a6b09537cd4f6972ac5181555f9525730ca816e776a5d723bf783958b65a387545797593c12324d51b1d4a2284597df95c7de7f20fadb431fad24edc8d9dde1e9feb4b59159545169bfb182cf0c8df845e98ccc58b2effa522a74b6af0d35270a2b390f158696ba109c42f6464f947ea6710a447811474bde0612574d5420e239b2dda453cc788184dc4c45c5ae33a788133d71f89df582a1d4fbb35dca3f908cecefac17c0f20291d2de1ed2edaa5643e9dc6047d74a74af26912caeb7fc5166671fc5da765d743ec704cf441df91828e590be69c79b19b561b9832d6b4f1c789295aa4abf72a843aba8a7224d1f58bac34de3f630f6f419eb3d8b745b671d30ee04255beb9f11aac12e66eab3558210a2cac58342ed3792ef456b4088dd793899e9ff3bfbb90431bf4ba561a3a25a43e103a7f3a820c08f81c9963295514e28f7a87b36827901cc2a7e40f2bfadcdc32ce07d5d3a54c30ce6855fde42712b30ca4442fb91c4477784e3942616d45fc15728352677b7d78d843d3a6000b5a44f7e8bb951364015621c1ed9ad14ddb083bb3b163ec410ca1012cc8660ff94764f41ec30c52e18b26bba1d670233d33e70d87392b201d7cfee0324215e9929d1792bd65f1ce4b17a7d433f69d7aeb0b55f9015e65e12c511fba91d387c47626b8bc7883b802f3937c8ac89164aacffb1bf9ee07484732e81;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'hf38c57d131963640c20680f09b1a7b0e3c4a2e33ceb4c078d3ceb0988955566a1076372a3408559aacd50a90f7a8219173ef60dafa94e3b00a71539f96f65ef2430e27bdeadec4daccc8509b4aae1d67209874102e09b822f5943dc06edf933131dc4701cf6dc301241b1568540cf9153440fa555d7c551d7a14f4c54fa2ab023a3d5fda95b5ee0aba60ff625f1a7b9ddcd09e1d037772fc47bad7181081075d7b07a32457814c179ec21b333621ab822ed64e1d0d47842b121af9371a729f72824ad6c0d67bab5e6c12ad77a229434300c3a9250a5bdb5827e25b63dd339a8cdd137ae6a349747ddddf83a9da2117cd31684db70fb7447c5bc2421f05c8e1623a08f59ccf32982b4349d342dc967b0a370310fb4b7b67ddf7c9a8de9d0453e4e74b2de82c89e6579dc24dda7617f41c4edb9e147c712acbe959e55b841a642ba24e481efab1513b2b593b4a0fae66087d0f6c16ee9ff8a0ea0fd363c4918114812331da207c0c97fa497df960a2269a02660cd9a5654f59023c7329dd53d34ec9f9db857e1ffb7eb748db5b0088b93044632eef13f3fd29f057d4f4a761b356bfaa3e6cd56149b2f7686dd8ace99caf15af8ab0c1999226dfb6f038278886f4c3091dc02444c8b2a46fec8458e4a95ecaa52b86c612b6db69b9ad1edb0a4da09d6bb47b107c7d7e4e2de2dce1dd5ef9b33d832fefda83ef187e5294b51ace9ae83e7bd1e5d7690ac35be2f7cdc21af891910d6b066fed06c3905dae23e0d85d11405ba91870c5acb2f8fbd140612a1955442b8af719d8cc5883fc3e85d393aea3c10faf6d8e9d2d1c6e90e698f4e360a519410f4b449ac8cddb8dac66145baf4bc594f7b3ad2d10554962d066e437695d4cc976de96b75eba97e73cd5a25d1fc5ceb5874ae01b4f4aeb30cb79f850b5238bb3973cc7a4afbbc549ac2ed19eb8b08a47173c294e9d75a600b7de2609ad2fe2e11a5a13122ac883345b0f378273c207a888b72b39769d847256bb167df1073c3cfe8aad0829ab223f6f26f95cf004fb5fed77740568412b4abef98c39dbbf3e455facd9eb6cba7827d18d43f0a294ca95d6511c550410ae6f7a96f3ba5be3eeaeeb2e853bc44b02787b8f6c61b69eb9f06ba1984b392c286c2d0a7279d344cec6f0ac918b6316eee8595415e9997175fc553e765aeecc611941b77525e37b542b7648d69222fde0d27e5e24c4050a841a6a4275392d7c3711c490fca2814eec31d7b7c08205c1b9189af59e7ae57bb8338003f408fa8c64cd41371c094f7d640496ab303912c3b107ef0ad6eacb1ff23a60bfde28cf497650cdc826589f2843087038ee4f55148b46f5e598ab2a0ffa4a8115dccb2d2c0d1606b777354210b156801da6d7208da705a3787e2b7e5d8a75e36991f759c94971f3fcf5f106db1ddda7d3a6a8dc7eb01e6f56fdcae2563e8af310783fba4d0a75c645de4ef5be277c9fca37b2a92754b7b5276baf4f66ef27a129cf90089ceda56c8119a48571964ce2114619013d2b15c7a8251e62cae8a21c96fbb83eb0cf8c4eb9aebbee2186387b2c2605e0969ea448ebd7e12d992fb6d001dfe9ecf2329de8778fb555db4b752543c420bb2c7d4e831b710f3b1af86c06c7f8dba0f3b3ebb50b2f73ea56b8b96accd218e9da9dfbee8bcadff614ea280cd0a8627bf962b82c202daea44400e4ac25a64a6b84f4533d5f49f19e1cb6d089e9bbae60bab578bc271ac9647872da01cab774f521c464dc3c33fb6ed5506c6063dcb2d2b12ee76bbd7e7955435251f488de64195ddd182322d66baf45a8a8fd677b2ac336fc4468f16bbdd54f54264a3f268dd4e724a05008b48dfb3a7872d95f2c2364e526b69301c91951484332188cf938b71c14070f75a8ab124155485aae4443f4b2d3300a8f61128205fbef28f0f47256e49a8e54dec515bac5716c4de4d7bdebc8af66c40c944546de59b7e50caacaccd6bf2116738b0f84da675f89aa03ec751ebb940c134b89f4fc79a8c6a2c68c71c1caf745ca8d3fce0388a06c2890d1a9406ff47941623ecc04fe9085d5d33989bbeb1dd4514050bfb872ab96ff2a46e71b244f8db74361819e26b477e3a64e8e81014ea64dd7ee1d189a2bab6ae30eb68ef53156e2761ccb0b7997aed3c927d7ea1a90fc396e9330da6126fb73f56ea2605b1ab8beebf74024622e148d7458b97610101e29699e4fc93ecb8062567a77a84b90b24b322a16d2ac61738f22fd5952a24828d7a02fa88986fe0de8cbad2e36f9255160ca96db00e4aa7586a9f05650c424233f21ad46b5bbe26d333576735156a8fe84d95be0c05d623ad3085606d6b4208394032a4cabeef34b67687bd5721138942b30c0ac1c28640f77fd8be9514efc5bfa3f3d8058a55b97a2ad277c61dbde9092e73cfc48d4a4708abbf3a0d3a90bd05368be3afcf67e0fbef2e7d31be94fff535d91d525b20ab3b80a7e4c906037ad9ff0daead8c0f4f8a816b1f73a78791ee3fbff2d8a2006ec781fee783c39f5b7ec9286d835c89c1ec8be5bc3ba406f5a38716f3b840464bc9cb167ed1656d758f2c5337eb39115da0a5495f36cf2a8a8278d4c1f145b9e13f36d5c6a0dac98eacb578229717e93629b9d5bae07dba24f600106353168bdb42d8decccf2d19823b8aef38bd7f980afaaede10f8ba0ecde38db3e2547d22f906cdb5477080083764a9b39b0bf018e2a92b4d4faa5fec36348b7c1ba43084ecb6b285b0e07c1b387f60204c4c78af0f30a2e0b58127368f1180a85f760a7d29b3ed32e708588c879609d93f467f3bdb52f44fc7cad96e10c3032df235271f161814849f5e15483e12d8c3d949699e25786cd000e2023180439ed8d4e6bc2fb3f14633ac8f6cfd563135e424f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'hc805686ef513610580b33772cfed0ec8ec077756e3b6956e7276cde9874bfb7af45978f1e94bf729c43abee71442fa1328f06ffeeacb37653277df2557d9de448e14190a0058b563274f9efc4f64f4f1b832ba59e5092293e53af2d10bc7c6d19b92c41cbe3da4876b67d27dc4175443c1354de86d47065409902354d1e56c4705046ce800fbf88e4ac01c319bb7de5d0ef4d1c398b331591bca188ca6e3528f7e04a582ad83797f78174528b278e3c8e53aec522ca03c7560ff7f2de5f9b8664a1b6e908dd470cc0947f88d57e71a565d602f544ef177876b80c456ef57b7c843d16acc0b883c601a7ddfd3323b76588aca4180b03ca98f21e1c535e091560dcddfeb819f6a864f083c60af62e10a5504abe08754c574a227584c94dd382fcf39ae0c889adf3447fdeae3a07b4b56d11e6f399c16d6c3c407e84dec597d4f262a9e9fc84f9ef0c5c35bf6c6438bad410f12c20c3ab4c27d79d6c7de73e7c96aa517a82599dbfa349d386eb4bbd1d0a1fb4cc6bcbae1085c328461fc32171d1cb21343b53708484bad250f028f7a79930a82d17ceb9a784c880418dc25c4894ae77029c9f20c7a260941a68a9e45c953bd3228883529cbde32481c8b23ed668cefda776fa8b74f160ad9d1529418fb6a02ad4f0b8cd3a71467cf3bf7ab8b07e6d2e1863d90ec39c8292200bd5e9ea97f48f070df72399e6c4fc192e2a1d88a3a83f7edacb5f51d5c81badc1e0ed03367fdefd5297c43c894601725dad2c44f07a5ac46ed1ed9a30f12bba00ebdf86220f0820418c8ccaae4a54abe10a7a334f2261182fe70816eff76314fe184e04a3dcd07ca24c31a9fe8125349f9c907b0574362e96085075965062af2685cd9826ca6c9028a8aa699994367e92bcec189300cc7ee207d2f372ed80b16c84612658cbbe4726de70a333017d1e73a15e205890dc0d4a4663c784083e6bc9bb98b0c1726e311c0e1c32f948d80b3225b76ee183f85d0714a0e9e555ae27e1964f9cf58fe632e3bbbf962077592ff7aa5625d1398cee68ec570d465f9fbc45b269f6b3ecfde89b882a2cf256bdaaabc763b99a6518510661d82a274a32163bf33cd4769f5aa46def41ad65a307a85afd5b50c11e71d5757f907cbace02797de9237b101d2a06220a3cb1d625f4a8110d0ac6b56fda933b9147db61b41a6bc15aa97b4f1713f307508b947bb3334d70de765556e48188f0722e2a5b37c5afa8b40b3b9dd42e7ffc92ed1e92772be9fe63e309d28bd430576884cce9c518ad58645c5a0832c9fceb873bd06d152bf98cae307f902d403814b2036b1ccdfade0cba46293f4de64d88f38e96d755c2d20c47ff783114a29eca20dae0b62be70f7cb4dbfbe2d9fa2709f43237db0a4afe85886713496ef2dc506c7f44509cddea90a85b3344f67b8e86234c7e4325b708439bc48f939cc36813e557127cd162fcc1ffca402be0150978ed65629268186de38ce726c8f062147854ab7b9fabba2266fbe8a666eaaf208911500f1546a3d6204094ac05bae84eae871b384b65f9d700fd7e0e2b72109032df83ebd1aa873e95de35501bd512a838456a0f400b0d482bbef16b2e0643181dfcff67abc673f3a24ae7e816acb9e9de0825c37e37bab679e55103aa39ec8a623ce499dcac9d660ca037d8cdcbe0604a97e395ac3d6a36a4075f13df68570cd0e5acd6de23bc635c76834c7c9864020f2a27a522893de8e3a9cf3656e56ecbe5bf8200284ccaaad296f47377614b7a7a5df30813b9017eefaa2366c0f445ae877edb8453441a95870d203a2ff9e7bb443234e748fc5122e17e006996c9b1a8c221ab703540648cd574a98c4e4f9585dc69fb6f87f8d8fe4767ba5cbe67657dd74f9b7ed23b5788f3b37ceb3f6ffe69751975309f496a4810aa9eb3cecc64e93d13341636498bb77c2e7f3619a710e21c3014cc5d5997a9aa47e1a75fdc92a6c03d68e3ed4f1fe4004901ce187b30a5b0a3d0b9152aee41d77460ce6ef5975e4d31904244fcf0735a393125b85891ef747c8a2fa5cf56fcdc7da8739b730fe16fa77f9697d06c4244cf414cf6c78f0551eff546b6d74ca81379973138fb7afa47cc38881fd561fdba4a8414adcc0b9af5849562ba8f38c5e7d3a7777984c095f671e7de1ecf8349f0f6f0f45c53584dff1c7b34d34ecc12f2f36ab32a264bcfc019341a8c712d9081b2d426923f654d97da7cc4e2ad9c37ca6732e568b426e1fcd564ac2ab9c5e947f9eccae78ed58fd6754e7c632e07cf4437fc0b18e9779862a7ae893dbe9b3a4b1db395a5ff892ff244593be37d1be27414f641030cbb43c7a572eda7d6263d50cc94e726b61ac9f55c713d10828492ebeeab3f010d91f5bd2100fe795e28326dcc3b66fcc3848fc62cab0c765282988a15c646dbb450710bb5030b0ab12e716f9482fd1c74e58c0a442f5c59ca3832cfe592117325fc823e21b0f38d9723069f769c5a585fb9dbe49d7848e53f7503aa6a0d683be65e60f2455a266a6445cf709af6c87769d05c8ad96016ac01e05d71a13ea5d4a71d400d855e6753941c151ab93718912ac652c013263d7afca2d8325fd50892dfc049a13bb58d5e0db2e990ce3ccf5107a44d8152858d9f1d3dcbbb66d4cd384d1ac277405ae072621540180525518755c5c95e42b852e3171dc206ad665efb64b0d706105088520a03bab7d05169e96f83ce0e221a9e9c92ced1dcf6f767c5e90918da8cd3ad2972123444c7e15695887fa769c59c80307a53d4b2663e4e3734455684477a0e0cfd8007bdfb41be23b171cbaa849c51a707c40df778a2fcb45a3a55e2f717f591c2524e6e2927a18b15c9f6be69a116ee6119e2e625879f44ea98b564452a204702158cfa970c2ea9f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'hdee1b5a56c6af3ebf3723f37a6aeb111372899eaccecaf788ec34c9e2146f28e80ddfb7dfc0628a3337857c2bda0af353bb7576c03bc73fb01a546ce6a1da237bcbc1d43f08f50f3e16a2d456e2290bb7b10972a78ecdd994aa90f92110a49b72dd462eb0159545a01733980fbbc97ddda9ca618b8bb75637b219d1194ea90958578dcd3f733e3c9f56fe69b96ecb06df4bea93d00e470e8579069172a4f19e56e5d9ecb0a361ed84203a3f67c994b5002b252cf7eb9c1aa698b9762e87b4b3bf0035a9eebed88fe2e71a11de0366c7c8b44b8a77772a890e4059ef163250fec72a958cdc7320adbd94a0611849a4845a683248c226cb20b663ea0a5c0dfc1ca67856586f057f36d17081e1de428a3fc655103865061b36c6f3996d4e3cbc78c8ac8f8836918830cc0b1cf3448aae1bb80c99e07c09d44871f4ba00139dc77f227049bd3429aaa7b6d1d61b34151c3e549bf001eb829b5dd063473c1d7970dd6d4bc0a163f8ef3b16282134efdfed8544ee9e7fb67b1258bbb594dc48c6afffc7b9cf0a31897cd2afa1ade6cfcf303b58eb6a1016bafdd9193dcd3c652531a9c4aa4094d36495b6b99669c84b3698dae035c2c87f6c3395b4c9fe826474a87e86f0cb9bc554092706cf99e21256d03f2a0af2f7bbec873e393d58b02526530b895910a84d8622f6ade6b016304b7163bb3571ecb41ca1087aa18345117b566651e50495a42e4956df67076ebc8ffad9e40ce694ef9cde06b2d47ab59ae02a282b993d2041069b947c5a942e28830fc8104b51d891fb39ed42313b7888e96001ad916c7ffbfd903f25443c65bc9474eb6f54a44761e0fb270e9125552053b5dc0ff7525afb2ed83db2abe8435cd0ce1b8871ea3d7a023ffc3a930c289f4cab793670643aefb481cb896e5e5482b53bd8614028f798e8777408febd3d1ce6dbeb5a17516d1f0b4dcc29aa19790a494cafbcd6b1cca4e8706e15afe62ed504bb0c7ca83486dcabd85ebd35a2800ef0665a2366b4b936390b2665b296bac87b1224df78a7e3261dbb3cd713175096740438697e76992b2384c84cec94d992e92c75332278158ee6d33d83ff109886e12dd555dc75eebe1cd054f0bc59b05e5dba2590f7a1cd6143b848ebc46a1ea8e94d06d47060f02bad5de1c4f127341de6e73992e62c4967722ffbdb1e4f25616aec8fccaff79944e259e31c1639f2107cbf9783a2c49749f3e7c6e91d57b5f3ea12d4331988411038b262408b0ed42498f7f5d0866e906f0ab4e34abaf681454d1bb65014cb710142924ed70ae8f850c4507c3224c37afafbf8b11cf18d640d624ab8878d70b5cea9e6cf01db8d50acc16a7f7fb6526a1c93a881171c6887997af46c78ddddac8b0a87e9469c0211394ec1ba445770b1fb0a8d0bb99a2e15f52a76351eccbea2c7dc670ee4143b237b5c692d78a180ae433794a523acbe2b651aa278ffab3ffedb09ebb932fd1328d2c30da211508f41845b8e86f99befe47f368b3396d50c38ae7a34f0bd81e022a9df0a12715269029c4e165a47d11aab019e935d4fd08a54ebc2bc20ade32ce8fca2edd518fe3acb0934f5d204f563d0928088e82fbf8cc98a7af0742d5fd3d3b3f9a547b86a3e20b2bc923e41c8f042c2f2d2f0d0f77a1876cc48b269df0ce61179a232492fba4308a7fbadda4096c40eff4954338619db720dc4f78c73edc824900ad6edb6ef77753c00a8dee81a1eafd96309bf82f4ec2ba1922f8a53ded746568d350ee3eb45c154627c767bad43a6f0f2c620ccceb965d2a8fec65e45de476aabe89e2ac7a436fbea6f0333b2ee09ce9b29f4dc68a80a33f8fc5b1735d1e955d398c88d4ea2c1e12bf61363ae40cf93c384bd984db0358508209e07d7a677a7bd009998b7f788d5a73ef74e9abc08274664fa0de1a0c2d9312e87e1862a85e74dc76bf7ed7f7614710a9946354eff475ed8fc439985d09050b145cb9d9d1ebb1ab62edff8ab56f553709a88889cd442795e0ce1b946d73c975d84dbaa88bec0ecedc036f8daba2c40b8bc59a8791aebf9effda8e94b28db36b8b7ce7c6cec57288cf872d8febc7514217c68053170230744d6295777443336317154431f71ad2fe5ae6a5021840ee4040a8f6742aaa107b9a8a8513c10230d9190aa8703ab1b37eb611cd865e23d0d867a27fdd3425f53ade3c4d6c3d871024988b5c6d68a57bbd9a0e164d03733c10932d5077f919e4a915301c285cf572634a9a5308d726c585af9bb71e7f8f375a7fa5ad0c178df490851f05f8bf9c6e0d8ea9b2f7fc44be63d5c0e401c14adebe10b0bbeca33f0bbdc48888ba11bb27cf515dca4b8b50148f9ac1b8e0a14f0f0f411f6dd78dd503e88ab0743bbc780e950f585f1554d3ab39569fff7a237e367ec087f885972cd57bfc297b144d941a8ff07349a9a1f8450d2490b1030d7402ac3c80739afae47f83d5af41ea13ebcbad3a009ee65e85a81128e60848855d7dd454b23c0ab9e21b085be2021880915d2eb591bc0dcd7c65c4ed36a77561929ce6b00fa5d6f086e3a2d54968cb4f6159f3b4c4fa017f115ee9858621aea4bafe29f9165d0ed6fb2f0548559d002acf25a88fa1cbb5308a2b8057c35d6f7d21afc56b0d8eefea78c3d1fc98ab4bfc377c077a701361691cded46f2597796ddb3bd56a50273a11a93cabbc4ea3a0d9ec9dd690d5d6eefeccf13f6c8cd55be85597ab206cddcb59d7c88767a7c4fb4025e9886f78242bb0aff250b6665495417a5673ae981e1f2caae5143284b959496e1a84dcf464f344e66420c1ea8c44cba319839991aa6dc840549574592a391c98400be5be969667da3d034cf163db95d41df713ee6ee2c306a401f74122644222746c35f14d0a363661ba5c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h1e0e9b8df7f9b53e25a788d3bcbf652e34935e3ac925b95fabf38bf2ceb691ebfe562abdafeabecc504fdc75bddfc3eb22b2726e9a2d69468569a93732e8a3144fb2ac86f27f2208cfff6260bc816ec12b98eee3de33185ce5bf49a4f4f70fda95fa743e7962ea62ba29ca57f241076ce43611559cdcf641ccec2c85dc96c1c7c9180991103e20a6d0e2039f6ea96d94b41a3ccdb475d1643c0e740b77b4837a914047c21f252547af0ca32875fddcc6fd4927fbf19fd7bb905ee446c880ee751fba809523fab0b4302a9f130b800ccef37aa6ab8d2518bae81c7d6507603ef8ab82c5e570d271809166101c422f088575784bb8df869784d33f497beac6ccf8b5ad9a91e82f88f818cda07f42c0362e625bf19ced667d7c7d31cce1d56b7de60a481c6feb9954d71087e4b323adc343f094d492edc624f9335e111e50d9d4fa5c2838f510fc9f174c4b876339a290879d00e9f06f19a453c34467395dba5ae858d4bd64d76cad689910a1027e96e921fd0cd200a76a88ce5225bf6d938cbb35fa786ad3fe95852450ff19e26e9162a3314d387c99c71c59842765c2a1645cec98ff07cb5a608c8fb9b8ac5a1e30c1cbbc1e12af96e57adc092f6a723e166e3d5972c9ec48ebc0190aa6687c28252e62a369f74a6c6e3519f3b2a9ce07529e144a54da71e4c3165ad3149feee458536830634c001327ee777443b13c1d17c4295c7eb3901fb38a0b7b0a322f011071f1e2513281ff75ffa5e957903e2b3cdd680033890f8358dbcfea7fc282f5a3708ae6b73630c144751553202d171ffeceaf620985c40813b7ac363865066048153c8b918c7ebac8337233b3c34b1a0ea77256a2936e412ad392eb8a55acf1754b2a1a19b2b0656661a566bff12ca15cfb37465d909dab67e654ae720dd40a3c0147ad4c44a3577a7335eb27c8d3abd312825d03ebe0d0cff4f3b10e3872291c7284c4d95b653bc59e95595603e4c351aab9b7747059f53bb11eda7065835c05cefaa6a7963e9395a7fec76ed6dabff06034e748d3da296ead107d1157f698d97e510ea0363ceec00c7ae4ae760818dc713d0f0713f1ab226e641262261b03e6f5733def10e9f5a8387c9842a5ff51a57962930c3e5a517e9e5be677c4594f9235b613bd19daa6cb13e23ff6529063a9a5829778c9b767449fce22989f15e000c9659529b34ba007d3f3544bc5ee3a481a9551ad8309916b0fb40499da54f358c4e94ebf0a0a24a8707eec40557a945091e6ca7760cb6d48b927615ab51b80eb21f4ff2f25dfeec303bcdea8a3723792f9b59ab920ac9628532c6443747753f38befddc81814adbd0cf92e28b72f36bc251879b39faafe90fe0fa23f4f527f4e6f5beb1220dee22baabb76e66bb2c77858e99cce8f731ec0e3cc4f2fca20a16e7c56b11609370dcdd4d776dd58ec155521806048722bde8d8f4f0b7ea1e840a57011ef904352a83adcbdee46daad35db85d840254bc3293004d6c9772af3e489fdf2dd5b9a1f0af81bec1ca949233dc87416df45a9b09275a1c4f7495aa234ae3a3b9815d35fda62b17659f3c4aedb8b85e696f7442e2aa334b6c99bbf76a7971635e287da0230785354fc2c4eb2d30cf6b9d116450666ab429f620d346aa599657cbe108f1405a8de4986b78d91be96280d022f515fa18c788a39f133012a1826011e61a039fd715f6fb9867cd479073314d33913ed4df04509929dd4eecf995e85f4f508e75149c7c22a51f5d3a06aadd9968ced1ee4de7bdb545b8b0ec9befd8d29ede3d62a27c24b3c848c2ceae18c46b8b7539411db657ae86180935140711fe8ed7772633533173f3aeffad24b9323aa7703de7e054356b360f2b1726743d8fbd0ad6f0adbfebdc98a44fc51a6ced45eddc167da9c276597b533ff95c601bf296cf62e9bed89284fa58b0d784b7d3d6baf02c8426caed8bd2779bafa45036b2d9d92e43b35f7789bcd743b473997dc3a078b7f34b853f689022a8ec89be69b9cf3096bd9be8abe237a1184368598f9083b3ae056ee0ecf4c921515bb1617fe8649c004560e703fd87ed4bce014ec8af4246af8f8277f90deea8ce5545160a100bc569d4ce1a248eeddb4dfd9476fc9e0bc655d8cd5a93b494340320dcbb0015c840066927267ffaa8341173fe30a9375987aab72cf78961675754c5a5c71823ae3b5d8cd4907aa396982dc1f461a92b4f7bb81ef1f509234e356870df8e39f1416c6a84a55910054458deb1e5a9ae2434637bcd84c9658f7b3eddc4789d944b6d61c22fbf9c4f034a605d970ae96b2ade5dec828a6fdcc58e7343afd0811cd4ac44352f3b59598c10cb485e6f4fe08eefaa3e2e74023ad22f32dd15b3b0118595691a7cf5c18820a86101c7e5a08e8369472cc24ed22f03c792ce3ad692a5725b0e6ed93311f680ac410280def0da42aece37be58b191d5ee7cf0249280c648e7e4998257152d2bc20e522017d0ec932eda1929826e64dc537b64f1153ae5e10a3b56bf94a7025d3455c957a60137c1b377d9bcc67a60be94de1ef4ec2299301a2409625d6997ce96dcac00007fde8b09503c05613b48117e01c6fa5798d0246405a03344614625479e7385f9308f0c6c3daef2942169c9829ff57e32796f9468eac063010c3bc354c0bfc4e1701a89eb86faba423d43612c691933707747aca1af9d5b4366e5eb6dff1ee4716720cb93e7743ecb1de76e2e8749560ecc33951f2b499ba5587fb2bea56aac4a57504ab1af65543a5c73475be78ec47fe79e60a0d9ca7ba9c32d84c32c321b7705f172ea57ff4b8eba083a350af73eeaa6dcab9d7e3886f9694c30b858c31c965a05f1b67856f151bfaca770ef96960261385b08fe95fca7bb94de999c3d1ac1cfeb2;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h79b3148948ac844c283b35a658064391fe061403335358c41ad1ed9820d409e95211bdc879a5d5f69ab266bd66df976d0720972e51a1a15b9439cf7f6b996aa138f350b5846767a324227b99980014fb4cc5c18415db8b1aad1146a465da8c3b4ff05642266bb227d425848f3c64f13d2608ed02790524771d2f6583c50e0d6102e8121802f6270637c9d5ede23a83f74d5dfb0e6fa082c7745411d01445c8d7d6f37d5d2c752f22af1d19542765b7736c38e5aae8bb999e0cab7a7f3e6430b3d682865c5fa61c8024406ed9bb61a38928a2e4989908bdc3013e39c94550f52af51e0a859640e469a434a095c17354a4acc50123102f59ed538019fbddfd0aec42e3689a419a744fbb37dbd33be394f3d610107a2d619e323f92387f60e2712fa7f05743ed878060110e1d270b703babd4740aa93707ba4ec18b20d3d25ae2d80f8e8655d9fe030e59078b9c7c2aaf2c2b028f91d2f4ce3b88a0a4a2d0e71c9e74bfc4025af2c6b0590cdd22f259a18adfb2bd3c0e36ebc64c701457ad1a620cf3153ab5a9cae21a1af5d0c903f4c42a206934832347ec5dbb98a6d49557d718939d6b671a586e05db7dac3edd55f438afa2386096cf971e487fa651eb7d212b90176b031f5673d9d53d8315bcb064e5cc08c45d6e97f743daa600190864d202287665d6c8529d8a1cd4609a5e1106eddd383ab76487e4b7edbe4c01cc76ac33fb6b108b34ac8bba2c5e29d07503e973623d9bccd3d013fcf5785f2d67fdc41b4e04719ac726774a42f6b105340989e3bd6e552ff62bad9807d6b0877b74ea70b917e1903bfcd1ea8d038fd2b466ff45476f38047f351ebfccf58a7dc90917580facf486e3abd991481295b201246492f55bc4b6dd0fada0be4ed9d5b6bf1b8e5b6a60aa34a6f20ac5a654d50e852f0752f86f0297b70b39ab025f601698ae2284d63d7f859b5e41b1a608571c8928eafbe42a32cadfd7d865a5e309c36990d80609bf52a1e3a8df8e40ad048a074a6263cc2ef4af8a5ca5f66108f0c0a11fcece506a58d64b913b7691bee52df23fe00a3d801631399ee3d91ca3b879b578f9385cea434baad903570783313e21b9a8a772f29ff5c7024c94689140a1ba04c8da82acc82c608be073a9554a65e8511a0993395f5ef3bca30b3927dacd6b8f7fc483e6e9a9a4cd73abdee47a2f6a96b802e3506c49b2c72442b793878e88778bd1d2737516059cb9f9ce580069ae4238a764a3d193ac3341c1f7b838c4e884944fb6fd065233ab834583237ee2aaaa13c59c2e958d93ca5dfa93aae5c77def3e1b862d4d86f49410482104558f2888976f093af45b04deeb667c5870c1d09bc7e1daa5faf503a674efc593699c79a681f055c2197e43ebcf52856c209f742f17bb6ed52d75b1058f28c3b6081236798f90acbd8571c609b66d7929ff260fe104683efe48e3444dde36229741e580b7a425bf1e7c1139963b653cc5ab9863da056fcfcdcb6fcae4fa9e8441ce166e362056fe3d38220a9dbb10e37a37d5b178a6b344491a89c28cbee1e7d36415989752deafd83b4b992063bf41458710843cfc98b119001f21a0ff45820be2d871fc531466455b873f7e077294a83d0f41dad3ba4c8a9d8e357a3667a12000f373d72f829665b3e8315599f247a1fb9a6d4f2ad2a2c4b6ae91537d75cb04616be7778674ca249ee89056442937105feb928d894abfe59a84799b2c824a9db9491bd8a1c35fabea1d081e87908d4a1ad44c748a69cffab04e3eab05ce7e5c33a9c83e21cf62359139331968c845eb0f249dd95ceb33d52ea5b1cdfda9f9ea1c3bf28a3300a39bbdaffc66b6e2239a9001693bda59f926498fab95d127927ad0a43db3f1d72d769b18c30fe04f8ce9b06a076d791d9b315d2714ad50b0a98b3d646579aad322263d8744fe695c2930b9b48128d005131cc5d9215dbba186657ce6a9fd44f9a80ad513c8e0dc65fbcf8df24d2b50421f9311b21915db1d42bb7ccde39f72cb027883d2c9725fad1bf76017976008f4df027b3ea0b11feccbd6c7bbb75733314ac6c39a33c31400c33ea60fb418e5221593d13e99f0ed4e9b65d9aa3d3337ccecbe4d0dbe63e8c8330526b9253bcd437badb0b452858f91c876f16ead04114302c92503625a0bc3c277e66e8c92ddd9d8afb41cce82d808856c29c334c1f98951b9c548a155ad7d8b8528f1d77d38a66c58c75774ce50147894ed70ebdd9904ffe69a3bbe0b91bf804fee0410420e2da205ef5f36143c3307d3e65423df445611e89eef9c285b08ddaa0eb9774327d387346289eab613751735f23a3b5915c1272a7d66bcb24d770c196bde4d83bd45c1411702bbdb884b41e89d2722c98695b60d6ea85c92ff12d4a4efc48bf74ca349d99e0a6658aebb1a8fa8d65ef4d5e8027d90816fd5ac0f2e53dd7510ed7312e6b0d7e6dca13590ba4cea8467035f1f81060522a4e1f1f681840d78919375405b8639275c89500c6cb65f54fa2f256b33c92566b04ef724443fa00c610b2dfe8a22a1a7c479f0b3f092de1a0123ed83e02aa075e1f00e8c0b1c938f02b3bb0789cb3c149d0755eecd667b644fc7cd9310493e7b24ac4500f311c93a669816ffcfc0edba6f363c48cadd52701418edd6fb69033084ce8f080b98f1ec27f0e2db9325a531b4034e5bba8145d41d96dc46d797fa3a25174681ce0dcb08ee61840393657e1218a36c993a445e2346404ed11f2acfe70cd4b23f2f658346a2fb9dffb38f4a5e9119d076a8b046218b41ee0850e099e813fb1bc167c76540185c79d0130444af6ffafeb2483829f56d75c229e35ec3b812a7bf2176013bfe36a97c8bb246a3979aca01b31cb2663dc902d410cf082c9d64db851f710d793ce8af67;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'had7e3309cef44c9b68135829ed7e2dac2ad517d7da1b08e27874a669dcfea5de70f3dfd8ec99c81908665036322c8681947086d2a84ea6b04bdcb395e7e390d034fb96c87ee8848f07c21221ea195874dfb5f9184a60c1307c872db01366fbec34ae3b6778e098db9ca90ab1b1ed7a8759c7e95b1b389ec3c88b344ec9cdde556f29dedc4814583b7561f19c599c86a97f81e0490d6efdae973fb2d8116912a7294c7c8b94ec5fa394bebbc238566c49436e097b483bb0d09dbdc8d155f653e232e8feffd2b3296be21e25807cf328e6ee62abacc5df8604f351b7712dd0a8f732dea0ac15475eed9605531af98932a86d36068e2b3411104ee6aedcee8c0897128a820f76f00f2a4e332d5d097bd6a51591ead47e895e75cf9b373c259318124aba969c57f22791e0e90ca048deaea103f0eb1f00641b15ca297fa0852e1282ffd38eeb0d0ad6ce736af88c3dc58f8ccd6d8d21e382e4b3b67e665556fb5df6d894dcd70b12820150eb5720e4f2f71d11be8d9b204b266c9b6cacb17d39720144e5f447157a0ff7694c8f55fb9d829b4083b52fcbd4a6143ffb6d5d106b83a0be108a64b24d67e057c0d021ea91913db4718d8ad8c7e3beea945047ee9a0b1e53b99e1ce496d74a64b453e9bbf2e8b874cfe059016db9069d4fe53f0cf5c05beb0ad594c7d32487f6a0901238c8ee7b7295fcffb64164735e909d114adff563e1a6e29a9adf1a7ce7e84886f72d72453b0c6b5bcdaea9f9c39e5a6b5d10e224e6518cafbdff4160f57d13e2dcc4122ab4478147f1b188c52e997e3064392cc83f8d0c156da0b751a3074078e70990a438d1f160f91a59832a8fe7ee9e7b2ea0d6371d74ef20a97f0584960aa6f5145c226d0d7c34a852edb8334636be5449ee63889022ac4e6eaf7cbcb0d9d44f258e74cd044d908d5bba2b5add2dd93a93fe08899b976a357f0a896329c39dcd85eaa38fe5595c6bc0e45456e44df1db75ded11b152ea463dd72020cbba12feab54e12f6b917b44ba12dd629b6e331cc924c3f303c6dcc2f23979488258c4867a389f37eededa6822476b287e373e4b4793889aa64981ca3c2dd67c15fcc7ef198c4aad94c87e8b7505162e84b44ec09705bb6b73e8de4c5658146677d1d5922f379e487589745a300a38493b01824d1a45042d494db9906a9f7dedceecb019e94e48e7e26936cf719206f480811bffbba5b42057066de548bc59ac2817ac6577e314fd12f9573fa833640a73d2f42d2b7b67566fe025f6a091c6fbb46eb6fa81d5645576c45014e3642c8b30f36027c00a3e08797180eb071bed33f764c96cdc544669aa680c1b8c87ac49a226ff3f3a083e93e6cac19fd0314c66412f070088b5261463932ac3fe75d7bb76d4f42c23c1ea6d0f7ec9a4b714e6adab7ea76869d2b310e0d10a44bcccbd7a24f59a9802222f28c37badb1d72a3913b91a16567eb9c6059fbf7910ff036e35e64f467291c6bba110f66ab33459e7a34b747a7bd245de657f8f11ee8a4bbe6a2b160e2a7bf6c2a8beae1719cf178fe073e2506bccb36ecde992f6b0df1e5714fad88bd9d71ccd358b8d8f99b88aade3aa5e91c766d886c3427236a895f435cebaf8185e154aa28f91c2ad1891272f455bf1b6aa308627837a1277b86a7e675173fff29b67734fffe4407602fe36a02737c493ebf9b8ba8cafc1a4eaf448e8c65585db7aa58497496c070c254ba87b9cad7b45f8c9c75199406324ba6cf656daeb0bc2bc49e9a9d5c47546a5ef0de7e590a8b1d29c0d8c10a1a75126a9d13ad55994c38882c23893493e9c1c4f665943d044d04cf939337f0e4ef56082a822e765e9136ac8735523c2713ab84ab9120f668b8a4b9c42dcc814b548113140f6f361db49f1403d03d052016fd091b36b1ecdf55eb837a68c028211e9edecbb7465e2e0b1dfaa79edd9263f6c06b3e341a988c8f381484bb0c3cad1b9962e5f11b8accc3c17dc558e7b451f01e6981626c524688ee369eadadc0b325ea1098f9930e985163f3cc28541f00eab22edc132eafa4805a01bb8e02d1bf5ae528fe93542df3918622e0ce055c031e7b6e0d4d75a04beeab998cd62b806a0947179b91bef1a7d28b37ae0ee6c289cc2e142f43a2e8df1b5970627b1f88ba217c3a46f01850d7f61f8aaf9457ebffda7c74b53ef19d1d1c2e1f93322981a3d7f5222041cc2d655c5682b2490db74ea2d4a66e036f2bc04430b6acee44aa70c88d857ca4bd4f579a0886cebb01f9f1eac5804cadbf4bdd449e34acb338911fab738e8916eb734e2bd906b2861f5832741db24f7af14bebbdbf6baa36e655940d232dffe703439af35ab5a0252a95151022b149a650624b286d77f98b09e022a8cdd3d28e8b0496eb6821d95349b94a095c9bef7f8483f5c5130ad29db888829b79f17a49c03506fc9c71335d0380dab0e0c9413132849de00741ed6f9433501e5f0f843c7fd8ce4064292a95c11babc879ed95e2bbdb2b0cc7ebb83dd24441e54c2cc9ae4f031f8ce6eae26b5dcc9acf61785e4ecfbb94bb19a77416fe5a45ff254fe29a782f65dfc74190f833a8f612922e0b5a960d589f3682886e022622337314bce334305e5d82a6ffb1cbd0ca46b1c691e3a4bc5443047a2e5bf9d2c345ff5cea4160e6dccba3d3cf660d495b3c0950086af09a0e5453c83973672bd899e8db29e908ce1fb59edd9f63cf470fe7914feb792957862f8315b17db5c2125b5ac0ff32096df56f2f2b4b083373a33d49c5225ab26d30e753c3e32fa386c2807ac77eb4181fb8965cb0c4a433ac653fa601ed1ff09d09edb5b0a4394b30ff2d1aeac046f54e85171e3926c33b67d799f9948e84ad7eec943843dc7dc9de8f989563f51ff8222bf71ddb904b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'hef23533a60210ebd6687db7cf596e569befbdbd6d8368decb82e6146e672e884d60b86861b4e1ee3a7a30a598cc0a4469fc5f31835910da8dab30dbe8b057506afcfdf94ba26b843dfbcb15ee791c5da1920dc099a38b6f8586dd2f3cfd1570a99fe6911dbe3ba8ee99e5dfe6a43898aa5e63073c77844beb5274f0b0a6ae86507e4e8f5caf221bfda4001daf7c56a4f0eec9cc3a571f3dff504d111ce3cca12015b676f8361798b65b751cb4d23515befbb6a57f88d68672f7c423b6b8067b359d48e419e0d969c492525be8bcabadeeabe81847f3f6bc1c55b4d8edb5f4d4b5244da6db172cfdd6f734c98b2a12b919e5681dbd4d868ef43b72ef3e4d3b187ad100951961f6f14b7a5ecdb42c35e3b0227f54eb5f32dda67d9b40a6241b1d440e6593a7d0b637c6b8356553f9c360270665804cdfc3ec8a52cc57e06d77d8ab974d65461e1b10231479d343eb65c60ab1a0b9aa5787fcfcc4425331c010319a561901ef6b431e7599e0ffcb57b3d3638c66215f5099941fe4da9cacefe8e95fc8cf202e6568c30acfe62a9a9d46a6fcc449a953196b26043f2f2440c03c1921de2b15a896653c315ebc5525794be1914e125eed1fc73c06199c490abcc719ca1a15e5bca62a3d114831a32acda4f91d12dcf90e5617f77338e23ab2541ce049ac8ecc7c702f1aadd4856548a07fbefef4e769465cf666c3f3316a9bbf55bfbd5d80258ffd962c2d0ae6779cb39ffa56f6139470585cd56b57e96e126c6057cd4e528ef67a13a37c3b478ab668929534fa1585a5298288f6799454131fcddbca7ce3e142815e62cd8180e313b97583786fa08dae988cee6c4105fbc384a5af01cb784d7a8d25ef0d49c9a1d3cb3e07f1364a286d4a568ce1a0aa047d8268126730b76e368ca2ea75a1521511285e6e568328f029a822685e0984122cfc8a73f78abfaa6bf959baa89f052bf4b35c635835042b0042005147579af12327dc8cc5480128487577e6c93f1225d6ff3440a0648e94c1358898a656da9d408733e2fee716a9a9affdbec2341659650d4d33fc2c3ffac53aeb6699d87df3fd4e1f9e838f9bc8aa3c5808c0ebc5070321462bd3d6bf7aec4912b3eea2ac6dddc29e6f48fa4b2988dd40def2ce2e8eb29699bafd87936c58a5259ea06c921bd4a688e2e349e2e29d4fec06cc5919e4a39ee9b6c77d51e909e7eb6460929310cfec4b04ae409a9254f9bed20fec25c4c92cef3446a94d3d72392c766a0c10d9a60d0550c707e8b9ce6e9c1dfebda2ae2936c50a70640c8671282ee5c53189d5bf8eed0d82e9885e40ec3008789d801222b4686892f3174f88f7bc8f3b269cba632f0d7d8e191590b6c06d3952c2ab43fb840afb192de1ae2b1c6724fbfd95c45dfffacca1af097d12d9bfa138355c044bc6badee4f424240ffa03808e289d11f22b1661a738f65c49e38182a1b3553140cdf0ffef609a18009b50572a1ad4341c3c7234b714f305d60760cb6fc52f595f798aaa50a240314e02d558103eaf49375404043c07854ff98fd6298441b0a04712243b98a57a9f391df9ffa0d0ea6114cea08101a841cd862b58a8a839daebde3cca66903335cdaee778c71647cb02d6e7e6c810d09c1647b6ac20268661fb8bf22914c786456f24a06aad9d2a0f36013dd8184f1230cff349fb2a86aadb6e4cd5b30723d65c4081a3e7eda5f31c7e279817b3babed6366def26ada438dc3f8e351f20f13d4be2ac418094d50e70eaf6b4010c9dd26ba1009bf3b36a88f3924eaffe38302d4435e063fcca3a22d219b2d4948121efd217b2fd85c9f839a75ff06df43d6eb6d9c2646a927b1179292c4de2f68f126c9d7c3c7f73b17ad56791f4476db7523f4cc76ce9de9754f7aa33c1fefa563c8f474a924fbb94a2186d53fc366420c20eb5e211046eacc87c54e88fa3857bc912f52d7eb3e8586e07737b091003deb3c4e9babc19f7d2dfdf9cc24eb60abff19b9a0a7a9b11183d449b267a8fc5164123d83548fba525ac4872044e5db6d2065e64fc37e718b63329fe4059fe4a320d2053e51d5f1f00694f0c97f593951236b2645768a0121df9a20218cd31e33677bdc4546cc6b103055af1fca6b8174e4f28f4c3d3157913dc154781364fdc2cb29b1b863134b37986a2529355b29c54649f5fde2e78b252e5da7927fee62756cf447169e0e6648ad00ca7b5c0f5ddb3b97cd056486801d5981e07d18c7463028dd57d23fb1a0eed8c252f0bb0567a29e11c2fce393d450626189142a54610ffd5cda2b1f35c94e719eac3eafe21de7458d0a8fbea8a54fc0792dad5731e6ed14242373283450053cf8adc9bd9c36d36f4870842cc031a4d6e029f9bd4f3a634705dfb9625a4fd4661ffb4680147542a23bd9504ef95edf00652fea16ce6ee13b46846a2b65fc6d466bbcf2a004d9ba44af4be9efd7b07368392718258d97361273db0104b870ac8aeadb8345d15cc50b4c5c1a86c918dc3f232423ac4e94a8bd9ca5b3f082fbcef0f34f80ea718cfeec4b01cd70f35dec4aee8d9f41e4e76e4e96db87839d0673f3b64f5a20b52c17dc000efaf06fd9efbd5fa829a8efdeaeeabf75eca4733cec6201f4516f37703b3458c0d22d23bd3a59c56f102fb54f08c166608ab13c79b068331b3b86ad66c2fa3abd0910d00445a01894dd378146a11efe1fa0dd3940713f4675f1522b69f8e0ac40e2f619ee49227504000ec19dd16e4a08da5a44b82e4de0febffe6a7fad8d15b48ff674eff71975818275b14b221b42ac96775e0961f57c75309cb100829fb0165ebca596e6f9a388a3303f58dbb978f11602ca66cfb08c77c088e897a9ff199666212b92c37834d90de418b8d07e31b111061705268599ec723d6378292f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'hab7c56086366f46eb9e1b59b88e7ea5913bed2571ae8cc00f0c9c56d978046b295e5dfc70065d11b8fd742d8b421eeaf91150d9b6c3cefbddf10c7abe71b9832a5526970f85e8fec3b176cd16df822da4677d3431343c9f9970760de7f3b69d92c4dcdb40a3a56541b8d25416ffda751e3072f808cd3efaad19df505a3ecb8f0e02c3b32e8a4211307709afb53da4bea2c5933bd8a22f796743e12e0366c97abeb24e93c96e7443de532356a9290b51f63222c8d21955a7afa4dfa5d51fd0f78278abbcf413d0f608c147e2ed0ab5693588e42a3caf101d98a1f3e05b45c7471521efb0150bf8ecc769adf33ecb26922a7579d115468d6ed15d444a6ed1905be3347481ac25f1c0e78fc352a87e999a92a5a381c4e08d70387082adfa5c92aec79bd750a978ea521ea165d3cbddf9e906f77c4040bd2bd0bbac12eadd3bdbd67c489826c1cd5ea1359da5c785737e06bee5f6934da2b2d25b3eaab0ca2a2151f8c805d27244674268a45037b8c77cfc6e3aeeb1fedb0de81b0891a17d1a2c5fa82296477ba2d69dad3ba0e6264c47f3af385d08de1ed05379d45c737697c571eef2eea70ed93d9d5599906aa984a29a534f0f95dd86c4f14af61766183339be150bb35e89a40b95e5894acd495430c85f7dff8d44039663b2b8df6e6dde41b7014843a9fb13b5830738245bad3a78fcafe6819fe29112fa0e5b49ba3cebf42c4b511837fc37beb06c045832f66a1407e9faf6a116315f40769ae7714061b88595c17807025865700ac47e1f0ffde521c7b42ae8ac1372f54fec2c2a0791463b9b5a9a3541a2e3f63f7c9b18f844a1e9561c8010b13b651805c6409103ddcb11d09f45e9a2adf165d1327ccc751ca49d083b8119d7c545cf2abb98dcc18f7abe028ffe1cca197e57965d4b8b124545f6c6389bc13b6209c2de54687e28d7974701d9402ea73e04c5fbf82bc52518499316d652ba679c569b6d0c90d777a2355e0c1c0c0fb6367471cdadce46cf6f0f8a13008730b80613107d00ffc4082cae89ace045e8b03d91b53e1d564bd0eee924f8b99d1c74b3dcf2b8913d3c5ac17443e21180c05022bf22f9203a54926d7be868c49ae4830ad3cce068038ffcc420535b9b057d006aaa7d65fb22b0d521bb3911cee23252a9648b2185b61729fa6523a71f95a1208adb2710f8b1ce1609d06c8819723e92bcd2a65aa8e721dbbb5e24e17707be03228f8c746d2708ed3bcb2ee8eb4ebb5606a344ae2f2a991af4906ef9808e543c056503b9ff578a733408fb4204df74db9555cbe20750e3442bc62101a57e18fe5bdc67ec8983c0698cdf25b20c0e700429d62bf73379438773eb0bb0a4af1c7a0aa7ae9dc6be68d85fefe707b1c4b92883cb5f882c460b77e434fd6cc2b5975f32065bf15678ef5f3b0ab21e6ba5f1f922d250124a1f77992eb3d5afa593186ba727a63960e50c442aa3e3b1b388b7b2e6ae717a15492003968ab4b6127e7591b59121c53476e5549c6f448bab7603924b58642be12081c98de373ffaedda3746b8fb92da9cca099fcef7f8a6e28776ccec3b1e95d7e3f5728c72160dce7234b51cc1b2a0a270f26e94b890579729fca2aa8ac1def10f5c262be3c804fab196c73967a6bcc9612b23e7dacf877323d41615572586b460367e2c0893269b7e0d1842c760fdfbc60c7fbdb864800b59cf55f63669adbb288b60cb75d7630d03fb87ab09151a35c78d9eb8da88a244b7ae1f464873f396ca3d7c690f4b3296325aa9b82ea16b34ab39e3257874b8a29077addb518cfcc87ba7008195dfcf54d9080c7f6b6deec649db417208d6516672399b5fdc26bd75afc5d0c2adb7514d5da3d2fb5bfadbb3a5f0a2f1fb358f5332b1f7bb648cb8a74fad98361d817a3150a7955f6feac3013ffea1376cd1dda441646e9bc5dc7940343428a20b3773f68dbcccff9c8e4182bb8a25cbfab93bec019e1899f1f5e8ea84ae59002e16c946357184b6bed296ab8d343cf71c7c87c871055124a4986e6496e1250fa91d68eb2b6d7f53009db5dbcd588c65f16638f08963e8542f9d70283ada39512a1f8bb9ba51ce17421b8e6c75f7a96ce91999d4f22bc786e8a4c6bfa3033b267d7fcf6e04f81377a659bc5de11078c5871e1b204ff7656c292ff5051d2e780dff77aee80ad1984d19d1af39a24c0da8cfdef68e80b9cceb656f5dd02cabb609cdf92d2855f2194cbbd49b3139826b24fdd738174ff39ac2a2cabac5fa4e4e168d3afb3da1487ddd4a12008824244440600514be6e81f581268d2c387c4be0433a8b8046d521a48daa3d61e04605227bcf482af23685c69db4dcdfda52e0e9447709c00fb05369a5a1f81594bcf9cf07eef6139a040d9e9d3e8d0c71c7141f9c8af2cfc099ca8cd5909da9a0521cd885d7b1d43593220de011572607a059ec7fcfac669e02520081a08a5c93cf0ec909283e2a9cf46d8b721bf6aed9ca184c7ea8c9c53486d538cfe1f092c00054a162ef62f74a2ed90b0180e7bad86378a07baecbf87e4101112b29af3f473c7d8e5e6fc3f669097cea04c178b73269955a734fad50caf0ef1b6dbc2db9f83e2ddd657b186866f00d024c7ecb9a1c4ca619cf402825466e8e98818b122f9e10557bbeebf3bcb968d02125ab9c273f81253a06f47e1246512f976cd702203a117998fac7f199d7d12d149773551d10bfe4bee6c41464b7eefa17e82d2e035c6e7de281cd3c4ad03dbd593696690e0b7f718aae073d04e0842f3cd0ace26fc8fb2b6f0261483f9f6f98c012c2e7195f0b26352799ea6ad10ee0ad705420b7fcfa34e1ed058c669feb636047844f6824bc647589c31fcc72880fa95aecab48c975206629abbe963e4a8d21e59c8c918a700ec933e55;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h534451fa752b016914f82508a6d1d5e3df076d9a98098a4f8c2b9dc5ae2c2e73f819f93b552a3fafe1903aac73651e579657935d00da775cb09be1372fd16742a83693ca7e29b497e7781503d214331b3c5fa4c07c7b2f033b88437573974a246963cd667b82ad18b5cf39d01a43c7b7f79d5cac3af4135735a3483c47412075882b4ae4435a94c05f3c3666aa0c413760c1ce3175ab4d126b06b1d665926007d3fea532ff3943a4d38f5d5094677e8709a2d65061b24d54eb0081bcac9ec6c5123b154be44e84fe0ac4e4c918911ea682df4cda9314d70f9b5225c0366de13021077de69fa5f2761a513a1a93affe870c50556e94333549f55637056fc6f9b8112ab3a16e54c10d8195f26975d9b4b2b68079cf4ca81918a7f357a2b7eb916b7a599628973ebe5df4f59fdf9bfc5352e5cb3673478d45f2f9b146d8877b680676930d549da27003331f162021fec76f283d194ccc36dea1adbc4ee67ef9dfdfb746a4ba7cf6c2afdb1ab9f4810cb47b13a47803f69c6e744923c3ab5a039a6bd1b5d2bb3c3fcf087864d7695cf14b505e1ce4fcc8e21b42e69a4fae13a68aa55958751cee8a935d098fd09d424cc4dcd0636a5682c1612f2380a39d57f8aca993b20ebd4a83a8f71640e6e9b197da7cfa92c052172517344a065137b7e221f646d8d130e152acb0397afa7397a52e63465828f41d81ac871bb9c82d81b5addfdc08a21bb615af410472341e9eb8c3da8c0d7c4624016d56cec00ba8f8748eefcd1b6d232b7a319426ed0ae7a9b195eb5d9ca202307fb5087eadd09a8071c19bca94ee56ddb28f1611f8f6c3748dd80860fdde10aef3e252903e906e658286a88f61a424a297ad34e6bb99686ad0c47c61f7bdf086d4ea910f200c1faaec643f79de49afdd9cb7fba2e5e98dfb0adb9047698118427de9b5e571c2861d123eb56bbb7f1b2cff7b52be692ccebf21e3f0579fc725a8f6be81952d29c52b632d8be9948b92fd21ab0ecb2f5628a64c2dfd8b95dabcc284c9acc803d1d9ec0d626d04947f81d6d4029427e7e746152119048b63fb866532bf8f1e9049224486d080c99e50bafc193c34244341020dcd1c0665d816df71376dcfd6aef3e10d6aaf7269c96e87a0c3f626cfaf4d6ae35bedcc3279577e7c3cfd635fa9bf9d5230b9d29531a1d9d2e8b0b71dcca9238318be0b1e037b2fc3fb8b40ae2093c28578c90c0a3a096360c69940b2408c2dbd401b45c38ab281ed110f243382376fbeb0647cb439867d18293858ff3a0ae6222a97e2a31117ea8a9fb69dec0125446b620d30a5bc3fa09abc15414cdd36a71ed6fd6513a2b8d3c51322645a73c59e1b5769a717f4f9ac42f5f269424f938d14a4c080a475e16e3db0e24b987cb70b444644672c0dafb16aeec94ee47cf035fdd7b1b31cedea901609f5f520f85af03618bb227f29960256bb91c46da8016b456cb8215ec2d74aee590b38b057332ea5b2c80763f762179916c403ba60a5d94a2a646cc518ac11e075132ec9dccfc664a8bf0c2f6e68f669d1bf1a05d9e94010c6fd685e15a923a82055b06f1265de8c9e892cb4541c35db14200aaa7e6a6b7cc0482cb15dc14eb5a6f90ee3d078dab4f749d7656edb92714df52912c5e11230817069c26c701382a2004346041a2c0008995826fc6547e9d5b5ae745a59f4986aef4f361fe8e38d81bacac83994682b72cf8d13d03048e16a4e4bf2c24f315580a7747ccce16ec39ee2fd1a827afa6daf11028afc1c00d0c5f3d22f67d92b229d60e85336b178b29a02e8a84368b55f7e0fe307a0985f278e13ea66454ea3ee07374f1b1b1b9ec5d00b174bf95f585ad53dad9d82fef7daaab736e8b4918a9d119fa72aa00c90d3b71840a938e94e793189e6d57337e8524086034926922bcf994cb1ca780a76dcb9709824a564c5bde807fddc4c8dc37fec735afe469bf347d7e8b7532673795f57a550e465b1f4d01f3187c684f456a4c0193112cee3e39f0cfa4155803a4b97be0e5a2b4d74e99dfa2f07b695c04682ea358113943c38f5b2b6be50e6db91e4f32ad790c6f5945d43e82d4e1f653bc13a92cd8411c34d5bcc7c8dcc72477ce28134caaf905e27267354b91b71080aae83c23ca18ee0a1f217051c72f0d0ea95b795a97db34207b734f599ac3da041c0465d98a2d3a768797feba64919e0c0b391cb34269ed7554c903d4e5c408cf2df6bd4e5e5f038f7792d59591e2b5497480e359f5257fa2ab6e42dcbe23fb9c4e13f46a56a499d084d5c8921ac00db36eff664d6fd33281670a9c8d52d504234206a193db09106f4276aabc58d6eb69d0f096584054709aac3149385db566bf2449ccffbb179ff467292bd610f2ebb67d15f05e8641aa7627eb6b13a641f47eb5f49017f1fb3d529740dedede44f3787aac826f7f832d52e57bef3d9fb2fd7a96fc440cc297dd12729e555ad9e989cb38638b4ad5d1c3c24d19dd826cebdb57b58b5ffb1e83a5ba94d3623e0d87b8d639bf1518bb0299d9dea23e453fbb9bea8ae7c2fec0e755ba9a49ba7080ab7f623522952fc227cdf19222bec718a39c0fc629f19801ebe66b072ca309b854383c2eb382d72be9d16eac104c36fc60ea6febdded6beb986505ce768bbc1878882cbbb45667f4dade0309ec023a10e96ea32fa609cdae4fdaae1e3b6fd5fc0f24229a33c1096e0b113ca7f53d0feb3c421524bdb199036299201c89fbcc1ae2ffcf122eea7a5b75aec8297a056557100ee7920199f3187fc0106cbc06cfbd6aaf3218849b6eb10617fc34dc65be0e9c95341a956443601c3d7dd29832642df8e93d80fbcb0b5d2bb2438c0000a3402e8a0d14561aad7636a586c7b91d342c94e9b516e3bc56586e5cd41612ee110;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h559621a749f9891afd7b945deb089c36411e248b30bef84f04192f59568947c1713186f22d0317c0daaee964911571b116464390315627dc1fe6c0e76954e192756bf6498ec5e12399d3a5a66ffa5101ae6cf0b018af61d7df5e2975a8a3665f84511c941c8b47434b999dda2ef7c3cd6ad291d0f3d96dd773323f45067c71331e54a0eebeee48a030f804aa872753343e8ad54642bd0e9596d8848fa58c4f11e348e0c9ae59c2e7379d7a2155f46d0a74ac7c76e65b112706513215a812b0bec92b1ab112c8b590b994d2a7fd701d0d37747d47d7687df6285c75e34f17f7f0cbff3e41b8bb27cd4c73f94fa0acb7a687035d6f027718a44717497856ebbb2844fa7f18794e6dca420c363b6b708e9caffc47ada89c67badf64f53b5b221cce2ac7922b153855308a4e1217a59ea1f3fdee58da2b19205d04307e7328c108bb2f6e89faa50a973c86c11a6a42eb32bc3502b5b43119ea4ed5d6493643fc6a2523d24efce60860d29823180e9b02ddf423897f4386eddb75f708557b32d3e3f943b08c28c9e38f49bce5d53b3c9e1d63ca7ed5bac2f01b6ad35066394352252987138277f8ba6282ca2ecb9ce909f8d2b65ae05f8ff45b0158ee060285c0d80fb454af69d4b1f2d4aa0711b84387b6d6740ab4ac1caa84b7fe0c2b1fdbdcb3c3eb98c3677aa933d28da813db18822b7c52cbf884ea23ac105dd63779b77affa7b27398d375288f000f8c22205a0ce0f8e6d106dedf95652064d783ae634a64e0cef955ada4c9eec5c1fd9382efef7d23e622d29f36090f1afb05b0a137968154c5a9247771978eac9423853ef985c106c87aa38c35603ed46917d256ef7a75bd69530f00dafd849ee9967496d9f23fc7a94a79bc2e61d148a16b3211823f1cf623e973f340be0d68e908594acefbb96c583ef4c0b6f976e7b47a6a88667e15887f130fa7d3d2e7ed2c23eb3ef8051ee90f0cfacb76442cc5b518a10e61e936720a4e02aba4f76f5d8e554ae9ccbe82791265e981e2063f76090becd5bac6e125c1aa35b19459c7041a22178bfef3c57cf29c55ac27c0644bc6a77fe62ded1b3e324f7eab64749bcc55661d38e16c9fe8c6aeccd4733311ae91d2a179209acc3ca38234f4d0a725d1ac2ee8b4c7180717a46c8a9836c92c80c3630d391ee4c590418043b2553187517a0188968239a6a06e33c07c6775747ae427ded19ced9c3a8b54e498c87b0bb20ee16d0857619cec550193f1d3b01b0d2900c9d57bdb9a358f9e592d5f2babf64196968e84c063414c4c23f1897a682293371dc0f38dc53873dc86c64e33a1a8f59ad850492a0eedf0f795a24cf6d256e0b5eb30360eadb0a0470428af5e01edb3fb530d32271274b842dc1c3706d758a785a6347215e3808d3ae592252714f913371683ca76fecd349b075fcee0acd04187179adff73c0ce6fcb36e5ad1b2b749ce3bbbb6f044eede88025e6612de9ab7bd5b9839b201042477574e7d6c93894580551b380b56bdcc89f229fc76342d2b533272f98e2b1d9bb15531aed945eda84a737f5864de6e060f05c5495268d15b8fe7308ce083fc4d60df79df74399b490736b28c63c0929f8ca4e86396e7ba877a9ca27a33018a525dfb2f7be4592082f7eb1aadc8303278b88bebc46b212820b795b7d61a720e807ff4f2dd318396ba9a0a8755e58eee5b7ddf4bb24f3e09b15d5b03235e41e6d8ceb75801dc38115e76cec0126f0c28289fa18ee42d1da807a1ee48ed7a54a21bbabc9b166da3be501492cc7dd593e22887ff5ece14dadfce5764a706c4fa08294c9b8dbaef7949b4cbce938a7bc520485c1164b44b08ef983606998c32e47139e5efb7d1b9a2bc86cd802ef8ba0f4006e456dd0e1afe35e842345eda8c2e6351a0b18371c4241b2249be915fc607d24deac5ec64486160b1e91a773098b39f10d13bb1e49ce338b8f4977217e07ebeeb0c84f65af1579132a8eee9e301484422dd13773b74c2e6b5f5d962c64b6288f9dea568c892288ce164fa3f5befba64802e6b3b33b8515ba315b6f2c67fa70f0093b06c197766d64181a23505302c1589ea279627e53e409bd18df756e7d09cc6f8039bc2cd311036ee16c4e48bd8064b4be8bf1802f0f478e292fbf73d304c5719040928245c3c6d4dfa979f3c2e6a57a68e00464988f84afa3f2fd1952ac18d3dc99514b0d6824ed540f8add1914f5c0cbf6ba63857aade3dd4359000a19e2eef843410a464d55758ae65e236034aefddda363d1b18f73d0a10987dda027c251d598c9d10b22f144a2ce0a505922ad1f50f53ad30ee92823bb541bcea6140bff11c48e51db4ae0c13287a73c262dd72ad261c8ffe5ea654e819979832ff7144aa2a6868ef3c0d8ffb2fe5938bd5def6b1f2d9fffdf0f0060e2ee5dd56faa9894224317cd06cd97a87a9cb24ec1ddbd96f19957964c685f9e9dc929edb491160b4f0febcfcb8f29e6cfbf66f8ca422e2b43212505eae269be88d0ea7a1b1f37fb6782b3945879e042d63fd557c567b10b26ee23a8ecc36128cad7e56a26540729fc92a90935f2d700b2265abefb8b6c9d5057a337ef49ff5bd263eb0f1e022c2f65858419aaad804e39fbe20573720bbc35e019eed2e20b9019112e515d3b37effe56d0ac94ab9ebae85b122ad22517c4c715ee71e962af1f95c7897f3da16327e04b45c78d71904f28a84e2365190443eabf00c3eef110b113e9f07c27b2f583bed9961e839a4c545a983dc7334186cdd0806822b89302f0539934f953ac8a9fc5fda20ca678ecedcd08b7ed88eebba7079f30331cd6924f64c50d885e30299621044cf08776f49688e464a1ecac1ab7511bbb4aee5e84c4db78ebdb722641b204d1aba663aafcc323816de390451;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h51bab2fe92d99a5b5386dad9b83bd2b692a0bfd32e31288013d6a64a9495f7f36552d0a9826112f794175c76df98509e5363d6a4a86516ee3d52e1a7b01844b3a5f374e67801d76d1ce333af97184c324632e06c6660b8e712ebfb320446780be95a6d444c146a9c580ba2cebea4ea3e807149171ac36ff30293c49ffc60c44281c221f6671ba6635a951bfb6f4f379e0816a7b792d3041049697a407c52de7df2012aee4ad5c4c87bead4d1bea45e6f6a3fdc7b5062f4c6e41fe3205c6b79e32481229041fb5ddcb62feddbc1e9c04d5ca38a1ff5689bce31875b54a93527bfb111500a4434a44d6a345086c95994926f626fc7077fdc2a328b78dd3585d0a1c1e5be7a338075779cdc3153ce75bafbdf415ad126c03b8eea8dadf2476959cc4aa3bac797dfcc61832a3bd1c19452683abd4f4a02195b406ed6115b54f22645b7f161b36c8b4cc3a9d044186aaf8524fdb7eb0bd3cb1f4c22a4b7eb28bf4a0cc1c0b2a40340a0f414a799aa651d04224dcb10502469de0a2ebe2437a06bdf676f0d03d24c8da9826899aa5e0cccb355ccb669e5c8ac6f2c03f7ff96c3ff1f2f6f6ea69f64bd8a49cbb2ca35b52dccf863bd7def85d81df66cc40ce67ab095065d0900237f9ebe3f1d2d1b6f243e45fc4de7024a28fb27323ddb9ddf3e483572c7c1143b18ce19351b5213b1184e95e5b268f424d1e691a42310e4785fca9b2187d8e38f020106af18cffd03908cec8b990231eecaefdb6f406e447c83341988c94dde947060d35e6537029dcf98755fb4f81a898dd084483fc91a9fbb60bebf058fde996d7826292e15b07b84fadde893866fad360c2cb8d10b39f8a8c230eb2d96d60c725d97b7d51c4ac68e379a20437801d1014720800080f7cc237eec273ce4604d2407e267265f273760994bc7e89f34eb6b215d832c5e1d1d576b6d2e7a89deb7ccf24ca11c4ee92d82854a0e855e3c52cdefdfb2527d14faa2fc0ae71c79e14c8a3cf107e17fea451a271b63e143d39c95288ec394a3a791d0f08e23d32cae31327645968721360691a9df87d25b1b06050a1170e10654fc68e3fd24d66552e30618a057efb1e01ca54f1b9bf58f3b347512c846fcdd6459d53cf263ff050bdb7a5c054a0473b4215924b6f52327236bef46508b7bd0564205deb337a0e74f4759769863d0f4f9d8ea92fbf434b9679df0020fe8645abd13d3b3433e650e09f9cf5f7746b09169787a1ada25fd367a021c222a42f7613191c8e575531241b92e882d78819fbe8707fbb894b7b08b448d3caa6c4407726290bd2db3069711faf6f4aae995b155226fb15c82a79c7f7f9be66151c41bc9f69b1e92ad17c4c505c5906834ceeeed99b39731dc38d816284341b06b304aff700bb2dda6eaf5704e79f176a27082e8c8abf3fe71372c916618ecbd00290d5bacf31e806363af60f7695bc125c61f140aa52b9343388a6b2de4d5fbab19b2aac2ec4add16a2385957fe510d0b59c6035da77772b596ff3b2e08457c6eed920deebabbd23f94f6798b1608a8b54de78d045bcfc3d9da1d60041f765a00cdb7bd2e83145cefc5ef7fc32ad9a2aed613e89e9dfbc2bf5b5bc3900591c3b9a535dd573d526fdf1ce71f6b69720934bd774f0646732558c0032083ba38360d08a060528d0def0eb8c2f8b223e883586227edefdb0c3fc91d4fd2248496e3349dd9df01ec26d04b386336c8c9228e833d3edfeb344438e1d9c5874efcf61076b748cd0c649866140e81dd978df6ade28ef84b2ee38f87bf9a1285073048e7c58aa8a2ca0f16a899ca83bf6f8eabe8a68e88ae8fbbd489e4a14e78b229888bc7e4cd8bc011d5db8b343956ed0d12108cce66f33d5ab098879da85866b01a1bc21c2e2f99af0f38dbd15fe97dd50dca438a9de8ea524804369e5d45de1473c1791fd30cd526628a74ec16505a218d99ec7dc7efcbff8cb2898c27fba1875edda859f98a3c4fb093892d110cb2f5e3ac6516708587fd51154703a4f58d199be17e806854ec8f6fc167ab782c10fd2781d6992bcc17eb31560ebcf9c62af08f6f0bffafa86f230c9acf43df7484c0be78587146c0f4295673d0da2beaaf61173bdcb27e506631d36d5744078f117f65d23284588f99836358d2617ac8ddeadac8c80f9fdf9fdaf9ccb2d3c0826e01a743cbd27ddc0567d6ac69141b91ae08e91a9c903c5407454488ee1fe99de30372a75bc9a158614cd14ea7e9ac7f689c800a22ef9996b08501df8a1f26e9167e108abb72877949d17a6db0ebd363e770a84af4cca0741af17d713d42504c8f2f5ad9275f8ef75b589e1708b22dd487e96cb6f515a554fff1fcd20966efccc39f221166654273de743307e1565a975f4a3cebb29829da844e81e875114c87db06eefb5043039bfc0766b1874274fe9ab2de6352f95784722a1d9f14c3b07eef92abaea2e4535c88138b387e3ce878311b07d341814804a71e79c425ee00ef0ad42ac7abd2593fc0e4e419c38199e9016db082cfc0ee0bdea78f6ced5874810b731692373d5ce181e0ee9358fbeb3f064e72316795c7516181c9e55da88a2b8b3e7bcd4cf6d50ea4c3b3296c6417f79291aca1ab422cc21bbcd52cc3f262546e85859774e6a57015680dc9530cf318a978cba087b070cbbda675d7656252e04d2c94a7a95c6224bba3a273406d63ddafea5a0564a95e22e7fd9dee318037cd1747a06e126d07d815e7b44a5474a4f9a89615ba4f20df04b7f94c07ca7ea325a749457468856c290b65ee4f7217809e8ce244521d601720927434fae984da1b6cbd77c53409f33f20227bc145fec11162b9de30d69e66c5d987e18fb50d7b294a57a0be4b0eaf05bc683a04ff0ea6dab31cd91d8425ce219b9e0ee47d31;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h7f9f5c321dc7cbb88bd3fe364649daa6400a795dd624ffea4bd760d3eddfb8b85eb30c63008ae5bc9acb418e7b1d2ff2e1669b7372c32357f81a233f9feb3780edcd37d876f7e23933a629dbf9da341844c3f052307c048b6835e21ecc73c4b34ac4df4948fb623b24316e6dfdd9960f7cb936f1b192abc88e8a104e4b42c90bc5e9c625ab2527ae54bd747112c0bf3b5f1399544399583845dcabd791e56306fa0dbc4e340f56fd4e08b7451d90f8636f56fd7c94395530177b0749d740ac13994b52e1ddd6b0934c3c8c0825f319e081bc79571be8d1237dde3d5286d061085545c6fdd2b16a121129ea40902ccc5d0aaddeef0ce402e66dd58072e7156f318f626747db5304808b5209da22ea9c1ebec8aabff4fd924f3e4f7882406b12350363e4cea40acf452304ebd2c8f748aceb0572d74b1015fe392e9bdef4a6ad66c9660708729c8ad578743b31627d635b1bf28d85885f74a3589de267b8a8a0f34a3c674520f4d5e920ad9b0bf5aab38d5326d6425b3fd0a383c7c476c852034496e7bc483b9350bc3e91e74236ede0c1d7d84143c6ff253ac09c753e508dfaddde650c74bdfa0cec4547a7f65cacb99126f06f09fac9dae8ecc02aa8c06c54e03ab8d61ba256aeb0cace4871a7c7933320f2d98db8739811f1b411dfba6c8b696327f89104a677b9158ef26df7a89389e354126aa92bab59ccfc954e68cf3c5dc93f2a040f220b5353189b5cfaec59a8c0ead34dbb4d01f81578e03bb22d4c0a7a27226f0f623504c6c4fa226fbd5a71ab5c49239639587c02eb7316387ba6217c15aa927c64acb211ef43735f9e3cb536cec780406f116a470b47e763da9fae395bf709991fca2b03e9e6b1360999bccbe10cb005d0063e3086ceb09132794932cfa55d00aa38c7ae6813095861e858fb296b792e213616207fd3b1e2705db6e54f51fcefb93b0deac36927cc27f52bf860ffcb6b73df6659029bcdd62085b71487b5568f042f423f2d992af0bf874a3f2b379e3dfe16d5ff559ee3e91b09038bbef090a7c5db840b5dace88b49028fe04b692a4f697898a0a6a00632bfad64aca7fc7c97d90d77dbdd6ede9803613492a6caf969c5bba453e0a4650b4b537fff8c9393a0942b44eae663f97c10e0e0a7b9bc3f6b95769b189982eec1106d807ca53a5366f75f95749a51f53b153ada762dc616c0674c15e3cc3ba15c704075ff81149c16a1b41ea7708bd14f5d3765eace72d44407facd9d67e068c990708de6e7e8d0e439fb9f79eb9bf8da07fe36d6cdd42fb1d8d60df3850670b6081686745a3885daf0a0c3072155813d4100c226031c2766d469e587b95ed8905ef4cf57391e520bfe8b50eb02f85d704a4be794dc881aff6e4795811c55b7e41a69fc7d385b8e2bda45fbe71c9acba13af6456f72063b52cc9471ec9aa47cf29cec90d16a9cea4204a03fca18228a651c1deeaeec572f3bbcfcccabbc27567f46313e6cbccd530f13188bda28d8e1e076508dac8069736561ab6b949457b2177d49bf903e14ee439e7b37eed0f3164295b3a95ae5df237651e829fb945703a4b61a0c019c260ed222a0cb309f4ab7ad3d262fd23c3e0282dfdebe4ae280608f7d8504bc4a4713217e29d39278944efb4dc33ea4b6cb1cbb85370f3d6b4773b61c904e041c5802c4fa17808a6ae07898be0f25aa9a6167d7c4a71f4e99f83bad734c645f406115072ab2de72e7886f8acdf9b517cff046cd852c39d17d4b3387243b485e48e842551882a4b0d188ec9b01a73d7a53e9d6536b1977a7abffa3aaaa5fff15276b32ecae22fddc2f677604f7445e1643c7a130a0dfb88fb18409c1b17b6bc902126d2f21220127ab53a932f944118e501a261da3405b1028d9f105ad9070471c9f0cd005a3b75020e39fe78d827b92eb8ce3972e391fa2b31fab85224dc40199d7071f95428995e8e8bf3f905a5353039d36d3efb5a54c20daf46ab0bb8ecd040c6328fff4451de8803a03f3d8c3a73aad85324f24733ce55540d72bd2f0d7da9b27092f2cc4d875eb7b80f58081b1ac3f90147d9e5e7c22ed899d91c191eefbc5e1962b78f15cf1b649933b0fcb735c8ddd11492142b6ac07abedd97abcfb09ee5d38f182266843bef2cd6279ed296c417ddf70d02a07568bafb72b8c516a8b594d0d75ede6b57df64aacef4b899f549ac1d844f5c6c0d3394ef5d19a1b073ac1c5d69e9e6add1cfd49d29084bd4b4e86900debb1d7b2298b7750707475cfc52b1786f1a7427746364443331d1e54e0bdb834d4ce4ac3ec3241e223c856aafb641916a9b9a56a069c4f42b1fad98bd006a0d1bb0b162bd88b0a00127f6527175647cb5c28098957624c103bd91fd1981ca139f73f563c9b685dec8ef2bbcd8cff1d660b86d8c10d28b77b22dd1ab57a12f40e54fda8f56d446dada7ffc9a3a0b66ba6f768fd2c20249c8c828ac0d81ef356c9c7a152b5ce42564ae4fbecce7be7931022cf080063015b933f5f832da6757ee3f86a1674a8b8749b46c5459c9200bc62bf0504fbce6f9e36511ceff1c2b72ee4c3f52c4346c41a3803c108cfb7de198b9358dec60634fb7ccd131207f9656fbb3e181ccbebbe258947cbf4bf1722c57c6d5d18e6fc9a59d0fac2bdc498df04404e711c523ce58d518101a368bd9a4272d8671d67fcf939d5562e58a2e338118175b9aa8cdc6ec00992550f7a50522b6d4e5b402da8464fcd8ea9f7d9ead9b699970aa737c6be260c0f9c5282ebb4f3e912f4b932f346a42eafa845a4471318b1c5ba1dc9b6e64cb455c096039ada4ebe53bde6e60607ffbaf53e4341f5c0b49b13e936e353bf10760ddd1162ef1bd0e047bc81fa79be1d05b0372dcc49b58f40fd36546ff6ed2de2c65231;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'he6c81340002ebbade210056291f529ef22358f78942da90a4bb50f9fa9eb41491cda61d3fcc8de2a9b9a3f07b125d7ed3b84a2be9286f0e6ba4e16828620edac05c186db7d9ab072491575012195fcfa0d27c72df9ddf293a8d3225a9647177b10f2985338f677aa537a0b736398732022d9e60b8f915aad7da75d9a17de6896271d76316710d3615bf9736e77be3aebafd0cb92a4020879acdebb703bab76b14c86644c1605d85cb183463f56b6cbe77e13a2f8c3a2b782cca6ce1d609efc609d128f2f59f9df647b9622e416fc3442cfeadb22891aeeef240d4b0550bd1ea94846a17c9fb051a6b099d655af7f0a30671f78976dd4d9aa8e8ea025a882febd14a161f03b559e6086eacf09d2c65739a6d2f6aebaea14fcce87527516c0b277564dfdbf4a264d41ba1d602fea6998ec3ceab1b0f51f253bd47efd331d5cbc36ccb53b99cec8e942d6f022642a6c859ea7b0f899b6dfdd951fa8204fe81c0ecab6d9d72bd44d4acccccf9ae544b938dfec7178fb322439437b179d266d6f45410e08688bb3556af890198862cbdcb0786ecff169bbc028ab2b6a43f7d5ab74ef37b8206d6047ec3317bad470189c209cb5644005ca62ea876d29e5c86079d971db69a6682979cd732505e3fde783fcaaa7d6ff00bb3efc960b97c9ec8fc32b8bf89af41967cbabaec4abb4de3744b1a18d37db221f2c03cd5b3e8c90e81e12d264e3021f7f48d39118824bfaa1368877bdc0a8290de0e650d05e00d8345fb172470e96b7ca741e0a463c55d75d02f02269bfdac8edbdddcc336a32915b6f6cb910fc05673b0278496b22e4cb4098aa34ef496bc895bf759b781f98c9ea0653f94ec43aa0ee6bd800e55d839ded52f575c46f11941fbac25ad023e201e4eae1b1011c021dccf30bebdc7f44680525ea98be93df7d0066854ca1af9d499957cfe4b767e66d58f127a812a6baacaf6e887d97ac44ca4d10530f812b2fa6541b6a7ced13e340374ff5e90ebf2a7a561ff0be567290f9477688864a459e3cdcb48489b5ef531e49e64ba32c4af250d3d24d8d3cd98af84e2524ca410de9cdcb35197e15342c5dbf49a68e100d7bbb1bc9eddd31ee5b1073593825c767117c8685c30ab555b93b0192b28c270c0c97ffd5128afeba7e554ce16688d625b7471002cb6a0268c18b49f61a7333d22cce472b88c8e1788e06e7a59c44247b58291d756ebe15f5961376a4f7d35ce8520f2e3494abbac1e30579bf2d7a63218fd04a3d238211eb5855c82e58c663a7dae0cfaf9326bbdc0b75f7e205b92c223a29e317006a13f3ce311e3e49450a24cf69716b5d1cd5dd20237dc817ff9745310434cc2a331609445c38ee6e0b8d35d53085f3fa85f469b9d52ba764d553a2f539bfcb308b2a8966a39d45d271a6cbbf682e7b1b261159b88649b54dc6601389a396417150dc36220c6b32d75175bcd92e7010731ee523ef67f54b328e9fc755754f8f638d8ae09c78ecf2bea2a62b647a32d7c75ea084434ea02688b1829596711a1667980d92934ad011a390c96de3aa0f4c67dc9ef3d5f3d62c207594aa9778d7f61cfd7525f71d1d46fc67a37778fa1ad0cd4625be3127cfefc331c55b05d46e4c843dcd270272eead06ccd90dc9373723ddd2a52f971148dc90347b348cbc6ace817ecc488d7cbd6bcf4567bce3b7bb79ad69a5ff504bc858352ff584896203f5eb946ab6ee45c5c0355b705fcdc93b2135d49fc416282a4f1af6b1d2ce9b5018e7e7e16a9933c4a1ec03ed3ee67cc1ef8e06e3a6ddf136602085a5955ecdd6a1de57fd2999d20302eccf799095784801a297fc284f63a31c166c5c1ef22fac38813c45044ad7e9832028cac66980cedd320196b103d0d35a4e66a8304de18a8dbabca25dcadc860ea5dec3e40123ea01a533e5b889cc2200bf259c2b075055706697ab5d5374ff7cf6cf822442bad7d97fcae2ba6fdba0daf06daf2632057849ba55f79aa5f13517e9a4eade23421f301cbf3eb3840646c470054f09400a57cfb019e8d99526ea8525edcf301a9f631fbd1b4a771a4f393fde1eb3356b7ee5af559b74836300559e4d65089281cc7febfbf010c7627ab3f3764bc19c6c77268d11ae9bc11465567c75c537ad81d9c5a28150c2a6d6f708ab618eba94317f644eac9d51a72dd6f571b3551a72845a02aee7113b588ec489b79eefadf81fe548805a8121d40bed3aa4b763854a60a1ecd787039b01e4cf592a82a65236e198e8fcbb57fc6424dd29a890a9ce7acea3d5f4bce3021af9f78b50ea76b604ac513a48030caad0d9e88e9d175c519e23d9ce0cf44c2c25232a6bd05e86639331948a0fedd1c978b844ba650f9cb05ebeed3ae1f8cc6cf21a98e78e2e74b71dd0ee26e161023bb4140782a50be3a4b959bfe2e9e6dd934d175a0e14cd3b6b45fb7ddd5a08308083943de17e8b1341b75b73c72bfff35114103a29c9532a26fbe2755c7fbf6bd68b9e1d9af88b3c9806eeacc6705b4415e64edd0d1e84dc8b3914731ec785334b74fc736eb61d07c7e20caabbd2d9e7b9e0fe355390c7b0859bc34963280dd60c0d8d0999067a49e3494a5db61193011f042e9ab92f3ad838b6d3afa444fa1ac1366a8533bc36276e9073120bf17004becad975071783a8d059b6f4a053d6b9ee5f1bfa88c4b4d13da8dfa0e99495ca4f88280b9e8c98702ac4e651cfa3156cc9e4a84c14a663354cffa31fb0b3082bdc12097dcd56a8968ef01b1317bfef7a4847dcfa53278a4d4b30c06208b7569f8208a08f12e0a9a04914f7a04596ffbd713becbb4df5c7acf868e0b08c7736cd2aa68d27c4a802e43840bb620314323a5f746010c7938648a5b14dac928230fddc4dddd952d5f7f0ea82624f24105be5;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h3b711af34959294758b7da915660988fb2b33e26487f07159bca218065eb83780552b8d705ab44572b6293335fc2710ddb9dfb497063283d721c7ba35a002ae6db48fa26d825be6b1c096deacf4da2af7a87c3ca3042e693a7b6962df057aaa8d26e3c1a9c7cd3eb7f10ef794d2cd5e34b985f810d176be5ab3b5e74ddb933267ccf5d79b4d69a7e1d673c03b5da174b49703798532873fc2ae8e2db229e2c786177da32e47cdc5cecb1f95973cdb6c72f99945ef05f8c0a18700366bcca73040b659b262ba88391828cb90b14db918a4d106036265a802d5ea885c63175301237f4701358027e06be5439e584f3e38a0a5d614cf65ff2a12b7d472989fcc98d9b0adcdd1ef4ea2c457cb6213a28980ad9d25a17ae2f985ea7695f8a1194bcf9678d840ffd3f41d3699cb75f3a03b8de0d6e6b9e1235eb8d13c6256987289a0b1033a46d1f4376136d9e9f3f23b16cff9dfcc33facceeb5464266c2e23268871c79b1498ecd53c5beb0a52e757cad2f41bd6d1256470db6cbe71329600e71c809757fced89216d352f88bc2da7feb1a39245c8346cc48d03372980df9cdd4c8b29e3ab414569b800631b6dda0b668fdd23cb893feac143f5b03857a866515351c6928c1d01aa24ca9111631546ac0acf51a94a87e07c0ed44f700ffc8e18a933c84cae184e3bbd18077c2a2f38881d721b3e06031088c0ba4df87350b12ceb330e1e5ec6ef51c51218e234a5ce128d13d7ab542a220e0e66ed3169c26d8f63c87720526c64917a11e604dffebac9d122d5e6ce04798636dcdabee180d0d5620f62d95f8949e8aae63517e08b33df23d1474df404fb1d24c22089130efb05a534dd6e7491504fa3d96cb2ac8f2706f1883cb88177f13b06ad4d909ef060d7bec094793307369a5690fd04c1bb4e2fb285aac8024fce8e228a87e3cb1bff844f64e614cbac1637f8a6c8002c2b7cc6af34b540eb4c6891dc56d47918090e2a8d1fc1162108df685867d4ea18f4cedc6a18479b7534c2d2303604f6fff485775d31ccf30276bccf2941b3b388b88f697d6f950c2e4fc4d0b723ae6c0046108b63dd9bcb4dd655b180e2b0d9556a195e92bc33e1f9a37f3d4cf4ef76df76bcab62a62e1831211b31277ee5bc4803950b9ce3acafeab46dff7f7cd754c5b447a0f21edb935f07492a69e42070dc275c18d29e3114e0b3c581dd7f880a82ad596ea3752d82124f4ef1bc1efcaa5234b37c23f78a710eadef56194a29fbbe492c2a5d8c49115ca7eef63cd97555f995c0a7fbc7d00c9665b55f053227fd0e3e6d3ed19bc64696be6d2bbf4b9c473536713b2009a00b008b45c0c04445156edfbdc2886d3def79662564ab8ad6d70a503928ba51061a5d87e13463bf451c03931c20880eec358d13426298b4e70840a2c43fe760aa77ec527332f2cbe279edbd349a766d116647c8da35aba46237e7540f3fbb29dfbb251497829f5f63e319c1a70b53c7c69dda51608f89869f7b4332793efb8e1a765e2b8f5a44223d343034a2fa8faa3fc325f4ca3173386f0d9d668e43a462890fc7bd8a46ae94374510c646e2a6b1f841c34a04757f5d8af3291948cbfdcda837fa93aff7601e04be3e5349b50ff44839e56b273cc9a04cab3d7423240c20feb0e4499ed1b8812c716d01d4bd4daf851bd906b2e1611af54e68ebc1a4629394e3be3f4b77ecde1d893c18fab17a48e7cd434666fb8b4179fd9b96ddf60a5b7c286299b7952c7c4432e4b178d429a977de948e561933d4e679e2d695164c6025c7f78a175e6b0c38047d3aa155a82f5052e852ead05b83dcb3fd4d1a83fa364145b550ca9081a396ceb8682cff2e4e9024eb736e260cf9150ef5695b1372a63da94a012f1f3ba51bdd37072fb2c5fbe32792d6184fd62f8f8440a7922e16beb23a24a1a1b03da39f97cdee8a456871112af3a73dee611a18e475a5cc520a861ccce97bd21eeb51bc752ba8302e1237bc7bcfece284526c0debc10476060aa3b4a05527c01c02bce36e6f1d398b7c959e6190c122d35cd4df5c202b3865651539754bdde84a4a2da3ccb0ba0d5707c52b0f8622ab93c2eaafea4f9c2219ceaa18e824c6820372c79a46ff70582474f783d49cb4396e02e9d78089b20924d9c1a1513e29d047399bf2aae3ac800b74a3d782b236ee91fa4712cf0b53bab903943b83d551fa2481e4acadf1a609f54b71076903344f7b31dad278e62d2eadb42b014ea9f8de3a1cc61892863a213a4f81222002cab9bbda1479155835ab43815cb18ab0c1a63a25545fd1a928a1b53b4cc8b7de22eb18daebb6613035c4c2a04b602b02dec3fcd21cdc39bc748f7394b501bedf2ad404ef4683b328cf90eee0970df6ce4efb95d084e8e6840775037574f43563f1fa2743c7361df1799fbfa0b65525154b64b940b607313e38aadee97122285bbe1c3bc1e31c104275dbe65987f8b238f47d67e9670572930355642c687dc42ee51f817272e91d4db53b3d2d74ed1c18353e4f2ac6f3a87baf3703b560ab45e515e7ae03e2a2b6ba3a3a302ad9e8c7d49ae6131ca1318a65ab158acb690d867d54f5ee9f22843ff9490d9720e7ce742bf0739bfad0eeb3276386cac1ab2c337226b65ad1bfd9de1cce91cf2f884b3953fe2ae55c97243b57259bda2b4d05f22bf76c97a4a4426fc2479c069db2cd5d110e2e42e178e4e9e4ba2eb1ad0accb7af8d372bbd49093e70256d88b7eaea442dc0ff73a25c4bb553c3defdc9f8dd18aa352f40890c6905c0df8ad2360376d22157202925a52ccb1f17fd597830262f3a630e9a5a703491a7ab1bff579650cf6ec0c6a6b35ade56826a08ef97269f4261c140129cd318e34ff09b46104fd990b17db82d4062a2cbeb28eef94250;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h32aa0a70c7538ddb2bcd8943c2a5e2e168cf216adde885c0311621b1e2c58b871e8fd6b9c7b87b66f849a4b63743349aca909fa226f15de0ae78f67ca6fa71b702ec7d845e652cac5e43a2966f7f53a4459b19da2acaa4128f0fe6e87a0d43f66e0553a079b8364e54d4924aeb9a084895f2aef763ee05361d5714301286f1efa50e17bf7141717f1da87797bdc34c3a169f05d3381978a8b4899cb86b5d9a68d878ac4312d78872464a26245d1956f4b9a2490ece973d50c77eca5a10b518a2387d1905c6fcbb73aeb3d1476c184d32e7f8914691532dcb1c1578528b20a12288b3dba8e457d40d50ed57a024e597561e038ba972c1ecc14e065ff67c4a32c9a8a2ff9d92510b9dd6c3629225495997fc51faea6e17d85ecd21328c43bc2a47b3b8fbf00e27040de8bb2f590fde3d99c960c1e8346f899d2a5ea9d0f6ee98f9b63adb404a0defadccdf124ee9fa93e109e7d05328742fc3e8311e9a4be8ddf7eeb4c6bfcd8443e236bdaa98186eedc0606b062be258a0ef29fe852e154ed6cc7a2ec3fbdf798d3cde16401df273488179f19e34c26a5d85813b641084e1108530a8eea05fc4c6e52922ee34a81a94d87907d6969372754bf07933e31df7f662901f6723b25d2dfa458ab5f6aa20270854af91d6b12417a375b3d0ac62b21116de559b26b11e1931d18ac1cfd9060b682236bb546b1f58b400d183b5f3cc811f4edbf833a57c70dd22eff7545b6cf74f9d4be8a2443c90660387f2e299810a59e74f75397d9831da930dc55dd1137c5fde7e6f98561ecde8e35254b38f477702f8cfa48458ee0fccca6874a7c78dcda1a07b2a1c29c56eb08af69ea5f7bd5d903ca055eac5b278ebbcf5692d2a1a549d01ddce22b07b1a236ad77901387d98fd3de2a3ddd8f2792439c821382ed813a5d97908af7b9706f6a57151a005e935f4bef2ee1966bd5860ff51e1f373d1fce82a6c6ddd670271e3576d060721b37b8cb3b671611ad73103e6c983cf6d3f3cfafa29594080eaf7be215ffd8c1c527c5b6df6b6d086433c3b10747bf52a02d80b7be7c50c60fe64bcb4210794acd9fa25e92c7686c92ae93c17c52fe22b90bb3993daf30cea4e81c4df96fa8277db83f29e1f9a1aea6dea71610de55a1f368338199df941f0dd40cfc1cd4151ccee6ef8d42d6d6158dcbdb4050723df901568160eb2d5ec2136dd90f50a0e28c60dda3d39cfb90230f101b7612ad02406d8eafb45d46c21c8647d67755755b4e7be0709aa27b3adcf573bf0b2b992a4c5dd63fea940227d489d5642205f354664d420cd2e2a38cba96664d2e80c57d96c35cc076924cd92b7820cc84981d9e1d58f24d450b11dd8c3c9093fd12dff4713d69514b8c72ab8a1cec395350b5e93bad8ef4dea9b1bc47cedcfb936ab4aed256b1cf53e1246788867ebb49b481def8c0a333fbb137d88ae9ced75c9750b44042fe8e921e81781cf898d40edbff422a9d7ad661d3daff2d8e5f5c156c0394d90a8afa8abcde3c79615435611eeeeacb33358bb8ab6603c11148cac055d4d202da23fb88985b3de379b58417c15fc631e34ecc858a58eb10f5e75be30683a6d9c983313d4a4e1330158c7d0d2143cbfbe518468571b9cf5a904d571d07ee67d4556e2e27e5ca7dd224ef31ef0ca16698e4054403a02a84cd49f6743622502e0e65181ae890782f3c79539fef4e249a6d214001fe2e41e2539443cd986f3e235842b976aa5b53a7c68a9c7c10ee4d428f79c0663d48c9701d4a59fd23ea5d0b0bd487d9c3172bb19c04d56fe5315d60ee0a447aee9c0e3d01b742c836c715a4290a4b929227b6b4e6ab2544cf80d1e49eeadfd3eb3f592679dfe28dab846cc636964a144730d0b891f3886e55aa7c26f411a7ed7bbc630f212c0645c5a2e26521c17b3fa9a3ef86854efdb575c4d9568fb05785cbeb4883098dca344921155055c14bd5f8f0646dd8858edec1bbc1ccf7dcc0c79d651d80430e1cef4cd867e5ec53f018740207f44f29d5d06f00d4d77928b2de06d4331bdd108c801c77d4c9fa46b8cd3ac7cd6e9ed7a044f66811cade07fd1e11477dacc54275e80af3529ddaf933302b661790a8bf0d400cbad687d8a615e7fbc89ae104648cd3edc24d2a07ccda92d0fbcd62abdfce1142ddcd4fe5fc152d3af7c3f424b94a5c30d75db458466ee404bbd9e34bfa294a0957a25de3bfefa1cd46a9270f9ac1ca1aeeead3eaf98d441fe744596230f7cc9f7f972c2ccbe98fbb5b8ef72b92c251108ba8cffeef9f1c575b4351e4e63fe5e9c578c1ea62c19a7cf58fe66c98b26425e921b7834cb36d1e437b8e63dd449f4fe8ff63035e49050f0df8000373c5e59f917e5de3d3157f584c4b47c7c14850c2bbfbac4bdb3b76b787ef25bf0635e3f9a3d7c07139b8ee5fe3a91aa9bc3365c307e0f43c69b7324c4dd101dc0f8a2a116bf7bc148f4ca43ee8d99d4aed5668889303304bb4125e061b0167a68989b8c33a30a5c996e8b075112f7372ad92cac9e4f9b6695a328a9373de8002c5c4ccab3f192ab42f56d61cb6978340cdd4df277d07f2a9fdb4ff87688b8d4fd912fe20f6d6104380be88688f9248c03084fae8cd72e06dd7bbc4b82caac9ac0d59c90924f2f4fb5397ee9e0ced6a959dc11829d3847c00b582fa93f0da734b5106352c2b2e4caa2cd53b264d56d0c4caffb8006057357f98101627946237a32daf54bb1ea29988958d837ab834a7abee71dd93382c5cc885bc3170fbc575b22feeb8c8888e89b2c8c972e8e0d39cdbb87b935747e690d7ff44929f58d56741e535b3d007d4764388fb7f817a12f11eed694e0b0b2a0cd96cf9eb5ba1e7474bcddb8808215ed36357fac88eebfa8403aa580299b3377b2975b411c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h1eff02244c0d00c75557ec3d941dc4e1d4181b3875784d39d39adeb5b7ae07639c2a7c1697fd3a27638a0a4d78356cb1fad5d1e42f5a2c8a0ec90c139ee81376a006baafe33df19b7076b9f3c114db4c60de4e69039eedddc4e4cb20dbfa9214d0734213c2f16b327dbd81773ce075f36da9d18ac6ab172dfe3442fed64381e81ca242549b6998e377448e55b8d2a38ee1375cf8ed4f8d79d1d1ce7c0dd1b37269b5b27b558096bcab26eef479b0489121bb4800e45f305dc10c6fb37b685de20d54d299e7db923cbdfac68f51346b78eef2b8d88b0af4223b27a498cd06ca819a9f6e00da04bdb58338e2446d4d21e1db99917f59c8de3464d05c0d4ea4c288873464f349563ded6b482a31a300cd1eaa7247056fc1de0d90e001ccbedcd796c6e5e7d75a6a2299348529d9be834307c850983cf13323ed33da50553919b9142efb0c61f22a61b730ab806860cbeb047f5f45d163e5541401a479cfd919b27e44824d57014d668ebfdc26f4e2a95a6460b06f510a22bc4b7fd402e879fc372c7dbfe6b9c632ceb871099a711ff2e3b9265e135fa7738b21f0dddea6f632dd1ceb7ce8c2771f9447ac0826d244c476c9ed257bab6fc16dd876e1e32ea1a9d3d750dcfb4e4f9f7a1e82cb92040b6e6eb661b6d9b6697f29ece040acf1bec8569fba984c5fb138600bcafd8e08b9df367b3d6de8ec708581f652d569ed38c5994ccfa8079d8bc012a70779b39935e3a89179bafa5b18417cb642d23bb121a043de06cb7c1a393e6b3fdfedab6b594de647f9e5b8a783dba28aaf621e25b868878dfba751fdc562c3b528498973db2df73fdc8e3d95f85305721710d44b26fdbc0d99d849f3e6f2d0c3d3dac273f847cc7334d60e73dd6eba2a73fb17048013f4244bf89e298a21817e198924095be6a6d861979e6464e04517986634636093ee044fb96f22c5aaa5eb2f0dea1d4bdc73cac2f2f63b0960c48e26e8652a8d55842221b3e035cf707220f563aa57fad0b8ef48ed2ac63b73c2b081d1ea4b2e9421854e163760c451871ca08a78ad32af63a014512be6563245a780f30109bf9c3b1054504de1ad34fec6da81a26fbee93e763ad24daff287d492d2d66202f46a99953b2586682569a66107cb1d2af2aed4c08c75da2a8f28bdb54f196fadc2afe367b8a52a44f88f5f0bc01735eaf85516b0b76baaa27d5ab3b64dadb70256274aab6b7a0012dbc8454b7eb375cc2966586a250b1d34bbfcfc1b208d800dd48e9ef2c858681a756c8b0b1b0ac7604f7b2f2a50dbf112446acbce04fcf6d1abc15d8377609cb5ffc5deea734aa29737aeade0c5b0c817a939cfeb7276d401de3db18b8129d3c4a8c9a2efed47aa01db3ca4d412d83b51f73b80bee2007475c9421a521a99c9ff48432a989cef90b26bf7894a0347afdd786329fa89ec2edeec3410f0f2c674d364f54cb40e0d3084de0ccf4dc07c730f78ac9368c12879d5a70a1315c808301a17ab85909bc0e4c1c49a0a123413879e149ba9d096c8b57817f7342b779299d7db30a678df616994a7fd4328fdbbcf77c0733a85881f059867ab8c8e80c1bf43b2ef2c7f7d5ab2fa0940c647676cae9dbf430ab182209a938db19c3583d1078c8acde19607977540b12301d464d24d68f9a65691464a2ef6bc80af2ef3ea7d10fd75d55c67dfad5764ee8d10d1b466ce6cf320657c03c93c6175c5ad0173afb84e0e19f54fce7d21fb436d2e805f53370fcdbb7878740a1a873661a78c4321e14cbb5241418dfc6668a1acee366a733a086a3c4f67743abbac8d1fc4fcf37839a05687b8cbec5dbcce2df43a6957e54e765b17df1583d94e1fa37c40e634b89c1cfd847ba83c8060c8017937a10a3b3b9f9e1e97ba46f45a4fd1966aee799449bb38ca8d0703f93fd8847150102736f47fca8f13025bd08617681d55a3d12882842e83ad6f2557aca70a80695964087eab31356536ae2a3ff16671dffe5e60fc6dc2c074c4b2552439e9750d3c3fc61688d27e1129de4912f7971a1f89d0b030d8461a6e9a8dbf634bb8d326577c2652b57fcc9a35a3616b56e86c6466bfee1dfc8975b128192069c818387b44e7129dc6d8ccf316847e1fb788b6ceb88063aebf83e42a705fcbe42a1fe01164ccbb2294ad58ee0652b71bd9fdde8b878fca8295c13ebcf4d381c70677b9a68c1e2ba80156bf89331297c80001f89964d8983dbb311006d1388401e5558a9df59f96086b047e8e5a0c317ac05ab579fa79a862f6d9dc33abd51abf8b9d54a580db8fdb6cfc397b8d82bbe7b031eef105e6cc9819d7d251bd48c30cfae6d5afb92702bf6774ccf7b60b93ee88b1416a0bdd16e49342240e06040227c15a3d47349848266818c36e20d7c187b329d199b3918b9d3bb94ef38c39461c6275786e86d0404ca1be51b890d4851f925d2e4d55c28f6ae59be340aac461bdd1a424fbb86aa0f05fbf1a6b78476cdb53c25d1e1066e69a68ac6051a96aa4aaa11cde64d62fb502747ae4cf3ce93b86ab173ac8ed6c7f5eac6b635d042d63e1a8ecdfa95642440b52639fb8eed3a68f3cbd8662c2499bea0862ccaa56555a4aa057d1c2c3fab7503373b9de03f29d7b5e6083ace4f4782f2e20978a287424b41ae922e9ba97cbe3e8613efbb808db9cec5b53625828bfa2eb3fcdb5302bcf9080a50dbd8bf1f8efc879a9a90ec757edf816089d1d8d8ad33e1eb8020fd8d961a6062fc5fca0be03a8f2b7a016fd9c1a9fa653905c38cfcfd79f5239dd5d2ab3897ba9136e70b2d9520e553152044515ffc661afad3a83d7e1dc7af03c8cc08e3d5b3eea164df2a5b3c323a7d8659dae4fccd6fea16f2dc7f64c7ab3d772e029bbc0e588213e2fe9c46aac2d0c4a1a79e857004e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'hed31ef4773186c38984ddbb8416a8eadc1e8f4f7b6f43e6226912046982063145d1dcd317efc707e8a05df314875491e70263bf1a73a33d05134eb09cc94837fd307a98d5b6bfdbd72cd1be5503e3c04beb76c3b8664c0d710e128db3b24f3cfe028c67d510420473b356cece45b91ffd770abc0dd71dae609a89d0be859d266a7ec67ad20e4b1ddb458d0438cd1ecb24f822e8a1c1b5e83cb665af095cee5a05f622dff35d98aa2b01702df27f43aff1f5be597ca64d685786f908751bd4a114725a0f1598573b73a7a774aa1abf037c184cece0e8afac3c7d18cb9c654b4b2194c24e3e8e9508eede196dc339eef0bde0da2cf059eea6d86fe4ce47ac4901a3a5ffd3add702e9825474814625190c0055d61a3ae03d6084c611ca4d1b61aba2687053077c5b9a639c601846ffd2ce71bd4117a31d26da040dc65adf2221183b9260b4688a372908149020388ed1cb1805941c251c22e9e28b7bfc2ca675a15f4ecb8690f1f0e73fd9debb6fcb358b8201a6578976437f4d4d79839d4db6af1072000cd96e9f69b623c3f36471aebf8d6068aa8b7ecfd310aa3969ecf6f6c4467b9db6d45eed2e24d883fed1a8cb7bebc24d4123dc45407e6f9ad3fddb2e73847d19f60e3981aea820beb0d61d863f41345df6d60a5db84a66bc815cbb691ebc6976504c32940a52ad14b48129eff83c219eb5de6caa3deb0345bfd3946691a9507ef73e3c7c013b0b63feb723cb8ec2b3538d7a82e7c7161369be3bcf2ee3176f84b51cdff2b593216dbf104fe736dab39b925ad639c2f86ebae0fdb4e257c45b6481068bd96f5f42a97a19de8b9dcdbfc83afb8e4ef4f7ed41e8f6b05f2b481e339dbbb2bcc8edc657ae9c11ae586fb8a159e72e487dae1190761cf4047a67c4730c3df19c3e3c4889ffc72a21df44e1d03032bfc3f9f9eed4a80bfb809ce778a031cc02ebfdc11fea04ed1ebc57b0e6376ec826e74da2c44c4b2a3d436dc298d6b2c9af366d7aa92f70bba7a032f0d1385f052ec5010cbd4739fbb08b39f6e7eee7fc9d8807bbd60735e2bd79c2f6fff8608167ded354550946fc33916d10f3d6566047887ebb4e15bee0f4134b487e696c0e281a9154462bf4800b0353e575e2b0a87db880774cf88df52aa132402e7818c8bb8d2d19d42a6accf8419261de2a78b6960f04085355e21ad17a3b0c359ff40065ad1eb53cea2aa35ba6738bedd7c010168587a9e6f61b515188641a6b1af7addac8d196eff1a14799611c6b35f6e0fd0ce1ef185c3a318b199f7ef31441978a99a0978bf8c8ce14c5023424c57daf5bc9e32e8fbec7bb71ba25be7b104c31f547dc5930bea4e9bd917c226ee5eac8fce48a784360ef3bbdb73413c793c43d66fd3ee10418b1582a97a812b458aafd10c06a5f154f8a9a2c64d6e6fe0bb4473386d6fa78b50e4850407a01c847de4e67b07774fc886d3266967c6f8959f8d88498bc8f441666aa027968d7fa01f3931b7de6d05d82432e933b31fcc4ff32271c3c868aa0ef5ec89d4b078268920f2ace55232a2bb239f07aab1b7a00934858b96c10fcf6a79bbf172879eb23ec186810c3588494ef04405352cef0fc418a8a24a16304741cbb99e5359d1bc0e7db54b0dc9d9e36039c04e8a9a160aeea78c16a730a8e57cc4ca9bcc1df9b4881fa862ad38a5ccc6b4e04c5c9f0620141a69084d6c179c286a334f4a602c90d74783403515066f3664f50e81caf8a74a085581305e1f7c782f0a843658b7e5238fcbeb5212e426abc29aa570ed6abb447c9a658c92eeacaeee223b13d606aeffd1612cc61dd8995f383af632ee8b4be1a8a6e48ee86a3c83cd22594ce4772705ed4ca3142ddbc80acfe6153fc8f24c60b0e9ed4a19d72634c31cf86a7099feaabb740138b90d14df4db7f5286b9c50c7c6c71c223cef063eddfe54c4973781b8389b90dc28b85e089b2c03f2a06a7eb0859b376a58629cc3185faf149065d409723dbca4825ead41c3cca9c12c6e7e4bf0281ce7fc6737aa575fd85ead6c50fd5bd1a8cf31f6519c56b1e97050a488749c1180477c554714f21e637759c0f0c1cad657bee3368bc387c03f05635737111715688793b7fee33599a64f3c8b9596a9a93b816991a1b929f05ebf978200c1de0fd1bd6d67a7c52b383776467bb5c7b92f5e69c6c49b52d28b39fa7b69a9351f1409c12a2504f7b88ca1ebbe944d6c758ed6850b457c192fa1678f60eb29d9522a311477c71c472551aa66ca8659c0a323a2540405c84aede662a0e330ba7c15f48220e1cf62da3d93ec0769347cb4ca9a57cab799a0427585bc7ed8ace412f1f736bd7d2b2ce7d8af25d3885b4572fa96c128faae94ff41256ae689b915705bdd52ed5436381816fc93ca70530520c54dfb55429fd98a14cb1238351b139e98b6e204d5dca8b7a12658380a5875172eca5ea3426b35e6b9ec4aa7861468684f73b85fc5aa5f12b792cefe7b632242506f71b414d558ae9a21dd9e7846f6261b8472b0d69b9a5ed0d15833dce6d60ceb71136971bb42ec40a142f5ae0216107b899353b014af40fa5c1f0a8d237cc64b983de1321f7083a295c7f159ccf7b7493d9a48d61f8bbef3df2918957609c5a528b9c9948d9e0232e632362b3911fc87393d5c7c6b1bce2168ea42fd7f2268fffae9ea3abfa2d20f4ded38ece87a39ae92af70ae2ddc852e800151e7d4c40826a6183650460ad3b6e11b876672e1dc8bc28aa8828937a8c2825105c8056ae798db0e04a493025b4648e08432606574ae8c06a00f6ba404b08769f0976fd85a009e1365af8317004a77f37b5f41fda53c3e8a8c4e1f2cf4f5899e709b5959709b13cd830a59732d2476fd3f745f23beb489ac4fec64073ec64210976200d2;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h93e4ba8941553389894639b63deeb86bec2d005550fdc5d450a92cd6d00afc370615a7f78fdf5a41a45ce8a9d4739cc4f0c58e67bdceaae8f96864f0c0099e28de75f86c224371589d712f27c271283d095a79bfb2ba97a419d41076ede64e58d94860b185148d1c13772b2b65d057c82c2203eed58bf2773bfbd556e598f3b5439bf0e352ef9c310822ebdbc196a4ca332a04b2a87b077c856c85c533f268007b96239804338e9adfbd4c8122d27dfe26e33088e0d257751e0f24a57ca80c8c3de46b42b1e260010976ad7f4814bf3692fc1aa0dcd16888464fb7222c20aed622eeb514e441dfecfc3891fc80d3d166abc8e5141e5d2f4447feaace2061eaf922ae2c415503f5daad2c03f1736a3f13b06ad3e18e67fb898933b10f5b63ec0e1aff051bb28d4ad93fb465279ce25b77c36a4ac76cc5696a712e0c21cf49d46e4c15a6c305fe3a8e518b9febfe8d2e4cac373b5f72cf31a23d8f31933c3fc6ec42c5fb27707e3935bc060250a0eaf776c76f9047ba858d224248b17c3c3345332ea8c22a6192e71cb392fe0aa8319d3280e1f60d7ab81abf988d143441c8c1ffba1aec98d461779b6b0d3d1b681134d6e6c1e4e6d871e0b4fd624cbe985edd1cd2c090cb182178b4181774b0a7f87c60d028b76bf0c03240aa076e9628eb566e682cbe9e5cb3448bc0d1d27f1b5f32798b0b23ff272e2f8a2360c6fce586683bf5f0ddb979d68de72a53600bd19724382dc63671c402dd7d928b5ef1390e5fd5c784741ab90a9615e8e8d281906ac4461bedbd7f05a824a9acc6a682d37a2bd5c996cae5421f07dd5762a674dfde207f6c0933bee4f8b2c63057a03a0f4b3a5a9cd4a0b8fae5f620a6173ee4e552d037aeaaffa1af936ae6272b0b853d251d8c99464976e634a80e23143474a9c71f628ad18e9c49c963eaa4c77530e7b4b53cef2d6c1b1a64f14288ac9a11bb8247969e98f181e67dfca2bc21f6140c87f56f8f488b843988ad3ac084d9f982b5c13eca4ca4433a4fb883672b3518884b3110eaf51f43f0a459acd3d6af5b1c69ebfe8856bce6dd008b6b7e3b96b37638c218cf5e6c90a932d2053aa0ee93ec0760768abfa8e42dca4a7878e67666a1eba011e66d9fac1ba224e3bf5e83b9d6e2c4f8d637094d68c0b958cdecf699fb259e28847a2e5f82f6327faaefa429e725bb38fd00edcbf8564ac1c74777d2531ca37bb3581aa25ce32b7e71aef5af33793fda8abbb4ef1059b8fbac42511491b9d3a66686cdc34482c04fffea42bc1e0f86ba77394338972e092f4323b7def5647749a7ec70189493484f024160335466d72543ed794e46af72055c39ea68dc805888b4ad496bc8ad04e56dcfe16fdbdc6bb75e282d27b99b1acd59cf1f6ad467e3da344309a28402aa8ee12d7ad7659db29abec4822e0de5cb7155ecde540e943df9aabf155ad1277ed441dc7cdf67697345673e041b557ead726c9e7d656f6a9b7e5f4b892a652966357c6293964a27b6a061965e893aaeb1d4edfeae174e68251b5648b57a3bd2b025473fe25122339ae4ae889529af34b2cf032eabe3a4ef75cb4e0519938aeff801f4490f35f8498ca9f39dc10bdb0aaacfe6940f95bc8b9e9c9a089691dccdbef1ecdec3b6c2de3b4cef6c295cf53401d971d3a7487b6f137e78fc9cb7a1b0803c98f223362bdaa42e453e4cdbbb0b46f8653f1d46da81633eb1faa1c86e1e98d6a7aac7ca9bc9bd6953a84c9d1e2537140c239994e62aa7337ff12516c4c8381e7f7253a5735ab468d86a4d399406027e808177d45399068c1eb61320f68e3197de1dfd2e0d9cf719a8ac04b9c7387ad0d2b7f29f49f7f7b78e232beab2f949ab8b48a6210549ac2021f4bf1c450ef2c02fb7012f13b0a6648a1301268ef073f848797de53bc0b7d7ac9fcfc3191ce19eb3f289caf7f6b2e132817a1d46b5376e55eb1d219c8292b410498f57a2e7834b0264be59a27b8f4c1c346e0bf60a04c01fb99ff283100b38ba2aaaa05547a50b9a41ac0f11e09f2d5d1338c9f7bcf8793e66ddfd2566631b249f4cc32d7c6534396a5437c11125c7253e2b3b4e1415587569df8f861a8e6ed03e43d255dfcd2e4fbed120cf34df7bc4d95cded1c480a02849fb512fd1ad45856d5a4697d5f78fa159ddcce71702f7d2cab42015ec0bfbd2df1e5e3203d93dc2a912651512bdce080e9a2224892c2d00252b5e6393a3cf461ce0e0eb60c47fde44f0cadc6df2b0eb2c1256304368e26bdabfe9293ef681c6e3335e35a1dd81c7cbfdd644a7169b97472d4a1df5b8c49e2c77842abdb062c274de0224df2e9c2e6b52cfdb6a5106d9a7bd4c461cbfc468019a21107a6feda5783022526bf77ed608d2cf6618f3fc2f5848fd8ddad0b672b0248c953ddb18431ce9d94a9b3f166f6f8d6098212be209bc76b7536b4570cd960b4dd4bce9f0ddee915e0b20bc0095c1025f77bedd5803c3e647060d5cdd4eb55881e7c01134999c01d132c693108a53fc1474e9f35b4ba20b04d61d78154d6569a2fa0a6c262a2aa2dbd35f1851714d014456db1b2e65175561b7616ff4646c3b13cace22da8e625a0cf14d10c89bf6348d9f9fad42a9ca2fadce33e46b0d05ab4d2d16682825fe5a52a52302fc7c56f0eab6536531262c2e4d2257c8148d0a15b34392e9c404241de743e1dfacb0bd93d5f7d860dca11024377a72c57d034564dec55620a07d0e275326869b724df8fef0ad901d9eb15973d938a70b5b9e060d5bba1b7c5bed477478363eee4b334efe489cafbce49148d10f90a25d87ed79deda9975102f356677ef5a4a4f84f5f76cf775dd4db1b5853db5e5628955f2c463e88ef580fb69b31dbbae3fddb367e2bc9396a458e26511146017ab6290;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h3593963ffd489c33937fa15595c513ac0277c7a9e22ea8b915cca9094c02b20e41c56f015405b4fc3cfea792ea75198e90d642b5fb0e2915932137fc7634d1c2e6bd736b9d9f740add528d6eb585a3464db13cfc0d87bc980c5071524ed7c830202ec31c97c61d93f4e092f8cc2d481c7f16413b1ceecf2a4772b3781628eabc33a26fa7389434a227e9f193e83e236fa2bed1c6f5d73673caa54812517001c85593d45703a05881f8409aac871db704607c186b3d539f7eef572650274c3e0ebd3ea947062208a459adf64d75fd973ceeb6e002c21fad53d054843aadd846968ef724d7c9b6dfccf0b267756552742ad33bd99ae262f0b61449834e6ba9c1421ccac43143d5d9a748d0b90275ac0c2a050786b8c4b77da4e0d7713a6911bf0ad9762740ddde349c32ddf5fb1ce907dd1e613be6c51c5a48cc019d09cf30a1e459a600ce45c75a2778b55c3f22bddf0c15f171c2b43dab52fadbe8f98b5f593e9d0c6522fcf5ffb334dedec1a15c53f8a259140fb74e15b542e6d997fdf458c3e617d3ab2a71563ab6dd1c26c660893f664550caf311413ec17961cc7537c9b7d640fb1e48b39049dbdc3cda1c0a2e3c0bbf91de57871321ea102a0ce957419adc0e9d8ea14da248ff98b4f727b52812477898ab431bfa352a4ab47c2571a485778008a601fe0193998a814d374ecfdf265368faba945e9fee47f9c6ba5c985c2bab87c55d25b534d878a7d30aab97434767b058b91c75fab24d76e913c04337c8f82ca6fa24b2cb0afe0654ec217ef4e30fa51286df3ecf7520ab541fd991166b8927a743b9b74070e338dd1c9c4e761dd5c6f30b764e9ac3b19b8981b1f3deeca7eae1a78569e0a2590cdd44c371e82affdcdde95df3dffc2768fb84b7918155670a978cee69a110e7a093fb03e10a2dcfc2f482fe3ebeca23488391f394d8676107548f98cd97bf55d169ec509f36b4e57db80fe7ccbfff28cb8d5b3583d7cfa1ec22867dd5c7ea2098fba3ba7d7e809d89b328f470532dd8b468ea590edcc77f115dc46e953a8ec5c55423e113e38117368ac226309b86671a6293dfd0f6e95fc2cf109843c12e9353b4d0da2cc88ef2d005b2afdaf1dfec151146e865a0838fee731f7506beadfac84cbbc373b5a081901a9bf158f083961b99cf6e337d74dd52847858f3ba568764544da5fa0f5a98d169388ed971cee2b92a0829bd6904943bd3de9548be94d3a3d59cbdb880634568324d4493761c0d8230fcef4a955bd0a57f3ee9a6f7bd0de28308c7184aeb6010f345c113a10722336677450c1e5c0d6038c69f16b046f7fe6493356946bb98dc7ef69d2e15122c804538420ab73f88618a218120511c8d8269f096dad19beda443967ed10fa3a450ae5c9de1a1c84cdef944ad76171ca7dd0c33bc62ddf8e0c8cb5ff24affd323b625866cd342f3b05083062ebd9edae5fb45942f89ec24ae442409eafd6d36bb626cee469a2d368b3d0b26dba8c54f456be9a0c2518ca8e5fbe7ae8545528ed4f426f5a2fcc547f7e9c35d192c8fa7e5172332b68603a67473758c004ea8f3b38e008f6279c7d8ecf796bea44f3567fd2ab89016cc8a4f5a37eaeac174efbd40db196308d9758758d57cdc9024b4d22222b47e4fb77a4fe231f9ab193b820c5db0845098373690b337ef46536c6f6a6e7794bd620cc6e0a21c36ba70224fdd2c0127c74e6d4ed61fd41786843d14991f3c98e04be38b13c37dda25fee6628705465c00299b478ed1fdafd224f709841bb14a812698231c2591e793936d293cd218a05e9953680b334ebba8554702facdadd34a0465d68ca1fb9ed29ae0473e5039e377f08bf124b1c4bc9124280793fe714fb158738a7290229e2bad124fbec2adee0ff3d8a5542300da1b42ca585a8aa383f3bd2ad9dfc1000ddf1d58adfc81b701efd534352e7a4547d5634d633263ee6051b1ff5b304f01dab9e1bd8c919e2d6b73e1ad7a30719702930bc9f1d08b16a207af424a353380cb58e49fce1d53127ceccbd62f63ea189904e08d1eb90def072aa9214153072db910c0192019e27f7e26b89a8745c3788124804302f1bf76b7b61955435fd1daca437bdeafb34a6ce636e530e3c805964c23a4b5047b15282c9e60ec7c929624d1270a79570b3b80276275b145ab32351c306a098b35256aefd3ab4e1593352830d8726c761528aec8b019eefca6ea9ae71a2a431ba7d89fcd9796d83c3bace01f90ee8b19c61a074aa62a6afd4342a20722b623af0988d30f2647f7951281feb84a0d6269b51a692b149d0efb909c45064aa699392abdd7ec38ccd20122fc64cd5416eaf0c53a733e6eb78e0e39bf7d07cff2b55555be2cd53394141d34729ce87e1f9d834dd5316217246908d47b069d08751b2049174c76bf4825adcbbf67d3b1cf74d0280ca1e8422901af8920f272e4b6356fc9038a23fae1496a0c67480a0959d758f9a841f1b75e3283066176089f74f329a4b022cad37ba53dc7374bd952ee424da13f063f9f32ce98ce7271c708a09b4876993adadc62b70a1a6014f5390c9be94a2b63ccafae26912ef745ffeedbab7d1f9e75cb02487f3fe219cbad95302881c9eb4dfea34e175e2930c924de2b441dc78b94737ce0d2946cff1fae9b4b43f6898c25a35bdb53ddb3696614f0803da44e21b04182bcc901ba832161689c03bbc4003a31835dd4bf70293d0136328ca61372990e7152f7a6cdb20dc2317c90523772539d09d69eb9910c206ce727e393fc7ac407935431f9f33013f073cf05a91365809f170f7d2c35277065964a0631992ccd2c95d369a14534f40f44cd542020bcd13107b4f177434b1b0303965dc231242b954fb663ad8fed76d733bdc4952c28f806e5b76868;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h18dd3222273663f241f2f38fec8e570f5024b2fb2f949118aa9f3a9bbd35aece8c073c09471d7499ddc27745e39a71f0b56d6fff6e4df843a37757596b57cd74f6d073f3708bccbf2a0b00f726e21583b9c5e1361d2d22a0db1fc6ab09f3bfa81d20e953658c3715a9ec35099ef3f2e55edd996eafbbdd29760e421dfc1c254e0eb6fcfef9c9c769765a63577d8c18d26bf56d45919be7f91196202ab8ed3b286d334dbd504661508ab98136bbf619688b24581ea0d8e2fed76a8e52c927ffbd1c09f3b7355f53457f71887de55ded9fabbc85c85cd5b302edaca9b8a3aad7a72dbae77c9c935315f5c77b256406479a8b0a56891a13d4c85044c2591fae712c216cac94e42eece907dd8fe58501ee693d324f705aa21715ef7ae8eb2b98597cfd51a6464a77815c6d773b1c23e5f2f476f77d4a848f5a8b470043d98c4e575bb56f585f2310033a598e62ee70fbb275903913cf0190b3cbfd20879c32884818ff6e1827355b7ff4c43c0a4997a75e53a53f411e0998fd23d3a288e0fa969cb0bcca7482cf218bbb826a28091870e18b0e9c492e69d205bf516d33c32389db0e6d74113880378552b083b5f4eab45804571be7d85e6a40fdd32e6ed558fe41c4b99407f1bacc1f8a4f37902a36f8ba6bdf65287b28d1975147e74ffa31000ccb9b1b87f7e8eca893b6648ab1544d5e0bc9a586e10324597551f4511cc02b3f72f4d5e9c549b3223addca463c39e6a95d3c5253767be2ff6000a7dd08bda5e8789a9794a85fe95159fb5c53b01ec9ee852a429d7af4946515d8a1d585df7dc06911d89b590c60b84b6749603573c322e9aa70c1802c7f5829eda9c38a492b9d39de6a49323b08981685c49b8f1b9588216ee9e9a809b5190ecabf08a4ce684f4f86154f060b05781d00f2acf67bc90b89aa92e41733260ad5b6ebcdbe814112447da2e091b0d6b4e536279a747f84205fc4534b5b8141d942c6a639734217a48b69c646dd8eaaceed17f8dc00e5d4ff450f86afbc0f6b9113faa5b3fe070ee3154c6c8a336fe89b1eba641463a1961911bb1ea3add278e8218237051f40d93596e2d96e6958666c315eba23868c4701324f592656a3c9e4269a3671fa0fd8cdb047df50de78418ffe11fde203304c519dcadf4b3a3e3ca536ceb4556782a73b4ffa5256b820a2bcb2da01c30ff9787a9890134205a4d6c2af23296e586705ddeff736ce610374bf5463cc430438918d231286eaec113ea68ae31aa399a9e320d712bf2d06399acb165416a335c3f6969ef4ff2809c9239e686df666c667cd00c0849b8cd89a538fe970e8e2a8322f0acdf65f8b7596e77e4bc842fe4a55bc52ac2c2e5d94bbb85fc5522a9d73558304fdadbba4fd35d8f207a109c69c093f7ca83b6fe201c339c9300417fc01156d5734551e4d0322038487b4552763358a697ad5fdfcd16a7b1e5c8c25fc1ef6f196c54a1f0bfe857a2a5cd8b1910799d974e39a6d82d72913f194fb2d13430ae87da49230e4547b426c70f905f5af0a0e69192005eee7c4b2562e57c9148f9bd2165a982d2274f8f6615a4ba8e96ab0728dd13421f99ee1b2828fc3cb97c0edd60e22745b0de9a838eb23714506cfe14603ab482ea450edd71a81d04741a606d581fd65b2d570287f1a3d3a9db1e8fc767cc95a7fa709a1b853d5ce4f5e0e9a5c20204c5535f8a5add80ec979cd5d251ebe38b4fdbcf3d195f3d403f4c358d1ee5ac57e86205a6000680cc7d29f5d13b04502636f43c715a7eb4a52dbf4fe0568e21d912540f510658dc8df965cc85bb10e3bb95315f9b75513ca4019a081ced1abc8daa77ac855171aaac29f6697298cc77e81add5de168e96eb138171e8667e76c2b05231736acfbc754de308595dab43bb213175f0a37203cb09caecf94819d946d7cb31359dfe1fb6d5b475a5a1c608402442fa3b69a9388ba455dbbcab492f8b3e582ac116f6842d476f78f8c55f2a35891a08a8439369de4bc47996ae94dd31b905a57b89d656cb59e02a427ea1b9d6282354be72d4e7e740b4d2a82e94080481a3b1d86df18406ac4fce2404c7502162ecd27db3791ba7be3a468fbdf647386921190f0c3a5e14b0fe3cbc0af97838c958abf3f9a82d062be96980db293a9f9638cfb9adb613145b4baafb9aaf2ec56724c38962dc7354f35054c53b33fad60bb229707628a7362182709a028c22536241f3ec28e21227e8362d0f32aab324eab446c69af9a24a47d781d5609aebc5bc6ff99ee597be0e3042fa852b2b3548ecc64898c0af9b8884f870e25787870f404e72148f172375bca26202aa758b79f08aa9f0788fe08ec4283f5f354d983b754364bcaaa504a26be7d7c80643cfc005df06ae62b26017aca19873dc7ccbd15d99eb5b3ef75086b615271edf56682bed50be027cb214aabcdc85d6ca08e386d951e6ebc19d622c2d0465352635d7c00fa24842c4808ef1f1aed4b60725e2d3e8c0c2e6fb71d9231a3420a6f5831e9ad8c1d510b9f1972abf6b5ded3af4d674a3ac083cae5f0aa9b4d7c2847edb51342435b4c3da4916332eb7fc9f51125beb1ac3ed4362b6a3a44097420169e88811eec8612661bbf29776840bbedb66a6bd0fc0dd84508c74b5153d62205c6c4e344a674f369f86e805004b94a94b007dadef8be529bd9d64673efb8238c6cfb3faa934176c4d16e6defe5613406d448f34b9d5163b462469ae353b89ecb74fe23b8be6c8e3a1f605f7a8147e8db79be0d093a71668edba05382827f2237e89be7e2e7ef8d398f299b56bf219c6e6f7d3d12dc99adf0df373c5cdb3d16ec83ad50a8ff0ce81b24f66028be27dc2bddd70685b16891b4aeca762aa2f615bf42011923298189e16e4286b04f0c4627ab708c0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h33f5348a31694173293eb7c1690077f4e4dce18889d9323c41d4df6d078a58b20bac2512dcc0dcc42c916acf03b8ca43db695c9eeff0d9ce0a32699e943a0cb1eaa728e0690a47249a3ee5bf34648b488a31eb55d27f8c37b0133cc312591f7e41a9014cc29701d6cd85bea6bb3e9c73636d726df445ce7192183b0a3821a4c0ed836e0f2df6f9912ceb265ea3b9f258f9845f5ab7aaa2ba798747f54d7c73e6860ef0f0b643ae535219291e4b3bbb71d958428f5a0bb145ce1cd06491dbde730de71986665d5dfd9630eb8c77243975c42202fd24e01abad1aeccc1cc043eef49453cd82895e26088a94e2e16a79a6885c1228b0d9b8793e0662caa4cc33280b195e849fb5e5e2f0a85ae7cccf58f8be833d33c29daadfcaa6b255c6e21458211c82dd84db646170c6879dd3133d0595d131032764e603676018d3ab433916b4555a07b7c814a0dd1e211622855d3ff4061c9aefda4e1ee548da0145a4a4d3661d07b95cc6a4ee311a051c36d9d97210637a7a2bfe48606f065efac1410ce3fce276a16103c2b40c366c6baff128fe4bbc63e562bbb0ef2ac0eef9283a6029831c5ff4fcf4c8d50d500051fca76b57595598254eea74dd93bdde07df011d6aad4d2a13a9d43828c3fd8abee6e82666de2a756d9af6bb16661ceefe46211ceaf09f79fe81cb9446484b08d61bcb92a55b55f4a40108be315737bb47d7ee7298f2fc1b862ee94848f8c90ce2ff59ac67f8233604a8d65dd426deaf9c1762281224207990fbdc27c99c37fa2570c3481a66b6045e0e0fddf6fd7e300aa4f6a4e7fb8a410ee0ea3b2e80f1855df4aa6f63980b07bc9d958aea80d93f6704233a4dc3ba240538492c5b32bd0ce2904d42e82eb766beed7e3df30903bae8a20e7073fd9c9d49bc3a5b7bd10f9faea6ebdbc7c995fdffe93b4eff3d55e224e2d6840116f518a9629b8557750527ba0ba5091e40cc9cf7b5f9b190c34f29d20b24aaa5ee9272fd6f7bbc0ff2053455b0cb515b6dc806877b387ae99a314983bceffc9b651f25050fbb6983536bb05dcdf180b8fcbd235c353b21e0a16b25ecddb07b83c8fde53f0693d329c43c6fa500c792c50896634bd8b40ccbd969e74acb297f786611a1f8bc3380fc2f6b51dd228a4af7011e92da46ea9ab2e638d6f8c5552187564ef5c8a266672f0c5e35fa699de31afc70aa6d0587b2aefae245394d6e4b9eda7803129843f8a4324056252313e626148d916fe4d558c2e4b699dfb83f54d15e46be0fbf6b2862230384587732ad97b9b7dc982cfcbffb6887a3b76388e4eafce3ff826f483c02090461ffa50026971d128df3bb137243731dea78e00e4a4a0e0c83b8c0e674786f68755c0695552ecd90e65d07f500a9c50701fe67b9a6b51cbba459da7e00f8e14240a2d35589aa095fe468db4e08df07e2dd3ef0017f0896ad9a5c46ee13741eee264216ac2f749bf054b76ace3f5422a602c0eb953aa5cec4ada47428879b8840970e9f3d829f5b92816f05d11e8c136350f11a272e9f38fd27251898be941fd5b30226162bf62965e4ad727dfa53f7781b1323e1e8fde2058ede9bbae6891d7123e24221602474eafb2ad6a79806f78cd2cd3a45fbc52cd26c5e33e134299211591fccd38c78fd0bc8f5015527b96fc4384c565173443209315ffaa1f462f9a8b74c5c2e5aa78316bc8821d7c790c0ad6a7d239c8fdb00500395f3cf354fa4d50ccac01259267b4dd82cac56c7fa7cdf4df83e4bcf28d245f6e411b1949316c3e4688e991dab700f50b6752c789cebcec120af26ba1c26c3e28fe68b9341d6e9f5cc9538a9bd1ad9cf05b30d4c740480809a63d9fa4c7096e15a44610931c9494c350d6aa84146abf4fbbb88ddbe3a4ceb15fd8c8e10bac092878273da123af0f814f4ba0be89cf511a9fb5ba80ab4cfb504bc70008a81968f71750e3f1fdf7bde09d00f2efb4259e7f3d70221b3affb04620ecfad2a9425d65038f8c68b1f5e50f7f0116c17a2b32c6c71c7ac49aed9145616f3f96fc92091717f06e88e0737f56c452cc5fd2c131105ff599b84a0def00af694f2fa060026fa75b68cbe31b90bc827ec9b9ce0dfa84322e32058bb56b7b2bb2cdfd1dec81df6b450a14aab744dc8046153122e4dca4e30e50d126b5db8b29a9d28d833cc09ff7acb0208d41ee0e2d0e007d1eab44fcc8f925df27343cd9ddc9a6363e57acef226d8266cf4347d8a0a787a563ea97b153fc985a10a5dc06ff295f8c4e9ca546a8b9a5fe83ede0612bee6553809e716eb9bc27d8e25bebed9bb1c15175d65ab283f9e538c0b79f8236a9cfc038ba20dcbab059992f19259e54d142c0e9676ec8ef8c2e2715c06fea5dbc9f152865d0c291b5a17e2f85afa1bd011aeb79c6c7104aa4acee541d86e544cc796bc75f1ea4f5209dc0d67c9d65afc1a32cdbca7c82789dad1a1377668050b4af344ca8461d9af1e98632a1b450337b4750406134f5821df5e110f913b96e535bab07a1de80f549ceceba12d9733c7e09e1cee1723080140c2818f54bb2598d97ca1dd2d331120e8f99f467db7945814ab88a2a6aa63757e94a78b3d3605c565a1b127df4de256b87305f70fee87e218dc74f9d87d9f7deaffb39680b9a5311220eee920ab5aca6f16d2a88d54fd86430d3a51b8898a9d703626ea5944b0d39046baf59d5febc83daad09a84494ce70bd1fdf1082ed7832f7b148cc815091931304ed738109d83b40d0e306620b9d9b9216934c041d504c3e10b37707268dcf4a0f4fa008089203ae549224054cb4b11f2c89fd9a7389624642d67337fdde8652532cb788ae3fee649c84e07ef2149e678dd8e7b26ba9c8e7ee251915f642f27fd99d93439a9b860582df9c2fd14f1974ec5a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h7f41bb0caa42634b02b8607f579361ff8221b38949b2dd53fcef03ba798bc73c739f6a15bea17cf9d4f3c952252f6f3588107f8f0d837124fc94afa34b43bf889020970171bf99b1df02177329c4b67b017389e8f1dc39160490f85f3e46f302ba4a6cba50017670410002cbc9ff00490f8c88b8fde942a34313495ca1ccc8a463ade17f9d3e258bed44cba4e119bb3a4d8b1dee75d2d7779b13e0d62a4b2dc31b0c8218bf4c1612ebd73d8eee403e2d2e6dda34a83a3e9a160e024c7d650f43ab11add4e454bebc720a0e466ec55bb5e784ce8236bc7766f5bc965e364a94bb279724821339ced2c58a81311cb3ccec1a69bb3b047b1da51bc28f2534819aea9297a914d241454e8157f30f1d73a2f6a47e63f00a6fbc44d9c3ac3dd596a4d750f11ced8bae1715ec5ffc5b381bdbf3621ebecd7c051b1ba8fa6161148e00da2276e24a1644e6828beb9c16503d647be3e879b3586f7d594c5e8b86e769d127e7f19ca6104c13d58b0f62819ce8ec830ca9a401577e565a380db743f0b6e5e79ff5a866021aec0fc6a49fb28a74ed1f941c3c460f58bd44254f0ced5f9d136858cd62cc202833d62c8db3e3f666d7013b64f5fe9de7d9e2cdd89ec167f0a81a2da1103eab21bbd30849c6b9875fd84a6594b80680260b45340d6840b02987c5172dcf8275c386d122d8a2d0e4a07728beabb2b868d5be704c25dd9805f57f72792a72b598ac8b89e25a2610fada91c4a56a779b5ea52ac434dd0476e29acfd83868c89563e3d66d1fc9b79b418f9e9b812df582f27665532cbbb70c5b695aed9bea51bcaae46e19e6c68c310c4a2c53abf4aa18fc6ab1068ee9e0d5b2a44a538e9405062564d44e6f92ce3b5b0d0b191e8c1becf9e54dc14719f5954c6b8288d9748aecea3ea66992eca74da22342498761732f2f886165c6d5e1d4ec74621963fd6768fb857dc441af67fb76158c9aac1f7704ed8740bad87a5b5a52bb543d8346a457400c44a9d8679ede753aa94a867b8db1946e6601e45a990c795923e89433505c80776ddb86b315a48de1bafc481860c4e1ca8db125242fb78af0ca03b34b3a103e9e097362670586e23a4fbe55e5c30fb97ab6748e6bcab9f79fd34bf92114634be1f509aabf1751461d9ede44b8c9086e8843b1697a65ac5faf175c361a3980661d3b3b6b17c40d0d4ab9a8c4daf84a8cfb68b52b3726034e8e616a78f1271e39c573c570fdf0ca198bdf4d992fc7cecc1fade895cf85a71292395ed8615f2a0467ba55f107fceec37a968e1809930e05a7ff76faafed5e7e7e0fdba2df5d67e7b57b1d543ef94606329c3c245e4cda308f7bc7502383538a731871021c59f70ff645300774e797e05f578fab9eeceb24b694d7897b5c08bb59b12771bf00c233ffb12e4b05e0d6adf4c181bfc22b5595d892bad031a2c72ea369b7e9bb0e2214bd3f2b8a11b0b2020fe277cd38561819e22d6784e02ae4e39cec6e659a506488ef45d2702f9fece578020f1af1f155cc67cab662dc6a815e076449c2377e024471528ab8892e15f4975e7704e44093b16902e3e432efa24668f9da70aee1cb06891e07f27050f33fac4d40d1587e66f6d5c08efe61bf9475702f6e6a75059e2d1b81bec7be19d067dc0c0184fd228741290c1f99081920a60b6143985917448ec4e397c0f17cb2adb993095fe42a0ab9a8177969cb7da2c812d9be179b2f98bdce0a77a2a411a314adba0c98d7ca5105cda65c8e5206009c911b7d6c18b663c1549ab69a75555f22e930ec7de58dee002312ecafe06b8e8931fdd15b8fa6c32a1987e0616ced9aa6edb11ee1b66f7d7df08ab6425a4fa99a9568422903cb3ea42e23bc360e8b3456d07805917d4ca91ff076516d4da0245b282c84a23c3dca6284077200bbd7fcc3b051236366927fc1e6406206ddc46da12d38e55b2f131f660b2b66d8776af0ad92b59995b26ac2dacae4091bcc233a5362ccff375aeb6b5797d28c6a372976c24355d3a84d04f4354b7f8bff2c1776ccabe19b3f399abfffa65ba158a56eba82b14a1776dba438704f3e4a38a55b2317a34bfac0875f94d5a0c43344093d51c2506da91af94e11e2cc0e0a3f14aab86c33f065799dbac75c166bf1ea23afcf11d9141ed2f2fee67d12cf713c80b7be73f8f084f05925ef47f3c572b367d6802eccc60550ee91aa9b2b11e7570cf253024388dd9c4287c32f60bc19c69e5b8e4f6b8ea452a9f6aa9c41aaf6f51693e7b8240ffaa076662710ccf874aa81bb0bf8181bf0ab92c5ac48a33c731cbc70e51f60fe2276e23482297b8a3bde8dd0b5cf95ce1fa4a066a454832e4c15440281250b3e3a4aba7a4d601de895f897083a81d91dc712320b39e8b81efe7937605733dc1c347d8947dff30a5f5f70913dbf300bb89f5dfdfddfa7da276a5a71b6b768cb785e1c14bbbf564ebb4cb7ac4b6a2ae5992ea1869071e8a4a159f6483cb1cb4c019806c061627659c48f0454be6febc66701db90f6806230770f17006cea38df7481e40047f9d70d7a9d55437703d1ad086fc92f8edbc8472f8381f76b5b901d454d674d89bcd7c2d72929bfc8c0ea2793a39ea8f4a7bdabcac5604df348996904e7b2e399d15438adf8d2ae415f5fef036d045c76d1997f1fdfe158f3aef4b2b6eaea477f7d48082a91c7e5aeca5c7c95f0e69e2e2f382c20966f9862ee7d244f68ae2b14ff406ae7513546e4d8c6f9f118fb6117ac56e9f59fb50a18237b0cea6f0b3432a58323ecfbb556df1f73abc290e3c0de4e69908e2f04da95daa07fd31eb0044c3dc03aac9bcb6304c94d2fbb2b4ac28a54d637b9502b7af155bed474b47a0e2af5f5bca48d8c8362571f6371985718e8c1e223ec8a1b01e63546c256b1;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h80dd20cc689e76eb700e6e97928c21f776ba1dcbc315f3f98f4e025382d1b12080f28c40345fb791e24a1d7c8f238fdbce879f311619c82e9bb045508a7f417337e626c7079eaf43389a35fcedf131306e0290616b66c168d4edbfc05ac956e94bd5ccf026d19aa4e5b888f9ffbef34fbe685b074c75de10b5ab1eb21411cf1128ddbbdcd1377bd582aa8f63e4ec73b77f87aec918c7aac51b261a0803dc0f427299b147d3be8d53a0f3a1279337404b72137399606fec74b9e5318ab8091a5af69f8cf27d3b064cddafd09a96b83ebbdd473501d23e79de3a7cb0179382919636af51f4a4d0a4e6811b2ee57879565984420870830147c63820b8ebbe66ab61308e3e147546054c8d1f23e834825ea3b0de1928726e25dbc71fa813dbdb832454d11fc680e320a3354accdfe41ccee20d3b0d6b21e827aa8036871331f9a35ac879c54913beef8d02d1955e800e1edbf08d937417530e0338fed21381b79bf4bd916f2b36735e5f1486872d04bd8a53505302a8153cbe8321c246a978dd6aafe4f627a133cf747ab7274859ee525b19a5a60b3d184fdd8d776448bf0fe633ba8bc7cc0780bd0df9498551db40bae89f2cc0c5eb03613e17f7dc89e3ae7e29771588bda7a66e653ee96e112028065188d7292941ec24f5280bc0a293e88aacbb52530cf017eda8d236241df756140d8a5cf09b91da0793273674478f4dc6ecd10a5eb797ea3cb647fa1ba50e826b85472861a083eb7437a17cef9cab00194fc77a9a7dd77343b227598dcc3ba46ff7e92b9a2730c7c8bbe422ef738dfa97b7f0aee2903add6cdac82108a24a9784004a707416123198e2ae87310b4105820379d1d1188f6f17746d948a6b54f908d1fb46e3caaeb0654dd50a81f3560fe392b084f9e03d6b5ebc8c994048689ef53732caa57780cc7553f1818b1a26d53452cdd024697dadcdead60a93cbdbf5b62aa34924b36d9a7226982f0c988624004b43a19263d5a847941fa09a86a6c69959493af2cd5d5f78872f4336909d53ec9f620a7e7b1ecbf540b6b432a25678fe77453c87542f36ee5e1e731655ce5c8dbdfd9bb8b046c9db8010afacacfba2971f8932fd2e83e3d61fd2c9b7ca04e63b76ad5d7ff8481aed21c5ec401abf8697ba4585f8e12d4570598eb05d745245c911c868c77ae1128bf87c773d64979cf78b3fe44492fb720bcaae0626ba110939cd31c6e41427b3c9e7337225cae842de3d82a3f301e4db764d9000331f4eb0eed3185eda98bc9474436e0a5947708d7638bd7f3f5270350672b7d8ff4a6f195939ef7b25647b6063c4a019d6060e93239f9c649ff2cf36f6fd3750403d93ca80d2830fc43c109d9c1b9bef2cbb452d751622f4b0d8063c67ca3559f52260e443497be5ede9f3dfea8221d488928fd136cbe12261bdb75042124999d008de66b48d44772c2bba1d2d8e376c56592ecbf580ce8553305e111114e7e2b67871e77cb23797e73ba4fb42ae6aad4e66e8188c33b530176f0db8d1bcbe1b7dbc5b68074a33729712a73bf82eeafad7df317be8bc0fb9da9b3d3b13bb2dfd7453bbff6c01f0380a333ad92ee93175a249d4d8e5ba1630f9ec6e0e92f70cc82567d531ae2f8a62e107b83eed3799d7cc8d6fbb207b5d1cefbbaf8d6d40376c739f03982ed6b7c45253562246bbdb8ba7277f458f9a556ea73d244bc73dd4a65bdc59c1e2a4597e9448fe1ac57d079f43579c340901e34e91815993840aea3863d3e30efe92ee9eda5bf9e7e6c6274be8edf62dd1022340379d9822443748afceda7e30f3f9ff1b0c0ee36e72e59f98d75a641f3a8f62cbfdc7ede0eb462979fe17e51fa7fad924a366027fb67335fb69eb9ccfa77af8e34a3c2048b78586d8e8c81842a135493d4fb4cbd0d231a2e9253b5f1ef25a131dd129aca800f9621d96d04aad73de40a3a274a822ed235e73b650bb86998d780bcc63b1d0efeaad127554a32545c3986a809dde607df4e208b7ea36f52ce26f2fa60317b994101c63b65a5fd534293a186a0de33b91ef72299c77dbbdf8e6a403e93db50c6e8b1c5b16429fa9e20e2cbaaa398bc5389423956a86e959b2764bab6f86ce945c0439af4e47333319c2524d8de49895f868d8893385538309a99e5ec9121eeb02c5fe7750cc90473d52ea4b58cfbb8c76a416540b315d0255204498629cee473f0c390ea8d76eea2b073105e284bdb5995f7703aefc77996becb049cbb7f7544eda9cfb4e3ac608c079aa45dc38e604bebb72ca9b37f1351c52b972246257196592d10e82923396f2df8285ebc6f0677c7453786f2ee81f27ec3069dd095534c59b0bc272e53cb6032400a3419e867e8214926b07c8569bf977be011cab7c9831fceabd669ebe3672a6ec83f3b18803671782dcacc25f74e385e590b3a93ebf772180e077ee4c7fa216da074bc0abb17d6dd8a3f64d7ccdf5bb5fc893b13d115aad1ede07d1f9db7d62dc23761be34361c4c8dc91c23e3991bcec8e6783a21b516d8afcb1cfcbab394d4dcd20329d20754bed7cb844d2269cf39f4334af5008c9e97f3ac59b31ab312d5331af12bad500f08af1661f2d0407edde5813be22b3630e008808ec6dd11f6899002f77f6bc7a48ca4ca643de9e9d8fabcb519eb2158b2ebb42814362f7471dc6f986392c09b8b8c097c52dff3fcb132d3d2b5f891dbfc3733e7dd217f8dae6d923f36271f4f17b98ce0f02069d26fb3d7fb5e0515a357b656ad671a26201ab6368a99c1ebbb9c3a524a1409596cfc1593ff912b0b20f4e21b0281ae69160297a55a2c29f78f2d515febcff8eb4885aef00724ab5aedd1a8f4fd87ac45f50beba24a562d20e18bca163f70149801fdfbefa23c1dd07d8c4aa57c247360a34ff89;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h8c08e735dda0dc8a70b2d24294935205cba2ef54e2f9b81a0cc29439ea42654ae08c4231342b8c7ac1f86abeb08d8b933405aaf1818bb25338b0f92175448e89d15a3d35bf72737446e0685f54131aca894406f7453f58b5c21029cf10a2cb1b39d9caae127c846b7a9942ae13ec46642122e827610367d1712840626c13910aa0ee6cb249031c60281eea1b0749c6304c9a3658b343b64a5a77077f47ca41b070818e3929010b812a16084c4c38d2e7a9319567ddb4607259a8bb2ffc1680eee65abd77465c99fd9ccd8ef2e2ae289e818a429adbbcedb178b171491246584fc17e2a3a284f70bddf0e27e7ad4611ba4cccc0876281e250dfa6a72b1f55837346dd574e8896e52fbed0508eb74755c5f5221aca4c6f4202d7db0583ea9584014a240986500427c163607b412d6dbdd8bb6754cd76824c97104dd3d10309251a873f226bdfa2b177a5e9f2d5acbed98d917864351d97b01e6cc5977eb19162594463e70c681fc1345e2043b1b859d3cb0c52a7f584ece46a0af4818890c7cc456325c85c68620dcdd48b726e047117971ba686144ddda3d1102e1270454e0d0ec5f1c79e50222f89c8415d0a4baeeac3cc61cc0cc2c19861822b1812755dd3026a6c805a200d246d3eea199c9fdbbb970545065febf73e273c73bf02c0c0154a94bf2f2d2b0bf64e36d92e7175db308eff74be5187d9224d4427549151cf9f1799bc0dc4eb061b3602e1f295fde3d9471f4fa723938fcf708142586b61ebcf2f8b80c6a96d7eb9330205fc4e28ba9ebcde91215e5362cc690ef9fb864a7a3ea303076bd8c90a65d86b11f51f326292fe8eacb3418b3bd0198a0335817ac246877bebe374090998f10f89d2a87d34ba2bbcee7137cb390a63f133e3547a92e30e83390ac6c4525df2338504cce62a3a2b51aaa9ab4051b2c4346cd2f80d7a73453d50dd72407c7204b364cf31f6c0e9ebf1c34025d9f03f7acf67b3fa4d752b89e6311a648d60baa62b9877d79ffde08e903c59a81fb772465ebebfa3b86df32f39771e8495b2e7c8bf22c3371740c2033a600b1e14f46bc5be1da4d65a81150ceea0a437723b9f68caedebc73c8037c69a55889ea5c2c2a1ec0c31b2e8f75aa7030dc4b52238e2687846446f95ec000dfa1bdcfefeea5b3cfaa0850c7b5cef967ba88527fcb68fe369b1715f483428c029139c8b4a18a12ed26857ea66766be38639a3ebbefff53854c05159541e4cbf9bf49a92b02278fb544a69430e579c6d5cdf87c2fc4e113ac1b9d640925c6ae3c227e21f51e2427d971f7df4b65c4c1fefd7039c8dabefaf0e7a131433141e2653eada86315ac3a47cded31a6152aa1be9d2858214c3bd2b9d01da8208362ae71b8c98d244f0a7127e17662fc4dbb854db102dd9d866fedfd81fa28ae232599c07d5a3e8cbc7f6482f8283c4ac4de719956d5c7a51122b075e90dd215d46a3c3daf78977ee2a339e91a1d183a8a38f1b86e9e1350d89e30e9904316795a5f63f16c3f474c298b8d294193b3b863c7156b5b194a6df26328710057a0c3fc8db21c092f5a3b8d907b607fd7627413449a96c389c9e917c54a7e65dec3f3aaf4da55162e87f379cbb30f42e7b3bf5627793183453d310158d553c7a5ff3c6fd9aed78491db0b130efa7388fa8b0bef57f7fd1c71d964eadcf27b3b21339601b57219cfc15735aed09a28ed71cd3350fb133e92b0340c742df5c55508557cb7e753e60bb7e5e45ba7cdc6425fe51e78a7e0120556df89521e050bbab1a84b5121f24eac82ed026e71a82b9fdc8d46b8c325cfb354e6c4464c6c5178e283749978adb0df2b874774cdef74bf3cf9869b9a7761f4461f6fbc1d0b72bfaf4b5ff7cf0f12ad9ab48414e0806a95867de56c4ec9c23a60eabad54c34145fa4684bf20bf61ec0fd575a36539fa10ad97b3fc08e37fbf698bb99a8ca8eb38a46928ba5e8ebd8b890df2c12d8255edfb01936f4ba6a3d5786b06d3e2fc945474c6bcdcfe4895aab186c36521acd5a612ecc5841f357944f5dc984462533627fea075bf6774deda97143c20f33cb71a14497389dc2e1bd27afaf9e2b073c33dc714207b0a9f47e6503c3aef04262b294cd8c23c43922771bd1b6185fd2b326222c02e7e8222096d3a6940e77287b10741c06bddbf037e4295820a51a03af421a21c07380b0d01638dd09c309356c11d4cc4b1d1401853c53f0aec5979e3d8a57bdbf1ab162259de07b70679707a615d3e2560f22092ca1c66348129b0bb2e7923a18114912c6b2417d94b2de2b9c91ec154500e52d234e21222a524c18f3fe455d9de9cbbd0382bbf485ce74c21c48e14383af2d10b30aa4b193895ef3c2cfb6616ee36cbec43067ae02873744f85f11a01b2e8fae85adc7397b4d441eb9fec676c4625e27f335ef3c1b2c977b28d2947f00137d4d10badc26bd496abc8cd4f58a93b2a417d922c88c4841aaab4c04e78a3dbdb61ff369116fabb667511ade35a0428a1af1f0af1058117c2d45e80e86b61ceb0a6fe2ca17fbc64ab1b686e5ac40a5cbbd9c992af3ecf568e1fa92c1cc82e0d15f012e12e603a8aa15606439e2c7732ef62d4afcc38950c3aaef5480649dfc3ce711b02a249048f64f76078617db5921c22c8285b7b5be10524e2b46f17d811c4397ff2f2ca7947b4336d591f0faddd51b8d7e3f8a3c5153e84c2906f283ad83e34fe4e57e2146524b2bb26461e6d0720324f806df1f65c5bc26aeca07c6232c411469e62addc252636da65a45b007bff7b2468910a06641b9eb6fc50a55d650730930e55acd9f81a44f37a77ddaa785abf438e772e051e2115b4f74903e5d695dd9256804058f1f284fecb5a54bc0a5dfa1ec5e6104e28b6b23eefc0f03b331b3aa1a7;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'hd62d46219cc355141151a860a9c6312b89266eac737dd58a22912b9716463b81aa61c3714cb5db9e5b1b44e0dcfe6a786ef2d18262203732ac32297050b663f6dcac2040c2f9e53e92b68eb29d15fbb0f295d8922b5f11e905eea02902cd3c025430906badd779276c28faf03d1029de22424d2bfae0baf9f8f8b17520a13165d0e57748a7d6a3ce6d01415b638fabd01a60a8347a03d05a552e5129e869a5f1563a9c12e3c9bf2314e18b3ec272152ae870398552db2a7ed605aff2d8f5c70a12692e3b1db5292be4fc54155d96ebe23a63563b6bca015288c6856ab4b84ff2bf1ab6100efa6729e418c51b1ab816d703affda3dc6742041587be8bb096c956e40a5956e45c88d03eee89bbfe0658027a034d79166a11525fde12cda7b55958d8f9c687d85c576cef645f6f31be358ec5cd2faf07790f0f7a0388cf96522e5278b8ca1e790dd605fe445615fb7a8a67750484ee3c9015253d70ca3465f420eec7c77cb6414906d8a3d956a662ae2f1fd5d8ff813b279d8f53cab89a294635bec9be1354a35e75e37d65a8bcd19314802a2a93a714b5b7e92a1c59f70ef60af40b37653b991c8c4284748574cf8c05e3b4c6703ce669dd2475d522f5d3248655a23a70ecceda2d5088790148c75fb7a3fdb8a78b169b83ae664da13df35f6c61b3a4444bb18ac8782f7a21779978114d4f490c65c8a7528307dd675b5f7a986be753ea79e73ee6fb4408a24dd3c11c6d1b4197cfd2183a490cae4c8e87ae76d29a68e3dbb33562f881534dc40fa610394c40545135bcf6410d232d85a85bc1efaad35c11163c7105209dd00cd6f21259ddad661d52f5e752fd9cb29209d76459e86899c354efc5a11ea0ee00b4940c15fc0dc34148fac9b6dac605709b459d9f8023c58cf43458144984b5c0dd045ee7c9f7656345b59e957ee0774310bafe8310291a826cff26dac5d945bf56480cb0ea3d381dbbd869d9d6acd5eda891d13d72e17e8e29d488a8931d4298ac4f335a9d4bd39af47e336f0598b50fa9c13f0356848aad2c5effe40b1b2fe6b3863ac584326d50e82188a20361b21f0e2e55080613743b3aa01fb0ed908c10e4ceca53e3b23ab863b06b426f43f9c7338ad4ac8a124692c81fe9cf5e67185005f682b8ed80050a4c9eaf43f02f5d30762ca87679bb971911081c5983201a023a163cea251260890afe0c19acc958b9bf2fc68635aad98c4516b046e661abe57bc861daac540f915b9ef32a228775464e0dcc4d3e2d4675ed7a3d6adc22fb0a898ee98554d56032a86ddb0f461450217a0d85bc5db5fd01aee51fc4ad41a3ad5322f5e723065b066d1119aac5f8b37fa960f50c80e43036b7910e5e4aa97d2526840d4fd6bd7c9d599d342459738792bac41ad09c4be2f30dd54e5fdd436fa164c859c1738fd05b86575742e19183815a8469f442fe2f7e725bf1695a8e4ff61fafb48662e37c94170c8e14de711eabf321e4003ed197dd36b7ec732f29788a4f3ca4daa7f87abdeb40fed8692f2b2d16c4be0d4b28273149e1a60d19ddb71fe4d16d50883e1a1c95f5081a56c3338d24b2fcd96877482d6f0e67719284a3151f76a93ac78349bac05679d272ca1906ec15cfb9ae630068527ef1562925aa39d041bc95bc4ee2f74459ababe876b9a856c9149376b0969cc32497a9409e9287c6924152e05dfaf685ec0ca8c77995242014a82f8c12cfb58742d4dcb791f817cf8056389debd2a383cc96318429f8897d453740f7ab021893bfc30bc48b29195d788648efdeb9b079229fa332f177fba62cd3c3fc0336347d735e084cda3f1a89f537947fd84a22c6254f8343868cab67b45999191b6deda554a0826e7df64b3e80d0a7d6656e6a71c695230428db8955ae521229c0ae1217cb88cc81c9a45735068a0298f05e6f550436645a757af4c01d5275d1a2885a7c04be2d592f4cbfa8e5c2421484b1fff7946671eaa92fd24d8c24114c4d6208649705b7828e6126a2086130806697ca2da14f15bbc12be9b68b32dc45f13346055e2daa4628c16d8c81323468b2c828c8c4376fc1c9a308b0cea0743e39802854f4cfbee3b3e840c02edef58760b3d7fab6e71fd9a97eee0d61e365758a904489a2d5b101d2b21b45e0109492d59f3ff012e1626361d0de91c69a20fb5d59742726b3ea4bb925d38a3065563d1e5672250e02879e5e1d16dafeffe7fe921bbcfa707564dd73ec7865f3c818a44e4104b94ea81b4ada0fe8af13ab821056a33dcd6151846012adb65b6a5bf4cf9f849f09f5ee0434fc5097265819212366878019c45b49de091bc417074d44ac4c4701411bf05511dbdd1456dbc60969e766806789764aead152b235b3bee09e1621ec8b509cec61736833df625d4d4120cd1f0d8a4e4d3eb98db94a3cd135572ab53382eb118cbc520a5db3949138969798f1659cbfa417835540478ab649813ef482778a97386429358b1a620cbf3deae003509a7a295b27025f7de07c2c217be698268a810c39d462f7c3dc8edfc153fb8e14bed5b78ea21045223cd2fc55a4d3c20431deaf551bafaa4fc4318b66f5a8bd187b78489ae75dd7d960a4b1c8ce5530e2855aadefd958b47cc3ca7e9241aba213ad802b4793123fb4bab917cb1d66ccee0b6f21c5ce48ab7700a02bf69f9df8ca504cadf55196bbc9753015c31fea52cd22c42bbbb793c0b53d00fb85b04eb196760b74ff820f79a79b4c5c6fbee926c4cfe3dc14bcea353e09470f9c00ad554a2850eaf9d190c983fc00d725fe9eb331bebd286c4ecd29572203589234635802630979cb593a55434b5c7d963dfafb2cd67aca963e43a5aba9f447d5b72c023c6af0d88fdfb7795b915da5646b8620f066bbf54f8b264674704098;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h7176c191e71c265b9c1765e51c7b7663f0b40367af20488302198ad6ee62cfc9dadb35e6f2829cafea5fb0b6bfc86e1d9cdbd3e3f7209a33360a1fe4197bd86591ae13811a1bb306988e6264611bb1cfdfd9946bbd3cf1330af0253ee0c8b36b1dcc89ad092b66a69806ca3eba8b564bdac1680512990691a644c7b31a6b6cf06ddfb3a139e7386dcd90d9e6d1cf7e699baeca8e001fac8d068b3b0abb1a459134d9ff5f173b9feca32dd7a7a74777e01a12f6cd82cdb85d6cf22905a06dcc7460733cca572f168d537959a2d523a829ea389b2fe938edf0312baef37dd4cc477d676ae9ca4a8d9e45cbce1801d5034b53ec39a6a0ebbb53fb8b66e47c2c947827f6e58a03d6e8384c08d5595b7530b232eb8f91bf4e1613f68ed2289dcd3c4aad2c768f7f142f100bbb2f108159f297af993e6b8e624cf9193c470deb6f557e5610a0125ec24981d7a2974e2bdaedad78c17b01d5bffa8a54ab6fbe2f773d03b1f136df09aeb58257072c301b1bef49603137ffbc5c8dae5d9c7d4a3e02e0755949ec1d6359784be6c6251cdfffb255dfcc4d432f66585ab082aaba8c557831f04e3472d22027563d7426c272cef872d16c0da733ccc61122d4eab2c86908c1c69c17b480ea41232653f634a2954045ab7bfb324f0a8f83975988638abe7c826966f498e79765cf674da4d354c6e00ab493a11c3b3a0fd251028dad65576d06a34eb75db12ea6de8e639f5d08d9e60b4bb55a52040e572a503fae22db4fac89a5cd7fad8559751f5b1776e6551068402a94ce8b9e929c2873a263a772b91da7027a5babfbea51352901c6b8b272aa5117f8d2ecd86735bcc1c2a30b6710226647258e308a24a2abfdeaa0bfe999837039f703256d0a4445b1fe67086563f942bd912830c9ede64c38f82b0ebbb4c7c5c18a102d391b66baffdf3a944ec5c26b592ce96e2471905412e70c4c73bdbfa9812ccf6d34d8a216959f5d810300c7eab0c82b90932775413f5045b628277b7ae65b04f80fc10f5e227b4f66a53f998aec6c8b7f35324911860b0432bb204b7c00cb60f8074e6fdfc5eae2f92ca34a5f6527bcb7bf5721854fc02bee9bd266b9fc2b106f66bb829b4e8528cf627452d71a2899d32f7ed592a1d2a50c6ea233edf95bdd4de85a106637e43bf7ae9b0071c0b5d3fbc2d2f11b90c8e0b81f9d675d2d1473163a3a08b5610ae1658b8ac30f115c3c426934a6e4dec222389385cedf4da329f038d8bbb824cbf0e6f666f72892ec21cc03d76367d202f19cdd2c15675eeed876ed90995421d468a4414323dce59ad435413ccbd114c3760cf8441958ef34753e1b8c62af7dc90d432958769b314264e07a9c00e64d82c0148ef3dd18651de3ba454a5f3eb212662ac181230acc6f7ca0f1f868d55cb923a7622e94f57e4fcb0103a719505598e66d21c08fb44952aa7799b3469a5a6f1c8af721e2949f6a87b2a4af7b9ae9e3286f19d4b123f279f9f4d63e9ea44d4d73001b7133863e85aef356f1cb4b172295bf957847f0200b90e11200d6a0fc9c018c94685e631ef0ee86ada0b282f315267f2d08a2d57c178f161636f8e9851b983aef7f908fb3f2bee346e6e65a2603554a7a84ccc1f7aa3b4e8961f87c39f25f4b7b03c6b6df212cbc6173fc6236d169e3eeb50685c9dc6dcd65ddc3ce88a80970c7287edb340acf692821b2eb7635d92231636bd9378a75a75623155d0d52bba538db9083cb3f27332c6e3c4d2f2b831e011f8957c58145886526dbfb1fa7cfc6e5b6c1f400453e51bfa95de56a61cb8f579155b289559e09e5b16618dc241e5a91360f61d27af0c982495d8875dda71b341cd7d5c02d8e23b71aed4d7760be33db5384a7ee25b02468e0b91a90447d49749c666101fade3475fe9f0f3c2858f1f8b592053d221eaac3d6a2f554db452cb48f5ba032d66db188d3b59bd4caa005d19ad090610a339a21889a35d00b454f11baba63c4cf6db2cb1a529d4f56b3b055e6071c09348db46891b7c9f029c9ad1a3ae3adbbad8b68368721a5b495563a8a78f7c0e0ff7e140ca02ab3ca95e2b4c9b887ad0da264934bf9302acf72e1f962099b83d99ab210be927a41ff66cb561412b25ffc41abc616a317356d7393717bc48a2e7d4aec2cd8a4d9b840215f6860c3c1ffe6f6cfa969b16ba1f7f210f642d40bca7c982d1b1e054bc4671c5b94fabd012f07691bf6297ed29f366db0bf25ba5a2bb171122f1405a31358a66cc544ee88bd797052efca3fb9041636cdde2c5c2a0bfc622960710c1e8c72d8ad090afb56a5eb0408943d78fbd758c8e7d3e2b246b74e3d08533297fdb71b2543a0571427ba20fbe33b010aad226b5a8009ec722d6b0c7f817dd07fd8569ae14ccb6777b98996bd6d40b2709905cae0ff3c73f4a6c38d23589d9f110e3ab6fda9efe744bc53506e199f07326ce48413986093e7739b8fe7845048df6b295e719172e4d6f36490a5a23ace77491e6a20354f1e5f4487e937ec2de6890dd8ee5ba3128a9a28b485044024205158dea470f438f5746092f4705d92e6d37589d585471baaa6e368dc761902480d08a141c61aed3ab3d430a69c834eea1042fd32c503ecf27c59b548ca1722904ea65315f8806c1622e14bae767f49c436b293764df622b5232105c8617a031be2f708253f9fb8ff821804cdfa3a54f01a8fa8b029b86399f1ff94d13fce9216504dfeb374a909b3ef6f8ac6d6323333a72ef857c31e67ac30690e16d53a5e614769c7afe4042cfbb69e46ce60b31f3df206488430a6ad8429e3a1b742b49ed8e7d17abdcadb824c0c52eb8d7d6903347af2e8f955f40fc0bcbef8f0f6352bf6a72c02cef808506cc9d39340e8e8865a55f6d47b1e9d9db86ca7d8;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h3f309fb0ddcd54fb78fd84f394098d24ba83e803280ef8534ad3bb32d2cda45f37b268d541b56a9c53b6359bd87c4654417e5da395293f5336242512c674385fbfc60a036706bd118bf7e086f1c2431b7d8b7c7aee6d69d613fefca1b91753d5dad02ec182e7dd3e76cdecb061a6946959188b1daf5c4aff6b5450ada6d254bf681287a216caa8cca1a03dc52121eacd36c20ec2fb4c82e23deb13f9c64572c3ae984c49f333dd88603505cd65c626d967ce5589f16288853aeb60ac4b025741b85dccb9cb366d5e134a4520913893b28b6b2e9bf45418c602bdeda08c4a7f7351e45792bef19fa042f46e3fb6615857d0e62ae62149cd9671d1fd99bb147f06ae1d3842db94db180e4573204077f682b3b051760414fab817471d175e43cb8ffe6f826379ff479ac1a578aa8f28e19f9831a93257b7e49c7ad6950a39c9baaade70ef11932c4a93aa68c7559adf9bac61a578cf73a9b178fcfd7762603815b90870965868c5797d0570e3f9f44432e0ab75867fff0ea6989c9e00f34dba8ab6390aa2e308146d7dca778baed91b9f0b2086930295376a4f87b3d0c23ca76933001b2ce4631d5c6ed32b82bda506ae0cb827af5377c3f96fd6c3cf837a399007c757adc5d167d641a0d437173cc011243865643eb6a6a8579aac47ad60556c9d47101ca423f9c1fe150042e1e084c61c9cfdc17f1380e50846d27f385a0e7a43e6827e58b4521950d22e113d866ed872d4bfcc925f8e47bca54099038e60d070c824dc13c0cfd856e6f650e4ef31e18d8df1e86aa89e7c569748e93bcb1a303b9280c0aab4f138e6be68808208f0f7e09e5df44520c716d49d310dff3336731e686e60ceb7e085b75c2c73737fa1a36389effa7f603743874f0beae7fd6c624091f4180073b3f87c94824108b8c4295e7b83e62dd2434427b7dc26473746fdf5b87c63f5d6b05670cf33fdc1172ecc9ac4b31a94d7d9ca4c9b7cede153285c4a1d5ef2ce58d33c88d25969a751a6fa7cf41579ce25fea44450ad0d13aaa0b26db17327777ffa2ce7e9e87c1dbf6634470c7c04a3f5b22f030b9c0cdc7ccee3b5c2bd622561bcb6fb74787cf639147c5016a176287614c2735c723cd45e7ce440787bfa46b8d3f3847fcad029e07562f9e04f4e702e9120f1b871b082357b0338e710bca19f5a2e93beac9b8588d7d06cca9018c45b981b1de4a0de454293b276667427ea1d2ef21a4bc267678e9339a4934d90efd8567ff4fb5a23f5e5c837621620fc97bf4f3af39d18d701781a3a05264f093cc0d48a4c7ca56dd66561efccb57f4a10a18967ee570b7147b3259f8826df3d2e2652ca074e3acdafe09c553865cbd940089d42c605ab98ed2852198ee71af5f0d595326f3260234593491dce6a66d2fa7ed9b055d2d17fda6cde9f2abd1815571d7dc13214f49b5bde7d82ccca9961617d72ad71dce1e38c596c43633af1108a0adc5db429e7e77bb75af3327773710d7358dca88cf35b697a3caf199baa41880099cd73dae07ceb9a9403d1a8e3c30d32cd189baa4add7fcaf3f4d00f4fdfd6e85957cc970cd365ec06f1f996434c6587d116aa9ba00843999805924d2570ddfbc8082cc38ea718faa0725be7849cd373b66647780393118ebd6ca480a5c1d0c32aca2517e7d1c2169639cfbfd9ae7a03b5387751b24e7890c6b7aff80079cbe54af40b6656ce6f2a9bfc43e9e53d7630c909263d296e1490615501dbef89f2791cb91fb3bce894a5cd04d474568a5e06059e324fa7f758a7d3b80cc9b44670ff7db24d838c77b943896b4596961ce1dc84fd546827f6644fefdac533541448a6e6ea2c418e2e5fc2bf14f0f9cb71334ce4234c82d57b4752b9b1da229e2e5c8c479715579c8065d73b99ac6641f2ef7f53863063a8d2d26c40e407193e9c6de61f31431a0d9292e7d5d5fce939928ba78b1e10530e9d77d2f8495a4b0ea82927878c2d8d96bd031eba401637e762325d14132d8282a923ca66d9b78d4ef8a42d7ce46e792dbaabe537c285456b31e367e59b043961a4ec83f6d98042207286eb277e726eb27b1d2a65056af4d07631c93c41bb18d0447d31372b5c7709bde4dabd98f46b35d964f98107190dc318c72a5286d6b00e8e3dfad386a077eb0cf23812a27ee63851fae461a6b724627cc053963a1faa0f2ad2185067059cfa3d083d0ce84ca972e236bf7a0fe094fd2f6460593f3a1bdec06ce942f01820f2ddf609fdbd2eb90bab3a1c6978ee142e047d7e4f2f6cb20a8b05a66581f716debb08194fdda90066023e0cdfcc9cbe96faddaa4152b4cc26b40737ae8f127bd0ddb998482dc724acbda490790d902748b26607226cb57bfdfd02ea5e1bd6115f3b0eb05f94821a6d201867981eedb477b169fc3c4211e630fc0287508d1f72f72aadb0503a481c96490424a2d4aeeb4609fd9c987ae56faf15b72a96a81a86383fbeb650358b38077cb5722da01ce81714dcdbb5d069838fcd668df9ee53d67dcd51929bc27532bc2aee89006758fd1ec8980b32eecfcca1feef6cc9f05ed710bed972f1ab80d1a829b041049faa05393d138656ac76575c1009313eb1b201630ed0dfd6fbdb10b953c419d9160b2d36aacbdcbb0a86d1e815bb740d67b421e330817e5b8bef306e37d84bb3bb6673300d52a7dd5dc6556d748b42cd054ef5b4f3ee9975be8083118a8365a4233c70dffe9f0fd45f662148d08ebec7153e06c107cab0a97e9362fd723d048d26be9d1100a63d2d4c3fdf380070c7fb0d16396fddd16131e06434665908ddf995ff59f6985147afce3b3030aac8fc9cb5593e01eeeb93bcb5dc5c6d4aa859f5bc736663a4b396bd0bf89afb560384dc706c5876fa35f511a63fc9f848db53ba56c1;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'hebda79b086165edb5943ef434f6b85d54ac0b33aff1819f7a02055785f0cf1444c3e97c59e70d0c91c2602fd1fdd22d5f4dbd2cf8edef1c6071a78557fce90453ffaf477c04e4d58e829fa7699d8b17990cd422926fff66c58f837e229f21fede28e37dd9352ffce922664989cf47ad4c04e44086de8ba7501e97d6afa76e3942e204353f76e9347f580b329c2f6c059c17989d980ad468319ff8eb14b21d9aab11ca34ead41e75437e72676e95307e6e4224db546449413dc3b902526560db80fd2e0c1cb8cfa8da2b9968d9a465cde1f0d448cf4930126b6ce7a3594766922fe8707ed5c792ea3267bfcf7237c00251380110d0205d88fc279ef7a88147c43e0220eca5199dd2c8676268484c5d0ca76d56965a5db818ee6f3f6b3a3db5da3b1b61ff162bd39c74745d5a6010e38ad50f42526700c297e94e00eccaf49feaa24e2158f11356cae7cdfc9564ebbcd01276b962e56af2fc08d02820c86868b6d7c840fa4014c6ecbd1b2fcc9be5031c97b24c74b9d9dc84b130a595a0d71fd12025d03acfb0bca4ee786d6b7191db8bd861e741a3079409e7eb2018054775c53233116cc5b0a3126d70ba599d09240ff0980de4980fdbcf6ce5ce7b47cfc52b4b84c5aeb12f7de996e330af8595d549d56db65a0757c76f09e8fd38198ae9f81cf484aa4bc8c72239f7f2ede016fd9c468944373dde991f64deee1241faadaea13398e49725f7c41905789749bc226d103ad87e18a79fc166bf2318ff98a816260bf9bc44f7a29c56813a750c4be6eb534208ebdafd0567d50e4f1861a0e9cbcb5e361ee56be2fba1c936bee5bfdde0c3b0b730eb3af9f06490bb802b48552d5438a505b56e3eade80b8a1125635a2b3028be14d53064beb8d3fdbf08d64f2254b66f513434274430ee5ab0565b7c0c259618f277d51b90a55306a5fa3a1a30f6ac71a2f2cdd473b4ca5874b1e8a6c06a014a1b7f383130226dd76f2e912c9c6e56093f721bd16e6e6ee67b0d152c7f4f225bf909f67b677f609c18142b21428ff781d6c691cd59d365017503b9ac8038e3e011e044a35aea9230085203b818a453342fb6cd72f09a9f462bd4a6e6db1842a50bc49125514d973ba5559126e85c6231f5d4641ff627e0f669d9939bff48be0347b59068981651d4065536aa4ade984566270b9c54331632f5bfae19a5b8ef568b13b7bbb2d914033255a86c323ad924dc82392b4fe7ca2fb7fd806598a58def2a204f7ce258c900c94502b73b33184b9da398a0ce087f92fcd836e30ef1bfb6c23ffe853319a661739c9d324608498058f664e8af382ae39c5afb4ade09e85620abb85226f363ec3d804c0efef250bd3cc7b7ea3794fae2c1e429d43407d670b9be2648d6bec0bd1165c67427a584c25aa7c8ac40116aad5ea632ee7c2f7951373655af894949e52fae7191de9c358675ef92dfe7f831eafe057650fe2eaacb3a21d3c45cec20c67abf5146249cd9100ae2d714abcf8be12edd3afb8e4548b763c1a8a504329d6418e8fb1e89e0c98a97d179e9c65fc65442a92bbfe56c43b89015e136aeb00d70063fa3bf288c7416003875987950580967bbd779844841a8351e8fe0a5038512c9adf9825e920fd9a65b2118fdb8e05227138355cada9b9319d9192edb7f83dd88a21182cb2431910d7f17969bf1d5de71f5b9f73dcb2392956bacb2419d1c4e0244e726a7b951d25ca111a962df0a1e35a716e3fb7a148fbd70a2b380c98d736fc17598159ad7511d2bb57beb8e72e8dbaba2c98a032b0a041ec53c96d57d0091ac7fffd442dae8810789e70f1b90d2bd5eca7adcfa8a415cd5eb0911b7ef5c74c830dd443d730ab4c408273e7237d45898ce23b81bd681b97b8f89580744bc256919f53280a975f9da838ed263d9d2c713d5f3e110963fd58537154e63c1401a514f8befa22baad789bd3325c62b7b315eb31eb58fc93d1715fba44b96d918b8e086bfd2a0476f4ab52e81810233bea545da5cd7e139f11f23b7c24e10dd0510028232052d6cc6b6d47461ab646bcb8f96ceec705cb374a580ebde77ca8cffbcc7e386d0f9e74343c5faa4a20a2245cf727f0087f830b151b0bf18905f5198d31aa277c5cd16c0ae8e27b0b3a72f2bbc7c0f1e73158fee9e867183da2609ef0ccec198acfedae95966e9debbd5d7100296b3ca7def8cb988accf677b0da5736e02c39afcae15e922789363dc8b6e220e9b4658431ea95c41b1e36b74ec18db34ad74bf1a14b06fde3482b8f77cdfa0c13f357f72090fae81ed0cc4daedda93ae3e0a600e97725a4478c8c0a53a17d351b14261401bc805e625ab74df47943e6fae0a02147303c3114f3b9571e9de9a9a9dc37da33263047ce91964ef4f08ea746af8c7678fb9026ae4b7f3101b453fb80f8c5db54a3f8b852c1e31d09322ce1063723d61b8cbdbe49c7fb4a56d07516d6004859ac06ab55a542d83d1319a4387c8f02540d6bd84046cc2104af72e7d6eb0fcc8ad026b183da883b9ff47325cc88cdc5405dff71bac775df054c8b74ffc19d730df5f3721bc049eef45d6f4260b19524aea93e06adb6b717993991c320f700bb661b6c553cd6917ac9032d8269638fcd63f96863578e2914217244a9147900fe4cc2cc94e6014a11237111e983c940dbb36b5ee0dfbf8119e7c1026db78fda7c152de22ed10794416ae5b8323275cee90ca97250aa57e0180d52e12f11083f983df0d4825c3eca782c512d0afdff298900229d35d8c93497c9c0008be5a15ca782f166feab56746d22a68103ac2a2d017e04d24ce68370ed77283b8c499f43fe5429c155705f557b89ec2735e416183f8d93e1453fd81edeb055e775452cdfd328f3d71544d4bb0f195c4404421e5e42f0f9;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h6dcadc676e02eab9c288b82e46d45fa09298ff18eff9db22b4989f6c12a536ce59824c160671e0e0270275dc4abb94193c0e088568ef56971c9c7b3b5d037286d5f46a0c47b0e4f2b15cb77a5b1106c8a4aa372645cfde74259cff28f4d60618d11809f8208238787db879eb1e576fe98d1be7f6eb9ef5856ceb0a9f3406ef3e83b979c47909e1e385a5a1173aadd14595560bb559f3a1af0ab8caf38dde8c578025186f837a7dc7b34a264f96e2fb58e92bd64abb196160072e914be1a895079fc057f689caf21a3612cc33bf2113a78807781024c71f605e7eee538ed8aa80e3b70b5559179c566f82ed0ef032c1821851f9a25fce9d166d066f69e854a00a658870100456282ba235bbe952a37650595268f5c08b3f4cfa842db94d49a3119a693c3d3ae7d480c167b377b467b73a6efead991fa86e1ff705d8132a02eeabbafa38036de85387ea8680934a2bf3fa36a3e53a8f8a24f275b5f627e4c7e96475494b56153638bd5aa5c42869c852b041aef7194d68a11bd2f8dc97ee05d837d4f952f90860dfb96f94cb51833ee9b8736bd5b5b4ee00ffc1ab704c56d5ed7260c228a11e04c7c81c9ddeb149a14e01fa52a4d551185bd926640bf35646eff06320072d6ac7243a30b89f330a54fd4da28ada1b36cc21d8161c2c94e54d4aa88bdb446aaa775691fe9c0de528e2b049dc74c44b485101dd437cdcefcfe79e66e8fe912a733f3c5035d9d40807adf82fc2ff1fe823526af158f0b7bb768871c2c18916313a777062d1cc13036cad6f1dfd4866b668fc1dfe270dd4b34b4e98aeb62ca89c2e291221ad0d4ca76135e7e96aa38eb734049aeb07e53d9228fa2df158cb14bf18dab0edae09db466000cdb199a50775bd60ff4df83d908035034e3d778b2e0a8e1d8c452e83d9827b1552fc5625fb310a3b9aebba435d27348ad8f7ba3d9567810c1777d12aa5b0304dd8c12867b45891edab218929a390c44eb2aef139756213613decd360150c59b57fb82954b914ba2cd0fcdd41925528dfe57991ede3ed7d8a794e07a7c9133e8403d949dbe6dce9b02a78b92e5b0ea99ddc0476536fd06e677dc7bd59cd70c1af906476a376c17efefafe359820d280a568fbcc0701ac736a1cde2eff2c3b157345d8b28c9ae642cba6c69d95dc505183263c9c61dd5595bb0c06378b0b05ba2f7731fa18576d8254591552eec87be82fa03a8dbcaec582469fc6664a4adbacb00642b552effee10bcac3339bfbff24b5708c97a969d0aa24ef25b553ce132db766512bf62c4ac2f7e5df08bc68f03787ad0d6678be03522d4f7a92c7d99e3b78573af803f3d82a9876c7f707be498b0bd2a492fcaefa5f4a358e4433be4c544d75f34b94b5787814014523312ac9f199ca3cf9e98d77e62f1e14d46bbc3d56faa3306d82c585407f02c4d6719543106fe9d18570602e09390fdeb42a6699fffddee7736c1e84b24f0dd311dad7c8a3da6d5e30411626a590570f974a936c48227e5f38eff002a78ef83b4ff372b7e47c0575afa8ae177f9913dfa59afcfd532894eee06d6b4c1ecdc6d3a464fece68ae8f9e28452b8f6779732038def9a9bea4a93161d2506e2dcd56b087d66a5356fd48f0eb105b6dc2be1250f45fd1571bdab6ca6062817fce2a2d29755dca8a2de2f2a9c6b04419e3d6151755a89a7c96011bc9a4de8b21e70ae14286aae72a421feb9a8c48726d6c3a49f7384fd81afcb917160d3c3dd83514f0c206b3fc61007088ca309fd3e5c7d55a48e61fca7ef84be2392adb19d0989104041b4746a2331f39ff376417b67a8060bbc0172f70448ce3d1fa150b7c5022432491f019e725372002312e82e7d8b8ea74441d1041695d38903439f851971b8faa47dcffc5f6c1de4110d2b3cbe341f9fa4b55818884baf9d0f016dbfc2fae8c6d6386d66e959a39e620b5d6d26ce5786b4a05c14a66490abff3b1408165afbeca0de62eabac2de5d11fdf1a29077b02e4fbb482fc7685a4349ea0aed94bac395dbd06b5798e85d0c202b89108a568b16e4f7931f6ca469e016953808a5a13ff0b2b97dc8eb69d1f467c60a85c35ca80e7051c0747b83f42e39984d865c96ddaa4c19975aeacb500ef44a0f63ba2ccb94f1a2968f03ed7a9c1b2c636a4280382e914498f5693650c0f51cd8e0a2e1a876ad649c39932083f44554ff13ef6bfd3bffb0544ec0fdd8dc03a6a70cba82908527709056fa4dbb761c25ce8fb03495c8ef570b2d51679dd8365279c34d7652c13d040129ac1c9209b06fd2bfd69bfcdb5a34358fe7625ffa1bc38ca5e66764a3ff3c0d1e05dccc4413dcb6fbaca1c5d21d6cfb8a38aa007942096dff19dd278207fd893c57e3a4c1e9ae79b747937649bbe61b7e2ed32ebce32378f50fe90566aff0d4e7b0272743360e47350c6f9e1c25b1c7b1c75e628074a0ede4796cc86e2ad69aebb6b28350141d2cd83a0e9391eeba30c100366c98c38e7e9e3181e691fa6c2413bc2e21411398f4836e37632369603332d64f422c12c2516003f3b265f61a7275bf3cf166a05d680596679e3dcbd0c09b7b4f96cc1300e182aaf0fff1819d526cc62b3777daba803e8240832c59659f33e8d1fd8294f7436e0fc9fb1b867b716613cf73dad397caffc55cc4af2fac2318b31a57b54d1434b813ff3a767f15255fb0659ee55a4349d3250b22e910e33fb02d921296c6ced4a961506b845ef5c2a4d5a4afa51890387f5682b06d7e12fa8c4262b4e5bb5a8668a7af806d6373777cf484fc28412c73a4cf0420c7a0a2a198e2e250610a9f3a162a2392f004bacbcb482533f4a6750026475e79237d1f2caf4a9affad29b9f368eb0b86f302ca3388f1f5fb7e66314b2483f17e604c41b2d9d3c1b9b6e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h29ad9cc4e7240cab8b3942d2361907d0cc49a1ce21efe9f4a4ebbd633c1e9ea172f2351675bd9bb65ed028ddf1c5d4a1dd71f3a0767bcddb73f4a864d600bb2f991fd07cd373980c3a8a290c44d73ae0aa34fc8e529cb0d2fccb9a11b6ed7f5d00d7773ba8fd88c638e83af717d0ebdb08a24051e837876f573d785e619411b248e35907d3dd701637ac432bef08e808a837469f140ac1e1c7f62e132c6aaf2864ed4065b846e41a9ab67c27122879a85ab27ca707bdd53356c39a4d9d531ca0d1422e286310c91e7387a9229097605700edd9c663b5c4b7affc01c47727afed2dfe3c94d0cd41b4ebf893a00c094a586826835738bfbbcaee06d0040b975c441e5ff62a346cb5a976c5b912a66de7cf2290d7e5f1698c6e4aed54d09f5d29dd92a0ae2803174280f4ace00159919728fa5724112cdc20a5c8d090709f6f3513541dc16cea05be633dbd4efc05f9daaf3ed4ce76863368fc72f2a0b024756bace06eccf713bbfe26d8c9ecf2bfead1140a16f8ff1d7078180310ac5f7393b5cdf1791257b7255d031b757304842e2594e61e97163988bdfb436a0e1567971307304b9b8066eead793ebc193d819dc47e5802fd25ed5ee525476738f155071be928a57f0dd509f3af85cfced198143e38f504533b5b4d1806b74c2e9d44dfcf2b68a0b1175b7ec5e14cb84c24e9c41585b35ecfbd2632c679fa88d074b6bcf3bf0104671277a5372bbcbe5f6a908f7fe342c5b3d80a4d0864e20df0a4e5db7c670e54207017f71057b6d95f3043729dc6d191158e04ca3bf8ac0b7992a80259e05ec7af1dbe226366a12a81a3bc4a071c07ec635e94b6d09fd8ba62726f33f9aa548053540d4b48fe5006612f88e3ff60023eea05bf7fecc3f38579720755f694b98ddd9e3791d725bf742fa85f346756a026d20ea9e1d16f226ff83e78299c26915110f962b5fbc0ff3fadb10dec2127f833a719722970f2eeacc2f5b2e134380322d4d91e8058d44f3acb9622bea6c2e72655594026a2a634285c2a66993412b983f47b95095d738525a1a9b3a9ac0c9d2bdd3a58b56ee510683bc656ad1ed3a8519325a583e8faf7820bc31453c661ac19f17f4973290c42ecc957db5a5a2f0d44e579c9963f00b49209da39b928def8845c94218819dcdb58d80a438511d902d6bb68cc389570306df48be60b4f13e7f980fa30963d3e8c83efd9246872e73f9fe56769d90935f051a88ba23418b321034383594f9c2e6a7dafc1f31e8303036ad302dc9690a1366adb94ec5e39b7d685a6204f7cba0916b7d1995a711b7eb328a9b96e7f286eda73a3760db5781b60e57dc9ed0b78350f44bb20b1bab34e0a2d7122e558646a20506e3e5887ad66ac6cb0c513813c1c4691dc4eabb8a2fdd464e369c5f033f7fdb232e62b4976c1ccaf83a1934ec2e760a8c0f80775cf4235495d6bad51501df02677c7ce32245b8b46a4248d773b0a9371e08a143a521758b612e5a68f552f99d47aaf34348598419b20519fc524eec9a55258f9d975033557298ffc0d7a76b74a43257bf4e11636490d6abb5daaca9ab6b8a807b3dcb766a592948bb88c244cebac1ab3e7ac9dc77a5912e5444cf62152733f7a4372bc76a859888d72090f283edec08abd78ab3d6f797038d24d1c04acf0cd95a78d9114f3ffa1387f9898de6f7c1ea65032992b08c1c73180f892841411988a1a46694f87cafefbdec761013515eb23e81c100c42d6d620dacb4d0d744eea763297564273c684f0648b72153d4907210557751308dd3c2cd01d4045d3301a89c048970f319ebdf6afdd9044c7ee9adfff5509761ad0a980f2b2e16655a749a3086abc9309df9c72020e6144518470f32a02dda14d4b9c6737b8f2df6c9479b27263991df4bb9fda5c9b52cf4d2fe8994e0bdf92c04c8a2fc59d825a97d1918e06e96698f6141429049d46d38beeb13bc8cc37a82e5ace7dfa1afb2ce4017b5660c31fb1d880a25aaf6bcb01fd8b393a9d00c3cdea25d10f6254269210bca1b8963452f623135202a387253fc72bcb5e99dfff56c8bd1e22243956ca78df90eefc02571c62c4a5916c51698801b647b3fb7ffe338327bf4f47da1e5b1991eaa0d846153fc77a24a642559b61a91fa563236114e5b6dfa6fda215fc9cd53f462e0c15a5deba1ee938c8f1f17978678aa39b81ddb10f916e7591f8162a714ea944bf2567c0ad946e4493e270dbd63b873ee1381964a5f5e2ac76d91f89e247c3dc1705138e507687d624e6e2bf7f43911b3d230ffb17e17af91a34d3e2d96e1b8d912279c27b9ac9411a9528312d8bbbaf901e9d5355ed483132e5045380b65e78f1bd5b6c1fed38ba79c6416de8ea00f3220f332d45bb640e742565830075b576a6b18ea12a808cabc8d778bdbf7b40150b6b2f292757b56cd2bd9f896b56599f93e8def9e1cb8492a41b24f81e70465abf5d309a8bcffe68df68e3612b2c173fed3ff71aa5072645c4a213632b79d8fc8d254def777cff4ba392238641790615c6024495aa2366db89a5b7b8e279ad46e2e7fb7753dcb7e08f87bdf62a5a8f198b5ac9f5f579634a5909257de8474cfce5617043b3fc44b5183e4bcaf08a7f1aabefcff855d7468bebacbc86f3d563fe0c61feee2e2b9dcb4cf0e1905ef713d54f53f20e791f3648aad0af6125f61f93b1c4a3ca61a68f595bc9c129cdd7baffa3956c6934a98c52801150348877f18827d5ac2bc7dfedc826c2347e79f9dcdb4fba09f028433974bb7b3b73acf8c137cc5d3de8f3babb136694002b6a057a09769ae253e4acd506be39aee152439b18598c7038117a1f30c7bbb9b77011ee52e1e8f0d0298df2599f89468c61cdf36ff38788fd6fa326ed3cbc2b563e21d84a938d9f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h6fc77c5a3b960ddf4011a8bde3658fe09891e81d49cce5daa910d3f49108a7829325846a251e02017ce0ca133bbf43c4a9e92f76a831342ef6a10783a0222eb5c5301ee10ef480f5fbda9523ddb58410b745eaa5421bf55197ca2f04fcedbf8d724779d0122d5a22d72c69a56cca4ebdf490b37c239018570f16ddb6d5be94779148ab7db74fa67cfdc3cc2072cd349ab43c3d69226c818c5b6b6c2c67f12041a1a0f999fdbc5628dc9f162c24a772922ea2a38ce7014701027aaa942d35eacd46b1a9d5b2f1dd5b165f833ee7492ed403f0bb0ce14e7ef8cadf2cbfcb2124ec70f2bf3a32883204ec7bd5d9dece8b730251d560c7021e08793d097ab8bd4ef6bce47ad8527ce3d38d09eddcf1ce3325bcf79012fe22ff57badff1abf68b3497138e26e6921c56d06cc0ccda28e96766d269b04f9ab164ef628c0f91317dbd8b63d8a52f1b53646919680c86daf2e6a27543805f763d596c5a5b969ad3c886dfe481289eaf3698cd9f1a9b7d87f85225c839f943aeaefb5bdf8773fce464435bd0ceff64bddd3dfeb1a67606f162ba672352a82a989503a197848a298108681ae02969bd893428c7849eabb302f181dcf32c85c408cddc280500c14036e6c1a317c75ab4bb9234ac8fcf0a15fa4d6fbb0e5ec5a3642f5c60ebab3c53600b62e41baae0a978cb78cd0fccff19003958f18f8b2bdaedebcb9bcdabad709c9f742adb2c19633eb69bd27ad97e30c9e8a73eb51be46d1d97c593ef26c81a31ce6b4712c421c000c56f62d8bca17c57f0793b544679343cbdb8a3ab2af5c5c3524012cabe9a05b2a30f965771eaa592bfe2c26a1e2200eeb23813bd56d62bbfcf6e786500bca1b064e7be60787b21baadeb239e3eec676742da55d530e7ab783516b504eb896c44644aee8f4b1fb40cfba6184f23ae32ea2f843ec7b9f0c9939ef3a8cb3dd2283a56fe6f346e8166bc2d59d7697e152b5f13ac10226f472b82b937c8649e3b6c1e82035dd1fa8b24e464974ec025d16c755488a3719b8c07d4fb7138f07eb6b656e8fa98cdda952750d330c3505b24525a8cbfa921929ec372f3647d41c8c13aab5f9ed38ffede2ecdd1a69593dbc4ff8b57f088c7074d4d38fa3bcb08e8c1067651f72823e0138c05daa2642c80017d007e51b416f7cb1555a678b95fa844bb65c53afa9e2758506d6cb4f666fa13693796822dd9a09143a3acfe30311bfbfb756f965b74c908c236fcf4438acde1e87a07a2519bee7aedc54443035feda4010b7ccf65aa65f7585e0de4270a2615f203e96a9a76965c642afadcd25cde7e8feafb771110a3ed5de397368bfdcc7a9953fe9e20ee42e0a838484798e2b515a93e7c8903b9eddb0dc65cf516f1773efcaa4ae188753a8fe5fea49345a7fe2cc2c5470f0fbd77d4ec1f92f1827bff08b84b97354e6f12dbfef118b1ab74a7c0f22002aacadd593a19af0b257389d8902092f4c87180c6bf803ce3622dcc683d680bbf23b36f15f2b669a2257c956dbf5a81bdbba4bd9ccb42fce580e428a1d80bd72ddad1b85548d7f0510df530721de3cdd50b50aa7ad496acdd6aaf0f5a08b63a9053fcc37ce49c49caeac70f7f6bfbf2024d6432bc4fc470a8b60ca3c86011df92aaef2de75e0c0226b3fc870cdfbc2f890492317a70a2087b18461a59b0ae87f3f69324d597bb17e5b76ee9c5925c4b2a08cda27cddc1cf6d4eb080a2188adea111fa49eb075fff522515dc5120fc9828fd8948a006ebfbb77b7df2a902227899620bec25617f0669af21b43362bb92a945b3d7b43414ebcf073fd9dbf7eea89634a7c2c29c18e44915e57331d21e5596e167803459df847180d3211465af481abf2781a2ecaaa82a0e1b827d14d6c94fb8bfbe0bcf5f0116bfdb5fdf966be93052c9b9e995dedb824ffdafae9392b6dd6838b7a1b71f5dc81f50fb3aebbca115aeee1ed01ff8f54ac111adce7540700490f50412a8356e086690f7cc3f5a9b55008243aaf1af7f4d48a2d654387d5c032366729e975b5aec4367ad390a9019cb1305ce68ea0e10481454aa808c7d411936e15803f6317722b4d049cb25e3b3177f3946c63229d8e8b7d55f75bbc9f7e25e2fa785c2d39a4e395b1afaeea50cf0098f4c8af0453f2d0822b6dea37014accb7b5624160c8dfa8c15e5ca39835a65d696cfde34724d934a013872a6f6d8ebe74b98cef0101d0b017e421b9beedf318a04084adbe32b41689305e25c7951c3c6313a5f5dceb6eff2179210e41babbd8a9ace333ec2900cba1bac20f972d5dbdb4f148acbd20e7945c7af0735f30e1c4606b247f56770bd6c691b3755ca2b36224031d5225ed498c7cdf612dbcf868ff5a76179d0a36ee2443e57751605ab4218137212cb5eefdf01e50763a634273316f2b1c8a4f9c58f6963b1396b3231dcd2004fdac54b37e8aae5026f8291d5efc4e3af58b512e89ed728fecd6fd6389e898b4153ebadd75bea9125247d2237ac3df0c00941389b26f6b1ac419fda109437e797e4aca71cb23f9a3021fb49dbdd04883c352b85b9f54c832ecfcd1595ca409373388daf65739aef804c855f489f8e28b41e028aa266dbbca55e5ec1f3a681d4874a65b9de191b203175ad75407ea98af3d63e92daa23aaac0c3bce0d56323289c665aa864ccb8d7780b6e57f7dbb3ddaafcf9499c9870d0597353e652ee42d8c71d41ffc3abb20f216a83d7879cbedb865cc3603ba214dcf3b8a30be690a306daafa8836fca03e768f9ff8e9619155e4c61d9e561d0800bba6d5723a60b23d11570763720ad758bbf401ad2b6e2ec639add934a83efc2200df4f61d3e030a7ec654618434f2ffd8f66398a39ef1cf581840fe7e32e11d90e513c065336cb38ab563ff522a001b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h60ccdb6dc1fb3974d8c04391433d1b81a7e7a10c3c4de850e5bb581f213c2f4e81f7c0084fefebcd219685569e82a099a41e5866abe574f2fdc19f4336040dad105384c0d32cf9d446b5db6eddc98bc75c11bb071d76a8c25af8496eeed759c86e950076e81269987b3148617e30d024b51a62621753d30c203ed78b5132c7af372914b060f5e1964225859fe007f4ea6b3d86ce3a686427c35317070f69d3d9934fbba3b68d6b4a8032999f46dfa7e59942a6ae83fd5c72cf2af6f84e9f63641bfa8b0f17f7aa8c43a3aafc113431f36970943dbb6ceeb5e795e5218d5308028049925da4895d77856cd05dc4f934a712cc1abd34f440dc1855a373f9866599f01492ad26f76fd34dd352b033551cdd283904cb72a5b99ac7d24bec59c8b5d75f2ff9aa458a119fa7da4e2c1493c4b35e621aae841e1092f4aafe4053521a1a9bb639412616fa50095dd76b312d2ead6ef144d60cb33f82a948bde06f4c63194d4370ad839a3bdfce75c150203e3f234d686603d6652138fab42269349b6281bb9fd33cb7f51d25660d860bef3aa91845df70d875a77eebb36aa4687c42391a7e1076a2d78a71c2b82794f8e2607775586e8bfd4d21dca279e822d3570ee5caa86f78c3fc707cb794038229f4745c871ee0a554ca615e1a7e5483be77dc0821eefedfa64de912f0545baec335db7a49b16a041bb09d921bc4d4d7f8ae43a02cd67d39708ffffd0b3596493b1b7321ce419e0bf3f8d0452b8040ec1d4a806285e881a9e4ead8c550afc842990a2abe4b4a4cf450a969f03845e2b40094578c817898f6bf4c4fb4f6ca1f5d7fd1a6449206f5431d6a3e9e8aa63eb5aabaa8b077613e6c3484f80d8173c53eab4e8317659c2d52e680ee3142a706660c94c1001d21c41d50eaf05fda70f8db72b74c8d2020a7292900fe6d2951ed7bddd2cd62ae7a618151f6ee33257d8cb89ce22d6fdfcaaf3755cdd68e0026758209c0b1086fd7ab839b7eeed60dbecffe2169de6d61f7b3754e6c55ff04d1b54e2b9cb223db2fac42648ee7043d9a3d8fa246c2edd9183d16afa81d815f1a291f165807be4714fba8780117b2fe6d32827e3fd5478c0c4aea530a6c9feb56d92490c62cd0187cca933bd5072427473ad90942c6f5799722b32baa087254c790bbe0216d90a827b52df8effc81472cc50e860a2c8bd586f81974851e7f73214e0a03a22654756abeee83fb36e2b0b92427302003ead466c13ff7f8f5466c21d735b57d57865aa604f52f4cc93727b665fc750ab6b5e6166e6d1e166e04efae2f58866651e0536fa2203141dbff9b218c65d095070ee62e38d9f181810b2e77aa4b0f7d543586a8d7eb47b4c421085872b7f56f6cbebfc612365e28a5d3662b5dc8dbd5d49c9a0c50a0a59d9e7b66146988bf61f4cad4d11115c059b29d536c9e4c1b5c63a699b1eee08adf5a9fbc1b84dc06f47e5c710a70c4064f7ec14892ba608adbecc9cbed5aab68adf79b0ff721b40563f79dd310b2011bc7e630bd735dee2e973234aadf293624dc031a231359e57f45b902d1650d38f9beeb1ebcf745d02e7ba950072c317f3cc3bb3293294e388163d109b74fa35e5f377d8227bce4f76ee278d6c4b3a364c62e88ac2a0b38e6e5651b774144c056af655dcd0ec06308c5b4d1f29d7352af96fea9b4f72b26c61072b04f251def55a108d2c72e1c816f455a58e5770ebf7e485a840fc0a036363acccd8cb4efa4533842748c03b1585e32399411908104476125ff8a16a47985b0f7071b9efad46ffc7c844621d0b035f4d7948ae15e81446cf5449e91f79aac9964ac17399e19977bf1c0226b062ce3ff79252ebfe3e30f508d7bbadf088574c93ce57045b4145fb1928d81a7685bd4e11b3b6f2c834321c09627f8c8ae9deda7c014a9a4064a543c281368edc9d30c8786b30846885eff375a1582b333e83d8b9e124ab6cab64f3c81b4951d02b8490cf277b8356af9ff00984fcb09139242482d5593ab69a8fbe8ceff35b7e961b10c74d086472cf88635a88a67bd1578572012118d8bc739404faf97a498c92891b0d3cc3b5a6431345055e6109825f83f19862819e87efdb1c59f5e173db22c37c10b897cf56478226782420e6870632e8deab085febac0af03f0cc9430ffc25f1324249dc135a527795255219fe4a90891fc81ccbe4810e89a163b4bb3a0f933ce254e04baafd10c332e1764ae29b629ca473fc0fecd7e13c51c041b25c480bf260a817c6c6d4417d4bfa43fe9785836af0343de555d91f1d3e0317febe46657ca88bd1fe3587dbb60e28de677be19a793df84ff7a729706d229c17eb961fdfea8c6f7380c7be1ce6e6d93e63e6f6aa85340dc562bbe4f640e54d097784c4e4d86dca7672203677a5a9beff2d7e711bf907914179eab702500db305ec08af9b876e08b999261855ad112d536bccd20ffc9f1804b5340b2a52620bfc439d94deb2011fa8fe13bc49e6460f5b9c748b1579a7c4f8b4e2d864de0c121448f2a40075a54c42f2682c670deb0a21b6107a315aa57b2b80a8b1002456c1649b84441652e49bccdee54725297cfd4f03ecd9ed80a155666f1fe354d560054e3c8ce7a9593c0c273d1d4b28eebb5cedf12788cc191888d0b2b933eec3636ad6339ce429d8c98fe53bffb542580ce369927a680a048825fd514b7cc1e07ac76c4658388f2d8ffc7f03f2161557c4a8bf4dc907210c9d8aeeb552b06c4c6dfbf19389149d229999abe09681dd5a5f57239548fedc579c3028f117338e0de48615aac501e2d228aa2cf3370698afa5f4b5fd65b3b950786c1fbf8fed2af08984e6356da893e110e4a504c8ba87a2a20ff16a78d63890d086fc733d19530e890cf5bd4b4b91bdc68098ccd;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h2d6ed6716d7c99532071a62ce7d47930ec0662d4d339c5dad7243cf6f94945419423a065aca086f4ef29519fe841a001c64ddd8d203751d15350d4d65b33decc416a59f61cc47d441e7aaab74b9f552b53b9ff0cef13a53d71db0a474bec0b5d137214f1ff2a9cd3de1034c2d05f9412ff50c0fff3cf2d9c3883fcbd0a7da9bc0cd4bc11d57779726a50554a156406ee0d249676abc3c54404d6250e1d65d3fdfa3c21ccbc5be0164c5464ee94c05df5b102e958679635e5f2f312ebced1fecadb380211b4ca100faf752af68480f06637852d48e3f65df92e5c4fba5b0fb01fd80932365060832c3f3d09e51e90f8518b7cde2b10fe7fb31195a2d9ead4e382c84c0f5831c43cf0c4c77a88f5835ccfb01e06066fe6e625b63884acdc021afdaa634c566f44264b28edd64a1d34a2e2ba8f4f70b5bf2e285eb5e2d0835ed129f475973ec985d0140df8f2a76b9f73a890b1e75a0a75c0d42877156b3d2396bba46ecf95c93d07e6531773cd5d8bcfaed0144ddd7168f42cf8e2bbe8cc304c7ce5619149ac2323ad0ef677841b6daca0acde4f62f22dcf98a415fbec21f35ea9e77d80aa98cf92dbe8711faf4313ac41518f69f8496c8d317e0ace586ca853dadc237cd45fc32ac40719f36f151ff0fae6af627fc4e021c97b17766c11ca001fc5f70663d5c99b49b0167cc1b1d39eca4848f3facad7f30dd0e243e407cf0228d40e910afa2ffa424b19708be9d5f5bb42b501070b324336167363881e08c826ed538439d2230bfddc74098cfbab79dd316d6b200aefa37b2af78e4e2a41178091e262fec750948202277d9a1d031228d770b604ace433b9f1a05f110add4f3c97aff2fce318922dbe13fdc18f6557cab523374f60066a9a54d424dc8764d5bd5470be2ab816889c844b980aee7ed227f53691beecf0528ed938088b12af95f4cbf910e1ed725ef91b56354583b0290fdb12f215fd88f24c520198a6266470c692e026f8be673ff9e19fe97fbb5c481b63001802a4b9e5506467b15947c31c3441d8d5b8f78f73c554d62d2ebfaa87f3a79195bee422f89a7a207f0ee501a1f4a7d9eea074a20259aefb323c041e9b964d531c374da561e6ec64093258eecb8bce529989fcb024578480780d22c686360ec75d2d2066e9c340f70d13ccfb4e09d7f8ed19933bee8963f000aae24aa7400468f0a3c73dea2eb1efb551f975a29833c0b2472a97f01c6a0de0c0dce1ff20d20341c954ae3a1e792281830bb5a605991df3e5217b1ff713e53478beea39f831bd7624050b0c80188fc0487c521d30c83eb08af9d3a796857b898321751f175ade7f0a09f6b3b4145d3fa0d00b4339b4f8b0bf80692fd73403097288a4adc5914ae1d5e28bddfe2eb728014fe8b52aab2fbd0f53d4f9d2278bc3fdd420e6599ee77416f43bab4dcd041f24e33b4bfd04f94fced828702664c725861a22e4b1a65105db6ab1171b5d6b4330195c7a2bb47a7bcc71a56ad8956e0364f877e5b5fe104fb46c95cdda379c8e7e024a81e5437c0c70a737a246844f4dc8e2b316b388bdbb12c34a0622758f1152f60f2f234e0c10640bd0390f8397b6771f7b05673fc9b2bda96d4ee68035cc24358019aecef732e0b7d93d2c983b18181981118445d3cf66bd79b9eecb729ac171c78037a38a316ffed599ce8c114797dcd541485a7a424cb1f17f03fa5e075ac340b10dc628d1e118eeeabf471f762f0e30fbf4ec0059c4bf5e380e3fe2c2d159efe16876603c1db3ceff6ebba5c605b1f85d0ce0c0c655787a25af57582a4970a4f50463ab2831610ca396432df24eab63c2468132d8cdb1da31e81b665d37e53248facf164424c67756ba75d25138ac00891f581c9f790b51bac4dc88ce7ab12a8baa064f2304477724c84d260c0e338d1d426768181ee234041f3b38bc3911389b532ed54c05956372df32334b8c005d9a18fa5c746192ce1a8bc85b24913b2ff022c7932ad726f844baf9667ef226697720616a8ae288b0425300fbf99b502cb4c9be56c9c699ee893e8d739888c6dcffd6e2b19b8e8b82dabf0e2ade7e126800173a4f6074a908b76f2c8a6a926f64c3ecef11d6470e18ec6dfc330c09279e5712bc1dd12ddc97a30f3f0a1a581c356f82e9310c9ae9ccaf0059705023c0c158c1cc24b56da6907510aec4fa37640789108570f2499274627f2ff1c96ba88ce3d2cf7a5e0d5dc631140e6495bce67038165e4ee3940630b587529fc903e66e0d8048e39368f5f04200e893bcc2d945f7bcc5986514f6b537aa631c029300c3a9f7406c1aaa14ba7048e95208fcda24cda0942284f31be42ce8e112b737cdca85e6ead7924acc53d34293416dfe04bb2b845ec822099e75bb654644a2476bc1220d108ba1188ed758875d51d6d1015bc69fe85c3e9f6a265bda30a5180db6ddc7ab929db795cacd567bd30c38ebfa5281ef5a414806c9990008dd597ea90f6652a0a29a23864f2d39eb91186ef0991909104af36d5416fac924b2ceae1a6e2b254610ed70d7a88c26a121246b4de2d500df6707b9716a4cfdd72de876480171fc8d2b338858d35204e3697ad17f3a561a8d8bbbfee6209a842c3a6fcd0b7b8fba6b7ab34e1190d8cc88a710d69d67037f6f995a092dfa0e958bcf00fba2361a373e0f3abf3e77e4367c383d987aa4d5fcd43665db15b8632060a7457e75fb9aafb1e3750119417bb1ce7b45a98b9fa319d7302a474828e22fa5970a5799abd81dd380f40c1f6b5b811905cf4aa56e2636cc3b4d53de0b6be60c8fccab90b360752e17e6714adc4ac4c1f1bdfa879691044fc60fd1dc7dcdea57d597e5932e5ab3c2284b7f9c3663745bde6f5861ffc2fadf73499cdd5a096d7ea01365bd76fa58e7;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h9efc5450851bde017b6fdfb23571cabbe8cef49b8ede27aa1ddb0e7778bde446e48d5abc5f8a09055fd5593db02dafcd9c8d1e9ca1e4a9cf65c5f36e07a0e2c523cda8a697157f98f7c5445bc3d375099e891cf7e54bf9864992416f536a5d52c5d77fa75510d5080dd4be60273d36d5a7279057d030d0be6730b1f1fe4b504938ea3d7441dd46e4700a66a3985e76b8b9cd68db79b05dfe38d2f20465ff094e8229c28a5f2766d4f088b4b771d74f45138195fd4c917657d61e732d9a19fd3996358c872ab3e3442971aa930ca8736fba8ab8d4a995514e332ab340275f6391f767e46244bd2e86df855ccba3ba13efab545d306eebd55fcf2f2cf0a280508a05c7c49bd4109ac447d9f26ed6c9f34bdaa5f6297fe45a533d9a1400be20db527b7a7061940377d007f5b47233933627abc561cda3974b025f9bd1c28f6cce152e72e4dffa3559c8e89ea2789b95210ec383e17456e9408efa03c0febbcc62ee96fd91f081f202d090ab11a6c57739a6d431422f4a3b8eff5831ef5718c7c7a7102395b46e296f6d591b3bc5e97aaececb4b0aa7ec4552f699a46f99b590b22d6d00760af9ecf20538d4c63b6ec39caed734b07f8c22e2f7cfbb1da341c039aafd75697c60b5c4873a3b5874181f5dfb7fdbeb87433833a044c2ebbadb6b22dad8a983889eba22aa3367956718802bb73dff73792a2f162b56c4a79570531189630e6283bd62cc0519bdc7b3b361232052b096f4d771282e8ecac35e1552f0ee3de70ecbdedc500e5b74dbc9734e841611f330fdf1639f15e117fb9ce941bb6178d38590d987951cc4744898eb2b64c7746f174558e70d52a979c6cbea9209fdcc068da367b9556e558b02653a222b361ba45bf3a94e997ab94aa6f25b77412636abed56e58606b855dcbaf01c85bf71367d80e1c74eb930abfddca95d080cda2a7fc100e5b308595aec7296abfb09ef2e2f994d61056489bedab1e70f8c2f17d620f2720ad1f903812e2cb49de4e9b4b824208e9ce8f995f9e5a21a763c811afa71e99d355bf0cb6873569f4ba10c217555284ac69d205dbc1decf15d05de0c23a73d812479b9e709ce92c367714c23f573702c09fb5b2386d5cdc8ef57dcb050327b0c8872bdbcbbab8023d35c3572d90b990ecd851ff9d0d072613d25d483e3650f427f011aa9565e3ccccb3e0dacdcf66774c3f0bafce51fa42fc333620eb44e3a0742b2c766444c243f7f245301dea68e2ae909335959d97f44ce23c56ec3767644fbe895000a4e2d10905566fcc43dc38a18f51e8933c6aa5f3e7187cc5ee9f25b65f6e337c9bad4e31fe9f13063397e62d6fc43c2e5ddb68e39b3dfa2bcbdd0862be2e9161212f7aeae988c244f6d893615d0d8761be327e82a5105b433970b56da3178b92d524feac84e94941817b50b5b14d7348abf59efabb986a6fcf8663a5d6b82249d7a88998a97327b3416cc6cbd1aa5ded0edd3dc593c07293a0bc7687a9138e73d391daa866a83c218232f5853c009bacf24401f43617eb8e92d6932cc96c90740db48074c3b036c0654c9291441ea29ec3f725d0ff6a4f02929486e5fe0b5bdafb57bcc8c17ecc648890459eb038ceaa4cf1209e41f73618b2cd03de4fcc068e77c366879cc1fafba05634ca7bcb5b582b92a85df5b659abf0a8b7fcbbad357c50ab252e3c7b467ce7fff85caede9df1c979973a227ac9140bda4bbd4fc900ef0ac6638d7f021f6760853cbc119f5cd178bd4d9fb4a5397ef02535cc26d5db28027e9e3b6e7f1e2a224f11fac6916dcca3be2268572c1e50e36361fb234ab72453cff52962d38ea6e5ee686074977c9050c5f528258bb0bf6480c1f18acf6be37f9da2cfb201964630a68c3416b244429972435aa755fa292e59a6d402729e68ffbf3569912d075e1cf690801cde80672fedcabea9ba9c76809edfcd2e8273f7c2db80c76a808b87bec939c3f68e2781d64c16e27b053afb64b600270a7520df7540f88919c314a4dd6f57386c894783aff0aca73171078a31a9e07416b734016d588c1048cecf7322f0230eba39e10cb699ba829c39ded001d1c4e4ceb504b90e8172c02f32a3177b6108a1bcea65fc8ee76e3f76191f7199e5abb759512bef679534f7c453c7bcb1ac8356b4bdef6d8eb4b0a9f3bfd56402913e09acc65c41bb57c989e2b92f0253366052da363d592c0d49b4ff84863bf031b3bf8e7548a1bbc339cc72df4d05731c1b3edaa8e80de12cc5e4adc2a5d23c4d7d8b0c64cb266a49d76ccf0aff2dcaa3a5d0686e12f99fe82ff08010d9dbdd3d08ec6d53fd436b363cfe326966b5edc0b65748dcfbb5a92cb749091777122b848aa57d7ae6153074666bf48fc326c96acaf216c47c300ea7dcf5e7f2bc857baea376829172db30a255edff8ed02af9b7f50b29ca9f1d5539de585bda671d8d6a25fd5e7a5877721512561a239439c7da5314154ee6822b48252ebb46b370d984b8e0a0239db36823f634997e0181fa6ba389490e66ae2d21b693eb1c88f3ed85588a6f7a780ef41f071b297b4c47e95ed43bcb846dfe1cfd8430f8e2000883a9f51c257d0e5bfe5db9451be0e5c766c17376ea6beb420d3a1504291cd33bcfa4ba864d8009dd09a2d182c22f6229725e6c15499683da8550646a2784575af3a4ba09d62b3e6ff17f6996b16cd8b05f2916b332e32f15ec1678e1c3dfd14e9095458ab4eab347e828c62a5d679038b7cfb45911b72c41a29faeb91c198fe1d9763b42caa8ac434b6159471ea1a2a70dced0ab3595dad40b6e2fad5a68a94ced0f5dfb846a13eddcf71da135dab611ac84ab72737ff7c2eb3bcaada6529ee1f25c4c0db89f193d21ab1b275fc8a3b89589083a85508f4268a75769139d45b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'he967a9b1853525814cfed005759a6a5e0c67ef5b62c0a10656bfedf9a143ad5cb99d711eae3de8fe2a77bb46f02f7b3f0080f8b6eaf3f958a4998668836415b1ffacf67a72d7213acb36e126e6fe59e0a603ee18dda5d8eab0cc465ac0fc135dc7acfc055cbd74d56f4b36f09c5fedd33eb7cf23c7f4f4128ff907e28a99d42e58de2cfd4589198eed0cdbe3138c7a47bf44f30109f033211cd596963fdec2de967d73cc5be5128df5d7ad092085ddb83c910ccc15b21021dc2a1ba37d58b4fda80adf42b1a092fb37bf2a3fe6d443db421fbc0cc935a802310242b4892b9841d6982d4632c88fb91450d006858e900563285143789e21b7d667f49609b1cfbda13acbbcd009e7597ed813484f48918b9f27f840bb8019521693ef0c5fe3d9fa339ddf97467944fc54cec616dbbe228fd21c5afca0c542eb6d83c8cde17245b81cd919a2a7732336b5a0c994ab1fbb7ec587fc4618152464e75bc73d2ab24d6bf4cad28e61f0d5baf58f2ec63641bb51436ab11c54ff1e53cc02a25aac7dcecd5773a053ebd9ff6d9b168df7a6494c8a24ef52731c3bc689a37a333c524f6d5f7da42ec474a3c954b610745bc30625e1669895cb6b55c684e293d026fd9be96b9d640414635b56a85907b911afec88e44022a4ba66d567f66dd16add958c864f72e62342efc9d793276f736b5804b2a00d90c7e2a3e1ac2edb073872d7fa6625f6bfdbd5a071ce5bcc0389b19d686c9443fea0d2e0833338d0fb9abbe9f15563b466721afafba1dd2dfe332185ee5ff5be4e7134317442fa9a1fe3385730de28f4430eeadb0c2850a55adf9f67aff01e6232c8f69cd228a4784f4c3ee8a5f736baff53a4a838c66af75209b3e1b17ded1fc958efd43c18545643dc67ec2aeb1ae9393e2455167cd872cc09966859351a632380758a06e1378cec9208dd778613928d4c54bda99edd1d526cdabce1d393b273326beae51b0ff6e0981507b1e97ed504379c1ceabb963b870ec75c8adaf69fcb12d0286ffbbc8022934f8c2c609d8ca4c79b5827d72329f2a720ac33eb2cbf4dcad7f1690514c3b4b950546a473a29d0b183b582d5abb7550162e59a708e636370c36b32f43da20ba19086ca2e4d39e3d2749405a922945df3a29c84c41e079166ed73d08bb97cbaa03dafb17eb0861ce25de235e159afe3a6fab0af1490ab04bc4b0720b9751736fff88f0c30a5761b62edef569e51b27b2a40cf4660d1623a93299300cc91b2bb2aee8ebea883d2cac1be06d559146af7c16d73d5cc9e0f2d8555216469788541bcb88532c7f79036a8e16246ab62226a9b151badc542dba5e594fc7aededbf5282db52622ac2635272d10891428a8cfe9570b21c77c4a8d91263f7c983d8b08368701c97db99bb7726b1183585e9637455251484b8af7e52faab25ebfae46a10922971916c921429a545795e29a503eaec5ac5ce55a0bda0cf39d6fb194437e61f009bff3690b7da313c03ba58c7faf93ff3ecdb3fc8053eecd8ee8cc1052bc88cb55b27ef292081d48844584a66962bc28efb209402a4ff403effec490618b4354ddaaf5bd7c070e1df3e8ecbac826983862f83a1dd47d6b5ab0aa1dc646a324622ed64fd0176e2e8f112995fcce140167d4eae4d75fd4c769f7ed86ab028428da86f6bbd9661c1f0bcc6684e805ade64d97464f092c200e1c4daca7d82084f2e8259e9b31c19ff7d983a5a3f566fe0dce68a56b3400a1e1a30c40069f232ac9f49b563a94a2c887d4c7a572481ce07151769ad745242dc43f0eba12dfec0c5ce6030f9771b90d7cfc28b15e2b02aef338454383dda93e63651cec079975bcda7c7d1704c65d654f18445987eccbc1b43a0906b963024536f0476d3ccb7f3fe266fc484e6b5848d6fd8c8f83d8fd442ae9e3c9104210629bddaa813f96b37527d67acc0042177ecf1c08fb157b3e43736bd3c3d91ffb735e9699a0811b41ec47829c4646a383857d973886f2fed2190f686775639b19079862883e6a083e5cefc74745f997138663b27faa140fdca805bac77aad647a943cc16e1a8530332f21634597b8eae9e87316b7d9eeee868f139df51029993699e24289f8a7d74cdd9e7ecbd82003ee0fb6ad22d008a78a7461f56766db26ffe19882371e5e965b94ac3c366f69e24b2f5f353e5a6e7a1e63fac36133f262ed7347ea201bafd7248d9e2751c1c07000e0c6c03b62d1703f284fd5734b081d2fa0289dad98bacd171653247b8a4c4d68bdff1c1cb36241a42964ea3f55ca62f8dfc272e2c73bb717da7fd504b90849cb8802f6433b46c34f751c7e1a49c78e760da2c687f118cdcabd2d5dd0fbec4a7d4206d0825facbb4f69649b2a846eb5c2ced1395b804639745da3e782b418f690211cd1eadffbfa1b23f134ca5df10945fb620ead112512f1905a9a20620b9fc99c16c8dccf2615f55a58c433a9708916a628f901e75578398d9dddd2042fe7953c51b73143085de0f90721d0fbf23a2f230628da33d8129248a3228adaccb717660f6460ca6c22ca95b3177f556bea5dc5087dbe5eeb23f3dc97d77aef16e1611859f175fcd87962411786df6faa25b44552283e60637f36c7b6dafba94f31d7c86531820982f0642cb0b9843dff9c866f55b393ab2d23fe876b1c3c63847f7fb4a18aea97930df88cc94ccc3eee68316a1920b348ddd4584870b5427e25d423b85a62a0cccca3f79065d03ec8efa2863346efe4d7d56b226cf8bf31c743dad8c0bc796fe21b1daf086e3f9885d7ab859b2ac1e03255033e6ef913feb79df0c2aca2cba44ae00eb605a3dcd664e4ac3e2689f27fa7d310f3aa2a958e9fe82be18e525f8c0b484926c3c3a9ec7291aa01bb006d062dab3ec21367b66e120cc00;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h5e13521100092fd101073d6fec72c5cabee574813fe26c2036775bbdce27c974e9039f8327c626c5b55aa79a9f3febc8353b02471cde78ff09b7ad9a3a6b8c247c4d17b54965c620193dc34bb0f601404cc8ef54e246ca6904d8c3b1563dc2ebed2d9a29cdf78a530e9564dbab060b33d17c2827477287dcf281cde6dff2845a19ce893b2a1c4e6fd06caa9f0f778d451bb187ad329b03f75159dc176abfe456b21fdb752c7fe2e4a834854031452f64d522177a37f7948b91648b72d6d9f13e5427dccca40b5b4c22787d05a6027f08e748e314c627b88e8729db0fb161f1c3795fafe51c1c753bc512af3fd7133c1a4e7c828ded299c6a00d658400ae562f2745074d61326d79c126484071c06cc0f33b7a779b15d86739171330c61b8d500a96230ba776d268433143f947878a57c4e25a0240c4bfa7411993156ad61d8aefada5c073ae75a0b0bd1304b8aba2632f115876f29022d91938cf0761369f86895aa4a2ab519490da0def5882a33719d01fba4fda5eb5ab46d73f706a9427458b2e2375d433f2f9e32cd8fa4b7663dad0c0ef9b0f0c74cac8c490b736c96ae922a55ee2214191d208f463b20d82affc880a58526cd0b2017963ff2362f5932139785f80530c1ab82a05f412b563e359189f6f9753737906888ca6a8740a844015c64ba4600b5ab02cac796a4861dee4edf38f72b0308c7f9d864f72bac945e009e01a9acfcc31b206dc9586d2c7804b2b6efadfe50f17f5e6adda0c1232d6a52b3867d131efb84bb309e4e802e55fbab944751fdc265435879c6964a9aa8662e60dc878f623ac7f62370aeb97dd85523a30840e2ca5bd6ba7ab9dd5f6469c56b35dec08e0ee938fb56a0be41558c304898dd53fe65f52dbbf36639ea6990d3b2f6de237a413d1c3964210e7112308f4ee29868d94888d4a9711144cde40152f37818d4780df6818024252a106688a17fe456378194b5f63fc7dd6a2a33b55b8c3dcf7b65d98173c84d9b039a6325d06fa78f0a0295ba88018bd5f7b7d5789ca73de79285a9b76f107039054f5bb608c5976718d3aa3ecf51553823a35c523dc288f1b36709b2f74dede3f233925f69642595e0bfb5a5c1b0343575888da2a1b0e53bb287a9ff765ec3cdf3cb814bf5a188da5bf7460563134c841d7546594c793321269a93b8c62188a795d1f65e6b4b4f4c5e218a3175105e234f9367585acba1840e59e52d77845bfaffee24ddf2eacacaec42fa2e17c052cadd5b39bcbe8a5430be41158f3d1bbe48f402229899f211f234a0fba46321970061a90e5f0e4e5461428ff225c9394190b0315c44970f812917e86fcfd202176ed2e584b56a35afd40e2df1a90517a5c65c247fb7499ba7fb55e3f49e179ee0a7d7b74bd0eac3ec0e48d5bf969c343e65cc384edb64d62dd7b55dccfbce48d316770f944c30c426f15432bf5df802d533a879361c2dd02a8f52b949b96997ca0862dae61306a85d4c64f13fb4b311bdff67078cb154882b4a6066a41a894fcef5aaf3be5a2e57e3174333c618812a1d99a18386d9514844a20f6e9ba4c9c719a1f427293fb35b8c087c839ea8c938ab382e470255857efed911e470b4fea4358a91a786a931b66b0b4b771608cf4c56e288a81ebea0b2dbb03570a2c3bc00627f718ee9b5186a369fb469dac326b8f0c995063115eb8d6e89b1ff4295a864e6932ad3a8739a1fc8ea234c1b91551f219636b41498bb402cddabdcf8760c99e83e877f62d83807f76d46fe566484881df945bd1fd63df5989b18527e9c2d1ee643ac50e45faec7a953908ca924c09e2f936f0aa741097cadf2eb8323184bf5ea73b302ae1557378be917b371048aac8f9e1207bf619b3578d656204689ce268210da84d46526f973a7b375e87e34fcb5f754d044585fd228a274451e148076c166b4573e94980cc2bd7dffe59642563f12033f4849dcf04bf8c64c5947cd322a6d1522d15b29fdaace441c35048dc4f4e2e8ed47c47dd3453c3ef22b7c88cb11c657432069e2b8b5b51b6e5731d39902abb5a6b153cb8e97376596b2a6f33863c98577264cf2caf774715b2f0a9ca6b390f02ffd4038b76600964a508286eb6083350c85e8c24303df173bccda61e6377dae1a9e1e2a0b9dc7adc73f204f8d06db20c9dab8b281d865bd20e7b1da9d109d9922394b627c48249a8ff063ed355d0aed38d334d630a5428a3e737b45def555a5d155429e9eeda18762c4d2ff4595b90b3d26d046e70fcb28be484cdb28f8eeb73c483d61cedb90d129d14a2e4a6aacf27133abc414f90a89c2b0c779dcb8d22987485aa036733c4edd6a4d13fd16d46090c64ef9672956d98e0a010dcf52a957e48070234fefb890b5d7e71881efca1ee10f87197de3941cdf1f42ab87e0c4aa10b9a241991f3d482ec2d0d13b20e745c04ab308efa9d5c3bb00a3561fd3cca7176dfa2f0dda58d5c2f01b23c5146e5bf419736fb8351a7bb017687c95f9eca4fc0bd0641f7904959b77fcb2a7aa7b8e16192c4768976c084cf0e09790603520a9d5e66235a85fc9ec89e7971da1c2f2bca39fe13544ffa83569ad41639d286fadafa39dafe5c46a408f970c247446c7a9c784ed9badc711f8716ad57f65fc047c6307b39c090eaba7aa8b388d6be062bc767126702223fc4a8c69c556ac585ad539007ed5a2c7959a620c5974a284d5abce1b2d61ad2a2fe3bdd15b54949a7d0587a5846aa4e9dbdeba1fdd1e24021050860865e0a46995833b14707a2a313d6be8e487563d2d24d19223fc86ff1544fd8d97861b83acff114bf8192250027f06c22479f7a97048350737e416fb80117a8731b916c79357fa4970bc642dca5ca1a80cbd63ad603140c61462ccc47109b35041f270;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h997f70bb5c6bae1fab95a1c283403b5821cf1d85c9d45656e1ca6cfa1526dc52c7363cabc0cbdc3fab49bd78766eaef4b2d6dfc73fefdbd50fe821bb1a1fa54bfb2d6e0912865769f316a25a2729062050c19bb797f47e54d5ecdd1435aba4d7448551d2c2ace0fdb3adb759970329c304fcac0c714e20dd43f45f171133f2c0ae9e8bd42130a4d9f7f9fb101c52e4c281721869115176ada47911e5b46264dcff17ab2ed379a5a8c296069181e96fb036fddaf2fc6764a8b47f87332ab25297d02f071ea93a278cd18cddc1840251d496da408ac87bcb564c3f8150889f805f0c317f1c053742389d5abf3fe8d7fd1b17c88495555917f660c897c774ad2fbc9ee461db5c29b799e4a440b654ad8dd35c02510f36930a562a4ad6da259fc790d69603fac7170cde35826d30804e0f8b5406e0afaf98676d07b07ea7d565f37d32a00a01859ce66555550b35b861698e330e3e7d327de7914cf61aec8ba117688f056b28f0090c316e82561a2c17fdadf5ffe50c7b471999d0236bd1147e9cf0c84aa9b2cef93c3a2cd787d54f1475735b5787f35c7a908a579fa159af7fc1d8d940bfc57f78b8b8e6101cecd089af64aa986bcc1dac281a633f556e1a5ceb3f3f2552e7a4d7279005b757ff14e5998a456ce91d4e86195fa3569c0cc7116237fc6d6fcbd32f56e8458875c1893f4dc406b27033078e85aede5e7d75e387b6c98701a0292699913bc6523af805b5d783a8002b2b61f9b0b63a01ca5a781d7e572c4d575519420a9a96a9727486932da1362958daa414c60f0782919271a20e6dfe91fb0095df7f51367f79220bfbc62f0bac78f64502b1bccd610f3c63bc52957799b5d22d1726f3031afda159c79fa7b723926bdc20975161dd4a2f4bb44e0e1b8a4effac1627c71d28def0bb676705ab935edddef9d9fd54e1effdb48fd5fd10bb51c9c016011f89d6b2c99321a3e951e03d639bf995292c9b96e8b199c218d6cd938968afb9bfab8c63061a7288b8d8a3712eb7128e4465585bfa175a75a445e6003f89d5ce7cc968b37cd1f50986b287c8e0e42cb44b95b399c0301502d416a5ba38b294b115c849e1cca6808880ea133565bf399cdb65172cba0c6cd3cda6de92f08eb47af3bfe5b0f754e9a761e92c9555112551526ee344d9f6b14e9d00e8a65a9df5e612cbd05fb9de6159d1596dfc85fbd441a43182d4e5c15006104cf6cc14a06af58387a502ac6603fbf75032817e1bd8a95f5a6b82063631ce24089046460d1224fdb6b1c63032fcfdc72ee47f1e4c540fc0777cb90e5e7ffbf76a066b2d468368acc0a1bbe8d0ec1047cd4008c1089363a89d47286988002638e9648c9a286d516896605c4008f4abafc752e48780aaa5eab95b62fd87606a105b6cf6ed152a1c473e814b2c658499295b06739b7f1505472ec7a7701d4a82f2d68e29fbd976fac139a6c40cf91c23a094da5da8981e167c2b660ffa46f343fb5c25a0d3d670e43e22616f0368573346d6f4a3fae7ef3573cd18442515300afc8066d4b4f2b6a96c1b31f51458404b5c36b51104a748de5610443a37f1417bd97c39d327daa964432b83cb1dcc143658a8d65530c1b605f21c3e4956d55994b48e8dbd646acb62444f838c7e863d9f43c26c96b18b01319d65d29e119de501410142ca71482d07f3cfb1d26c42934993cba5074e7e791979d687108e4508180cfd5ea181b3c18dbe5e20038a4f15175a52d526152859a81b7e879fae57826672c1ac215c797a97e2a8f228d9a1b308ced7d3a5e25c021a5780fd858eccba9388f9a15a5065f42a040087d14e1a985a6557aeed580c96db2545911775d70fd65039f89784b4c016beb5d5dcf5e29f39ff2dd1e8dc3ade34c353f3ec54ead34b56bcdda8e82143c3c0409999eb2eda6a2c2f004457cb9c40932133c18a53d1303335ef1a2fae1ab231d1e1396f167a9a7379aeaee4e55266b521b624771ed8c60a415604de9a2d4a71aefe1d2f12dc7608ad4a870af3845161d97e014f5f66591841f70e0edde4bda4636bb4dff3d9f2ffcd52bb0c7dd4d189a8d42b98649430ac9f7efe2c4cc35456b2209db6016d40d34a0bc2c66dfb75cd51d7bb478682f867a5ce792d316f4dfb9dc959fd8989b67a880a0c6b12d4a883d102dee8664a1e0d48c6b5f315409a1b609ef1e9439bc5dc670c90e8ca4c2b5279e5f3bab55e935cc8f8598207ec30d4f8b12dac3195442c40b16df5d0771e68953bf1a613542fca4a04ee2a02b91ec9c1dbaf0ceb1c16962cf625a77abcb2d05f3dcd0c02744d136a6f5a9cc12ac361c4a7a703a6c83d75cac1bb3363fc34be118364d635cc70a8a239f363a2c874707dc208c875ae83c83c556a646e6e4837043c551210e9d5ba088122cfcdae1b683beee66f48f87e888b6bb2d510c79aa48ae7bc2a0337cb3b4444590a19b60e7f15d36359dd512bd480465e96e5786836b63bf625f7da8996a74defd4c439417d980f8857658fb24cbd066001b349e5730280b0e19ada067d3ff6b62bde187719f07e7175283de6240a10d4cdb4fd746d4a21fc414dac925acfc4ec0fb7a68f4e6839e95f60cbff5069c160e8677eb5fe5ce9621fb0b8d84b4b6a79eea8f763dcb6d669b599745302662284ee9efc60f0c77fd94ffb210178ed1280151a7dc5e33d6cd5d00ec453d7a6c3382511942e612ea688c273fae222107899f1c507dc241a187de746698240d7e925c368e002d7c0383f5b79d7cd073240b391243c3b49b17a27bc3c78b21bbba8e2940b3f9fb2d096001e14dcc69bdf5b5c9879bb549fa83ee19470de05e5e004135eb8aaa16761231db55ec8a4d9333e44dca00d73e6e8d9fc693cdd77eab326121eb05c30949033cdd1aef86cb0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h4887f693fe0d0c4134e95ed6f191bb7e3075f1b1bbec7e8f0f5b914f7cbfb1b0305614772ea6b246359455ce44df4e3ff836b4cf76b7ca8dbd3cd4913700619e47abb3a7faac477d5ee133ee620171f1ccfd3776da50d613590b1df47adfff5a10d5ed1f540c9e0632bbd7ed0083c4188d3a2cc52c796bc77b77d29e9ef064c973ab2e69d769c4cccc8075d92bba8a0ed3574595e10667cb1564fdb07c271ff6f2d30cfe2fd79f21e5585e2340cd48f8ec3da23d51ae06fe0618e3f53b4b0e99bc7fb20c14979af3149fe97657af94113a6ad00efd1b18bbe4ab14f589716ef34f8bde9436d1b965e3529dbc6f492eded82e97638128d2c9e713224e622ef7c3e94557e649edea38af23da6f9779afbfbd88006ba888db72a028eb68d9a6a051fd802704dcb52709d828d7460850d5dae5bf45d4823134bcfcc54ddfb3f2016df32f5b9cb002e5d26eea6e1ed4f799ee98532afba44170359b4ba8e81ce34a3f1d2dc83be160ae5ac9b4f359fa40db42014de8cb0f4ce3591668b9711cc8f18741b7b5ed5adab48acda49fddc15c03480b36a4e99063305dd55df84241419b7fd16586130a7660b98cc815c32a0ab1f2d9d0a28df110717d32edbfbab68fab298caa10a31f55b722dffb71e2d7ab984b04482a8045124ab52736d1a85bff4b841566cc0b76e224d8bd92e7146ff8395650f1aa56203d7835ebc16dbb41572a4fe3770803cb2a17d740050f71b014dc1027a1fb31249f89764da5d140436b2b353a5b857f0d519137bd9da56b55f566d19b3c7689ac8b895af2db822abc81a76871bcbeb3d8cd50c2599f51ef704e66a14e626a6edffb8ad4af8a71bc5b3ed5814a737726364b6290e93f330f2a063f86320a92bc88bd787b457805dddcfb31327fd56228a76702fbe544d82988c6d16b9b9defc2291f8f37f87ad770086c597a09671a406d39b6cd393b849c6ea22850c0c78dab2726891b5e28b7fc0bf496e554a3eb30e657335db1547612bf19b406385527e5fbd0f1dd6ec28cbe8aab4fe5cf9f0f79dd5b6d7b74baaa30b8c04baf2fd13124918e74f9938d7e6c7b22bcc6de36c9c1a6c7bb7909556e25a9209cd7110565b944e984170c6b0b852d131ce0f6cf6e06a128a52ff9a17240c4c4b0328020a5694d4f943f015175644d5a2a7323a2f461eac3657354c25a5d0dcdf8bef45d31360d60e63f1d402a7f9713155b803fa067c66f7ef7f4a0a219f0b921e72ba98371a5f7b550dfd00de05e17a1c2e90ab5f756bc87bcacec3bc76735c6a674b6e57260bf799d2151015cc9d5955973d08e19e99ec55d860bb7e25bee95fce35a7400148ec1e08e173015168ab5f1e34dcdbf5390923580e1ea49caf15849b25a4f1da6699578dddd424151574caa2e54ecac90c4929bb2a6fc69f806d48f3d1620686cce7fd3fa471905939c204a2aabcd311e7f3574cb1793fc7e8e799957b619f0cf566b37238e2c902a42198782f85c554bbdf248b1a494a1816897223bc076d06b2471efeeb1983cde53a9d5ad055df65ed4b79ea8f09b527812eb7283a85cc48dd5ce6a1d5eb04c50b8cae7e1901b3e94714bd65bf048fbb2e80dee2b5177ea01f65626e78e50e2da50f2a25417991f4b2aac44b3089ae847dbc326b9c9e9c720b6f35e602cf3e93aea8948f21283c678a03f49402862bb5e0507b3695bfb827f8d72c57b07ca02cbfd921e0da5d5648ab947699551cb2c216598588cb9ac9da72912afffa3b1e3033a904e1d2146fdeb7fbe1c93dd00739d432f1f781bd5ef94b71d337ed25600e9d45cea764410f6f50646ec5e81fa1125d3ae4d2119aaeba3671a1465cfb31b3042389b05c64719923bfc3de2322d0230a8062bc6408cdf7186f80d4ca182d44184b133ac637f933018a93ed361adc6e602e5471ddaeb1c01eb7cd7e886c81c751fa61b42cfbab713aa3a5535f24b2dd54b6f619c67f04d9ea76b4608b5084a0dbb08e4a4d9837ba44f27d092201a1dd852cd560a2e298a0d6082c072fbe89b662076f4b0244958c2e0ecf88739fd88360c28ff4c5c01d925c92bac7bfb0094ffc239b99261d6c4298cd2d2557130d5a6554d69f2f8709f07c9891f31e5e0cc081a2782638127b0459787bd2d7a39a4e81035efdff3c01d8dee501fb176190ba6d195cef4d75241f17b523e96215089158eee865cc157ca837167fb4e15fa7fc99ea3e76f2ce11d4c9da914a3c169531d0e09c91e369cc39305604788cea0ff38930e00d5ae171e1e5f2c6a93c2efe70732ecb8acab8993d4ce649ee104f7336b4b996d29d52b3ae90323921ca143c043c7169db53a3d364d2e3c4cde7571b75e9668fc430881030f3e8a5372e0f14c653bc91c949f378147b2d23e3f3eed3e785d756eb50e3fe1ac3192c3a206cf63b7ea4ac11c920241c2b5cc9724717488646f510139f1e48800c26dc2c88c786d764faacb6ed0e8edb106dd304d238d7972605487f7c9337d80d6a8cabd7da689de74c5f4c434cb687a9d64a2fe358b4a0a4b13c9bc3c678ef6309e4c97f7938022ee8613133556af24505a8e7a85954b1466bda90e3e36706f39a584f906bd574e82142ebe888672d9eeabf803bb57bb02627a4c7130ce39ae0161971991c18742c722196ff190f35c3d02b2c481d1282a91566709e55f4ddfde00ed40bf1e1083f84d0623cd8979321cbaf75df3addca98f2745ad9f5d8a0648762a4aee9921667742d9af8098c6fc76ae1d48a95b6a61cb0170d9c8eed4da32ebdd4341b85e92f5c34f19b00ea1130954ec2c7f74b72d5fcdf0ecc49e1bae2ea76f4f5ed60d4f063822b68b1ecfad4bb95d365712cfd4244c4019ec4d79cbaaa9a4d9b4b4042d388e352dbbcf283b3cdd5fcb4f62d09fa6665e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'he2325fea99899eb5c404e41944b07535089db6d0ba060bdca9d37a56ed187e901c3b14ecff111c236e798c30b79083cd5eb9655a35a8a91c50a7755edd9373dfbab2ae8a4fc9c89f53050921fc4df3ef5c6120070cebf357b28cdebac39a0440ed1f01b339b4b4666ad05702683d2ae336fae6bd7b7dc7854b633381b8c05afffbb831460b3f689c5ab7d0db8b35520efe405ec365dbc8eda5f40f64a1b3d3e034f3306be26a7733c35e2d7622fc5c6f6ed2b6b0a7ec086dc1eb7bb58f57bfaab523164a685e59e76416b2ab23497661479aaa51b614c03bfcbfaa1a44e53b99e44c2322370c5a0432e32d7c25a167fc0d3297edc465a226587b77125578b0617e1dcaf6b083f0fe387670343989ab31e099fcbca5612263eeab0045bdd09e4c01d7f072f14d4fd78ecdbb5d060be6eca750384e5096ece9d08d6a9f21cdcd1e9e729f1bdf9bb2641081a20baa0f4f572332e9d1236de02f370dccfbab9f7222706fa5236b8c3f035a8c3b585043b7da038fad7c0a126abfc8ecfdef80a603a53e35ece6f74f844f6ee7eaeeae0ce904041acfdc378a2569d586c2357563099ed26ed5af9c023cde58ee8f3000e227efacb40b61c22d1c94325b2445e10e2581be6be4c46f80efeb9a9e0fc689f4e63acfdeff152fba84863acfd7418ef0ccfb6ceb37d15c214756047fdc26f0b99725c87d176df4eae77d2ba59b09e435e59664e75023f196fd96997d77cc335832943147d7dad3178db730b7144729aba6f354a1a90e2819638845b9bc96c0ab84ed446c12d802de01cd2b74c2826fe2bf5188dfda04bc925e0c71ca0ada95ccaeec61c43a2fcdf6ec3d132b0e5781a399d2f37f3d0d24f0f91233f05385035c9cab0bcf6d3c11a978b66c4f23c688f5e21fa83421bb403ae15fb348891e6634e6ad56ac4b36e0d9f2d1520a01c86466aee7b6e296a2b0499943a67c010c24439b960b7cb123287a542082721339a01685ecdf41aa9399e52c45ff3cd923352d02539914bbcb6f59141fdadb65890939b510c3a6c7d80831683117d746d28e6e8e8b630af8b70bdaafc125d05deb1fa2aac49ca51071ceb060513bdcb5d1f690aa1bcae4cde544df16ef4f7aa69c7176e43e3c9ef623636a66e4bfaceb60bb072d34588d2c80fab9f306fe49a7e1caee0884458689688a8a1d79c665821adb30f6c22b33ee0c2361ce31f5d950dac68a7258c8b377f943688be740d9ee5dcd807941ec4f34d976873801a496fc477270be52b7d8e1b290b3bf0af7b60511027cde39ea81b4fb3bf98262f6c849599862e1a8d6c65b353c1efb25deb0d68bd3037250c5b715be8a34850af96bd4c32759d6538f6cbef9e8bd9ced95d9d550e4126247f2a47e49a64b999d0ed26dcf6cf22ad2375375ba64480627a2fe3d38237a2e37beea51865b7fc6dd72e5dda41188fe2ee9a633e55ba40e132d21b2bb72d53c1ae7c252ce4ce364698af0280e4eb864703f851aeacbbd80c434ac60b2437ec06e750462cf5f83d41cd60b96534e58bf7b23a987762696d5bceb81cbfca968ce902b351e72eac37ab04a38b12ceb9b78a4e8142fdfc15a28b17fceabebbc8a1824a3afff951d595b9716e02864c87957567e173c0feb5934dee7a03d7717649d131bca4169b0067c6dbd87ea1f8ce72e0907f7b72628280c54188d6d86ffc810bbc2db8455f6f51e9cd4ba835f32e8032fcd1469cfb8cc0cae157919b72c58ca5f6be3cffdd2b629e9f3fca04fe38673c42eb0bdd7a534f1c0bad2d5a776bd251837231fb32ac9169a2de4974157dac33459005e3ad85b167ba03f447c6a1eda3d14e61c3e0b3b58d4249734837a675bfcc077b430c52dbd0655ba0adb580a5d280e6685c8d451742b4a4ecbf231d20fe0fcc418c36d5666c2dcd918eb888cf177b9ede5daa70bdf70db414a171195fdf9654a014f117b9443afd4cda24849fa7db875319cca096ac4071f4c9805d8f7346aece0bfb970791ee1aa9650a8c75baa02b078ffb0750b71449c784d868ef619e758289ee8fd86198352bff5e985a4151b4ddee27ab7ac894491d636a828a4e037165878de6c81120c2dadd29e412969617d6261c54b80f72684d6c2d6647e522865eac47b67370a4075681fdffbcd9cc104ac2464f660f16fd37e1b440f12a81aa6a880bcb523e83dab66129fef4ccc0e3ed8f7eebf28f8d726b23c092a88a92e25e655371afa52b37cdd27c2b1b4fbae903498f5f850c04086d00b5f587fa0bb9ce03a3985cedbe829880ed204fd02ce2f83656846eb394c6b62c58bf0ece75238c62f4ab53a41eb848cc6d3f2cebcff986aa277ab84a52eb91b070f22d6a5e794104b25f8d80b62a89fdc2af6c744d4d97bb2d5b0914515bd71f30472157c4355ff4d00f7eb2f45f90defc7b52f2cc8f8f10951013d51bbef2ae6de52be75125ca991d449c59c77ed6b0231df08ed1e82dbbdfd8326d9729f7d7693f2afed4c346a38385cbbadeb0724546bf6921cee366f7cf23d2c993fdc70065030a5c869c91a928f520c98d802fff8d40299f3d31dabc848e8550ab55ced6df75e3a83f9b4181bfcdf2569462c612d46b7fe3e9fa18e2d257c3c7a7ca69e6f95ca16c9dbc0c5e7e472b866dd668222416d318a1c9244a3ab19ebcff8dff2d5dc0cbaa02d90964a655702ee09561777448fba1f59d8b6b4b777abfb0d305b85de9a6370e27ca723dcbaced4c2116e270a999c9ffdd514ebdfb3b778989ab3d89ecd4b40cbe4cad60819d3ad415fbabf7f60f1c9cf9627459efd54c783beda7be24d62e06f76525db3fdf9d795a93c7c744808ec27981742757506fbd0477feba4ba32187e00a67b793c21104c629b096a508733ea92dfca4e1fef7492b2e273faa8d48c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'hcbe11b74065a970b63e57251e2b59e5111bc76643d9fc36bc3fe0a4d03cd441d6b4521239d59b01f9fbf2e8939039e32bee07fa40be29000553efa40423de36af59529bc7590b18db60a8b44e7039931188487f7a3e3f3697ceeb5a7014e5444a2d793e5f746fc24651621d291e3f366588bc11896ba5dfe87327f7ac0a0757369c02b368ac95a0383086a7e7e7417fec04e7f35700fa824287ea8672ff0139e7212178abdd2197663c7ea6f9b6973cdb5fb74f7e6bbf58e1d7dcc963455c18fda2ec450a21be9846dbb3b2ed58e14955cab6b3a156bc075e19577e353851b0376b694bef09c06f709154bca43fa4ea7bcd5097d62474ddf0de06a24f6310c834f10aad68cf870e37492c2928a978de7d8156f00c021890571400bbae833fe4c8b69ef85717a549c9738cec4a1704b8630c5a26828e8854661558a259455814f0b301d9df6581b6bc121f1fe22aa15eb454e105658b917800c5ede2c9c1a7d6cfc328837e87f00f6a3c4fe9c40c3215c112ffc55f3fb817c432d3c60545bed92ca731f703296bd5f18d937332229e0f7a2773ea9e744a15fc9aa851246f0c31febc627a5ac66b7a13eca3857a698d10b4a94ce623e04cac7e0959811412a3c14aa85b3880051ed3a116ac628fb94dbc9e397f48db94425dbe222261213d1a8e97346e0bdf62e97c5ef353bb9fbaec9e0368a6eb43e7e32945528b6e41947cc8370002f431053b7043309aa0a72f6ba11d77c370cdd34f97a2e35fb82a1b0126ff8ebd95f0cf1abaf09c82f7f09626dada7572dc7cc36a23666d284dcdb541d97f2a951edcb88386def85e5beadc187b3b71e6d54dc17b416926d55f7d774d73413df3049a9e846b58da2b9e927e83914ef45157d2b03128cf81ae676814736b5ad5af1a821a5ac4987f9e089d47cb835f0a1ab62b048fbc84a10279e54039571ba3f84e7165629e64784a014979dd03d291a42f86a961f683e66d43b3ad2d5bdaf7a1981379ddfd0d2c12f0d94e109da633a0d80d074a0fb4881132ad1e027fad63d4446455f9a5178ba298d3e43bfa14bb58f24e0f77893d7bb143b8665f5241d9a390ad3d5277e0be1f146fa738b0510e949e4f75b2400c881e57eca4ac745e6b133d22009a84da5e6a205f23492edfc6a107e11fb276130d8e4b545d7e9c56d1f1f9a5f582ee8e09e535539190bdb9685629fadcda2db9ac366f2c4edbf8f2f27ddaa648b056f2ed66e3bbc8d6f568d38109caa723b06954c35abdfb414ca879555bb9acaed59a5993389d72a9cef4e2ffb77d427ef8e348224507c6101e3700483eec644809b422d9e98b07b52dcc1d57416ed20bc9bce461e4c63e61f705dcc30ce78dbea498f3c5980e3c04990784b8d3f23a74e22321c904f9dd19fe2ab05fef1979f227eb0bc2d48cdd1c9d84182d6d0fcba05636f8419b88c495ed4222ebb7830f3d6e20594cd4a898a9782882fd5e7b116636999ad5e9cfb1352b69fa693c1704e6f8d67b13e2e51bf4a2643dd96a877841b16fef7ce747c92c0183e3a90902b6127363eae485faaae515a5b8eea398dd66b6ef9a8c63da6167673e0d41fc3b7639d19fab2cdfdb673feaa247215b32e825b22edeacbcb238d3e2276bfa0226c4356b262d30b241c173bcc11e68c599ed7932b576a3286d91df07d85268e810e993b0bf5bd2e8b47c918f2168bc34fb3d8056d3967f5ddd8e75033d379a92a78ea147954d85f7eb232c91b69b5f64f6f7f15c56ac7734e26cb1ca494b4229cc813c591d2c9993495f04d2faab981ff7ba7204f7da91c990ca999b113dd65cfcf965f960d057511d6b63df174a94946fda062292b157cdcd49a6f5a9baddfe2a22c88daf2cfc06d179e122c5a58021ab42eed4449841f5b160dcbf80bcecae543d792ed7b461d16853e8a577c3892c7c1b5853d6cb1af5a4ff3feea94a6bd39dd14da3270ad8631e1cd33e3ca9397326662dae7fe51ba0e9d2488452fc464fb60173d02e514e1949023e647f2ec212946d5b16c6f6f8bdfa9760c5450f7876b66d025826b6cd91f85db18a71f71ce38d6babd14b4cef555295e900fa2bc67e93130a33a4d8405ebedf6d3f4a9e8999aaeed90221b6d9ae528571ff6118bcbaf4d531a27958108616d46d37fd34ec33a0ea7a62432d918c4a2baa1c7a5b78070a9f3ac4bb99c7134b2db73e0868acab422326b355299d3c0bc5c05d373bc89d0c9ef80fe9f65d2e19dec610b394b938031651688b8d3ce5d72c6df4adc1a68c85344794ca9444f78fcaabbd24a26f7536fad245ab7478637838f3222ee0306ca4a07a1cf957207e8740bd3f433a24d76451a3c01671abf58155fb145539ee6e48e89158f02072decc9e4be242f8e5ae26e09e5f994a751f7d477eef7ca573ba7dbd96a6a330d73ff61c6a51ee749d54f0b553b1ddd2a21653272eff8885d45dade02bfb746b16f08accb6df3ac7549c22ad78c3304a5adc29054e9d26499091a5cf4ef752939f83e819701553231cb33d85cb8cfd5288259ecd59f34cc329aca4dc374e050d9fa4e768fa844a09687047a8f6b355d76c57344643b4b6f5cfdfa186e82fb59b70a06cad702f96781312498805434eb73a950555217dcb7f0b291705efe4ae52e56282784fd3304d84ba1f6793bd3afb7f4e5fcef22c235a762e6a20abca30d75a434068e6cefca83e72d808faca9a3cc05cc4f0627e87cc0220e5893016c7cbbb2faf212287efcbd9a043ca2a49950232fa5e5a8d8e3f618e9962044c07909a82ac3b48e8e7ae20e3e381b0111654ee28dd869bd20b15f83f4a6d64eb32883d56766c4b5904df98eda98f84f06b352402d0a495ad37992796197799e02c5c40b47d6b6c214fcd4ab0d130eaf731479e406cccdc82b21;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'hc252e43a46d3ab195417dfbea63ad23d46ed174401f70d8cd4710ceb743f0aa9098f82c0cd6399bcd4d9d9638abad96fd2b09ff80b1dbdd1a2b1458d5c041a979a0def7ea63918cdef6b89ebeee76d377b146591809edf5702520a27e533cef670ad976530345ee81db6fbef1000abf595c5390b923b7fd21afaac04dc0fbe362027d912e767e2bc39b62a45a45adbd4c9543639db19807b179e712ccec1479b14beb95879282b8f8d1b8aa1f8d02d5004e6e8471112b3d78f8d58cd0e8af9dce450c45e01d2a6cf1321df17b82c7f86684c72c59c066a6e560017193cfa386e0433b5768faaa3c394877e0d676fa0c746091b8d6b39e3360ff744aa9ab859647a647103fc0087eb18fbc50ae231c1c8637949d8afcd20173d305d39f0d704b68d00f99a59baac7a7cd9de8ca5722980f27ba4056758e8cea898cafaf0aeb8a24a516bb075ce6a4eb2c50dfe4f1a2953aa99bcf17f15363136099c8627ab3aeb8edbbbce34538e173eaff538eb99cc00fd9a66c4557c3204f4dd861d79ee92fdddc79e0cc4ff00047398f5c31f292c3d95664de825e12794100f88288fd186fe30ddc9dbc323212aedf62dc7dcb5d48fd63601ed68189875b0ab47bc7bac2bd54fb43576b5db24d6c894115b79f0958a6a996b8a5be6d77a931eb2499105619566b0ab6398b76a390492af3a0e3ed2b37dcd936d15fa28a68a2c367c0995aff6b82790c41cd1c962be7efba8e5fa1355c38ac6a1a6a90d94f9352ffde05106a605de4776e8f72f3b58a8e687f68b4ef9ea5d5695d1735ae3edf45b303ba7709558392c214a44766ae0ab84cd6eaace2be49680ca85230143410e4614699837af9edd92f3b78cb7e5934c7ee62b5274ea720859c2d357cd843c13b979dbe89e56434c6f6473ca6e1dc4e7b46cdc817ef72a017c92ce7d1d8f49dda9601b12cd43fb82949cc74e98bfb9df21f4efe80fe67c919f34acec9901ea633583eb251a39aa7aea7687d8a8ae3da4c737cfd91787b6f0ad818902cbfe0f59cd15d1422aab94abaffea633ad8cba2361e9c60a3dcabecde82bbb5e0324932360600dc3ff33de23f9a70359d7aa8a3488cd3a6507637be27d007bd0c58460a8d402c48550242e9ad3d8ae45d17e5ab2ec64628dbf513d28a7c7ce6c80494b86fb2623b00042954914ac6db9f72fbebf1a2866388f68e31abf48a84f0db1ce43870410c5e8bbc92b5e21b1d87ee5b6bee11fcdb546dabb5883d24a55fd8c266f5bd0a80b1f50c09770e395fb966198cbfb9f7f3516791c166b4ea46747768c6167bc7e3bb181860c17e4809732aff7789a74e8689174a023a4ebecc9b051ccd1591ba82f1c6534bd7c35412909604476b787f75f1934cac307534ba41cf0a0f536728f1f6ebef77cb8f95a17dcd6dfce8a928741a6106bb675c9856a572a593e693355adab9e2335392b2402f07ae67f41beefecfc543a8790e5f7a1dea32962295467f1c77f4cb3633009ed5239b9a12a43c506b9c93e15863d8c013d38fa570a566f226aff419786018d8b33532f1fb9d6bb7c76e488c836fbe3d4669c67d6926841dde5da435a53ac8138b9f29f9a0fdb0877e86a97888cfa76ad5efa0205462d16ce0a06bc2c8dd7199548ed975209b8af02944279547e339893c9ff520dfc552c3e9a97d858464a2164010b91b46f1d880038df5732c699f3f715e3f136b892f0cef7b926c50cf108d7a904d23c39d1d12188c65a7653f7c414c3357a073858942c2703513f767efc85a8030d6e1c7897e603aed9344f2cbf2798ac827be2d6d6c674ad94db98143b6bfb420cc67bf89af9fb42c20504ab9db2596748c268d8ad60ff994c40fa72ab1048f042b2cc3b8ff383f859d538849d1a3744226b545ebdbc484817cccfb37ed4cc034f614aab492600ae4bcfb6495f0b9b130847b4d25ca927f899c0da213386531147526dca23e027c668e1c591bb4c43b36deb070a1cad68fce6b24edc25868767c5418beafcabc2493315545e00225fe81872ebc8d55fcff3cdc6a2b6b2a19dce3972834b05c2391595df1cf35a1e003209e8b6ade5cdf94b95074ae1332ef697056153425f70cdd6c7944f34c47088c2d083ec07b537db7509e9d5c81d0706a93c1f9911a8e3eb8ee544dca750371c2c69983817cb3741a5a20a4eb7818060f23d4fb944b0382e5445a39450478a4bf191dd579ea464d4b8050b9ba3a3dcd90d20a816295031f79bbeaad4bda8c04bc80c4e2a66cff36b4dabbfe98738b106a04013ed7cbe844e18873623b585efa3ea34853248e325553c2a34b85e9108a69196f4c489700405325cc97caf892a4acf25f2456b81bdc24c6bb8f39dd5f78be3f849925c42849705996597e9b008e0f1275de0851b9c503b4c1cff7c749ffad766f4fb35ae061ac0357aedf3a1c49d21ee1922fe0588cbe57d457923ffe477d60298bedbd1f1d8bbc73cc14ae3d224a6953db95074843587f20cdf46ab062d63d11f862d7e3239e23d9db883024250e4a700ed566b6fa979b97a9a62ca724b91166ab466bb8cf1718593498619d3ba52f2ed254a76c3f491f1c196dab2e0abf1bbc50e56f639cc52cc9192a5c7120b2ff6859db425849946428eaf4129da025b32f326ad68c1cd679807fce43ec6de2ed41237ed4ac08a32a4c322870562a01794e67925effda2925634ec9a34cff9306b668e82610967842021b6d0d31a03012c2edd2377a159bdeb0b9a94f3e5e7b2288412fc34aa6de218c0917f5b8e141fdb8971ed906a9799cab96594e5605e9ca0ee8d839dcf580bb9595df9dff7f5c350f8f68ffe20ea1cf46c11de527317433f78b93e6e4054309566811b23fb66213970866dd667ccd0e7b2517bfca6e502df96d0d94891d8e9;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'hd6ae76bcbc2ab4f39167fe62909d92c5105fde8dd765d41b3f2d196ebacac2f48dbbf6523a0d0efa7f762508b39c59b20499461fb4dc9807c7f84fe890710adafe37dcb8a25b3b7fdce8b1c40c35ea8155cdf551858d5f83ada3b5baa937f8c5dabc748c56338a1f800d3bc66337ec285d03072604ba4949dcbcc0e0bbbafd063c58115a3ab103f1bcb0ac83be6cf23cafd19cdd361d0a380360348a85ef6b2d7f5707f839d34fa1c87a8fd543080a72d2c326a52081aac15eaef74a0c0ceada1ab1fe320aabfb6aeb035fd8c560c272b78e9919ad54beb76c9573694d24325d03d7966cb620f0a571c437db1610df038579b3d26ceeab09b0531f792d8b2f69daa8c2e9f809c21577a732821edb626396669a2114bb28dee8edc96d539a4f4d62beb88f385eb918ac354bb3598d4a28d615df6691ab16ebde9933b15602b866633038eede3f8f2c395a730b9d8b29d7c61d656afa63c7d0622595e477cc63b32dc01fa3f0773dfef274092ae83f15ed7f7a18098b177b7dd70fbcad4ebd2914069e945f1835c8b5d66e61b91f7ab3e5b5b06e7bc02f2ecb2d881a4052b107bb721f6d2c4a892e123323aa1f1261717adcc84003106d53c275b2893c5eec99130c73d3a05e64628c574cd8eeeb4a899612888dced236691c6dcc5942b4540b8fcfd3dd8294767e8af9b87d85325c34a0746ba080c7fe48da7f12548ef3de05722fe2653dc3421ecfe2c76b4303aac32e09f498761ba19c5dcbd00a6dc11e43bb9f11977f85efe1c26da2966a1f9f8dc43e4993f54b117a6ade371cb730478cc5cf98796cf70a7d21e9702a66f52fdd191a0507b3720c3eb51913603dc0ceda763a1a309d58e16c8f6c25cd39f4dd66de1e43735059e5e348987a72255c18d7b4966d68ecc50bf63a81996fd88b3b3f44098a5fdbdefe157cdf40c019c048c0f5fa176ca07da83fecff10e93aaba580daab5d00b0c558325ea320973eb7368f1816147331467199c79aebdba6ff2ed137ffa9db85c392e53b5c5ebb68426b478892d877fb71b2e7c0a1dd31b4873b25250d8fd99d25ce5bd234488bcd9cab67f8d7d302412d10ec4903be543e96675da1bb2a6c1a4128584956c2e6c7112f1a5c2f582eaf49bcf8a147931805dd415397feac4bbc999f74e56299084404619511b3599dc247cda3c24747d0abf96d64640c3b7b6f0467209dd741b5c9cdb17f92aedaa7d4ffa765da49e3c79362806f2bf12c255ff3c5bbf29344451af2d823266855276eb0c30960830db92b61ab20e0d872f5b3effe2e9f62ce8aba995c6838a14d89bd8305d7955d9a79ca319b1d6b148db8a5f8795a076060e5b6429d165eb78b2d767b45cea47c85fc4675705610cd25b86216e61317ab37310e90e9ac3680e8ce68b12fe6e0320dfe19f418f37185bb4f69b549e1707b4cb75e92f0105811fd9a8b619c2938584a7c6fc5f7c89b3c32472e2ffc4f73e512ad461da4339bb00a80a47537a78521887f44002e68f2bce852f10a26228b9a149031373ddc6a6ea84a9738a76e591012865f27dc8ef2f51b7c6d3e2352b895bb5287b6d0f708b6e2d7df03a23c1f07d6cbd89a8e780e919df879b7834d917a403dfb99143b9471374613ecc450ab3ea8d699b1cc1310bcb5cc64874b5c3f278642e12546fc64decf773241399b768f0310a6a81319fd1980b75bda10c838b17d4f8ae1e61b75140f76aa70a2874d79f0fc8bfb67effa1334a35a5d670596367b9c93505c047d29e25f239ceeaec56538fcb3f7bd9ba1353b554f674cca571988388cba6b6a1c13ae71c8483dd9126f52fcdc198556dd8cf23f035790e9cb8f6e07ffbca489c01bd9ade0b318f81ab4c4ccfc08632a866c30344ab6dcb50db1e43b3190dab759ff763d284ae99b78ff6b0581e6eea9c98fd680f82d5781c603038f9b421d2b21c5fd329a5ad1fa0b47959dfccc9e5c8c3b4c7e333d65d6e9efbc5707597c05b151247b57d6180ac66ba2334893a523f1a1f7ba74362a036705ed099a39365a5fe93a65cb5f7846fd1fb1b8a88519bf6116376049b4cea9a42e6fbb3d56003124498d59a4c61fe39d18174d1bcf9861f8c9db8aad810ee4d12d4028595fa00bf2ca7bac7680fb867bd333b1a729dbdf9eaa17d7cf96397e3ec0b2fc4eb8d695fe697f01024d2bad11c3ab12edc2820375ec4425e0f13d1a6726e477a5daa00d79e62d2740e7a423d2a85babd8d41c60e05f200f9a8690e43ceaeb3842ffd9a5d73b8f3056a2714c01ca8c80b071895e4b8d8a266f68e07644d1314f5671d5bb2878361c4034bb34e397471e1271021d2ae0d34a0784e2a74c5bdc6dc0a30dbfcd38eb9e5d09d403d5ac5c788373864b70de47dfae12bc07e02b56ec1f6291da6e1463ccc77bc0aeee5fb36ad47544229e3a4f160deac0986530dfd892dce40e9c7e07ef6b21a1c80f956121b93e4ac50be7260fee27604e086a1d15875ca9be685518bdbfc674e501920bf811fc3fd94e2514874789886a520146fbf768545285df36d9acf48a7fcff569055df8adbec6f1cf8260f307294fced6cf73c9abccfa3c013c1c08e02139bd60aea4cf66ecaba15afeeed16622d5093d300d8b33d9326167ac2406467a7a8709b05ad76f1d73b6890c8db8d27bd8b58270f25e84304f2c6ac77dd1e5cf852fc381e28d9af421212c8c6710830a6963415b3e6e1f9156e6bdbe04c585c9a80aa011c15f98a34517c717d55aff476088faaeb8f831851cedf3c011b8ce4d9582acbadc68aa88e7524f5991d48aaa59ad133a115bbc8773b4638a262376d7a277f87e8edac9ec8ee300a77e9e0abee47a4d19b3aced3a572cf1d4ed78aac4a5141d59f3356ed90de84b5c3aeca8100134041cbf198caec4;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'hbef66f0888e83d9ba1a951810bbbeda044b7dedfcd37e9b6227d771d9914cbb16b8b9e2d01a062f51746de2f11c2db82b3164c3051e1629c17bffa2f837a2a4a09036f7e007dc04c713ebffe3e4845d5f17f57d851b365db53fa71635a09d7db3a9bc41f11187acca284c0a5312fb1ca557421fe75e76831b4f990704ab386a51096ae3711f31d7b28fa0b4bb3a01ae19e20fb1ba93a2a37650b12aa17d0ff03900908e2e60d40d99ce48633e61686a8d3dfe2755ed16ebfb73c2d4c00a862da25f8e8e6e6022948bc5f86912e55db5233ed63e745fe642e8cccaa925004169f0603d36f9314fc21391cff4494d54f4828a3c1e27602831e3dbef02e049308200538a0b0a796d3ea1329778291a1627f2da89ba3ed3767a2a969e75f8698bc9f63f20b95d7cfbc84235526c050c87608fa947a1ef9aba733b6d29ec02881efa84fa9863c74868e99ca938c7713d98dcc01c004e541c3f84c8e0e13eb5a3bb3065724d113392c749a82c3d383bb8a08cf15bf90a8099fc17922b14a1b1d3df95217906b59e867ab76174a664b05580bb9e18747282687f335253ec6e73f5471772b2a0329045d45c951abb52b5fdbfc79005863fb73c4c3f67df5a595462d4940dded2fc395209b0f9090eb320b23a930fd51688316d40870983cda9e4094d9de3151a4e2f884fb0c1439bb4b6f3e067ab06de41cb1b2b6298f90790dc150fede908eaef8d980238ffaef7c0e98b37f68ae2a924905b95f3f3bc940d2b8de6cb96527761700c900aad7b33489145556fdf3313b8f12f0fb6dd18ba8751add37de3381d943f9b334cebc3624ef6539e0e00d57f7e723eadffd34c297cb126851b49ef86cd4bd172560e6b724e3246a9787301b83d06bd39b0054203791e42821ca2c6471fc727014ddc32c5355780fe1cf2992560a654d839f3153605525b6f225fb1133678063b2251134b1bd67f871ed7abd8ff0f5c7b30564761c45500cf5ce6f4609e39530d51dba85337b36388959dc5d298d4b867bc828b0b0849599a0cf9ab20076ff5b2f6c6dbc7ca828a0110e5c0972501465dcf0db5d5a018cfddedfbc53e2769dbc588d353f657b1b6a978b08577d1ac97aa0332ba36948534815931b0f3b41f7c278e0a6a55e0a3e2c08f4bc0754013051ab17de39bd7399de52fbb7da4863e5a932a4fdd38741a935ae0719c182a0e4a9cbcdf63e12d12d92b37a9ce514001bcb32a819cd314396e5e6378b9347c476e0c24e492206c2d33fc4825c3b4945b43036c05f8b6db6c8832cbd1c1ba2bab01590b0898c92e772a90dcff6ac3abbfd85881cee2e69be5a699f0d91f6712d75502c116f06ac38e2ba216eae0fb9f5b9c3beb4b491a72bf4c7f0639139b99f337c894cffa9922bbff891000470b500bae5f3a8fe49eb98d355e660abadc5d67648210b1bdb8222bcd0c8df3eda972fce31ac7825580088e8dc9c710245ecfccd5437e580dd2e8f434b1d950659e5468945e5a0219bee0a379b7b333a56e6e44f3f890811110bf276f12c261f858b5e6ab5904ec376c4f52c01ec4574d5946de7b99e5a336463a2514eb110b091b73016203bfcc204e6f7e024140b9ff64be32b09aedaceefbd4c66f951c2eba65daec2dcb64cefa0a621e7ffba7a2b88b4c72d91bb3f9270472f0e6a28ddd12722d8bd43fceb8e8481b760bdb5f0aab999990730773f009276c88610b91e63de1b1bbdd24cff57490403e6572fa548a8c0323548b052c6e77f0ccfa309550166587921a0f82129edab329aa8e60bb36cfcc1e273a5535c1f75cdb34bb0ec89d197803c3587386e85b934463b1a8b3d6f7470ce5418cfbb82d1571047122c25e9a678b0a167f014de8a57d7b6d8426ee2c4999f2cd83b76ce77e5e7ee3d6a29fcae7d1dfb21550ebff8259aa08b7c35e50dbfed73c37edf598fcf43c5f3d2faf38fbc394b0f9d3274429f1086c5d307fe0f6ca4ce3e019b8995fd120bd2d33679ab54fd8ddac9706844dc666a515fe2e2b26b8f081174aa34a6b3d996d29c931a0e313e21ecfdf75c5d8eb4c94a04de96f23b12b16660338f67d79ae4297e3393a9ce4c9519f1c103efb8252cc96e74f234ec06482d434d3552c5996a0fdfcb4db5ee479672c6d3bf6287ee913a4f9a2edf1e67617b45896351a15e86ea6452ed683aba2e6237a8f3227d00e4d9cf4effba6c3be2fdf1b1c07f8410f0f8f6c19a88680089713f77aed172d674db8a77931ace353129068b599c370062085801a47d42c1580bc8a5de918be136430a9b03597021567869c5a331bb3267125a5badcdfaf855d010a0874a3e077497ce025507f5affc3971948562d2bf418ab1b3c830a746769c5f6ffab440eb47c6502b51f0f99180bdc04e88b6015a6dd066d5212774d97443f6898d6eccf58ba9263f3b8f22df981e28e513d20ded8e6fdd89e647dd552613f4db794a90a96d6939aa7da292f15303793c0c0b8739476c4c90d986c69c0ffecb9a31c945784ce37193915b8a2946ad6afef376159b77b712c2b18bdce4eebedbf390793d0456d1b3c7a41a525302a7e7b83251b98beffbe32419344332d68cf7a6c4f95d59d3a209e2f07b92db6e6915ab5e58dfb5029a5cc072ab05e1808fe974995177d8f3aa3e7b0cfe705dc33a39005657ae9b52c7d51ca245377de25bfd42d165354aa43a85f3a2cf70d5f05abd5ea1854cfdc18ba673b7c6a7cffea18099e55350a63440c78197518a157a2dea99276d82830ef9e8f9cd164c22f6cea8b897b0e26de98e6e5c4c0f2670abd87be157ace246a096e564521127497766879cc3d7729ab101eb9514a28376c1c43f486a1eb2614ef4817655f68b8b605e9ba5d817212afcaba530c1aea516e7992350a819f5e00ae57b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'he26accda54ee06ace1e7ebb011d836f1b18b1c4712da17af5599c8605d63a51f071d637b4137b8fd82c6579c8b6a18e60340861111b1f40fcd8877cc5694444d8e81c89185972162d4e541f3cab150d8bf929255ab365ac6f3512b2fef60cc9966548be0d1ba738ee538335de4439132da7782c016124e9c54afc52e6c19a2a2d8a6b7065e4ec02979e63a828c910437c140f3513bccb485a356a92d825880d88e21702bd4d53a776035e8af9b42b9defa11dc88246c8d42193c4e6a89dd234e17886fafb13a69ec7377f700e0b90ed775abb6922495169706f923311636cc7831f27d2498e421a718c1780cef6e859b3eb6f213a6ee3186959b7b6a972cc6c12782dda19c1a496296bc590f50a5c24c868b34063a567de560a6a103334f89a38394b84798706fc664ec1e9263e168174a231a73ec24631854029715d70aaccd729c2b15ab17325305196210b961ce49a6a18aa74906aa3e95932795b619472a1f5a20fbd8d774f4f188ec85d5e2194fcdb94e6ae02b03ea12b2adb81ca1c8d3774f6326d509f0f3f1e09a7adbfe7baa0a661cb59fec597ad2976578dd1d787f04f14dbaa5ae842c3aedc60d6c06eaebb46b3a0603b9d25587b2b3b896a904ddc0af9c4431efa6a23a3306fac2349af8a14f1108bdb7009fcff7eda54d533139df039a6dd35a808de0d3a0bc9401fb54773c4a243cac9ad99ff0be3ea80e30842f0df958f3585480b4fc55160b54f840c8fd8e8d0eb62c751585bb92f006523faaa36d801eb5c0f863ff3e7f1618ebfd98a8ff43b6a147a54001f9c0def0f97b88166781ac15be30b1c78228397fabe05e7a97b358057dee987edade938a859da66105a581fcf984adde785db1e107be1df69daa2b649fff505f1b2d60880328610ee1b9687f560821a3c60fe847646c3a95792e239e170f36b129c7bfdbe219ce2ee3f42a1e024640561b815bc337551d2f6a444470d5ec8022950972f92ced54794e20bfe0570a70131137ad1d707df2c4db494692d15ee5b6fa5955c2fb9f3c38b103080573280771f7600b0c6cf1e466c0265baa7e648f74ff3b9a9c63d8e420196cf0c8c65551cad12e40a568f8691968c8eef73cdc98ece40fb42db954c7888104fe92ff9d2e9d8121e92d17651cadba21c805d56e8854227ea24eab124e3bc5ad70f2c9eac21c5abf3c68d964920ae9c998272c4d3717861a7321a9a2853f5a23e91a5d9728196db456d04fa402d3ea2806b5020ca0fd26b5628acbfdbc220209381000afe5086f5088c6bdf67b98b472b8efe2e6d949074638e8c81f4c44f222f02037c6acb7e4e743ab1f586956810550b0137d43d9568e5bc0ffde6f67b1c27614cff9d1a26355b1ab2bad2f7014e02a879b9e6fe6c0fb2b1f202e445ffa60e385f687e00492df744354ef910bf33824c2c400f348dd12e3a4ef6dc7cfed3a7dddd5bae5abc39bfb04f9179e5d1959748ae22fe269791e6dcee183db7e6de3e228da6f97347248979868a8b30de916ef4a7786f0799131c6d04dfb897cec0ab48532771da842de7aa4d4892b31e4e14d7167ee5df6ed543c312244e612f5e1c438fe1c02fc3afe614d74602911f974279d1bffc3add82b07a2148eb4556315b8776a339cdc4068190b5b9c53a56b2a252b114d18ce27888707ea54e3df7d3838ee8b4f20a7ce61d662051597c0b96ff070cd6986c8d43017f357134ddb8c4dbae045bd222769c13e4c88244fdfdbfd86afd7b3316206f19269b04c8c1aa431eab3f91dba21458be1a89cc629997d29f822bbb86dfeb6f280c1eaa35f5e8c1746b27196a93503f1e973221c06f412b6079cd5994295738ed73a1bbba7bf36cf6da0199794356c8d6fee24125ae7869536755055a424175c410bc8419957822508038e4cda00cee156fe6e5af5a4da5e16638c4323b957401d69a8f1c99a134bef86a65d2f054c9215bf2664f422f31613f0ced9bcd1010efc33f6bd508e0e285f21a1df13b1309706651c0f685fca581872e4b1064cb177141f08868f6b00a4bedc885aece4509fb141f8596ec7843833bb9d6941da28452c90e4d407459d7f5c7ac5538890269bd54ce06fa88eced5546032622849758348933e495be8b80baf7c9fa5ca06e72845b9e6713712a33aa5f650d74706120c1c6d04ee7cdf53eb87b88234458d2dbeb5737d0d9798001502f5615a6c435f7565f31622c3230a13443249f59052e7db5faeedcfe463b9473d187a840450856b25f1306da2e450752d4262a25cf41b2f52774497fffa4d72f97b59e89e2637149818e9452a43d3e2e36721374fe11f5b8716de9ef07f25118c59a7fd8c509e7e4f1eeee39eb2b6ec6185f86e70ee0e3656f3e967af1dd64cf19f66fd0e05ff635cd6a78c3232ad959cf078bd7d8c54de1fbba844f1e79349a365e9792d2aa3b84db6a1366b3062ca461bf923e84746c6d62c84ecbb45719dd479162d2c127a0f910088fe6d6fbe81761c63394caf0265a28045005c0cdc7256301cb42813735aa302087e5e96344279677fa46bee904da4e15d18069b083883f6c30849accbe54d6cd2f0dfc7afa5ec8ff4513d1733c30a278831c65855f787359ce493bab285745947785296502b50fd38f645ca611ad55aa0e2be446694ceadc40b455d782eb1adaf6b2db1fda8c597fc89d262740c2513b6d6c9639e2951863a64dff325a51e1ea2edf74b7a1ab7c98bf72f7b76c5cfaa62b062218848bafc82df31e41026c8fe531c502824407c4ffb7468c9e4919eae46a29763e8d1fa882962b37930428be6ea359e6a95722eebcf9b4c8eee747c5cefefeac06b389a722ab7b5d04adf99c7ddadf7d6c6d1a84a349b08413b45623401a536141cd64caf8a702209454b2646485e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h89691b8711f4c51ab5436cdea16ae6c1cb506a93c7f1e1352f8c81abe509f2f2b8eee31441444e2c7156e492d3119b3ff8bb1e5538c117ba029bdb334f5e205c1ee2c7f500c17d357dde1b168c6badcb998415c5d6924b090eb341003309dd36a4c3904d451c39a445366fcfa6641a0895a461b3b147ca4db9e6661495a3109e62a2a84fbd1411576e64be08bb9eef9cdd9f477069d6c2050e1d51dc71b26ff529a4b7f8db582df9d2c72847305038d9ceff1c5733f75b9c4d5f5b76e36711e104e260db98a703c53ded054963da2f7873eb67a9e5ecb740b6aa4e64c8c3ef214d877dd64c7aa321b05b4917b80bd8766d64984e4cf9e87c148f033a8c3ccbf9dc19a42bd0d55be1aa60fedafec5b01eeb884e06d33405e5eefe198d93cb649a514a058cba0984ee798d50add6854e8aa9acdbf941de3ddd77bf79836c79dca061ebd9515867c3564e28f7768764ac8642fb2934ace7897d7ce7a272b08aea315b023c686f6c89ed8fdca4e3dd513c80cb72ccd8bc8678ed35a5d1ff89c63408c75881d73ca682b30befd31415b44dd3c999d45c81b35b02db8cc27c3d4695fb0b03976ab6d95e85443afaddb511432657a634a20a56afab567da4a0efe862375a1752f91d771e88c30355f01e7b2cbae412bb4291803e3b5c1de9f97b1c3922301058a915bf2c784fd0a624666787ba37a3ad01802f6bf0b2f3dfaf5cf198882d52ef40a4adf68ea78e4b687f215ceecf5e85b4af0eaf088ddb014e19fec05be35c91cb7b3df91988927ecbe6d1962f099766d5dc7111fd67b1a42bbf30a26dc973f054abb56a554eeb7e13740e2c7de9f341c7e71a6b77afe3bf1c24bede2d5d3fb0caa4d42df482eb498b713dbcacbc59b810ea75cc8b58c7c55cd9ed997f68edecdc3618fabc419ec1f7e1e566e9e23ca16b679686e1e476eeba5cefc6218d96d68aaab4263194d2cb1f57f6d5aa3d319b4c20e00ae74b6c266e20cc7dbaa9d4b1531357b017b6c718349b648ed78aa519aa572d015c8cfb886c6825cf73314820b49b02d31ef9eecdbee54ad5833f0c8adf1890c8dcba45c4c7d7cc8098c5e52b4cd779a99880f069a004640e529a7988a501f28986a89e0cfdc4c956567110dfe7fef7224bb054dc17367a72a9b0bfcfd3aff941d2fc48ca1ba167ba33f945bfb700547fb5d014f75eedbf7fec42814bb851939e6108e25a672cd2a97a49efbec31d03a23540f95bcaab711c3c670373aecdfff6feb98320134cb011454637bfc2bd1613bd4788230634d154141104b1822430b226bb9667a387420ca1ef468bf42fe710439fed8ee742de44fada12baed0c59305f54da7f0a081588b9cac8eb93112ef83d0aca0d92c95b1326d6946dec51c562898d0f907b0e3bfabd7f53fab2d806da8ef082f142a81396c106db6b3651d0734c801fe1ce3dadfc42bc5d71bebd256cf99d74b5204a40bdf2c0f04a9ed46820a57d7a2a9a4dba9e6bfda745c1541f2e555bbab64f42515ae11d92d03844089415a9f983a0fdba68bb4e57e398c9079e2dd544ccd5c38d58686d8584349ac6d224eebbc82c5e0493217fe4891b5a55d636e80cd1c2b1605f22167c1acb38def82e0f35bafde428b9f19f46919dcad911e8fd8a455188b52c012ab9a2cc475262a7ad05edd0f19be21e2b70b973557829c8923d6f063b3b49faf12bbcb43ff3ed2aa38bf4a3b7146046c0a8f663ae05daefde95fe2a0644ea16f57e9cc19bb4781a3d334b5d00c1793fb1a1eb9369ed03f21d572bbed6450595402f8d51c13eb76a736ab98b110ace64ba1e9168832f45b4b78bb1ec03c728554820fc2bec5373fce1555905dff3d3185e38e7029c24d79b03c103962cb62e72f7e719e02b9674989712be58d88658f48ed8817a10688d6a22f9bf1ece27b8678ce5ed3f6b0a0d86f98a40c88d8bf20443240fe6ece86b67cd2b34c102bf3f16c0921478d1d63d4c6a17a6d4cbcdcabbf38d54d8f7da38a59ddc0eab8134bda900bf622e6089a8801e41a243fb80d94d4909f75177a2a22e8f6041fa80541c0725a002555c0c6352868aef45bb1d8b4ff6c1ca9419315a20d46653f67eda6d4e3601f785e9a7ab2bbba912b6071c3cf4cbded406d44905e8b88e9ac04972f6ebd56286f47a46f62db3b1a949a964c8b6dfbcce74f08cc0a67ecc50a82595dd6d905e843ae16841fb1ed8f625adcff6f024273f410e41e14ffef38365c0ea85d610e4001ed1bbf85eab06f6d14962fa0d4594eee6932d367a26a7260038e6dc08d4c19f247ceea46c06e4b2fda175e7dbb61e564421e5d865f16b9b6ccf194b9494d2a6164087237cdc5fb828cfe0c4d1c982a1f6be278d00728f05cac3896105402dd7701156e976452857964bfc0a0cb7ce9f0b40713111bd8a6ab919bd5510d915e5e566b16216aab4bce1c7b50cfd936d78bb6a51f8bd5540980296d724c8b37c244ae08388b34e7b004fa5f2e20856487fc16af963086a938fd03c9c945d9faa8a1bbf3c6625c9abe2a27dba6f70cb3bc8c5d6be33dd244e29876dd2c1a1e2acd5a855c30089ef88e17c00d414d374b011ad1719b3078aa624c7fc17e2eb97caf83ed70fd9a297cc95307452a63705343862956d3b09b819e158fc3da5762df1b75236e5bfde0bde266e6cb36a70c9fd6b2da2715d069e5827707cdcd605a40c32ed49e057146e66f362bfd9ba9ee2a0b0ea67ba3b010e5da5542822856922a63c3ac7b0c00c072707f013d25ee34c1d5baf3ae6e0c72c9e8d228ecadd18dfeb43d9dd7db89ed7b509620c4bf397809279fa2f9359719d11c82a89bc18def6ece05bc58650eebfe42806ce7a47676ade200a09437109518b912972f018fffd5b1511c91dd273cf3e729a628f22f9;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h146c96d1569f79067422c9632b2df5300f60894d9be9c0e0ac91ea5e611f858ff174fc400fdaba5474b81117d0e76b7b39f4b4f385eb608430656368ec41fd409c22e7eb25b2555f7d30e3c30056174f3dc6c59f636ad7bbb7d439c95ee4649f5b12e69b76a477fe3901fe453a64417b703a6601ee86dc7370be8c6c611a796f02aa9ad47fe0d585058258520e33829988292d1e38e8b42208108af36c5faab865f6b30c3e868c259800be6ca053ed95788836cf38dd267d4b57f3f3925958285990c0d6df2459d4f148843ddb231a39f2bcec9c07f862ce07cff0282d06be05a1ea3a8e9bbef98c5a84571d502725496e146f2f2af7a199a053b8acd8d545dc094795d36f2334909a5fac6cc3d2c7307d06b2d5af4b5b79a277292d812237d0a10288a4b0320af6e6538d45ce27f5ba4979ab173da216373d1895cdf349ad08ce547c9701f0945172c6496576f93154d102433cd5e72af0a22925369c6feb89d242d1ee32350d3685773c8c3eaccde789ef60fc397a76fb8e98b4ab85d45b4400d21bd4ad1f6fc955bf227b36a233aa9f2c204954e6a3af24d73987f37823d477528201efa4719cff2efd921685c1000f9f77cd7fafbb84191f75b8a16cf90454683f617ee7a500855d628b4f8e496978ca58c3feaaf6f44ad2dd12b86cbe190cf2933453bdb7f0f5ee33a89f7a4a4859212662f7b76f21243a18cd7775f58a67368b52a107854b9c3247813d2e7ff040ed153426ef9dc1210982a35dc299b7c7a957910e11ce42d3a6a53497d13266103d94c751d8825cfb67b4723f3d1d78a04c3244187fe92102355e7a52943815c2ac035aa00eda332c651dd75d90f7623a0e5812dba27ab7598f17d2143b3bbe8d47617bd771e3ce06eb5be159d95b2158f3b57ec980c32b36a38a15a957663992ddee081919072fa7f20e01050f9a550a712e462952635eb86a36c7c9133a4a4a4706b722f55d5a635c35bdb01195a076eb61d17e22d6b8c0a057befb1f6cc7f1444664d5471ac390c6d60a2a9c3e6a1a0e3d260a5ebd43db94bf81b573f00c55baef2dfe030ec9a4e4f086214a968cefdd69592fad4e4938fdd5b6ca21a2f1637ae663886e0b859e90fe8d0a7888123369caceab78299ef116a01424990b02af58038f7115b9f25c4d5351df72fb9ea0554735864d1b22350ba15a6d17d84db0a3b718c7ac01e7ff4951c4d44cdffe584ab43123c71bd4e3d1e92bf10281dfd515d73c02b39b3ec1448652164e708a4e7d589e9dd23aa74f33720d0727275c1958175101b46b384d31351dd27d4092695f20dfd271a5452189ac47da35346fc77dc2cf6d89344df6ef93b27e008be6dcbd44497834b948fd37d569a9bf77c5d04a17b21bbb58228a84462024f9f2552aab2dd8438b672f93a3056b78eca6314575c4513588ece95c280bca46178974f7a04937874efa81379d32b738a6ce3dede52add5e1c7af82552d15453e6e579622ae7adc61f486d1f6e936c3a9e57a45921becd0d1609ab858e238becec1e47550bf5b9db8d888f9089735e5d5a5112c9f9cae12cf084a9f95b25ba8f602a6a19bb3b5f08c2c619c2f95e31d897d38ba9aa8c4df8965cae9242369ed400cb368ee1dd777ceb4582bd579d5a5f4b420339ea8eef7ede915f0da91e4fb7538e8bfb921bc80d7fffae7dd987651299256b7e5c8f50051b4f2d58f40a28fa807a021a917dd3c6b3aca9770fd76591098beb5866a0417cbc3fe88426d240d9c2d58bd01089a10bf421d58adf03112c6e1cc18adf1cf79baf122bd5bfd111242ae645b11fd3f04edddd0d9e33e1abd7de34d39bd36686c244bef6703da09473d5db5321c91c654f1e1fb09e0adccac17b632d56b3ca376ed8f6fa4626af9b2a5b730f6a271d9606da0bb74e9cb531457f80ddad307dc8a3b58dd606bb7958f3a08f22c1d01dbab118e9c17c814f7e137534bf1f1d1b695ff4687c11e85df82ff8aa5ade597e3c87814e57444910a103c4aa70301a4952a0e3992c5bd9d0bff00a769d4e519e1fd141a2d5e30c3178298af98574e240a73069e3bdc8968779e91941f62cc58770593fdced0056b8770ad3a847c6169a26cf21ca2bd7b501cc162b4205b64cd092efe0edaee85e4847e40a04711ecc6c2eeaf6ae5826652b49f81a243c41c18b51f59f5992a137971816cfd2d71de8889b9b217833f4e86b29bce32d0c093a62ebbd0fb254eb6e0b8eab734a0eefd7ede6cec0589cc9f607abe6c4dd7ee786dc72d2654359a6d2cf5c25c030ca137291512735f13451a9570c524f7f7f2c817fedfe67d45a2bf17b488b90fe49d0b2ad8d19fa4a442e2f38590101caced50bea917d33ee45e876602827ba8520eac2cc5a391653e1e95a0b18d7fcbb0cb31731588cf2cf5a334a61ac85ebb46fbfc424bf049222483545c3f1a6198f6afba1d714ad23206ea0c31be9295c439f65ac9a00a5505632a4daf008111a85b8b26b748d043330cb82508344b56bbe981ab7defa7b5343040cc3372f5423fa0b48a23b9c202b084550026367f16b5f9589b1c8dc4f4e1274303532202234aa5add7ce07d0b30c21ecf791d711f782a83ea451a7ba140ea22234c175fd20804972fef2201152bac6d19e22f8b6d00824edce87c5b5bbf64166a863162c10ca744673270f2efc41b79f472e3efbd585b44d152790fb1dc4ef434ee9b52720a2556edecc079eee74fa7058a42b243a9cfcf1a47ba4e5a5b4e1d92b286c7afb8c5b430d5643661711c1e8cd54a94076ea09bedc730c2538a3a2455c6e88f16a6ef9d0be5a2c586ae1395b2d785debad245dda7f12a6eea9e809fd798d9e92d4665caa8024f91e9c558cb80ee5d19521cc0f62aff6097d262d133327dd8d7165d699c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'hd47f77b437a9c62da2efda0755eb864dc8adc67696c993b9b0c562d905853c4d6cbb7966ab39e7d2ca8530a32892ecf012cc5b54e9217f4f2a214657e577f64b3cf2cdfd7eb97bb330b8cc510431206a7abbf05509f4a9a2d316e284608195e81afa967731f54b28736c16c9c1aaf749d63ae6d1b2016dacaf799565252aac04a31f08b18252caf23c1aa227d7113e8b50c1b863ab07ef63789f6c08d70e94d3860c7a0557dad8a7b21e424132c56713f3d2da5bbb957099ea74deceebebfe30d9a97e08d36f74ab9103f7725c501798675ea3586f7d47ae9836f49bf83dabd90d83022530939473c973bbcf5a183e800d7e0a462bf9e130b8f431f281ebba9cc517528a896b1d86a436426d95e3c67b91632b8dc82a6f00fecebc5d924713394885a323ded786389a3ed35b6649f70b92e79aecd4434b177faa819664048022f9e19d8b1f1a694f726d988d379aa154a7e8a9fb924969cc36f66bf835decdb99066a8acf67c77ecf64cc033712856fa6a1de224e1f8f3470b9c49e8d4312cfdecccff99a509cff1077cce4d0acfd5e6e5c9db8028a112df28fc7359733a71a7fade6d55175ead2fd4e989342c56e49e13960d3f102dcded48e9b1bf9fd5275519717a03c43b0923e77ea97ccb3ba34ba04e8b8a57bb740eee8d270bab98e8fe41af48ceaab3bfc59a638bdbc4b647bf2f0aa271d8a06be46c416c16ad0f45b49277cb68bc01353a32512371bf57f02347e6bb642a58e87ab1d26c9d39de850ece02289bd2768d936ebfae8c36d82f3689c0829417157fe046572a5afe1245fca7f062d335c5851db03549e2f7ff2a0788bd91f03aa7cace1052916ebf1967b6be0e7ccea0bb5b7341aaa9e1d23a220267cce94c1b89ab8110dd972d25143a67ff9471d14e35c0f49f5d4cddd2a45d4a1c833fbe542267fde17336ff045d013fbba836e72febb3040e9aa3100f4cdee8a996c90712d9261997c6936d7c41359a384ed32d66a168af4607ae6358d5b1a5c39ba3949c1f2f581be67b4140c903fd957b4a5e5d5c65cc0f45ddb3d6461b42771cf4f926d29193a99babf4af723d6a22c533ae314253a200b274e08cf839afba318a0200da38696bb6ca057214cd5dc5bd0f5f14beae08f8d0f199a1a036238ec8f67b127f06422e9e6008a2ef5651fdbc6353e4c8e75bf1f678e86d059a70f7582691832bcd98884c3df75de4836598fd302869207b5e8663a5b6d03572db74fa2e250aa9839ec4fd5a0e0bb73768026532488814c3cbe0e619b0fc0d9997cd7ae5f62012060c65165b6e72263c3ab4e496f7288baebb3cb0d666c086897318f856eaa5c3b63f97a6a23b20dd447921e4cb7c4bf9ceb4ae92a99dd60faf63fdf34fc393e6a809c7c753db7913c1b99b9fb9a58131154a158d8b5fade3b3c896d73443f9636efe2fe15bb8476cdf2a9d95890005e892ec20393b9cdd66daba8ca14dd54cf453be70d9ad666533d2ed9e73d866a8ed1dac1ab5d2a5de47d6f0e16b84882cad4ae541db683b68b1301bac36c629d098aca93ab8f0a42e8d0f6528534c46b70daa99b56ff0fb4d822771b04dcf54c60f0b8a233eb0a48540bbe2ee64fe8c74aae31da263749b5bec06ccf1248749328945b7d77f894381f30d8668709012e316001921d316a625c985a5a03ddc05f2fc7a426c8d0a8b8e0ac75d1bb0bc47970551ceff6e2ee16b916c4ae344fc7e849df2bac202940e5cc495dd3ff7ced217ea013bbbbb9d44ca841f2486fa4dd55fdc03aca6814d682f0483a00fc4f88d9552ebb76003d6591a20844333bd4fc436b1b386d1f6b297b72d8e89434280c2b94c1e5185c7673c4d7df6e8ee9a82d56d9436d218e572564c25f260ac6befd4203ccdd0cc2c3c52a5bc48d36ef41c1d8cd09884af5a823fe2ab3f3461987e8798dda61dac34e0a1a76f6ae20b8df50916787075594d94a11bbc2c6b4f8c1dcc99e1e336be1510f2cd60b4f0d05505615a540952f790ad44c825fff10b684b53eb56f5035ce33f65d951b5921d6d23e2754f246a3ca01a37c67018871cffee0ddd264d5372acd48df8f94edb76013b20b84b6b12cb86789c10d6717af2d7b1a80e9049e49aa608780be2afc63541ac3d8799554e23500bdb2f153488f6c8562f0f54ac0dd6dfe74ed32956a77604fca31fd994a73c6c00ce9f7485d4f4d174ba32048b36c2d64a2969d2d4540e89963c1fd0f0d831220eea17213c7a37b208022fd959980885954e529141416ac47600b17d3559ccfa2831183106fca941fc85d724648c4899e1a3c3c15b45f7991e58fd09d2b948ababd8f0b4b4ffb508fbb6590d93b7806fecf0e411edba18bf5fae656b1422b535a40ea03fed13b4f5ad577ebdab18881a9755417d78020ac37032edb671e09f23f7b38f99c17b73144f96134409a7e4c5aba7665e350d2ebc761ffb7bda51c41f30c4419ea3e4403ec801fb311d0ba7b2b649543f11d2e3d2497d73ee6aef5c2228ae8132399fe383d3a584d20ad1b96d5376f5d2f68286d075f9b1e5390c9ae83499570fa9d2e78720a349b700e212655204c9f64757e7759f94cb30afecb11767e2325636a01c945f9082b44bc9fe53a5c5ffedd280c3aefa5c4b5332d171152f8be2ed62b6701cf99fcf43a8f58627943b432c79241a0edf73675f0c57ab50bdeaf95b7270035cc01712e70c803ddd888ceea0b70acb7f424ae16f0314620368621d7ba6951842445e14f6158671333c7e58603c544c539a2ed38f4deb196ebc82022e98688401f490d3262b48db5d7c54ac476fa23b762d6a338a0421aad486f938304640d6c479ead1fdbaecd7f79e01d877daa52d4cebf21699c7b6f0f36ed94c75ff93326c6fc16b1a9bbf7d382eb7684eb2ec;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'hc435a0da75651b25fb827994313c3cba0b6249e7d4ecc7c11ec2e7444d019ba520e23f55374e675363075a85a57b126ee7bd036f25d466aef5bef41fc60154b952c425e7ccd28d75ca034ef2ec676ade1a58c38a207ca6703e9daef057ceaf9a27f4a15a0f78d7c25d6ac0d771f548c0562a4f9862fa1f2a58e122d73796a33895570a27298712ae16d940ebaf2a72873ccc76eb5f2731896100da1e7856f26edd3b3bd912dc332aa900e359127a9cae8d8fcaaaa93f815462e6909c0874554cf5a0822f4555dbf8ed13bc0c1477ca654bb7e00c23489656b0fca332f1a064546451b4e869f7dcbc8ce70880635b3e79e2e44dc23e4030bc180e464945658fd5c2fc85122fdd9aae7cc97e275ac3d42b07480ed1cb2cc5c7280fb666e0c40d2ba952d77b2adc1f101b099cf5afb19e72bc44d8a9592940809b54de49f7d0c88114d7321b683a52cba524ef5ed1a84e0b9471ea5676fffedb2302dd4454c527b51436e2a21811b3476b2c59bcc56e0bd51a7d27d3e2ea3995a7f3b50e355133328c0a47eb5bead5e070acaf93a774357562b5e07f2b08792be3ce1a97704fd47c2ddc704f08baf50013395dc2525c0c4d50d0b9a4686de8096043269f7d4dae846e5b110d2d3d5c8c0c0b7d212257f991ca5c54a82309e9ab0e5970ef065adf3e8a603996bade9ced7a982ed6cd54a5fd8fa4129ddeb11359ca78550350c1ad1ebc1075ae6236b94df7f0371f1441d81cc280c5d158250cee48b205d603f4899c086df973b31f8d39bfb9db956b49fa40f3bfa8fe93fb7434c81aa0c99fcb2fd8922624ff89a705c87c91c1f1f59b0ec59e57c2732c0d57b638838b9a9356e76d0de812bf47fadaac4ea1ff342c87295c38e957f3c5e3b9f09d9fc7f152f5257f1bba5ba55d9fb0d3ba473fe9d2246152beeecafd9545318d97f5c8ea81ba5bd05bca8d7adf2af1bd501f6a7e0a4a56003863cf1721eccce26fa748efbc32f67deb4ce4d233f25ac477eb5bd591f855ac174c26d397fdf02cfcd036ea96db92251ccff0631b623c59689eea8614b406c1fcd4b2105a4b9a4d3e7cba888d0a7b75a29fb303c7cbeb13dc71c49a16e4d16906ea67c382569c1322de42577b05f504f5d93dfb63db80e32fa057e9ce08fc01cc7132306adfe80018602ed242018de9f476be05f2c81947579da37d2443a0c70fa9647cdf935b3efe8c6b9a75d867c8cdd6e9383aeb554e25050eab745c9e308a5ea3aa851616b0cdc430101a85d9acfa5fe375fa8e634de6210ea92cce0b14fd03c68c644b1c22aea31e7feccdb633f17dd52d5e85589b53f4f47ac4c234930c3c79974fdb233730062b37e85982726375e6878cf8ad2b673919a77cb05eddbd53c088c5d3877bea7b962a70f3021b5fc2224788cb9fa43d9a69d5d6ab7f1c67907d7f816f7a52726ac8099fffa2c8ba87197d1e97f0a689288dee405460eb58b82b201a327e54da9a8f80071364bd68e75af15184462c157c8ea0f9f927104f056e2e3652a90ee18821af842d029cac62727769fe91acf4b983ce1c2c189e7bea8210e6dc672e2b62822de34e2c9ccd97deec78d1e9ee889e981b8f37d28ecd2405dfd8400a9bc1065dd16a6f1f86699e357db2474f2dc0431f1bb0075f1d9e6a8cf8099b56fc45a2272f68807f9c26176dc4ff72f242ce698750de94059ea35b8e2d400239a6d5363a0082add4cd48eda4a9780f8dcb4db6948b124c02f9675aaeaa8313d65ec928a37cc42f1cfc2f5aff4372208f934ada5ac4e7cd829c9093e5ccf74ced62e8ecd0cb0823f12a846ea34908409ea18d5f6067dadc26a92b2b60a03f3b6848a7ecbcee4848d75e0708262260124d151cb64358fb26fce7224d7e20f58ce8f52fc0058b34f4203f39e8ee7f84ba479921d43162a3e4dccd1ef01d2cda93c103a4728ea5c488eb3ecfe78f6f6e198e92deba59bfdb1113bd1ff50a29860e3c3290257db02247b6fccf79ab93ca6efd7eef10c5f3d93b6be01b994adf1076024544893963cac57f899b26718e1801fbde9d796e1e1298f800892698f23d742ab23d66fb294ef9046e39bad82903dfbd1d3922dbf1c5a6e874dd5c166ce007215f6bd89bf7e2890591a51ca8d98232434cbc8bcdf43e73ce19c4dcb63cf76b23ea3a7f7bf4137c6385bff4f3362044f475966c76e0de7db4853be6343d3a25ccbed3750b25b16e24d7740b01ccb94cec9e9813d02a06621e19f90e6076f1d2b848863e1ab9366242c4909b3ab0df17e3e27c06bd0e3737a0c65381b9844912fe2ad1087492d000142be9624746c7e33a554f567e41a3c913f7be89f8387e7b473617d198bf628a67f613387ca12e66e15d8e74f995d58df2be5b6662efb532a46671a12d404e6507b0617564aa0522a7f1c2448abeedc24d6e84f1c0ce66dd71afe467fe18aa4fab7004d493739052b299e5f789fdc83af0bdb331719e46f0aa1ab83e617deeb876f43acf9f96edc2ea879deea58dd7469b7142a7442db24c45fe537f9df7c9151b0067d3195e10ab4e4baa6239c05da3d9839baacde52f209d7fb6ee738abc105e7c245bcc6a8758c92b8b24fd86c36074fc39722847900008ed8561e29f86f2c61307f1ddbf90aa95168102fa9ef89e6eb3134cb55c9c35a1cd63a6ff8a065c9688777b18bc1eb4c479ca45476c02bb0d9ae98c3737fe34235c7447e51411a83ee7b593f98761cca2f5bdfe9d100e6f5c07c71aaa0b1c7ad70b4d67ef1f8d70faf31a77587d5177e9c5fdcaad13cb21b26d97fd73a111e78613589f8d8248897a120fdd3e5e3a1d6bd2b6bd373559203d3be6e8c59db7ab82c3e3f325228344e1eb7cb3c8fa63a5ca759de1e17d7853fd779d3b4c25790b88e2e4c09dbc21bfec78;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h65e90bfdf5078cd6e1afca7c4d0af73a9627518aeb9f01e734cba16349aa0479b102a9af833bfc36fd67df46234d0e9c77d8fd5bde0332b8c774ddb396869b6f9e6d5227dbb989404f48a21ccf3ca2e4c40245fe4206b0cb6c74428aa9d77024f34ac27ffefcb441da6451093a62a0f9e0c388577bd67d3a5ec3a70412f32b96cafbf56aa1147020655c21be9a787495ba855b9492fe68f61cea904632b6ad10f3123b23fc5419bbe5f8e903f4c5ce9915881454d7144bc4ddca79526cf498880a9f27e94553312da7a763645b331149183881d5412f456436ede8150dc3024d11a7f3aac023166946c7795ae7da21c91b3f1998390cc2ac7d4adc4eaead791ad01b3865731849447473b9b5706483da059f5bcec3a8ffe6728d4ec6f1e61696ce0634ea0d1306f7c325069a924052c2e405a64d4bfaa81fa6e43d0664650a5dfd103f4ba9d7e7fdf2c194a5c3728f999dedb2785ecc4ec28226d91c81807343cebda31e7921fad2756f0c0fffaea0e3d725934abf8b1b3706f409574d75c6bd9ccd6f90d159b8bce89f6b0062bca1ab6965e65a40b8f66cb2c910e4ca7ef8698e41bbec7fd82ebec00544663780e91fd58a494c7e513c1b67741e998a883e2cef6d41dfd8b7bf0356462469c1cbdebe0db5a5aeea3feef4524ddb661bdd02aa48478b2862bbc003069bc9486512a570455dfebbc2a9ab8dd5c401f82c9f52e55b1aaa4fc34e116b157503e9dff6b19f435a4e6575c125c74853de6278b61c2a43dca98da1e9918bd40e5cf7e3a4e726a1a09055c7897725c37cb57cf9c25b8665a3e84617061fe949a304cc7b9b7eae690edc983d2ba6618d05b69638c46528757193ac0b3cf4f8aa134d94bb6aecfad29fe37e164832c65adf5530da846e2a0fecea5e909d7b85fde41e51f765d552569bba2c720ef46a44ad53191c8bca9c3f1bbde947e4d6d3564a4ef95d205fcb4ec8f73fbd967f2890823c247405bea87cd05606ba701c6e0be43936c935c4c1d7f924cada44f3efa2f50d17a5aa8e1f286afe9eba62cd257eb53a5e89c7020e4c5411146069bb966f271bd475762e0cba974821f324349471dfd323c3d53f9414789b46c13be10deb01e1897ef56e1bb89c23ccf9c8e6f0b67242c9e3f5a3eebbef40f5ff38ca4790a800afd10866898063a72d39e54e9b01adbe1b9cca07b4d331c60468fb5a36d859d45673fbd773cbb8281cfcc2ef43df1780590e2bde02a54739498eb9174966e4f433249bb0d0a1e8b26b6011c000b9125708db2bbaca967bcc6bd6644603f2e423e08fe8c028af9a7c2d9ba0946653915f4a532254dbac0b65e78a148e9dd651ab3f8a90c6313cb96942a7ab803e2df33a88f8f3e8470fb22955112ab051712878c87490746b6e1d144bc58fbb45a339336552784807bbab4cadfd60fd7c6ba7ccbe50ecb7e8963e92895a3f9d3a42eea774f737a2bebe3bfb7ea18a0d30a103a1db734d468552d389ec6408050d9e10f06a641065f7c17b1b2cf1b260fafac6fc30f8d7fc4d3f5508e3bd849de53408bfbaf30a190e8b59eace56b0014434f6612bc508b76c00492b10f0fc2ffb4f54ad864aada36aac115d3af527ad2f683d898226be9584eecdf995409a527d90d8c5c21011e06496af60d1ff600178509e79b17fa3cf96f938bd2b78bcc8837bd35f7ba48e8a6e562d5a78106948a8d45b5e445bdaf9aa0106171f1422eb2c4187d08a5d5b2812fe9df3f4551d1980bb0d64b6499c1f274cba143742d7e65c70efe5923de757f1da2fa3fa72355996a76b8ad1d7ff9d3c0142c6cd2d521f615b50e2e62a18b389dc6b0d049a9fa745476a322da660ff1f355e6a3ea3e717ad635150cf1b944d8c67cced2d17d2f8bc6dcdfa3fc3e762ebb506269d94ee0fa17fae45dfb69f2e5366d61e5d2b3c780f936f9d60a822aa52ad81d6c80a4f4080a1eb37f62ffb5dece2f766905c5377c3c191b2048b6969fc7cb71b5298f40bf8f54d39f8aed4c9276049fc9825b1e47532223de94341235e67ad5de45ae28d6981a6d8a9c7e9a693f6dcf7dc2f9de041b6819c6df191bbc06b3bd4d2bbc89ddc86601c6370d556db2f0cbeb09aca0bb175a733291489fd2bcb6c9e0f3785127875737e2949405cfa07a6ec6b02c8f7c6b73e22c0736ed33d90ffc65c26b178550a712cda7d947e2f2fee80527981bf762b5cf375bfd5670fb0a85b00091de3c978dbf884a325c3dc6e92e769e78c01459004e3efb9bf4fb5377200b915f2f6fa924f99bf36fd1645bfd2fac8a872979728b3207e359d3e5ffada0746d82a1e91181cfaf632fd079159907f4e42a162727a2ee8f22a38e26a7be05de043d90a1f2e8445a3799f0e052103e3aedafd0622fddd5cbb37ed7c992ec2140f579e1d590827792b3c6507e997afe31b05d5c463c5065256d15462e2053285fb8dfe4a47812dc3d118841d25810cd1b060e126a85be47467c895f83ca947b29f2389925eb818e2812b7b3fe6094834ce52341da8f4397b078c06f92a21d354049021ab52c787521554c96197c221be8d2fcf23fd578ba779845164e3f63cec46c23dd3d78e78725f2eb896b095442a98c62254a4c203ff195ad84b1b7c1788a8c9038a48c3a643adad0a78fb1da49d82aceb32e1e157d09ce35d40b5df5c449b2ae2e466dcb09c060b4ba97ec1f350c66ff48f7c7a3fc9799e05b1667f6f8a2c0e6d511896a8180771a6181e177771807c4d2776eb9dd6a8853ed323b2fe0023b1f1d9ba90167235d10789d97c1af150825c077ffb36d69721643289e485117c2ed0ea7012ec45dbc4a2f46b6af11a5c74a8d137e31b7a386823876d737558711121917577e08244b05a31a15167f792a9aa2bde7685090f79e99ad3;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h91b0d6613161e533a6867792465c0b70d2e9b9023ee5af2da62b81800df1fe7d30d2542749251bac7ec5b1db9261730f830af99f76448500fb02ff5630101789e7f83b387d2c6fdffa4b87aa838efe731a12d766ac1ec76b9321717aa84e69c7975bfb3058520475b40aee0f963a2a713e6598b043943080fd212c41d3631a4ed03973a7a187864377b914eb0275da1a28e473f2c35eb3ed415e1b2f9a10f462ba226d19f9549fc940ba851974a22e297f27c622378d0f346f7f5d7569939bd27a2b3d90eee92da3b254876259209a9ea89bad99fc1cc5fd3afa94c5f470d367f69ea6b49e0e1669cae87b2f51fbe2d07e05096b899aaf6628d72de994533282830e6c3ac1f10f85d309a0a15fbd3e422387927e3488162c354e4edde37ee367b327b79a1b39b1120f044d0af4225e330071fbc85826cb9c24549fb66a0dd1fd02f628226e3d6659d23a0d24349ef0259c633cb63717de6ddc4ef332758ad1d344e5bb8341c5333acfecb7da42c3498dda4a94371551ffdc83552cfeb2349a505b44f5d6e476212685bc32cb72089447b78eae60514520fe98c8b91cd24f29aec66103fb1d4a89d457695cdcd2c0d8507f4aba4eda5417c5fa101bb2310f5d869934ea2448d885af072488bb3d2a913d54cb9549c48ac75b540383d5efa197b064f589bdaa4eeb8e2571d970ea516586615db1d1eaf32a25ea8c49b8520153465adf042c30b899ad5236598dab549e75c9c60b7ee735cdf8e4747bea35066a35afbccec6046b69601d5494aa9730dbf3308e061a10c9342a8f8156bf3782125b9a2fafd956d80a9daeb8efe2e6e1fe1243800b6402c5019a42ddfa725420d7efdbb9ec432109ba25ab199e1c47be51bdf8c2c161661f96805e8b731ed0f5cb0c34da429b7c272116e5f7f58017ae2b681bea4a2de5b4703ca32736867e5d8c830ad547434acd51e52e900ead20778eb5fff739f284d87e8e3ebc31e47e491f618bf5c88df90ad1f8b0a6be4df88712d90c988d634ab128e46ac02030fe0d303db169691f721032101c588da9aa358f4b6361ee755b7d5cc99878410fd2ae358402432dd339924e1cb54ed6dc4aec66ef690fac356a8144b3e9bc01249bc64c8a20a7c22f24b0907ce3edd39cef025da034ef585f86588e3d8f33cacb83a4283f096baabcae6c6b84a98eeb8f3a199ed9c3519c988cf0a1e941019f258e4b8b7efae7d9a5f19161dfcea6d116eedeeb46b63044d361c8b63310db92ca963f1db3c3c226a12680b757a61f78283fd8be0ad0f647c552857f7a2978678d5930a2be4108f748d516f57d25f3aa488f8f07c1a3f6d00d377129afaad654856edbc1e6d0beb230b424da6e4d1f6390b9263f0f3d8494b3c4f42f7260ffec372136a3cd659c5b60336dfbf2ec9e95f347d91ebc6612b209ef944996df6bb6a08c3cea0033f62ff0567fa8b22b2801a70b10fcfd140449d567238b3597ae7bda69b0046e5c931c7f60afeffb222e065212a90b5c8faaa90302169750afcb5366ddc4d5f23a232c4899160d989138f4513f29166d8e0b598901dcb6d87500c4ee10d5ef152425ee13f0233862a0a7980ff1f8f2d21de1102569769d55e6a43b9f242454f6e499398aceb6ca5ba61651c0e34891115fda85988bc15ddd7f0d8d339ce8281a4b97ed5ab58968a8070feda0a161b5da86dd8a3c314a589fd8878a2cd9e09e4c7439c5f5be7fe00954b0c71d9734624630b545052407e158b8d9235b17ba2234790a3641d960cbed9ff353473c215f3141ef425d2af519d3f7b164fa66765470ef85296eb9eb6b9eff98dece736426ca413cfce578e2290e67639c9fad7697eb0516827e7d40f6f31c93adbee9aa8264c346a3c6b417ef6ee46b674f95719e16c2a2885b52fb352b09b6a816d3f9fea3da92242897aa8ce15269afd7f125294ea1b1ec08eb86d0b699e20a3036397f69479755a1a13f4603b99745834cf96ab33286017533c5992dbe3939976f6c8da390f2cfc0bce5033d7cc59193ecf2ba0093e3447eabbac89cc9406a7cdc087099099583834cc7ef9bf422b96d3cfd8876d5d9b75ed0c8837a73ce56afa6490f4feffab4f6a3057ee89a244d7e945c3ac41425bf368b35f3851ef2ae44734711147a1548a9338d1db46dea310c2141a1f1e6684028f50a44fe782bf24664ced32285f0cd3616c26575efb790051afc4a03fbb78ec009e6ebb43aaddde504f98416253d1fba3f140cf769c7a41abcab66e69ce353f9815ec4af77e647136995d4e9de5c1ae9da5d7d0919cfe23dd2648431645b58c793858c3c1687c057382e06811191942c492d642f8245f8fe778158071412d0b16b915e92c0dc1fd1fa292ee36f33fca2b061f08f63a22e7ad70817e2ebe1fd0024fd105338608af617ed5fb20b1426245ff1cb0699418cdb1a72b97ae4a695eb033ce3e06044b61356883fe887cd875593da0e2f67ae4924ee49297be6d02223c67c308470203f15f4425d6ddbd265099778606ac88fee4afc327489a13f38d1bd9ec65b74a1249b1e43016bb309802d8ba3027930700e76a5f835c8d7b512d93f9a56b08912f3e17de4b795e6cc437dd7737cc2542e482679a637e16cda56f6cb862bfc3a1586fbc4b5e3b9bfebeb42f822059c9b47b184b69c821a271f0735022bcaab8aab10ff5994d321696614ab59a530edaffe039cda7d7e1acd05170d825e4d720e0a329e9190bac22cb0a7ecaf27d7b35f53de9e8110ee45fff5bcb4d5bda1b26deb4a21ee4340bb7d0eca8eed270801400cbc9199fb92f1ff7f26bd9e767444b7fb63ac3bbe9100c8c0533c47f88ef0d307b1246b5a478684c146931bc90a3488e251098a96f43090aac535fcfab596dc85b051e93333cc;
        #1
        $finish();
    end
endmodule
