module testbench();
    reg [0:0] src0;
    reg [1:0] src1;
    reg [2:0] src2;
    reg [3:0] src3;
    reg [4:0] src4;
    reg [5:0] src5;
    reg [6:0] src6;
    reg [7:0] src7;
    reg [8:0] src8;
    reg [9:0] src9;
    reg [8:0] src10;
    reg [7:0] src11;
    reg [6:0] src12;
    reg [5:0] src13;
    reg [4:0] src14;
    reg [3:0] src15;
    reg [2:0] src16;
    reg [1:0] src17;
    reg [0:0] src18;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [19:0] srcsum;
    wire [19:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19));
    assign srcsum = ((src0[0])<<0) + ((src1[0] + src1[1])<<1) + ((src2[0] + src2[1] + src2[2])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3])<<15) + ((src16[0] + src16[1] + src16[2])<<16) + ((src17[0] + src17[1])<<17) + ((src18[0])<<18);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfffffffffffffffffffffffff;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5da1d7c94a4a07f1ab3c6fc00;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hac2114521dd04010d37e72aa5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc586a3a01e5d6e483ba5c6646;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he0e0f163bbf3f7ca0c654a867;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf0bc2768ee8410bc5509c6491;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h127f7804426912947613b90d5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfe46687c7968584fd65fab297;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6e0cc0b6ee70ca2747e306b4e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdabc12cad15f25b197fce7d1e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h81227fa492b431e7b41232eee;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3069060e89eea9963a8685eee;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdfff2ebd8b3edd8616303342b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h19f24afa96a4dc53b5df26a22;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8655c2715ae7b9c9cf0455673;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hcc25181802c930f3ccb08f86c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1875f961a528930477afbe9ec;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4f31ebaedfbe90ee9fb1306e0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc6b7e5663743275d088ca350d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc9522c0a732407cf06ba46b85;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4b2994059e0051312cdf0ae13;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h541d707b741d546e5cc6f9c13;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc58940084c60e01fbd8415ec0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h58eb175d177b66be927cb241d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3bdd381e1a803c0591a2bde75;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hcb8e6ad9d0d8ece2f1f827641;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h308c748edc21eaf828567e167;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdc06293ce5bba5e14814ff9be;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6991878bb51c0ed2da2b5e392;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h77e0d261fc6b7480e97984ece;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6ee7d57b6c19234132f9b58a1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h465c736a62715119039540971;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5c1b2ad96ecdf33781c577db5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he23c78adb8b7425b6ec200ee4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2c8b1dfc51abb52691e086f01;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7fbefba241eaba7bbffb3f65b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbe50679a9b86906edae738a93;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h56b10e09e9a0953ac97f2d402;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h93087b212b3195a4f94ad55bb;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfe0833ad222fdb767a7097c35;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hafb907339658909ebf5742771;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb36eddeae27d4e39838f6a23;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf7e79b93bd92b7673ed5fc83f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h855ff31350f28f0024e8f57c4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4b0703149478bda42f2d5e41a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1a4c52ffa037dff975f01e830;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h600ebd91f103b63e73b503e85;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hcd7cb62f1ef40b39a9226f21b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hab7378fdbb48f812a636be95b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hcb000682853f8de2801ca974b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbc3b7d29f425fc41744e3c4ae;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2b77fff0ec5d373cab286c396;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hed8cb6a9955b9988838dc724;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hadc0c37dbb80ad7aa07434e4b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3131ffc3ac9f6d6a1bf81c724;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5c84e9b719e9de6164301519d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h429d248aa2ee4917bc4e4fb1a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9c3b8e5e247d87f1be1bd0fb9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd3dc60339569f10e219108d50;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf45a3d898a77a0b43e6c6c299;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf452f7f94f63c43199dd307bc;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hac5abf5462ee51ddd0d51723a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h24b34549c282296e5f2abe6a3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdbfd203a232bf878e1b9f8f8c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc1b585a3acef5126edec29e8e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h754275a8bc20b0390d8740994;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha6f23bb45b44bbaf63f83024d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha4fe16f7dea84b9e7f661ff59;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3af9c14b1231ac83494819551;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he52471afea5d3e43a6faac6c3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h99fdfa0f51df853df2215ec4e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hebacfd2bc70a55e1cd9089128;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he3ed2ab02b42c6da377948645;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6714c66663ba1f702b706b7db;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hca89748f96721666e7847183b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h36a51c79db43e42e7e7d74030;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1a788fda53577a6a2f1de0812;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he017c294015fd006a74e1ddd9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7276a16bb8209858b409559c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8c41d5f58e6937577b72fd47b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'heeac260003c699959708523e6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hea5b467c56aabadc55cf5d8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbea2fbeae8f93a6cd79406059;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc214c3227908ed16c04df423d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h15983438a3c2533c24e9b93d7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5f9a1701d629a5c425e2df3d5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h335cb4360e31a8ae5aeb0faa5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h44a475e58c35c32e60f6aa81e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3ec5c2c5e58f473dfd8d25c43;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h90fc39a460f5671975708c09d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6cd884a51d7a467174b3f0ae1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h96426f0186d318dd67870c1ed;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5f285af50d94b79d4139ef176;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdd8421d74832f6ffecd60b940;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1f54bcfa278cba8b7ef1c39a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf3e9908ceea0403bdb09db070;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h66e0ce54a1454af08a1611590;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h146a17cae9ce41035c4631b6e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h30805c3ed9a96114441e0e346;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8ed7a0c0a8a36ff4f23ca6892;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h50f31c2c1690fa78ebba25048;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2a7c2a7318daab3ef34ff57d4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he9d31c0d415f564b140aa6bb0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9e52128b351482ff9937122e8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9d76176d78b190c0f847c4c87;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbd68a48035a095fc281d268c4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf69bfdbdd5060f7444caad3ff;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb541b6614928dd33590707124;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfe6f7f01ab08daa16d4599bd8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6be54776ce1abfd0265a67c6c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'haeeaa248f5363bf52b187e600;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd3fb555b7c6f17b8881a07446;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfb726ee347073227f314fcc8f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hba74edfb87a235886940e1940;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h60bba62b1dcd0119caf6ca5e1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7c7040eb7215e26407d819808;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h20e4b928efb15bd8dbdc9e22d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'heae99cbfa24461025143a2eaa;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h77342a7b15435e8c4c76e3592;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h75cbcb219b294f59798122bc;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hcbe08ef5bfd736f412daf64cd;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1b1ec56c50a99ba8334d0088d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha97f2571c9c7b32798b6be37f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdaebd3032226a15da041a5966;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h62f94f31e50400174287a5c81;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3c37ccb66be0f519d5d757c5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he4325fccd412282f2ed4125dd;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5851d3ecb3422acef45e2fdf2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h48b357b77b6bdd6fc4c4e4d5d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbc78cb1ee8d012fbb61b3750e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf6532d2f7966b263872353e68;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf136b1e571e3937d490758bd1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf979a4a6a3103cc41c52c3564;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h26ea8456db3554416e61a88c7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h882a79661b6f8164eb7eb7cf9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdbb37213ca5606c104aa5644;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6d8d0d18ee7547740c7c39ef5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h37f409d220bd17ef3cadb57c0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h961f2487675b31e3148876bd3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd9613f3115f7b410641aa738b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h937d6a31aa45b690c0ba93350;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd7cc39f611ce887100fd49903;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9946db12663f9cfed422bc29a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7d8416a369498ad96f9f1d8a6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2ab73cb9606dd00b339077fb5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfafaf9c2481d36b36ad6ae51a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'haf791770d11e538433ea465f9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h48087f4de1271956267809fae;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h68d2bea30101698217ab960e2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc64913656e0b924a3179d668a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h745ceb5f8df375caf348ed0e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9cc04c37e6dd2b61f2a9c4c8c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3713ef4329574d6b478129e2c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd03becfc32cea57c76babe844;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha5cb3613f5c20e6f691c0e791;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7c80c1162536d997034f10d8e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4f60c5231976ea657f33b1c4b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h67d7c562183374fc0da7bce3e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h11a5251bc7e28b991fb1b6e34;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7122f2a511022b177915e5bc3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8214a980fba61bd89f0a57b3c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd4c68b6a40114a195f50a97ff;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h25f8ede20d631dd6f01e745e2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2de072860f6ea051554abf5f7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb861d132b9a0a3b03f06726b7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he5bbcbd5277db2d227c61f577;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he91ba9bfcc37a9bd6d44cb15c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb8155fb6ab70e4e2fbe3f523c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h65e68025e13be8f51d521b2c2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h159d1cea6d2d031466814e083;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha00013ec7a0f2c97e863bddc9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7b2285c6e9fb0d7a9bf81d944;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h78c51e76f90d69667b7f298b8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h10ebcd87288dd32ae6c7bd01e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb0a8c85401bf935478277a7a1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hcce1156763d773b5b2f5d192b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6811cb543b807a610c13a0bfb;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hcde93afab2dc8857f1f20a841;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hec7964b92fe51849bbf0bcace;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf85f18e1a45ba4c97104d5863;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h722bbd7435af19a1788381f6a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he363ce64a5dd8b82ef869994b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd1d61c256b9f760913382ae5c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h463e257ea138bb8057207157e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'had71dc9589801cf4b6b98678f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdcae1add8a68e5619c88d9ae0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h824c7f7b5bfc36ed02d6edf86;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h161c218574dd9ab99b70bb93;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h91e32150e6975a3f522cd5a4e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'haf160baf7ca1c21442ebb4f15;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc09f4ac64fb5cac99a31e3994;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5a3f8e81e8ef3b03e41e3c80f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6017b3de6356a28b40a56bd9a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9bfa6fa47e7135814c53f64cf;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h231ee1a8119c548e217777493;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf08b9ec85b9fd379a4ef9065e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9b3020e62636d03cd6fa21ea5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc0ff140517fe326c5641eed16;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfb626e9a9427ecc29ffdf1bc0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hed1bb2011d6117f6f9fce4bff;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hcfe056ab61b3c126749d913ab;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'habae5a50311edded63c39ece4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h77d2359d91e195facb659cfc4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2f413130371ccafc3026d8e04;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h65fa1e7f4814a4715da61af9d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h907205275211f52e0ca9a3bf2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf1b38cf68c13f485cd65e1379;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h853717e22270d66f8ec8aefb2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf479dc061ef1907834476417e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hcfbd4ab377b069e1f48c6c573;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbdacae78aad7989258fc5f057;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hebf7b58f1534c6d75eda7fbb9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb746afaec9460189fc1966ae5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h98c3c2d18e7cc7e3331b627a4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h44b1e80057e568451b810f685;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h83d234682cf086161bd2e520a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h91fabb5cc9d8384b0e972cc78;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h45ab832e878fb0dad9ea42638;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h500e1dd41784eaafc2a6a8a6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2e3eed4e1ec643bd8d8e231c5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9bb47750c1987ce2db82cde92;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h673d0a5882264b024260e7b10;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3bfa1795f1261a0654890ff06;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd5cc8a0c74045e2397d400da7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hde3fda2321a0d03bf5eb17b57;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'haf3093e472c944f83a756e753;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h581f8e3c32baf6e6754cef9f7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hab6f9ccdcf746b531545f9e44;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h87f3d38598e687bea1635406f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h44fb9208eeec4e4442583b3ba;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8b28f52ff132d187aff1118ed;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h93e4f4e21939c6fa081dc6e90;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc8851a7d38561b81ba11e52ac;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd1ddaa4b33091b546017f93e5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd129e7a082c13780a895fd886;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h93bde3c5942804e6b206d821e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h193bedeb569cac2335a49ac4d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'heb465ccf4182fb6c75b7075e4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd2a14d95d36bd604d8c7bcc6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h233ddbd583e4404342dc1416c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hcb7b20526a3df672471e47df;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6d152462d639acc24463f9a1f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hce3cb9290283b28ae76a9a5c7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h49c860997c16fe1b4ed8f988f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2b9011b6c19c0de3bbf27d16a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h52e66aa1715c761a3663f4fca;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc4e1b1c8df15633d3ba18a732;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h96ead31ed69bb056163ec1eec;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8c87f37d6d001ba9023afc499;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h30a3ddab0c730785f608b2380;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h10655d83de353c5ff30084dfe;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc3d32a08c30e5847371792043;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdc94342fbc731fa4da682befc;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h52d0be08b45b5047a54394ed9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h10c256ef28b0f3b7772d358c7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1085140b9d756df3569f372d4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he55359600d68ffff27020f777;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h579f15432de44dcd462dea8df;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h26210a96e7995e99304f84902;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hcc44b5a4c2cda26660ab507ed;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3a588f73eb06afcf84d9ba89c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h219eb2f0fb1e1c8afcaebaf9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h16fa40b0ffe0767e940c7e64;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h77d4340e59b79bad0e760c288;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4e0312da31d0ff4cab8aefc57;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h557fee9c784b13c8ac88253d4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h38605ef64518343d64f9a73c0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9a21f102c25bb4d982dcf8cac;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbd0c6bcce2fa2c98bae02183d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h38a838d9f03114b78d303cdc5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb3364e73fb3b0ad278207e6d5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he53ffec3821a2c7aed48a4d55;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h57996ad4d8af0529e88c51bc1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf8f89783c322c827a80a59576;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2c14bf934eecc1263f26527b1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he59c7a4954e12828a3a6ca06a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h531f4bcd36e37e99f4d929885;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha170b228c4e121aa73e23b510;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5b18ead15c49f4d36020ca3f8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7d63c620583c1695df6efd66;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf942b4443caf2fca5c6a76e79;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfefdd9f4e1794380855ffca73;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb4968f863d114cd8ed37b923f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdae0afd237229d7f3950d4e3d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha5d13f92edad16bbe144725de;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbaf9babbde617e570de67ad77;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3740731a5fc8374ef6371d04;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2b54dc10dbd934182f5f2689b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hac106519962c09b5ad8aa3d95;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2aa5e4991624341157b9cc529;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4613fff4e24637e60c913ea46;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4e74bc3c0b690341b21c11df5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9f0b9097755196d764121b02c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1dfe8b71feb2bdc0a7ce4ff80;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hadd2f54821ef7dc83967bc906;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc7032c9d9cdb73b5e1ea3bb71;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h22f8afc9e9a738c8296ddd7b8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'heb1935e30d2c31ce46368a7bd;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc67de9b5278c45b54d2f0592d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h564b4565b2effcf4108fe0763;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2e08405f9742792962b8bc2af;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h390f86e7c7a3baf9e7402be0c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7005e9d79caa6b37c7cb80c7a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h367389c66c4fde9a7ae84c86f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf121981bc80e44326e192e9c2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h31741702558825b1b298606da;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he3ccaf7652591d7e3459d7823;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7763ea8277931280c11cf8bba;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfa441fd53c50787d8c508f540;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha613626dd6075d2deb7d81c8c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2ab10a4f920d42a829237ac32;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfe6126781f0a735926f0c13e3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'haf739e2ace61a040601e3aa71;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hed5c0748fead29b1258861718;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h191df42f092959638f475ec7f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbc9081edd77b419cc7441e68f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h442fa43d86213daa0aef05193;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h618fb4ceb0c87707fe8dbf39d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8ad635d8f8f795355676f4278;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5816b07836f0519f293d76ca5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h39bfff6cc54500927bb8aedfc;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc5286d1f5443a415f12c7d5f0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd814af5ef543d0d6bff8d5bc9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he4d27d9e22f91547ef58a7e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he227019dc22d647238412de7d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h15f881b687f7f57c1b946596f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h25b77419eccce36d6028d5e6f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hde600e390e578aafbc830bd0d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfd23b91078b83c1bc686584b6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h37becb1cb2adb7efc0fb286af;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd176e853ba4b3f69d4f205ef9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h498672690f20472c440541820;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha6fe5f755ec33574913fbc87d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb17d8effa8c770ca1377b7a12;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha883debf626f79772d41c2de7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2dafabef915ddee0ffe4dfedb;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h43f1047cec59891609f52e942;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hae82cbb8d4537d0c579aef505;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6778074c152256fad43f2f694;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h15f369b40191d356beeb774b7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc37f2f8baa1f83fc5a9e9071f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hee39cd0efac28f700f9a23b2c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5260a611f0e3bbb11ee92ec32;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hef3aa9fe471ae4a59f5a4cb6e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h945a0111f15c4f2476fed5069;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7e9b071f1c009d2d141d91a0a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb11db8712b5f717102b071afc;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h78670fb357d007803fcc6aa62;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1ecf205d47d0775147b4a5149;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h921fd669dacc8d484d682b9e2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h93f6db32ff68d0de294b03018;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h79f0161c851e1b0127adafb5b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6224ef4434f6f0e38c7122561;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb1a875f0dd60026b97aa570c4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd6c957fd8f78c4214a3be6ef;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdfdae6734a10ae7ffb8382bae;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4fb164f28aab1e04a3b2d550a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h50611c4fe631118239db4bed9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h81ed6c2a61b1a0d1af67ae124;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd4e35dbba320edd3ea02f3eb5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb416a82bc1080b0c5a3abe41b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'haefa553312893e279e1f480c1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1c5e0bda1120c570fb0616bff;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha87865ac6dd70f8ce7bbedabb;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1da11838b72fb8df7aee4f4ce;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h23f05a6decd35266309fd199f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7da0fbfdaceef75b3bdc56344;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6de8719cc8ff97979e61efbe3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd2286fffed8c2ba3c1846e70e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4ce4935642197a25c6c8d59ef;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h52d72a681b0682ca60d454191;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h27a6682d577abb8306629f368;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h52b305b75439bc1882981b5a6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbfd6bc560e0039bb32e643a3e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9352c47490251da048ce077a5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5bb5e94799df88adba9cfbaf0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5e1f582f89c2f54a242582874;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h93462f9a7b87652133771c9e6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5276dd7a0005be73d0b7e02a5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hcce5f487dbed68d1a0ec4ee54;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7443dfefafdcb66c3f01e0c11;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc786d7a66e9faa8c34170fbc5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc12feb9ebc62b42ba8e657d8e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc0e1a6288376088c072c77009;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha4f2ec397eae81c9db5ed38a4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h739b7e3b8f784d170c2079e04;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb1d2f2b94228756aed6472d04;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc0e457ff3af64d6f53c3ae03b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h756c56ef382b4dd00ba236f0b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hee38bcaa8f31321bda94b8248;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h39616d3ec7e3b0b9e60b594f2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1a9bd3ae18a76d8d06cc579fd;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7fe58622df080f5a58ee3c5bd;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1d53333c7f33d07e2010dbc60;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h731f74dbd43d6c208e96e42b9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h212f3c12e208925c896eacfcc;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h17f1eb9599a0943541f2c82fc;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h36ecc077f969ccf1388188f11;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdd8d4603dcc987a7537c28ed9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1b143750fbcb35f1e99836ddf;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd23df6d7198b7177163917bfc;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb2918e96466d546bfeeea7b7d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb97683e932aa9759e11705bdc;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf528ba51b9c1fb14148a39c07;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h22068bb4f074fc4a16b165aa8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdcafbd11815fe5f49263efde3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hcfa5870034b2736ae8e246bfd;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4e788f69b330b3eb0cd019f01;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6c2f180aee9c25433e5afbcff;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1a0fba919ecd3125102261e0f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2b699c3226d7399c82c048806;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf8509730e99d2cd2561fce059;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf78b73594ff21c6d04022ffa8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc85f48b6fdb3237ef18a21518;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h758137e6594012eb111fae34f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h712920903f3f9593b080d7add;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5c403d8362f264297feaf1916;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2bd94228d494653c6f798c998;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc4f1fc7bf1c55caa8daa31dba;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8ce96b4dbd9238ed482c29608;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h64c1502492f37caf414ef5cd;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8a1fa75a71d3bd3a7db9f24bd;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hcecd22891a5f9247346c1365;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'heabcd1e887ab5d028e6e421bd;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h94ce4258ee01628f743add654;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb3d5788e3a6dd0d6333894837;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdf9d9dd429ea710060c85aea1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h92347966746e3d84361aa96b0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'had35ba1024ffa39019255b308;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hac6bba82cbafd2b3fb699a99a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3c1bd0a932b2ea9e07ce01cc6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfbf683546bc6edcc4eb21ee57;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf247ce14b85c7d109e2dd00d5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h332b142676fb5357551425427;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbbfcf9b9f66998d82d0665b2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h771594756aa9d6e5c90bf1f95;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h85efa8b1c984c01bfc69778a6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc733c6716cf11a031916f7dbf;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h958b8cb7a63c63f2300a61d96;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h33aac9d4aef90180b84e470e9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb6b398943f674a60a6048d6dd;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6096554b13495a9f5d9bf1d23;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h32fd588c2ffa9e2f673566751;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3210e2c82d02f37e0c829f8c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he5c2b548f0fb6b5d8e35c924d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7d1281f742698570b6e95f8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf61ac10167a34856884c25e5d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbb6210f5222732a6619f281c1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h41d54107d48dc8299e80d4a53;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1ccfa56fb4c19f464c074c48d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h27dea84ecbef46a06236ff096;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he1b52700a429c9a27e3c80f2b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd2a65200713e532bc5dcedbe6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hcaece77c4d07d0e1c026c5037;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha970d12704d2a7e486e734382;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha27c3a5190f9a114f1662af2e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3c062b5085cfcd2d2ba265667;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb1d8694c66f2d76c213c3a230;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h548287d030e8657094443c90;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2d34cb1b1535d9652384dfcab;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h76dd0a739ed5ea0350cd1bf8d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h23a8dd6a9eb8156f1ddf7a65;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he7e14b2bd1b0f4c41162fca74;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h27612416aee3db61f3a8ad0dc;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4c003fd4b5bbbc71c9fa419fe;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h15a2a007eddd682f0e52e5d51;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3ff265fc46e994e905a5bead2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7060f29e6515f4f0dc9e131d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h87e73bae2fb12a25fb9ad8f9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h19a8f4c6a6bb65dd291538b54;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h549f5421516be6ccee8e46ca3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbfdf3c5b390e05c77e16d488a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'haf97326f2cddd9e2071b22001;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3f8fcce85115e10190c824981;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hade0940ce5fc8e7f2bd668e9c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf25d8822464e95143f9abd73b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h36632a9314a4baca465d2f497;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h21c85d15695138be0196852b0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9341f915ed25affa578ac0e3f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb006043330599e0bead2b4253;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1fba06682cc38bce44d50ac6c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6f57fd48f690f7f98e1fe2dad;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd6480201db9cad45c95795bdb;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbb271fceff07485fc05b7bbe0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2f1b030e81d5053be85225c02;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he4bdc809174439c587ad104a7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h86373aa4ec30f96deb53fddb;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3dce7929d747c0d81a78f8a5e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7c6329d856871bd06c0218b5f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hed07ca14f010f4e25ca1e1bd6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc7b02075d689e5629a9e699;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h91aaa456945d9fef94b66d2bf;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7934c4ca247246d1a65d5130f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he30b39c429d40b6832dd0ab33;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf5827619f25481373e0e7e079;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6cc0d2aad5f3056921ee44850;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2b657454828f4b53294c3759d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8c7c922d05b1f6aeb00de8c6d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h12efe173151666c7c5e682cf4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h405e1abf0189290b98233fca5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8233a4883c73f0621a2d2d563;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'haa2577b91ce37361e50b52646;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8e4ff8953bf90746f6097dc0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h385c6fd83daeb4bd41fd4e412;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5046aff8887cd530e797e487;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h86a223e73f9162f6de4c82bf4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he82e956a60c79c90f4b465ed3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf6cc27035014901c3ad1e845e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9f4d80ad93292326e2681ad8e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h388b6da2215a63410a4f872cb;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7b0ec9ad240ebdc6d774a47db;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6addcab3af1e3d91da9751e44;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hec6316b9634484262a9c47aa7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he4c5bf9ad0b2e7ce8009a8539;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb42322351943c404e2187d2ff;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h781297005bc90c8a46d2a9c1f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h816859a269470a27f529461f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h59cb226f6864df2dc0214ef29;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9c77716ab166a7a7c2f79342b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5b64e62964fe1106413b3287b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4338a2d7123bb8d0069aa945e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdefb87674ce6acf5b7108ff0d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6ebe0d5fa7b76b3e4ce765d35;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdc46868486f0338b1229bd5cd;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfe413b28b3ab8d563163c6169;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8e133574b86c6d5f187eecd89;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc0ba312423f3a14a782478ab2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha9f988ee8731ac6ea485f2977;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h704f4ed0325b129c356ad51b1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf59853e8bf17f747f4f227eb8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3791176ce85f36b537cdc038e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h34d53ce79990115a88a00ffaf;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h423f337e50479930e6f6aa1c3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5585d602d2554824bdde8463f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7df512869caefa2baae8c4a3c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4289259857a1b8058e66618de;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he79bd7d28d392926f3ce0ff49;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h55104a8da3ab1330eacfef654;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h622656498f5611ba3af88f36c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf2c638760ba2b7ed6f00c0d47;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h761a421a32faa37d68adf1449;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h252d33ae5660248670582beee;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h70e1ed8464a23b4f9b23b35d8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7d4d3a8f4f8104d071c6b3b22;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h81465d29dee01a1f53bc8b88;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4758e0b5b0c48c7572997bb48;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he5de2343c20af2857feff3f80;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5b1b7a82a163949bf8143651a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1c8bf51da177c7c46bf49695c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc9a064f3ccb2a9ff1426321aa;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hefd3d24f173875c924c6e212b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb373828ee8179f4256afa517d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6c5669734ef686455260b66d4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h34aed4fad109894b461d0b5e5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdd6433713b5eabf1e0cd782e4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'haae3dc73d1d63d5c5dfd9a129;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hcb360fc0b2a07deb90fa28b84;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5a0679f47b8011213ae378721;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfab541c621e5002d49b22fc9d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h524d7addedc47398ab2d894b4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h82da68d40030e6ea098f1c2aa;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h85657ae0767e7d934c8b4b992;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h63724e7c4bbc6a9a9262b93e4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he9b57cb3e8b9dee34efa51745;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h47b1fe1647c3e0b55a90c6bda;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf83b2b6b5cc52cf21ff883846;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf4cff5fe15fe91166478810e2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h954f9ff65889fe434706a4949;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbe29addc58cf00bbd0110f29f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfeb41e851bf7b5cf27c5173f6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfafbeebf4d9da04fe7d1ecc44;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h61f28facd2391b5107586e69a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd91743e39fed1b2f8ca2ea459;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h900f3c2987b15062e518e0611;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7e03c4ec9b508b7b70fb087a7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha9c1ef0926b9af69384375c9c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h143b97ccc4b487feb8374e381;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfb7994865fe3ceb36e8169656;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2a39c469ea8d8a7223cd76ab8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h40cbe7285ea02126077cae7bc;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he16c396396cb8dd162659be77;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h80d60ff57f5ed9d95d9507e97;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h593aff7a123883ced34311560;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9f61f9bb403616be74ac30ae2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h103dfb13eff5705f8c8fc539d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h13e80eb2ce7fdd1a5755bf8e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdcca1c02fbb5a9a7c2b356cc3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h90c4fa1c10385c48f6394068d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc5dd9ec455d2145b666fc7d42;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb4271e1a9408f1163ef59da8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h17a43d96d94d121e913d2c58d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h429fbe66fcd980d9de178b8e9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hffc27a410788bbb2f04ca7931;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7ab2d52ec3ae4b8854c7e82e2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb69290ca905f7a6608a7c2447;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8ada93cb271d29402e08c6d51;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h902caa878b1982fdbe5189b8c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4dd9c2f70af8964e9c389c75e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfb9ed33de9b84fcd2492524ac;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he21e4d6bbe8fc796fd13781a6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbfc4678ed736c2ffa8be8b59e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf2840da8ca369c313b878b98;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd5b205c427dab89a6fd6af46d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5e9f07f2a4b0d426516f52b9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h84f12dc96a4aad2f9153b04a2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4cc3891bd3b571f47f03c337;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h16d7b9a861790091630e49e88;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb675dc2ef4472b611800bed21;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfe655ff02f2baf5686781de64;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hcb789eddb8bbf44e0780b7c5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4da4f82ff68467cfde98803f6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf7a81b81d6ae3e4121252a2da;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h42ff1b673b7c5f2586488b5ba;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc65985b3e9641a87ff70f97f8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdc8dc01ca38bbdb6f9aeef095;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1678785c411ba6df711eed75d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb551b29198bb3e365b15b5fa6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha584cda3bd41af39c90433cde;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h531ad3a1732f41b309a654663;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h92b1cb7c614a9784a730c30dd;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbe00195910fb329b0e08f56fc;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8f67d2899dc217e62b276460c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h94a0cb90a16d1134c67a96ed6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h356c5a75f4fed72b645d55bb;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd398644c7e3998f6002aa1eee;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h85f89904ad6e3a0572b9bade7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2d0aba34d75d495d8ea5546e0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h53ec6dc4c8bd0e3cac131f091;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd2af6633c495335f0ddf31406;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4d76c34ca249219327639c611;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdbecae62697fcfb4c76985b60;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7054c37e3cdcb16103ccaae6b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he0f24510e97bac574a1a488;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4df5adf5a005798c864176546;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdada9aee62445ffc6de6cb035;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6fd0cdf2dce7fd93a127278b2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h65e2cbd0d4ecab37a877255b0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2a76926412defc72b905218ea;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2d28652cd45bb68eb61b9f2c4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha59d34fca13558765e180630c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7df96d0613a2b22349e6c5120;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha39323458e94d4352c54aca57;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc609ff4bc03e3f4f5d1c4b404;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h10fc4005093a4376be90679a8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2389c1ae1d83f2ef9509648d2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hec063370174f5f2de43d4a877;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfdb65fdcad8b7a327b7892c05;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7765990e8e8d0b43fa968e63a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h82c7615c37a451bb95bdccf1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfb9be4c12909545f2b5ece8f6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h633a0efcec253f8bcd655da26;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfd6427d0222e715508b7b4384;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd4aa02a09a6672d11996ae30;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3ff10cd3f49870e9997776df6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha228e9e79385e69bfd817e139;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h31d1f28ca49ce1c4910cba11f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbf5971c8a0b3768b3ec528fff;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd9b7a3d7982b7f3f41670db49;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h18926ebe92662eebf925c6b2d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd3763c6138b477a9d8be64cdd;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf083d584dd202f40c5c6ee0cc;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h13e3cdc52e858fb0ced82ae46;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h41605a6ea4c78825a64450adc;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h216ee085c66a1500aa714a5ef;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3d6d71ec6d0b6755f95510a27;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h678587334a7b002416b82e758;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h203d3f61ff9f5745a5d9ef467;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h52fed8b4ba25d69c9195a4ea7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf2d8862664c7e20a718834b3e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5282b87b515ce3b9335a6849b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'had33a09c18937a0cabc316d56;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb77898beb8e866ec27d73e4d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h94857a3a83119c8750c085159;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha59966e9bd90fa8b8f6eb3bab;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4a7ae5241694bc2155a94aab2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1ee7b828b5eae3a5eedf7ae52;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h702c61d48ddfb0b15e7587ad4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h61f388f81f9e8ae3524b45e2a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf1e84e75fdff01aa5bd4dd274;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9ffabb4759b56a2c8db81ab57;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he37417fd510566957c928d649;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h802e0f68b98723661482aec5c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc594edb6b4b839186ccd85d87;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha9e5c3059f190161833fb7ae6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6984cfff13b6f8c8fdb070287;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hce77dc6f708d929136f460e8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h89184b821577ff3308ff0f835;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h44b3fc361b8cf7dc33681928d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3a6a4abde759064e6a72f371a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he9e203e46f905f1bcc0fa5556;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he63499a0763b145fbab9bcfb9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he440b3c18c6d6d03a94757d31;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd48dc19d856890e7a129c1a7c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h17d273d5fd2c3e72d0e5b8f1b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h150226fbf61755c64128c3022;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd36e5de3efebc99a746e0f89e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h445b4f89a3bcb4b9501e0d38e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'had459a3cf7b4f9490d7662026;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb55eb2bfd7242adba82343fcd;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1a44add4e1f0d993948807a02;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2239a5d83ee530175270e4729;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha62ad409d3b39b7e41c8558c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb6449adb5cc2572e7772979f8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5241eb5b3e80fc86f46646129;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4d2a6571cdca329234c549e8f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7b28d1cadd8da475b7e750c85;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h41d66642bf8f8284c5b583be3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd8c594e960a06fa817aa0579a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h122004779b7aaa14d095bf095;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h431b557514c520ea36e3e3242;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3043eeb9a167744bbb461afc9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h60ac1c9d73637507742a361af;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4c05ee9baabaf9dc7f7a368c4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h503562c52420627da1568f31d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5335ec356dffbc6aaed7ac366;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9ad8d1b4f73d1f2e3d8972582;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1732c1ceb87d1daac3f6446de;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h74b33307ff13a51f1403f274f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2611f04b7bf2e3cfcb21736bb;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1f747f7e287fc50eaf36719ab;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he23215a31cbd3935f80f1173b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1458eb71523eee4bfb5aa3bd9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hef7dba0d0e4015f545f032d41;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hefef8edcb9e40d6d063880289;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h427125e3538d1cdfa4f20e965;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1129c0f5a020fd1ee73318ab;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2c6dea4b5f52e1db1d2d0390f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb47f65a7f852a9db74b2aacc8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h900b4cb1909527a2546a3815c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd094ff959ec9948c4dfe06aec;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7ef83d834139dac3a4b7bc7ee;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9875f1038f2ac59887fdd1939;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5ee6018a1d869e51399f49ea4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he2944ef1ea52b4700a13a3d02;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7da95c539c42784e4d5a8d1b4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc8e3c44d520bd28077afe5bc0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h66352aa1b6154b9612d70e516;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he8f95b5eda1df153d51bca6aa;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf4b2d2fa78d075a554c2373fc;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb7b8301dd3df72b81c2d98fb3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h45aae2ef6eb0036b3407af62;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he8a205d52b58458dad862a90f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h74d5d99a8450c1d681214075b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h17a75119ea97faf6d72616837;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf2c5cdc1da66407b96422b0d0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h92743ba22dca708cd964b5906;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8b0d5f2a67d547e70d80bde8d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdf2e7314b881d9ccd2b9e6459;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb488faf235b27b3416d0a9402;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h205020feda202f3884c9591c7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hcbcf748e715cc3e2162f605a5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he3f1ccdec1f1c006b0c0aaa03;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfeb7c9c804d868d795acb1a6e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hde0fe5db30f6849197d3159a9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h588a542ea89c2e0aba6823c24;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4be79b5ce2d218501933cf4d2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h42eb585c007876002f230a24a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdaa446ccbe4a108cdc77a5054;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc2ac99cacc0ce3f28c1d8548c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfa426e4823486a2354952b44e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h68012caae59d5481435388de9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1cd0915292e0e7e62395cb317;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2767e52d1e8a65a78b742019f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h14f4c79313d51844cf5da38f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5835caf12bc3266b8471870af;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he31f6ee0f4edd98015b944bde;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3dce2a9267751c75c413aeba9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9964488e80267f3e89c537955;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7e80579a17be45224d1481dd9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5847d605b10726c3d2a0b362c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf159301d09533692fb11e33c2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h678e9eaec43e2576944607a4f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb968f71a9a6e142a4792de57b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf409cbbda13661e3fb9a4a10f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h891700fa3ff89cac5af6d92a1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf9c29f619337dea3b5ded167b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf75dec33a4e8b33d78470b3dc;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd7eaa3c615b2992ab8dd7a5c5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hcefe9c094c3f0388b90eef30d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha6560729907521b6229470c18;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h434114b94af3ac1dd5d489d4c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he2a25669ba4247a2241cbb7a5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'haf7700942bbac2f05b9d08743;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdbe8be12db10ef1bf51c79c42;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdc5412326db7f705ea8d72ee6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h238f8274f1e53e48db6dc2008;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd85043892fa6f2ce678b2fd8e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h75464f90a2032053e6ab5cb89;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7f403f07bdfff33f1ea8d94c4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc93d6858793a6ebd566a3d55f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6ddcc2b796f48c4a99eb1be63;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h984fce3ce4ca62de95b5f13c5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h14698d2c3b545973b63999985;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h90edb557fc99fce0b22eb4061;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbfb3cc2ff9d434f9e9b713e6e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9d0776e139aeefe235e9aeba9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'haeb08bfc6176669c23417a54d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h91e6be9c1aebf06e5fa76c3d0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd4f21f22b889934e3a686c01a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'haa7842389c43cc0d77f31e203;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6414ed80388fe92ff73e79bca;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h237036822f4b1772382770bdc;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5f4e7689b7e3804c68bb24032;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7267a4ff38609745db3f8666b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5baf579dce5d63905f166aaac;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h26d552ccbda1f32db64fa712;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he76f32f807b4b6a06e7c73ec3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h721b1920a5132ff9fa48e3d4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8c71b3b418b5226d432573b60;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc1d4add30cc35e5c9e9e134f6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1a641de943002508291137199;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h85f3a60a3e40128ceed38e1a1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hea34de85c4f4a8719e0528605;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd38cc5650e11324d997df4fcf;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf9206bbbacb6941cd175253f6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h25a6ae880207f9469dc335058;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb31baa7ee80abf958fe52b730;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h61210c54ff90e356f3ae43007;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h31c81113a44e3252ef19df344;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1c62131f64f50d2cc04547b49;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2d286a3520b3a0c03fa749cd1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf52eb5c4741156dc82feafab;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h786e60fe1291d1009ef7a2bcb;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3f616b1ed502f326a1db96c98;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2ca1eafb7b7fd2f83d47342c2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9bd7dd3f0d8e56d4f2c194ccd;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h82159e39c878dceeeb59c51e0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha739abfce4f70b236d32f2ee2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h589acb98fb956fd2fc6889a1b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc146997e6969eca3636e3cc15;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h65b120b9457f39464ead01c18;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc81a06632effbfd351b03b7dd;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he6b0765a734010fda26f75876;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h144c9ba7bcaeb1ae6bb0d5335;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9ce75dd3a599a16342b2a91ea;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdbf23ec00df66016bfa7459e1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha425b2041a826b6846974926c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd37f0bd33342b09ad79102b95;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he0f0250bc096352042707591f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6d31aff840c75eb9fecf21aa1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb0f316f40cdd59d39cca7361;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd05b456f6fcd648070a6d6c98;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h57451ce3150cc0102861ec9a2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd302beca88776940256161de7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hcdb1b3e45b83b796b0e32594a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h11ab58139af9a1477a46e82b7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h12c3fd43586e2c8a4922186be;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc4a913fb1651fd65d7afd8b22;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h71ceb2411d6d7e4521b013428;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4420c844c76a10d0e61d05100;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h87e190ea9c13af70a0ac21cf;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb0204a81372e2e81662f4ce75;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc3ffadd6d75454ef7a2533eb0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd2a51069fe4bca1bfb6f363e6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'haf01f7ff153d15a43c0b6673;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he335aa40be785024da9c3d5cd;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6069150f64e07beee25df5d3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8352e50cc0b373ac013e99edc;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h787a131dd138230db4d6ad6c8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he5897c9fe90f9a73fc5232611;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6359a83ec33f46b6b36c784dd;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb01fbe49ef42a634fb5668c16;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hba85fc343bbc5d463d2e5547d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf945debb3ddfca5813f9a0e4d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h912a6e2cb121949208ba469ae;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h728df2084ff213bca1342996d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he9afe4407eec38ce0ad231ffe;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd512c63ec33408ebb3ca30ce2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6bfa3e1aef7486ab8b6964219;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8b5c58b4f9d2287755d650c65;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he7ebfb71a90e964b19b015204;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h18c7dcc3eb019bc347da989e9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf935149e8580052ae4fe4b8d9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h424f9bd0fb8fa8462ad937fb4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h42c03ba5355180ee986a98ef5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h98cead6e730324150cfbc2415;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfc0781b30a9dfd4d5a847838;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf08abf6fe7ff4f8a9efe32232;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h93c4509bc8439b7c920a9bd98;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha2f9b2ef33b95b24716c0f16e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h53e7668ed8e5f2b5fe9e6628b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9807cb9f1db9fe8ca065d00d7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h14f3387cbd1b6bfef7c6c8177;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6a9d02c582e9a35b0fb8990a3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfb0d5ea9015fe52d3b4a712de;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6bb29cb15e5abedaf17b1c276;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'habfd67c5acbde3b4ef62663a6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1d6013e4c860a5569c5c63a26;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h17143ea1f56555789a15d5fdb;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha3861bafa439e4e8d8dd26066;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h229205d21256ba469b9907797;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfc46c56ed39765e1bf01b6fe0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h98fa7ad3b75281c44c6c2207;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h35fb505b1832fc94d240cea83;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h455ba661478d9f9fa1ab54d4e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfc89ddd65ced785fbaaf4f1dd;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h16c807ab574e1a5b4b39b58e4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3a49c6e8d813361ebff25cc6f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h18b8482d0f66c1f6d0cbf3c4f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h901467bfec578aa912f0a2bed;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3a3f3aa00c2c3e11be43caf9a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h812650f6700f3abb0545eb2fc;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb5bc0e5d934c59dea54f7ca8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h244580ad9bc0684a5ad647e9b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hcec695a3c9cede7b40b49c0e9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdbe7b0c670ac432b66df40f30;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6252bbc7ff59a98a1e2efe2c1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1688873a553606276b06a24de;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc7858226d84accb46896b72b6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7e98f596a97d47fca0424c55f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hcd9c4940277c437c69be4ab4c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd9a1af608b1e0f93ece570f3e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf362f6f9a7ab59800dce7c795;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf37f08abbc8b07cfa601cf8ba;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4ecfc2b54eecc1e60341b646c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8b3bb6559eb4a564933cec3fa;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h466d9ab46ad7c1f536cce2775;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hce243da0bb616edd3b10308c4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h99d38125fee71ab5ec2442300;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hab0a21910fdafcb14fd89c08c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc7c9c7319d6444d3ea7e637e2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h619d1e9ca49254457125ff740;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h53294c9987069cfa7d22c7e35;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h792fe5ebd71ca4e1b232fd27;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9c193f191e7c255459a5ca409;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h13ef1a10604888677c1634b9d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdf888a1bd29a965eae1894564;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2a6d9c9c59be7effa080a2aba;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd8bbd40e3ca2348b6507a057;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha5659c151f66479a5e8535c58;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h87087141dc2e43cb10739e7b0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h43716908ca9ab366dba14562c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha10b08985f62e479544931cc1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf82c15fe77e16566d4d10ad5e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h104dbbfe0535c1da0a3e9f5e9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hac8ce846bacaed0a345651575;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h16943fdfd17583683a185ba92;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbb3a8bcb6a0a45f456b76096;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'heae9655b24f06799c0521cbaf;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3f186b48d519bd66fab2e59e8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he7c950a8e7d96a1c608ef43fb;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h805bd41034bbe9e36fae16e62;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hefa718f4870fd5e1d593e9494;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha61824397cd6ec5419dd51328;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2677b37f2a02957abe5cf0995;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h19dca5f1f7dd34f4bf3b26fdd;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha84334012e385432a2ca1eba;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h74e7dc51dcf30b3ad0e3cfee4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5fb0421259feedbd5d1c70fb7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he8776d2dcabed0fee1b368ea2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5dd0e19df7de320a268786f44;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h75afcbcdd19f20e05f1102a17;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h84c94366eb9dcf5a1819abf30;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3aff400691ff0346f6a11d9e2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb38ee6159bf36a3f4011071c0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9c5ae1b8e3f21a308146275a6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he9a9a650a9ccaa5dcb168c3bc;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he4fe890536377b9c8b1a066a9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h75aec65f166d004a60175c72a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h969ddbf00e2d79f5c66cf386d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7e7df678be7b5d2710e320566;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h527e82389240f4c23dceddda3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h149bd4ee7ad6f1ada537cf2e3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf783a51e663403c0b6dac1674;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9a88e9211d2bbea63d9e344da;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h998b560529896423ac66890c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h608cc7535353e8a62f3cfd84c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h948d7d0f079b482d2be1c5bcf;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h61530f122ca64bfe1ecb11f68;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h57cdcb98ec3e711042dd0e586;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h78d53f902cb5a28c693a05cad;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2478d3b7ff9e699f027488a94;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5e1aff4bef9a13d72365c13b9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9a7e0f3b3b2ab635b1ba434a4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9e1b296a5d3aa9dc844bdcae3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hae01c2401a315b207131d9c8e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h45d6b47b58c656260ee965802;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h70874d6b8116a13892c63a5d8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hce217d456385103e5373282d6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h789a5d3f99e3e5102341dacb3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h79a6eb7754657acea3aa8eb02;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc21c3d5a61420900b0d19fd30;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9148c497735c1fc0b01d5052e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h396511c445221ece6c2388763;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2e90434e05f38ada88217eaf4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc0ba721fab8282e1188f31058;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h175e964d3c46129084b304507;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3c5c8e1e0d65dbf730da9fc00;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7fd2686d1879fde35a8b0db73;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hcd5e3b0afcb4298409768cf4e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he4f82573d1c114121a0a2927;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he0b71757f5980851b5518dc87;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3dd5ca2b8e6dfae6370d48510;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfe21e3327935908c54fedbad3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2d8567b343f501da94393f386;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8b978cdeb9eb418a22d480296;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6ed4fe5d4c50756ada10c0949;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h400a8aae7763c8ea82e86802f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h78f66df11ee0e52d39d7044b0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9496fda792c468d5b33a6d3a4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6f1c50841e1daa45cfd263d91;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h98c141284c97702bf9cfc0ac6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha94df92fc386c5c616408fd7c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd2cdcb815f5e1ebcff9cb3f15;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h191da22dffa0c96e2d212674d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1f9757e39ad8e829cd149f573;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4e9b75f3abb37e58241ea56bf;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h42dfb60492a366749d870c635;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3ee072b95f388b64fe5842fa4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hae5990c1c3af6c7f53590543c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h56cd5f50357c9c26d2dda0781;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h95022ed8a610e1e480e777b58;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2639a036b93baa683554231f7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h193d3087b4e3c40f92160a5d7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1588ebaa38bedf0d4edc216ea;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc97bc8d50fb406196cf55686a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd7cd872db5393a756b7d57c97;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd9701e61f3ba39aa57f813e0a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hde34e606941a53ad07aacc7d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h688751e7188ca052a128af57f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6966131028d04081409047c46;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc70b679d228ec21593dc676c0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h502f50a77d7ff2c56acc207d3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1eba8abac5fc9503013dc2cbf;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6952610c34b760bfdf22a4206;
        #1
        $finish();
    end
endmodule
