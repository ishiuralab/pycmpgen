module testbench();
    reg [17:0] src0;
    reg [17:0] src1;
    reg [17:0] src2;
    reg [17:0] src3;
    reg [17:0] src4;
    reg [17:0] src5;
    reg [17:0] src6;
    reg [17:0] src7;
    reg [17:0] src8;
    reg [17:0] src9;
    reg [17:0] src10;
    reg [17:0] src11;
    reg [17:0] src12;
    reg [17:0] src13;
    reg [17:0] src14;
    reg [17:0] src15;
    reg [17:0] src16;
    reg [17:0] src17;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [22:0] srcsum;
    wire [22:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13] + src0[14] + src0[15] + src0[16] + src0[17])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13] + src1[14] + src1[15] + src1[16] + src1[17])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13] + src2[14] + src2[15] + src2[16] + src2[17])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13] + src3[14] + src3[15] + src3[16] + src3[17])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13] + src4[14] + src4[15] + src4[16] + src4[17])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13] + src5[14] + src5[15] + src5[16] + src5[17])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13] + src6[14] + src6[15] + src6[16] + src6[17])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13] + src7[14] + src7[15] + src7[16] + src7[17])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13] + src8[14] + src8[15] + src8[16] + src8[17])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13] + src9[14] + src9[15] + src9[16] + src9[17])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13] + src10[14] + src10[15] + src10[16] + src10[17])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13] + src11[14] + src11[15] + src11[16] + src11[17])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12] + src12[13] + src12[14] + src12[15] + src12[16] + src12[17])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13] + src13[14] + src13[15] + src13[16] + src13[17])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14] + src14[15] + src14[16] + src14[17])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15] + src15[16] + src15[17])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16] + src16[17])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17])<<17);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h0;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h65c90701a33e882eef8e329e88ab8aa7fcb16e4ee706535c9a0c79c43768601d86fa3cdc6817a5959;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf2b9d5d7e5e56cbc7563c26058beb13a25e39c4b08193ea9bc697c2e664b3cdf25fb944ab17fd53fc;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3aa35bf5dd7e2c9f0ae526b56663df66d977b77113fa33271ac38ceb40498fae5652e62e0916574e1;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h99dd4a5fd25c5e48397c89d004d5959ba9bea71ceabf07be7874807a4dce4d890606a0a263b9610a8;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h47814adc81b97707ce8a5e43ae095e354c916d341440cfd1c3def6d293439e60a328042d261dae90;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h48f9970ddb5070a1ccf3145c13d2aca49029bc0cceb2c49eea2cb8337fc7174cbf3c88543d68c73b8;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h173901b6229f71ead4d1fcde5f47494d82d4890c6fbec276592b390252726f93503d0da3ccb219b26;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcbdf0ad7f36a0f127769d8741748930a7b4b395dd73af6279d832870244fabcbea5bbde83ddc68be0;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h37c61946b18433da3ba4c44c78cf79473f990d2eeec1adbc68a937de6b37a9cc37219f79ed9f0817f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc99ec6748a883527c79fd9523cee09773d18a93fd0cb4c2e303f14543dbfb752f3964bc6a114a8beb;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1cf70297248ce2aaceddbf0fc0d044184348dbeb4fd0292dc0330dfb781f533b1eb100bc1b3bbbcfb;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcb0d866515a839391db9154f5b0db84816b7d95e7a6f41f1766a06f3a1bd472302a383d33d3f45aad;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he0ec92b6199a3d0726274f61438ff3101c7398ab27331c4f2ef1e990689c48d39b7d025667e1510c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1e409e9f4589b720c5892f45c5f6a9835c3ed3df3d34a2bd1ae577c3b41e22318bc277fe9edfa81a9;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd185d9f5364214866cfa3a0aee9320f97e9314e8b114d7b21bb903598276deadfe65f5bc218da6fdc;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4bc0a48e429d8bda195df5f084e53d1255dc03dcf0e3283fdbbc1d4a8ab6df020c21db43fb9146ec2;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h318c05ed4290f74ab6bd5d60a02795cda438d1626f1eb7f95894e885816c0c8d0a49ec9e6455f923a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hba5718cbb3fc5be8812b997521847f41a79c8d1cc3cf0255396ea7b8de653f1893227e4205c355c92;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h74342ce101fa2462fbac4d3a302a450f6f8b3e4645caff79dc75344fd684c11510093b13804e1c697;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h213debe02a89d4c8fd79de223cc6d6265681281412d2767e57cc6720215a2802e45fe15fd22de136c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9136d42edbdd8ea1f7809711838a9071cdac0b7f9c9907233fad7006037065483054d7906b5ccfc4e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h969aa266ecb12fc245b4c3276d7a8798410758558320c591261a86b5c44ca6b3edd54f20fca25541f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcb78e809fe7a036a9605fbaeb720f07263af31b1a0bd08e5d3ded80710221db22a5973542c6b12784;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7d958ea65f07f8da4591e8034968eea20af9a6a7277824d03d2fde37d6431ae132da121bd0669ccdc;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7f0c54e32ad875a8fbf930d496fef235faa67d190658b860a0b4360bbe1f757bfef7e8a9c8f461626;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h725756b005ee959d9e8ea7cc08f113ea8e5ad6dda37f591bda017b4dd31b414035b66cf98aa70bbd2;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6877e2d0744794d26f25bd5bc76421fd2afa6dd509d07dd1d2d4b1a83ac155ce8a8c7a080285bc279;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbd37f8fdc0b139baa1cb991091895eec6ebdcafd73fcb7018a3aaec8e68794e918ef0c651d7fd457;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6943f3f7113adb094c59fd5cb939acb05733d5da568de854481faedd7f730dbe46ffb9c61092cb761;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc3d35bca6365821b622d41bc7a379e6a7380d33576c5cc49da20d174e7c14f8a9e0c4d928d953f21;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hefd98326d9d7ec4b1c5d7b8e6d29f34f74470293531038b2368c48ac35e6c9bccd13423982d0b7eb4;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcd94bb436feae5aad90bbc6e4df8f6b789cebd5147f8e3bbf8637daf6e531b523fa7f55c11e32acc0;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb8356b97a5518b66b1fc27bf9b3151bc8bf3b786b6e51ab705485216580fce32078a6f2826be440ad;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd195f4d84d5165efc8faa751fedeccb18d3aa899de844d49a2933298fd69eb31b7c65ed5ec33e2c61;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h797154138e75ae739d5dd1ec118709ef95b855135accc5c6087f3b8a8909eeb98efaeaea336b9e7e6;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5122bc6e702d68590419fb626d21099acf104957fe669140cc1943caa8995596664e9790e468e1e6e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6d2fe41d0dd8e7f9d7a0302b6d170917f5534139fe7e0d8b497c1e118dee7ad0c479a906c990ad20e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd5f6d83bf198b2e650a3e90e81889a3cca8b3825c72a2754c1ce4ad1d9f4df3c6589ab6ded8d7f9e4;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb0aae07096b1e0a41a64dd2722012d3c9f65f646be5ec0f934e390a8db223e598eec5f32a366b18;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6b443e56b4bf26dc5e3d8bf64bdf2ef2c41be21d2b9d17d66a5b00adac3c4917229c46b29beaa460c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6b263d954ffd7b23fec9d5f882d23c242a5c39272af43c1808a2d6df156bab826a073ff89ffd8543b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfe4358e44670d349f19dd56006b86f8f296253420635cc903b656f45482f02b7e2d81b2df9a9174be;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h29bed977ac8646d0b45447ebaafcead701d0712b265c122de7365b614f414fa58dd88118a4dff014a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h388454de4684f17660c100c1763fff709a24900ed7145cd57198f164a1d37d3da4e91dd4e4390e7c6;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5a33c110c3bbae2bf241e8f3ac3754d82b58fa55a831b61d1a9c4b46d131975a89ae2d40f5280383d;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9528ebed75d0c066174a16e5c3eb4e965f14cc127d528214fe272b601c0063c230978218b93228384;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h341759ae3a96c717a9b7508938972213b6318e199281b25de5ce5a4ac190dd08b696cf62c443c8565;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5906d676e8f9ec0e1af95af8603c54ba3125859c1cee86dfdb420deff1f3a92b7138bb543175b8171;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcd1febacdab8c8234aef8eab4c997cb72890f64271694c75f3beb539be341f01ea4c2abb374ea12e7;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2126b400b4c59f3a8a0b98e49f8956d751f714e1f0ed80ba69773c3ae0a6cdb05f1c4396a1fc5a079;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha39bc38acfb309b9a0367672362dfd95f6033422384623ea0faebecfa273a426a4e450821d0be7e2b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5e79d2ee59ca087c880e133c03926ad4d8174e7066a400ab61813c0123eb2b7c45f5c90b5fe4e784a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hded32a6c9538d96dfea4a10b609543af0fa7ceae3ebc5f0ea3cea9c1c34c4389679421a50403a5e0e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcf7e01525366b7ddc9d88cfbb79f562b0f3823ed0e1f91837f9c877bbf0ea1694b0b5ac72c7eb0c60;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8c2aa0f5cdc3952a14d6d9ad033902cc8f7601d010d696f528631d34b388c1e78dfdab6dc1065e57c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h893e49c4f7d3f635c2cad2907e9444d5ebf9562de7eff2b5fc890f1c015bde803b8a0599d2ac2b77f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha763909e7b7172a86935e1f9b4ed0aa4382214e5fa591740a95588c565c5a8816722d1c5e2b2d3ae3;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcfee2ece1d2733764a5bd80ab49bcf7a008e1b9f0bba7dd8af9c1ed5c78e5da1495af44994bab57dd;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb6b3e2eb1fd811a0fa265b44d10c36472c916fb2a166f225b2faf232b94505c465d6b8ae4786805a2;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3393b27f5b1ddacb9693925924786fb3275eb70e10f46faeccaaaa0f15404d28efa57b0d6cdb821d1;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3f4ea8e64f269e595b38e330f12df9a71fe95a6780a773f04b3395f83697ec8e480268167af44b4ea;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h40b054ad7ea5721bb650835a3a9f437334ef329b9ee5629cb2ef6f4086e6f1005593605965095115c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h49631f0e4f7dec49f1a4860eb5ef66779eb243bae3f65ddd1b4608560aa1583addabf8759bcdec117;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4b6ad49a92fb1954ac37be33515666e5ecb31ed07f404f9836179b746fe27c1e1c633924f2d7cfa5e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h90c27c959e5a2dd4715179aaa34e9dba7d8a09ddc3297c523277728c3636b793cbff1c64d341871ad;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb4b69a3c49065c96e2f07351050fdc5281780282a4b418f09a27c0b4b70f94f7c8aaec20992c8e589;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcbfc984be2689406b2609cf3045b00c9d3be0aab9036cf14642fe4416fa1b4c4de1d0f0df61b37905;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h600ba121423df65e61d338aeebbf8085d36f3c363e193f11e4205af30020e605efb4a3d70a0113389;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6df904faa45d920d6ca8d0f00cfc6f3fd185b119e10410eb456ab1a946c77392087e56f618fdd587e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he50c863398991086aac8efc7203c86c0c954e617699885f30f1ff43119ba8a1dc4c7c70899290eb25;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5837de75440a09f8f37166af0f6d1362b61362a48fe97af09d2140debd3412aace27eec8188954817;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h54c5af03cf479bba1cb692d3d7d55195291a29fb8eae6205fd483bda834c0d40e8001ca1ea9f115ba;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc7ff6c874e31629f8d665d0054d5ff21d5586f8b5d3efdcd4f401d11d066abdec6a064db15d0696f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5c1ceaedb1a45bf7b4aa3bbc523be886c099d17d0c90a0b24d540da43acd4222e6deac93dd6175c1b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3d78521fd93fdba60a467c6a02b346615fe61e744c23e4f724bf053cc742cccaef35e682ebd4ec51b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8ecb2656c902bc39fb16070d4b9402d067165368dd4b2e9c88b23e9cc34cb482f048705b04c324125;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h54c116670d0671bfb6269279dce0fb8b6d8182ca943af98aa42d056a4c1d6dbf23403125ffeafe6c3;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3ddd39535ba9a392a437ac82f127f65650a80bcf35cb9fef3752ba3bff086e41ba869bdd82092fe1a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h80c6b3cdc8e35b416c4bbc3c4727cdf37f7c447be442fad4ca596f0ea95aa473ee6c6ae72e05ea12;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he9e509c91e14caa128c213a2352786433e0aa0a0eeef2301d482c6fae7bd21d23a29964bb08bbe3b1;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5526e388b4babc2c023a321d47eee162d11c58b386a193786917e4d471a3db6016a6af7ff31893b13;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb58a3f079c35bd93ade2347f51c54b0c44f8f650782d8f9d85c538354c59e3653c1bb68da51a08d91;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h94db88b08c5bb2d51ef13f0bfb73bda460e415549d5cc434b7839af2a193a74aef58ae36883267cde;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2f9ebecd4a4ea324d9004abc7437aa2fe162202a2f4e328324009e2142368327a7b5170729edd41fa;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9fa3d06b4dbee42a48ad2e7f8b7ffce03e3ad8e403d35c340e6ce96d227f1058b7e1dfa651c4804d2;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4a94ec22f7fb3565c784f8f18368591b9ae5a3ea4b28eced610225ed440fdd3c1872cf40fa5d2f6ed;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6d5b1975d491f72711b454f783dcba1f8501ab2bf1cfcdc164a75b7988858ac04279431701d9fc4e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h831f4aeb89e0cc6db5330edd584586b7a1cb31023970af137279db2e5d8cea4109e13ec4e8f011d85;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h69d3781167e394733914382eeabec267a64e91fe99ecbaaf79d2d67ac489c299a64046d0fe07673b0;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc44f31970d7817a972954996eb81db74cabce6f4dc33d4c8240e68888298c4ecf8edd490050742f7a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfe01af5ae494ebddccc9bc9efeb12286f752cc6bfaf6832a53354b259ec2b9243a4e51dfa75d348da;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd0181c8e1b1357960e134c3c0acda7fdcedbbcb3c4340e7453f2c2b1cc772ad6fe9db50dffe1f5bac;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7f8448ba12a3aa34354622d5b9a0dcd7f35c7d1f3f9d521b221573b06a6878ae82e9976fdf615276;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb3e85d1d3a47094d53acc4980f89782486c7609cb193615ff19f4731b75f338e527984f61698f7a60;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb6e87dddf97fa08f97d8677ce7da5ae706295e89256c3b3710000c36544ae9a0332068a4298723eb3;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h538b4bc5f05753e9e6a517f6ad89cd9ac051075b9c98f205e2f1f184bbf0c9c1af86557440fba4166;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfe48c6ea4856e54e884a4a933ad3d34c2253db0cb7f5254483718aba890c3d20548cc9512c94f0988;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4ee46d407352c55170fdad032aab3e68d356fba50c0464406fef24161bb3714e657b383f153c298eb;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5f4703c5820cb372e781fff82099e05af4900b27ae9712dde41f5df17b9963f3691e8572dbb205611;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5223a8f6dca47109a5aaaa083d54d7abaf0659b41d9fad0a76a7b4dd66f539f605d1df2e7a5a290e9;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7fbbd45974e0ce7b176775473d50a48265a3b483b32eda4d634f8a8d8b62195464974ff4aab47de8f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha7299902a7b1af5b2949b9879cd6b3ec5f7c78fe2a86d5d8000e148fd5c60ef43d2c73dde697bdcb2;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd97f7c832a00b9ec4b9695ede99615bfb0ac6b9b6d545801bfb99c751d65b65ea4a137aa43c82b366;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb8f7c92a3f09b814ed185c55d2da690811b65786f469268b27c70a7f178418fd6d7f2fdf8f3d5c1b7;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc861d23246919de11e54b9f83203da9ed9bbb522fda91cf59bb7245ae5a8f6d74128a81e8ce67288e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9943d8380fa9cee1fe8c987569f65209fba1b407d0b5de96d623b67426e371fb0eff820d493e80415;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6eb2d7372a693aded8ef884d51f5d244a359dffb0850052389ff44bc3d0b2d2227f44d777d74005ca;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h18d26bf320d8a68275d7bbb248712c7139e8e12191aab2403094cac88436c20c7ba021f21e3d13f94;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4cd05ea7045583fbb5184c49bdaab026cd383a10bbc6aed845963aca6f052c7ffbf22ea3d396beb4a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcab70760a71d2165be9274b51c49017480c427b2632638a679cec72f873763fd325e60120ada4bfd8;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6e772b335dcc397fd945b7a5385338d47f24537a99629aa03af7cffc5ed7c2f55344a7188dfdd1ea;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hdc6608459e7df87d729686c3d5aaa8951099ee65496975cff1011fa7387f5fce24c399341cb53768f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h76aa83665eda74680f9370d985645246fe06d6a376d2eba74e7f60eed14ede0404b21ec05a047f135;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h83a96956b0edecd67470888b382408ddb5cb47aa4d36090a428db0c55d7c2438cf966f73204336eb3;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h37bc41c36b87d87e7eb4bc073ac5c4694ed29f93efc245e6c951ab5f4e5b71cd67362230c2db7eddc;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7fa770cb699d8855b7d3ec6628561a026d722d78bfbaeee202557edb3f5c1549336bf97317073c050;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h689c3dc1f2f24931141a386ddfa6566d294d7076c25013981efac5d022a2e2ed0eb16711755836a31;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd1fd14ce9291cd99ddfacc35ef93bf814251e58bc2e2417594df00634f9ba48e23666909e670aa848;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6f4efc80edd7bc3244a056a290b1683114642cc7b024a149ab9a0ef79d2378c694cd6957b2000282d;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h804c5e2ebf3d50f66a83aeffc27aef9873263a1aa9f865a3b386d4bae8e9fd7853ea7d6ba7989d708;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc50015155968e4d207dca73442892d9fd5261c26a221cf0e6a5a8fbf9571d4734cbc41a23808a7523;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2255022299615e992882d0e6c1242676e67a3f82ce390cc60f37bd2b452c1a00b1c7dc0370e0d4e8c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hafe973a6788f2f1d28389612eac6d907395dc3329adfe0bd7e76ff77685abf0dc00ea7062d8923acc;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hac694df1b2be84849854c32105d7377a0add6600b6d660773e2cfb60af2d3cacadd26d3e887e14ecb;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5cb17d008879bc9a6f41cce4cef68f314d9d40b049ee79dc9449be6cd656ea67a36f3e5c0750e4782;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3ecda855aafd538ba2772054ecb1509e3bc6ce6166d8ead4cd19d9066be1dfaf0a42c5e151dacb230;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9e580e556a64c880a35f366b469ba8eaf2ba741681ae868a53e07f67344c0a75ebd2f76fde2980ad1;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc65ae941041af17d272b29e989f52bfac090cf76ae6ce76f9865ae05943925fcaf165655f5648da92;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfe656c9645f9b95a695dce8fcc385ebf77da6a270ab7ff7d89ae29eccf00d706a69040fb34e89caf7;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6b4f9b655822c7b8e8cc3a85c188964b9660bca70dfefd684dd8278e2df40b4d4fcc8b105de572515;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h681a4a1416619d478bad58670963d746e29867589576eb098e1ebc4f19ab2520db3230a60d8f612d2;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h51a39aba4318d2d0a125dd66025e77763ef9a3f7a8770efbc04806fbda1fc1b1c107c54e48b53754a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h14f3221484fc0527ba7bfe6043fab6c42bd3b2c4675ef76411af31251a11d3bda3437ab53f67bff17;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1f181629ae6963f779d62f4fe96c3a4cb6a21f8faaccd7c1afd5fca239958039e536e2b230049a71f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6c0502c165917f125e2d4fcc5819872d307b3f67ad62815a4fa5afc87c2312e40597140857e178af9;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc138bd77be9dee405f8ce54b5899d8597d2cb088b2c35d8ab8603b571511f73d1ccba06a46d194b78;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h54883c4c5cd79fd88ae3706487ca6a8e49a9a0bfb4568031b25d3e755dcf1705b39febea1a966bbe5;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h27a0be2040633d4b8688c196c24d8d6039058d30a89edcafbcefe709c600f4ca4146821b5f012ade1;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5018163d4f017468c6fa48c76ce1b8104a720f6d0a7fde692c618e9b8767cd496444fc0c9eb7be512;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9a781af1f723a19ef55bb96f59d4e2af07e4fbfa0ff5f07835fce4af248b2b42184f792dfd8b089d;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hed11dd2885c57aa137b1a84b0f41814b1ef780787b8d7811cc462ecbf0220c30000fc9e3ff7d4f48f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h77cf41150af68c8db328ea691a81682f2243da5d1ccff7bd52175ba3dfb770dbfc49e682d533ee0e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h157bbb3df8bc4937c14c974733e6cfc33b66ed0be4b43ebdd340049137cd49de839aa68f90245ecab;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbaaa612c1cd8d3d41a715e803d4f4edd5f7e47273b6b419cd32d258fdb774760a2078466db90580f4;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he9bb07a6621498444ac2f55d6ee8acbe0fbedb7b3e342533cd6846d53ad6f89d051b647b8ff69c7b9;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb67e4a799538f8b3bc495411331f7c089df0e990f4e9e9a7afe22322ccc784fb4b0b900b34ddc50f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h57d83072dfa283d574771ba9bc60501a9521cc434c739d5923b5b0fc4bff6a63801eea5c4248b51e2;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h26b60f7b7cf18b6f24d49c9a1daa802b27cb8083bd9ee9d66d30f92538acc5720e0dde88f5b281095;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2bba8081000e119d6925201f155f29dcb09002ba8737648af1790f6c738b50d5ab99fa05944d9d8db;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2b1d0a4cf47af85764f8ed67bbdbadae606c770a48d89ad90d3323aeef491f430308b064ed2ed44df;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc5586fb0f7973a58f335f3deba4b6dc02488366e8072e5252c56e5896bda200f21b3d6d73cc72bcce;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfa73477c1018f2ea43ddbe3e8060a4a6b06343b4676aff2411227fed46929ff0e8090b85775986d76;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h18b71ed56edd3f580936bebf176968589ad4a3fc5b9665391f8280e182e81d1500bcfd5e89e2728b2;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha56db963897a4f8fe73c4aa80b4d3339767636593d203914deea7b266a6b417b49ec9a02cc617e3ae;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h51f5bd089271910ba1c663a0f08f79954472a6ba5d36f0c894711557a30e8b97c61d6d9f26199294;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h87224cf459809b2902157a7ad4a6a3a3ef42f5b29c4f07a4122b5995d8f25daf7be98bf5b536ecd5b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h70d6c68079e286b0b2829baa37d11061a972e0c7f155291e9353d2ba5215e82a9767d2a025bcc124d;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h90e54588ec1b35603f3db91c18efceb09891de4f54c82786f7884a89116db4dd367f6a9ddaec13df;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h467743743d1dfa62fc1b468c8fd06032ba69ae4d4b838af25d40d3da2816150b8b254b599df864c7e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h217c823a58bf3cfc072c728d65dc586f2ee84df85685f9a6a766d852e3e3789b55c94b1167d1653ff;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hffd5c0e30c121d06b50dc0324eeb03b05b1f9a12dbe0de67531834a25db98b7739dee705e14fc235d;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h64212427a060abf5ea29c6d9287ec76f99d5a093899a2a4f9cb3bd289f5d445723c616104eb394cdd;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha1b4052f51e3454f45251224952717eab1aec4fce1477ad2317a8f499fe6412729b060d4d2c65f259;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h75b01f5d4c3cb9de15a48ad0db8cfa79e414d099909acfda8f20a74747c8ac0ee500b09a333defbe9;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h682b5a70db20e02450a8dc075768c6f43523917eb51741ac237cd56b36c54e2a7b1969929960f8f07;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8d0404d40ad2ac7870f2f3f1b542b7991159ac89717a7c98e47abfd277497eab1a350ffa6c6c91d8c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h72c6fa6c3bd6feeb6f66ef806dcc055a89fb0e1eea435a75a1cbfa07b4d4e4a0e52673da874df30d6;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he9d491a493bf3266e21c67fc57a7037cdb2b94819e3151ea276848f65d7d06799fed70c82ec117f6a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6a73f50e8dc3706fa143fbbc34c5b84e43c8a2120afbd8541abdf5d0cfd9e5b752c0f105d9fcfd724;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc38d3549907525ff753eedcc9dcd2040bfd2d640c1715b7f07ce946003c5540056da8cf226792c701;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h777e67cf2ee9cc0c82d4d6598bdf523296957ab1395143d7e83aa3881fabc20b0ffb1a7a224d324a3;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h853a4ed3953ac7ff850a6a98982636b52829f4885a5354f66bca297f4dda5d36a05a007c6508a6d29;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6794e512a77df44d9ca9c45a71a7ee503bebe89ed555ddea23684c537f60b4366d576d7fc2d85f828;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9e1d552d61c5151d8d83ccd16f73b94c48c5b47fb5e26b1ad2f0354366261ead59eabeee13af95704;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h511d7a7b86e1a3d80ddfc7a8c9106758a702c9642a22d8b6e59d7718ad80b24970b00ff3617ffaa6f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb921124a81d8ca7cf15237c086be1b32641b15575a8c7bfdd98351da5e329f0ae87b16da60203da66;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4d071373e3a7a2d64e250ecbb49b00bf9b3bd3736f62ae5a7bb1af761ae82ccaf11b2b6b2b91bb8ed;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h25b84aa13707a62cd5393efa70951cb98818df510a5ac010d3742f95a37374c11c2beeae46712d38d;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd5602036e5fc3a2750d3ad10d764b7ce8b40bf85c414af68fadad4123ecf547aaafa985b0adda936a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7dd54075b22610a8c1ac4573068c6075793d599bd49ecf0a4240a416c621c67293527efa6dac42bb8;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfcbb4b181fdff0c3c0975e84167df152d1c3517b3bd56ba165a3aa23933cafe7e33eaae61129c6dde;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4bdf953734419c4f4f59dbab92b1203b69a69df96be91c352fe3047c4d5c90d69a72c38c197810a84;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4c5eb3b5d3b2fa515b975a96f2f16083b7f205d03e41a1060cbaf6fb7a2429e9e703eacdb11ce7b39;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h914f5ac5f09ecefc6225196ce5fff7fe765e01e9c068d9783f740995593bc08fe50586f9e8ccf133f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h34b095b6ff4a39387847f828ab59eea59d000ca868a7d6f6f155d954161bea839f1c694eb6e968e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h443518c89cb2dbe082aafc57e1e81ec8c78eec19cbfea88cfdac71a12d38563a482bb7bc1c08c5b52;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hef71ab7825bd5c69c9df1363245e5fa643f3919e7989e55540936b5e18a8a75974e55339ed00b89f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8c97f5b235fe00a9b68506085749283dedab68004e07e86d123e4bdc26dc8fd99bfefa10919c2630b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6e46622e1376eba0a3d66cbd97641b0866d3b5d80e649317ab76315c8d4701aaa4a6dca161f7a089a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hec3dd830f0c52505f08b5e3286111af3f30d0f19502a6393d91660b6d3edffacab0122add79047129;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9e58c915650a9191aa78f6c82e12c594b0465aba4b8a6569041af35deb87ac6414417c54e5f07b6d8;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc586f24f9854ed23ccbb54b498d05a8c6bf1fa8e3de5b38a52b533b13d24f03cdd66cf3521ec9ead3;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2fdfa6f32cd3fa23c2f4b5686f92c803ea7faf7d81230396b1ff62f1faf7757d60655912f458d9fd5;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5fee38c79b5585a1548bb1d73657c6b91f387df8ac645c1aa6fd214dd4aed1e5fd153abfffba0b76d;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd1939e68bcdc98f5cdf66372c92127911fea55455d8c07281f52be75e3675d0771ee17a57f41a7472;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1284e4113ad8bf9bf514d042c1186ec09cee23963607d20c4d11631415055e5c0c436ab00915ea105;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8badc327103f0b9e37da7ef87337aa878847b2a1a2997e01d55b4a866b72fba782a249ce0ab2601c3;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf4ed3c3d678b09db83f67524031538100bcdc47e8ed0056d58be8d8a0fbf8632747c840972dc7052b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h861efff5d035a4cf48e41218b7dd387f2e8b485c34b9a77af1267a88023fdd1b6afe6b15418612fe3;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1f157d382ef21101dcb80cfbc3d91d438e516624f79b79ec9f1a86c4d0d2a5ea7e042482bfda70f9a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hab04baf79867362982ed604ab1791cd580d761bc94610095aa487e70f5104674b89dc73a06790361e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1b98650eeb7dd40da6f241d70f66a7000636827426ffd0ace22b705301d6476fea62d262e4a49285;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfd5dfc576a49abae71c73ef2b7a18667bc9bd38c2e840681fe31b94b4f962de2b3589ea71230c824e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1de7981e684e806186f8632e0ed572c1e2b0f0f60f4f3beccfbcb199f1b5fc08790d68f773227b9dc;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h59ad2ed5e72c83abfb4e56729f008ff5f8a1e0fa952d4f83b5f28a1bd1646e8761e691843bd801dd2;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb72500c519871e03f5623b59c030547d5a04b9188f9939d8fcf273b60e14ed88abe0c5766ffbae93;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha1bf4f78fbc8be8cabe7dffa91d3114521b2b51c96516fb371e10ed40ce9a1d4b4cd1e98e9a608af5;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h93c023b688ad35122cd2c974c6385993c17da2c0f8648d8e64f668ec753babc298dd76a9e0c7fe33e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h15890cc9bbf68f73b0e35c0c6d0955f8c53e87d0b005ee594d69a8d9444e5464d6776d236fa476ec3;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd482619f832b1d081b420e4c75c670b0c026f96040b9f7835e7a29507926258a874a76778ab88a5a8;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1917e3fe4b2f54e9adbac77cb8a77d40e4168d3787e5f7475585943f953c22d4a5ffdee01cd3f7100;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf260f66857dc4a8cd680704f25366d565008db895650c6f6f8de19a3226d10370df7713b84d1543dd;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha65fb27bde5e1b5268c2b21c13d78d895c45e8b193a4c3231e7b6b29e87df58817251d43e800bce7f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb6abf8e0a6718a0247b3cf4c889fe1883c8533d4ebd9a57fc2390dc5731f074cc15bf6709467eca51;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h61a25d154b6b1701653adaca9e64d4b47171e36a52611efd5e597065c0ce754b9f1e96fbea9544450;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h32b4c1f543fd80d85a5a6c06dca1c39872c551b359f040b2a1980d695a035c942bead35d0e0b54a04;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha5692377b5af58881a50e27cdf4caa04c6826d94c6f00491c87e5f3be841348e5d37e0290ceb2df61;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2a9a0d1a6730271bd9a8f1314334d40bf7b8260eafdcc3d730106814a54d2ed96540b3b5d01df8cc9;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h18642a69a82c3b88b23f76ae060420ddde13fd793f0f008b23ada54d7364f0da32b356b87cf300cf0;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he6f3d82653d679977e446ef0a573b3778df943604c5b3874a4cea4f0a2f1ad26aaf09a28f89b1d5b2;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h986f40e8e9baf12636bd9149d9dcc63b9d9122b998e23ddef6ee56b87d7bf1181ad7b8c2be47b9adc;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf403f51471e01c7383984b422ca6f4382a4215b5df2ab41a9f75a180db828ae43ba06177fce2af273;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2ea12797a3ec654fc59702f116aeda25feff4b8944838c4821435e0542fc7a8375483cb0523e0ecae;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb622a0a0119d4e306b0322709e413fba340bad30844acbb45c1e370327c88f8b6367edb1fad55bd75;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hdc22dc0047ad10be2a38541ea0db419b58dd9eb3ad9f4c4fef3fe24166b2928d17de74c1f14dca970;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8496df3128e25fbbc55dfa6faee5c4cc7a6540c7ff96ac8b45a09d2bde12d07d3df4712f9b55b738d;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2998429539fc95f348141db5b787ed1a564dc8362ced5a3ec11098aa163630fb617609c2ca8be7e8d;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc8d1fa2f895ee23ed6d85119f479d076711980c8022ef2f132f4564259f7be952c60824aeb9877a54;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h52ab598e2b887a23d3f06a455e3ad98207540ce43013203ea0501c38ef7250f5457ebc244da66252a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8e105a5b0bec30933e1efeef5ca35b39c1f1133f31a7d7be47b9fac9bae8119581b5337d20476bf96;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h83d933bbde9b501b83975f85a5e15f7ac218d8b363f7cab2b1945c5f6340a9d4d0d6b7d5683ba310;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h51691b4ab867b4bd76d895fe19eb51f988e60b0613893f1ddcc59ce3982198bc59cbbb8d6b9c2db9e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1f5a0e2c49421be198fe881a35b90b5138e31b718b3756f314af382c6f4e849dc7e8b47df951eb0ea;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h564f6bbf294d850a1260fb2062877d8c8a43641596314dcccd983a823c634805d1ce28fb5e19c3128;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb514395f7ac02f004e5d9a7832371a4e4e770a0d4f4cce42bc4c587e04dcb961ceb4b11d841c265b4;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4f508591f2ecb9bda54981a97fc1fd250ab1ef070ffa1e8dda8568018dba535e9d6e97cc24a1a3a66;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1a1a4871b265ed08a7ecc9938defc745b8a803c2d0eda0d3f3621465afdedfb9e6b143bad52144085;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h801c9f1cd225468274657f98ef67fef4212e4e7c433a10896c6a724aea193ca9a8b174f939b79f18a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5e64dd312ea0dedefc7a2051798ab36f62ecdb4fcb378e2af726da951b8722900dcf34dcb65c911d2;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h80fa4228315bffe62ce1003a5b0d4b80cc270f254c117a451ac857f8fe3e0c56f7d29314e3c1ffa24;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf9ce63e38e2dbc454fd146ed59dedc275fbe1fe92a75e6bdfe93c736c5ab9459432362d502e7a5165;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h801218af685dfa96d898bcc4626c50a0a38ef580247e8369b20270b75c97caac4902ff0f11474bad3;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc45ceec647664ba264cb44aae4fab7379a44d47a8f51feacb600e2094e4c9cc6aafd141e0af89b6f6;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h41b5a112940cc512238f666ef4f35716d2dc15e48f2cd22034ec7d866e130dd388dea5bb36e94ed12;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h550321f6d058af598d4ef51868bb514a2b8ae1d3aedb03e05f686dac0083822c2c1325c86627200d8;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9bc3bd55786497d4174e7ca4d5183d15da8f4c66601a1ee0c8600f795370aae81ceae64e8cb381d6d;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6f34683142588cbd3da28c8fcd56343e11cf1dab97af669db5aef94160ef63cdef0532a79e1f7dd27;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5771da6cc0c6ad7e9f1efe9deb67483a3d737671ae848026d7bded66b2b9ceeb99d4c7951dbf1b36b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb003529d1aa554c7b271f7d70762e6f3cbb3df428dd4dea86f276291ebdbf82359bf3dd9c6e5ba783;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3c2d45edc62f9573e4155ca7c761a2556824c277ee2a6583d996ce4c98531ae103fdbea8b6cb1ef94;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd88fe541f9d29a7b4a8f27e7effb81408b665caee918100893862d671239d9766bd3c2ea193323f7a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc3b4e362b6fcd095b796e137718d28a120261e93dd240d167a7a41598d65e0c558363b99127c195b9;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb0f2185244dc80c23f082131421dee8ae23520b5ccba0335de9bf6ce4ef37084db52d4286d86a8e74;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he0c1735de256e280fd69cbeeadc1d8b57fb80285e71fe2558d37cdc5bcaf7f5894773659699065a4c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7a16fa5ab605f45a48c1e671a465883482133fcdedbea9f3c3136310c7b7396dcb4e96b92acb5655f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4fd366f173865b121fc9441ac89791be8761df3ff3f7e44acd476898a50d94ffaa516895b7bf8ac86;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h57b5ab13a5f988a08431fe1d365385cd1bead5516977cb856cc1ea9bcff2e4017dda6b147aed58726;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h72227b5da92c58eb646899d75219b2d6dc6d81f211f2900a7a75cc5e2b1df0c75387f9b6d1300ab26;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6126ff215ab9395dff60d24896080432197500253c0ecf01727ca5d665fa075aa2ef02e1c18ba0466;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h70fbf252e0e0939e834754ac2974a980ac24a1373f281858f0de254baa6aba82a91df4c1558f42a3e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9eb24c020e72bc17d2072f1dc095464f719c1c13e4463548b24f5f6db65fcde47ae8b1d4397a3e836;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h837c40873a210b94ea7d3f820ce7b1604925c43f98a0ea08bc93c991026429d838489c198b36a14bc;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h69af0e0c9f130bb4981dafd083094fd61a91f5adc409c71a6adabacf8a41ae5dc90735a79b4475745;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he10b562471465b555b3c3eb8026e66ea2b281aa5faf0dafda48d210f68a6058b34c02bcd9f790e300;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7eb604542496af4875a96df9ead27d4ef7c7cd0a5d3deb5c09145d0c17e0d737bd7fa43bd47e113ce;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h16bbe84086430a4a42fc4f073a4c5f36d821a2ca418082a13d3f6b727207196e654a0402d755c8022;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he07fa7d38081126c978b148e801c3323b05bc6e6d49af054c38ebefa871277944740ab26e68e076b7;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha9a20ba0970a4e94d162c4d9238fafb41a9d44e3baaa5ed4e056e10b858e55ca1d5eb9a1da2e052a4;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hed276a5361f19c73600928b983fc9adca0b5df36f079c5f3431765bbdbd0a0bce31ab7f6ffacff84a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfabb296515fb7704c1fa46b6f5f98f883d9112f0d14ee8905c1f886df13f6ab658e24c7544933fdd3;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5d2ae96b9e7f352f569795d7d1e3b0ba3304e065f7592c29cffd48209e0ffa803b0fd6db8acee045b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha931b3fd02bfa2ccc682d8d0a60ba56e757786316cbbe3bfdc4604364f32d795e632ca8a1d94d77d;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h44cf41bfe8c39da3f6d447866d94916054c07adfb356fd8c669ee388784da34edafac3f45781fb2c4;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h993f685ef9f80e48c708369f619d5fdc54fefbef6f9f4ac734312e823ea743896c01a3f4e91f7396f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h756050a35c653c30675049e9ccaf777ed6db0e53d1c3d80d0bef63aac4662a5dc5169b021fc54933d;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hab7046e8bdf0a2002ac7c5185435ca7125d7ffbfcf4392b695b0c0da9fc3bde0254bd178fbba1dc90;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h612c4bc69a10edeb365c9cdd4990831c5f94a1df0c0462e495e359ad4269889656074a89402ecd81c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hce3071a2b484232822f236452562839dcb3f8c54b3da86f2caf4968aac715cbc55ae857115816d200;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he246690bbe35116fc5a803488136e2a83df0d9138f0d00a70a3ae6e326970007f162ce5764dc6c455;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc5abe603f2b45c6654951fd37fddf103318231c620ad55fa9e8ed5f1531304a10fc32bba57c7c6ba5;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hae529c3b61fd724ca96eb78d2586178bc27bdf363b7be802ac911b97cea8f54a13ec4f319c64f4aab;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6aa514c8512d1983cd83e09a4fc85c9d0a19a00020bb55d4318f6ed5f3ba2e6b54f91127dddc24f70;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7be7ca03c5e94c44afc9901d5b7eff4292b04d9cd5f66926173b1a26d33e99f707bdb0c3f64576501;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h57f2983954ccb98eaae240405f8d365194e9071aa9320b1dc1cb053d6b5e2c69bd989c859020ff696;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4d7c472321b5e4aef2b2439a887732b9917c83826e660d3534d7646ce14b01f20667fe4266ab10a7a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1f25bdce90bd5a96ee3c01c13173c180361a6c1aeb0deb65fcff15abb357446a1f11ee73eeb71c0e4;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6b19d65a4d581349e14204614ec7ee3c68f445478fabebefb7a56ad29a8b66ecb24177fd5b6cd1279;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc2ca61be329178ccc7296f7c02761f6f9b91bdd719fd714e7f5509e67d89e9a33c679ba531e6322bf;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h37cfba0132d0fc1a4489491ef4f29742e9b58bdc2ca93a50cab1278199f3e47043c5e6ae7bffd43c6;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h699d68e9829cd18e306a26d875642a6f785548ecc7590b0a16b347f370f9f0c06b594361ada668c7e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h269c300f982c0bbf9a0244a74a997020904ee2d19fc55fe452f73f5a1d7c51d551c859de7ad6f53b0;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcc345493e99e41775b8765e9f1cd51e714f3c8997f52ed996948752a91e25dad612b16350ae30ac1a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he863b3acce3cc94cea38bcea114571c42bf6d84e64eabf12063bcec12bfbc3f2baf21d62a9b17974;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hca394fef56d2aac6a81381430ea1de828851f8e1f6c897be88f79933050defe64307d6fbd42221233;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9d16d7dc6554cd6317a63d6ab2f47a6d9a08246a83c9f47fa64faf617d881240abe9f2365fa3b56a7;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf8ad89eace8cc8702269d374edf608ca6f858fb979a2d0d3fe109d0389ecd924065a312a1c73f8a6;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7282b0744e5b666a7cee11485f1eac45d20b6a07433dc75e5b3f649e02c76764df8110a5e4fd0c52d;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h647139ab5b73677f4b3306714316a0a2a27d06a7185d7bc3ab0ffc0d4cc69d6f81bfe04e035c4a551;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h30e140e4fc1b96f61ca055e063c61a332323a20e9b56ad5bc4a61b335e15f03035c8ab1aaef8198ea;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4ba7d6a3ddf76aacc6dc3ff5b97ace50755ba092754ee93b76d925bd9395ffe827912eb349a0ae199;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h78e5c7873d00554448309a22be7b9f768435bb5131867da4a80e4cc8996fbb5748b7fc70e5be3dce9;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h909803a93491dbccb8b9a15bd8539c96a9920ced41ecfb4608a47caf1c013b52a70ab23c85658cb46;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6b8ed6c53c1caf5327deb5f8a334c01de1e4c2bad27dc0443501e9974174be3e00c2c0de5f67af402;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h89a8d47f102b48b200a9b8509f196dba4f98a86ba4efa648a65d82fb61d040af2513f97ebdf6a1f22;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3898c717686b7734aa832cc5704ce257e2bcb9169a48b1cacfd29392908e656b35baceebdbef8ca4e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9e8a8e14cd83c69d3f312513200067bb4988b693294c29c32ecec4b5f3688fc3d6b9643d6312fa2db;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h33b90e4bc8f844d7adeb5964e67f973d78ff15f978c14d266792ef5f2cfda143a56db437eb90630e9;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9e6782a833a191552e8b40f2cb152804c31f83a2a18a2ce20d39dbcec0d8f4f10f3852635fc72b97f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he8cc03dd36cb1d221fccd73c5e80bd652a611a727a044ab13549eab341fc001be6ff64748f49b5024;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd1d8dd6c71b9b27bbfa90c8b50d6789f1593562122f38c6e145d754d359946b7e1a10664680e6e3d1;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h378058c94a1e6934b509baee7b137087c9178e8f225e852322e6b0b2f1aef2f05a88a579cf8de2433;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7af1e7d3fa1d8b1539c90de6fec7d6987501f19dadc0edf72e86900db1f381ace702eb721675c81d;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h933936b850ede5a552251db3337a19869deb395b526bf3a11d70ba166cf72be4ecda7a6ee64b52c4a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5ba60e59bfc86e212164fc70c1db50f8fbc5aeebefbccaccd82b2ce3eb7b80ace0f9ed489c41aff68;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h52dcb9142b69c8fd03e7bd0424878af8e0dabd97ed415be37d765f1de5ffba8654cded2fe5194516a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4e1db3d0b7ddded758c293553ddf14e4d01af7216af95513411378698ed6f673aaec616f7507174b8;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h791a585e65becd49588eec7c04975125d4f4f86a9715070dfc93501aa7070dd5131d257787e7121d0;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h70875449746187b2d1182c6b02700a0933f3cd9137f90b94c846408868e59bea9c6db88d7f004c665;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5b8b1ab1e5788e683cf75d37bd9beaec2a910746f69c3acecb126069f6e8a97c99c5402cda9fe309c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha46bd19f95b86a83c73b93ce2594e2e1268d46d97ed820c9dd74897d2455ee8c4c357701c9fe21b9e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hebabca60012e278b2065038b8d700f860d5c0b08ce7c6348bc0f4699b31cfcf998db17f617c8a57f8;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha31c9d0b25fc4aa6c23e58471adb7d844041833f3e5a7cdfe85bf83d981f4b2069c03813c20939479;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2020d52585aaf0043d8047fabe7e0edd2ce791cca47ed308ca4381fa6c2e4f78d126e80f1d9778627;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha368a0324fd0f34bee4baa58dd3c52deadda91f626e53f5cb9297203f9eeff5773ddaa43d6cee9634;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5e60e1acd9a2ea8bf674a7fddad1f740e9bab55f26d422715dfc7436219a3a1cc1d695ad45c7cfd74;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7693b800bc823e959b07d88a937c0b28bd0024946bd52fcac3dd92b00f2902603990088b9d254d218;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hca8371a962651a49dc88ae110beec6db1fd5124882e1d45d72dddefba98e0e9d98849053e8fb1833e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcd505dd5f50bb6430bfadf69e3b8f1806e0b14ba86f70e95ca34121de54ac6ec65a47268177a3ee0d;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4d6d8687cfda648a52da232b9d6a8d3de6fe3db08b59c4700192ddb322fa8f76c198ddfe08363dd7c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfb60888d016995701e7eb8f26564894aa84c4e38ef4462e597e0998c49649897fcb55310e2c4b1df;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h95cbd168235b6987ade71c10ada703355462d996fd4b5c8407d9dee92e810b54f7bdde58800831c97;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h20a8331fbf1a813214a38747e9bd90199bfd2e004edbde366c5e6d7090ebe374dd0a4aa4c422bfe61;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he240a79915b5013c4c739fc11c3e95c7903e3ba1b0b2ceff278a00aba92a475af208c7397e3a6038e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hce8dfd72fb918e9f3f353a6399df956461845999a23b37ec3117ab7583c0ebf6f525ab7cc768281a3;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc6e5497788b5d99c49a3fe3508dedc1ea71fb5f5b78ea7439b609cc749a8b31979d97d0952e04a820;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'heca2cf4123156054213be5a036cb12cfc1d39f7f97fc02a9b179cce99b40d37371aec263c5b85c077;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7d28e14a40db1ed4d4c26c3b1f487c6b23c550c5e949f5940cba2ebcf31fabcd3ce39ef7ffaaf3b4b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h70781c15cf4a4ef447055bfb48532754ad9553d91496367527cb54b262bb9991c6c9fb74686127102;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1aec9b7dd55c573334ac691320425283b7e2bf673cf7d75af39973f74ea8eea704e9a503de56e0016;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4206b162be039d4db589bcc4dfca215f5c79e32a29be256055cbeaf77d498d3fd22a1505e98d3681a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h58f858c0eb6c45639a43751e8f96a8e939948b596ff303bd18d8272ead7473eb911dd48976b98f985;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hedb87c2f0d68ae31be319ec7dcbc5c7c8dc8d13117049338d1151d12ae64e3775427e7ba594e920a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7f081b5dd583caebba25a0215293001ec6c7b9031a0e500f89697fd603bd01dab41fdbdb940b2643e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hed3f388eb2f9512adb99601533a7cb5a06e283aa7100799d0edeb6a55814971e8d509f10aa478beb3;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8d4ec7011048d75fb897468fe1b0eaaf4b4e389e1e7c8b232e8404103f9df708e2facf43bfecba25d;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h161d955884340d27f16faabf77cf64abfa86ef5aac8832c2728ee90ffd3bc88b39fdb5b0490f21e69;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc0e27136fee4303d321584cc1011b1da40f450d7f4c19d32a1a5843d607adcdc0c676d3c5519223f2;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc3db960fd42d1d4d3f7df49289ed77130e2ee115f9009850c252e2d490a48e19f3a5996e35141e21d;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hac40553c91e3b2e60b6fa7571426d8c24dce44fc1ecd3d1b9d6e856e66676cbad894ad7d7facbd4de;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd6ba5e75f707c704ee2f35b04f3ff79205125938d0db0a3f17040eac29d01814ca3d26feb87ecb473;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h911696c7b03d72368c6da70c4f25e8b37d634c0b1ac0cab38c60ad7dfe9a342bd4cbc01cfc4583ef3;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7436e2e667429b5d0a7c895d2de51e3e01806ff2123332b875f13ad6a9f632430641be0324058b678;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3b3bdc53e4d9fc6ac9f07aee7bd89ef4d2cd533c75f8ef6c1c79b78559a81317959df547f54bb7275;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc5b2c68dc2b2e1257e93e8b9851b8dd4d4721891b6ddc86b5c35df434bb24bf979cc30667ae50341f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h48aace34c66df62a1bd143439ebe4e2c677ffb43b8043e7818c3b3ff1f5b443634fc4ebb887c73321;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h99c209d6dd77534d38f9777274fa7b81d3d1033aee5f3875b57780c30185c5d3ff10eaa223106feef;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h36b6385fb09b563c8f16f06fb64f809675204e7444d57702eb5ece2048b5c70029cd6c630560d05aa;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1fa0cdbd66b54ba6693fa98402101723e903425f40f9a90dd71cc9b13fd1105083a803d91c1bcf0fb;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbc73e6db0bc102bf5c862a31ad117d2895a72bdc25f8ac40e05878765bcea3468e7e9bc70f3a25193;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1e2ff80fe37655648f44d9c55eb27db5669c01dbd9fe65b3ceda8fb26ca4449dbc809839d5e1efe28;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he37a66b00a37f8e52ea56053c4bbe85dd598be7a4dc708d1cbcb6c4f8678191c488552ffbed1ef7ff;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h99deff5542140ddfd543cce457a290c7c5bea7a4f4b8affa6b322d5eae54d4d77f06a101c5220ae30;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3eddd50524c5f59f31576ad68b26d9c891075f8cad9f37707bff49b1df549812d2c2de78ab95f68cd;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1a38af88a3e9dfe9456e364f2be66d89c6b44cf89a8ac6c21ee53d4d4c30f466d2ce6f67a613ee3b1;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h86b26d99c858e1318300fb31c47525ba102f5cc2611b7326b581c73e6c8c7dac7ec492cc4db53ec88;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h67aced6f0d5acd2b3ee4608cdaaf1108d35fb3c8914c085c7cf0c7cb5939d2625a9feb1ce0a3506e0;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha8e652e1f06e34cb08f42916c05126886c10caec7677c5dd35af4c0b42f4ca72e1909e7c5e76fa11b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc03945f874fe215ea13baa91ce0c4ba1471580bc5ae42b61a1dccd9c0e24f303ed58d08ddc207a6b8;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hdd96fadc8f2d70a83398790a3f59532ef988d6426ad5892d18a072437106080a8e1a7cd1100da3c1;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4b156bb65b9d6bddf870635f569ecb923e703fc471017c943fe80d2d1e32b6efd917b44eb74fd9c67;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4ee0661fd0c7dde5ebacb32ac23a86cc80537a764c4f6ed4641406a3f6cfe22f217ea28511a9a5ec0;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h182794765e150d8d34a11c7507a24e3f7025efdd537b828623a4ffef4f5416cadea3a1adcfe6483ee;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h43139574e3d89433d5c6466e9155886c219cbc822f8f153ce02ea74097d462ba91b01a4a6bf35a37f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hed56f35c16992e213d90d8c97a96caf71a9e2e0a09370c3e7f25febe04ef00b629e8cf46aa0a2dbc6;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc115da036e61309e327acdae93d798b9605ede13beb2e677ae8a178ad11a6d2325b0faee4c9f6df41;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcb957cf0216d0b134e3df823253be194b2808709ea848aa901d68e9e5dfd781da5936b341d3767b42;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8653c406a4442bd2fe5046e49866cb775ae7a1754d84a3c46c6f57c8ee2937021b70fe14be2adc02d;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5f0b134f309677413f8c6247a34ac08067e12220d1864bdba9fc754f9bb352b84f1e7fca5d7f63c3;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h12933ec2a97d8ab88892b4f24e9b4c398d0abdfd3242c819be41d360ddd1414f6d2d3642f8db021f3;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4419167e52b2af7afdd76da622c7fd7f66debd86702307e51008029b3c99552a260c808803ee536f9;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h67f0f1a32e2300e2ed1e088934f368cd4766e337a3396fa9f4f9b3a4c64628612b3409730eace6f50;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h383aca4ef025a26acf93206ddf44881d0fadcb99e0209200380c5ae9e80b0ede9f3f2f1aa4eb6d2d2;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7841d45f7b7b65f5b4dcd916c64200a0eb2779336d80a729f11d0a7dc0042de9d19f7075aadcb3356;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7008ba13c6ad8e9d5be2e6e562b2e6b66f3781b94b5994d3349b115737d663e73fb35fbdcab21286f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha80918b3f21b4b3e09926775c02a1b7221b9e928b11fc36a3058b9fd28b7b17dc32bfd5d5f454bcf0;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he895edb45f695e524b421c0edceec66f10deb7ff1831b95a16697fdbc269555cefb3e398a135f1389;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he800a0a9b907d82e90686ac4b931896613bc16a8ead0ec81eb5301d3b7ee2d47ef635febf38ebb558;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbf99a4a79cf940857906a50f28e2fdd1a2904a813007241a5f819f4447cfdcd99eb09d803674d8529;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h802237557f5a9ece048a22b08807b5d40471ed0c9bd50c4eebad6df9f52ddf162636d30a4b54d033e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h23ee19a71b5fa142d5645e1ac39c46f23317a799bfa8d491167de98703fa48a329167e15db590f89b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7d4e3a08bfb228eec28793b136146198f37e1340615c9f4271a4fdfb1bab26ac97d7cf60e7515f317;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfc378936fdb20dac0dba308c3cb10102b2c59a6059c82a85a27eb9aa31de737642af7544c717854c9;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc47bfcb410e75808cb595daa8ee2f0335ff97c417e97342a2e6cc6a6c3fa6d1ea3326e79bc74d65c0;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd7d21179b9dbfca6e58d999b631bb7684f8cb03183ae7a17db8c4ec47f992c46cd9bba8795907bd19;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfee3a6d80f9bb81752db9108f5971829c57d1c526acb251656afb863cd06e15d61dec210c64a647cd;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h22fa8a4aedbf698f984224066cf7bb5f5f77af94030fbcf687d12ebe415a3a91c9d78c63b804464e9;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd178faa661d558f6ace5459e59502f44ab695e2e63b73e1d64de36b621318fa69c1c219a3011f5e12;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he08be75235555c3d7efdc8c072e58f6d796da18f1a7b681103a2d3297ff5ea77d131c5852c3693b47;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfc92e15671eef1016ea275598a7c74a8ec8a0d9c7794d9e87d3494fea07c937a8e34aac301c84f143;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h222e279910b2afede7757d688bc9cd58d0c2a8ace19bbad0222af44dde650c40580555ed951a7192c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h189f1ae0fc451c98ab4898cf1abef321506004ccd3fb317de7a3b7fb60c62feb410f387861fdc782;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hed46fe8e230110b9a31338765ef93a0497530a9a486fae1553888e8579ac38bdd4473631d658c7cfc;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1afedcb1937bf9e6a70eccc3874ef0feed5f7da0baf33a6d48c305200dfbf0417cb3a1bd943fbaea;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2eef04f22ba9928bc272da2300f23324b97bf20ca1db2bd0fa9e429d98c33ab4cebe58ab32b784a54;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h646c2ca37a297da55c4e58eb2ec42c6e1f094c115fb27101d0413644f621ac00635472b47ce52291d;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7da4d7ae8d73b5d167f2daef18fa510c44644221c60fb763f46c2d5b28f3733280a14eb3f125caf4b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6883ce5d3b788893079f9dce4b7854230bc99ce94636e403b21c0a0a96b100683e6f7c9b0e1855aef;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h585a2b1c1fee0ff384471ca5b16a4070fe13e5ea064930f91f6b3b8a9e244e6c9f8febbb98713ac8b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h99a257a1ddf0c82368d482565b43ab454763f16946d839bdd42fa5183cc07ac257ad82754dae1c7e4;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h37874acb646e2282c5f7c6ff353c1952c09b466cf66b627b99333b193068027038e592dfbb57064d9;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3a2e644feca1ded9f8a1bc2283ccc622f3b77776dfba18c937f38f90d74ff0827480289f674c527ac;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h97a6f0d6952acfbc41be49b4492c9dbc2b65b342a3b7ae7bb81a28534bc5ee429131acad81e4716dd;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd4ebce83d478a56d85a127c77043395b01b84142c0c9cf1b3431435c9bf3c5a47b24e2dbf8f679288;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h41f99b769f036bb5ae46658d21d6c5155e1a70f069865988a2824bf2b640a6f7ef03ac211b26f1393;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hec51008dda974324e7e23c6dd681a4b44071e2710d993553242267f139232f4617b377d8454294f77;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9110b577ee82212f608009544f6d65c4f7a3186cf6f0a0bfff19390f51ada2e336f3a91acb142f85b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h390602aa0add6409359b9df175f07ba81fd6afd57d3c679ec21813a776284d4d2d104a5ec8865a4b5;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h57ea159d4240b73cf2f9089a94f8b7481eda2010926587ef0a6c8819615d328042d25fcdd5099680a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3f6c46c009f0fc0129fe9923151271221a87cce0d17904ece3c3ae28283a782f1b0c5e0508e1c8282;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hab507ea182fb5db404400d23f910ca1432ec0eb7deb4db86f5434cc9ee6218e00ee1af369e4dea9f0;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1c6fd3e732e4c05f66a0a3d5b34f7fc042ce58468c2c9d83f2a73a6e8c15f1a6d456cc5159c0f6828;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h57ddedb638368dfb58ef45262892f28b3c6ac47890f1db8f1b6798d3ac846f5ee6c7b24dfbd37b626;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3104cae81143b93112681b787dc54aa61e810d2b2cb5763d940593bc4d2eecd0e4d3de5c35927b282;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8eafe0c0d2c77ead02e14039aacbbdf1e27818a58260174b376880f8707032f10faf2d3be20405cb6;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hda2cd059edd53177c5368ec340307549920997db4d7c4feb4b56ada1b603d351e2eea18bfff03b6c0;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8d1eabf3bdd45e97dda21d8edd18e93d4c7a6361fb7dce7c3f6bc10e412b51767940f33d550d53ca3;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6fb30cacb2bb496e4ca83bbba43a204197dcf9f424f9f702694981f1454490d54bf9cc2c7df965ab7;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hdcda7014501ad47f392a23a9887c0f9c0346ab43c28fb49b1edcff171e04ba4d4615a44c16a78fe1f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h53052a7a91ff9597452dd075ecb578d4e16e9252874e4a0ec0c61506aa0307b3ec41efa35924b68d0;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha13a8c9f08809ae430ab184c5dbae717173d270a9274cb7a1c3d8b20c8c4626fdf74eb3a1bddb8dcd;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h45d95244f1881d21c1cb2538ee2edfebd7cf20e83cf8d573ad3b7c2293cc10866c257c0257c5097e9;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h858fa9e5553c00559a2e2fdf1c69b2b066a330489f43c5ab2081b23d0c07313eb1be86f27d2f03d9f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h586ca9fc061121e2e33e970934fd809da11ac4bb3c13c7e6a59ce7880924b28319c8b82c42625671e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3840b509267060b78445411a9415cdee92013ba6a582e5b454ab92fa7ae4e6a4d12a44889a3429aa0;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h975b54a2ade9bff14b266dfdff2f97efd93fb050d8b22eb0456e752d5ef3d5dcd3d0c1527bd0f8a4b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h799c4a549a93fe39b374904f8ec0d8d941c8ebf240e027e39553cb407d5da2bdd3d9a2d1128f48e3b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcefa826a783958144ffa8ae459096c4a8e8b7b97ad2cb43a06258b7556be3bfed5941139f1328534b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfe3205c5429d38f39209030231923777233a832e833e9dcb7a435d19574d1a19533b92e87cfab399b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h652545c629fc8dcbb2106dc0d45bc2e82ed300a80f478b54e3872fcb39fdf1145258812a0c96727a5;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hdb65d0ecd81577a08de0402b82e70b619c76b404ffa11a7ee1246d6806ba865995ff8dee791dd8863;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7667721e0d28a34ed05d9e61881e0063f4d7c690666a68152c424e9d3ce201167b352e8cd4c0a9649;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h80e82adddbacc65910b5396b8737793570d4adada236239de70cf3040318904f7c9a324d3365b0a50;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha0f4bfd927aef5ba4c3c6c88a486e20bb0f634c96737735ecb3cc240d9aaa4b36f923b32a5a8e56a1;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h32e6535fccd17949837d42e7de2440725b2726caefcf4d70f55c17edfbf852acf4b0b724fb076209a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf5ddc0849396699d278ab8ed41cfdb0b92333d913bfb4802fe5ea12fc9121adf22b13d7fdc237513f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7d6dc9f3ca3ea81485bac47cf92f8ddf4bd45d6805fa86047a7120798a06684b95a2524f7bb139954;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hee4b0c526a480796141a767ca0412d586d5b9afe7f34c20a43662ad63689d38f40ab47ce9c71a770c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc833f5be21938c3b15be5b0f5b648b5211e422dcac6f4e977cdc7993a7bc7b2d1fba203acbc8c389b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h68157d7b69b85e9c19eaa466a1efaf880cd0be51973e2cc7e267869d508f343c62dd7c0dffd527cf2;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb9563c76600a2e82c0dfb3b4aba682def704de2649394dac7f66af2d17bfa07929af33415ecc459d8;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbe2dc7eb1d42d2a317009a3e5140a26c299048708ca6d3a0fe87e1a6b918f5833705ffdea0ed68e2c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h92ee414e753d0a475358da07ac5cfa54e3e42f0953135d348bc9121696c7e94ab52343df456ff356d;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfa4423a4002abae8e19cf96ca0594f56fff832e8a9af731610c0b4cb9beca7f263636238da9941f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9f630148e60661336e8fc523a1a183ef58b299d7d2c634c98c4a79f6b9b456e7ac42e87b27948135e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2d24897828c41d5a2578cd3185cc5f40e0d98c8fe64d1f6734e6a90097c12fa944a8025a4ff909fb1;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h56634e4fd6fc0bae24f6705339236b820738e93cb67039cce0ce34597982bf19406edc57762a78225;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8fc22573bd5a290e7f2c4024414e56800dec026ac6404cc9e3977c047ae315d331d06f8c6321e8c21;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hff99e17cfe97463ceb0f27750637bd8e6d78035225918aeadd9eb9e9edf6b5a6fd1da5b8450de93fc;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h97e687a3391e88ce20e19636b184d993806bb1bbcab90852faad059410574f270cc06ea70cf76dbc8;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb1db0a36d5362acef051698fa02a026dfc7dd170184f809006e8cadfb126acc6e6e085d8f101072ae;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha08fddbccc600ddc9649cf1b403bad0c2c90efde7bab5053509b393a4d8211e7066343e6328b2d355;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7747635f019bb51bb6bfaa10b031466f7e528f5090bbb3ba479ca7c03d31dbdc9429196caa54806e9;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1d9427c8ef323ccb6f27d2f63b72094ac79d68e22882d134e7e9c9acf51cb43caa3fbb22c0b14611;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hacb70015c28d3410d93db3ddb2db57f4ec7fa1f626ef82f4182284b04fc4360e9a28c974ddba85d61;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hed59bf1f3482354542f50433221a12b9255569848fdba3b1b9060d4026d84670b1a1602ee6091f917;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hade48499ac70b8809817c47d545973faa1282546b781fcc47cbf26ec2a4f8845f6e163cf57d99b9fc;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1a81f13f1a6e7c1d6650a6cea7d1174e7a61135808da9624b6bc65b7a044c4ec941efdd42f6066dea;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2486a9c225ea9b73f5e9f5ee0789c832fe687c4c50402092166d58884585a355db38ef8108ff369e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9182b8e0b3dee3be5df1bab52799a97eaca173573adec6f811a2c11128361fd3ef511e2fd4aa09cca;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4183e500989b97ddd6fb9918d3fd79abf3f7eac33a12bcd7431fea21a60837122b6a18b84933b5492;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h77a285ba752556fedeb83b2a0815498af8891c26e027f2bafc45752313dc81c17d7829f3de1298fef;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h60c9f414b000b20a95c6166a6bb11396981ef4c0c331c1d78182cb15d56121dccb521fc8bd18f5085;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hce824909f8f30b716a145e0967fba813c9c1dbfc3330700ad347a9d0b1f376138098ec6e3e3b16ee9;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h236407a3d5a2cc163f06575702affe26192ac3539a5369c88aa4cce5e2cb901dce10f5446a48c755;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hdcea2a123ce4fc9a822fef832728dcb71bb252f2cc8a7352fb7e1b84faf27a177ffa038ed76f22d0c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h832f1cd56f435ba44376d022247cc1df314ffaa484dce94dd6bf30222d6336d2cc751cf2ef9b5f83;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb5d65664535a0720435d1e3bd89d15f12327cb9ad71d5dd7fc0a8507e699d76e9d3c59120a6e51ee0;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8e90b8a03a01e51c9ae34b3e7d21201c4a28479d09f270ad6279a7601985b2809767bf56913dfb532;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4eb901d124b6a77a3103af61cf24adb3a86388fb31d59bb166d08569a6a440946dbfd8a57b22d8971;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'haf569c733b8985888423a667a85b6aee81496a4e9f87e77f8da69ef8379fd3f9ca95b7c177abd8f92;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'had62919d160300d594e34781446793ef3205acb32fd74a6e81c83b695774b2a86c7a31acd5185c61e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb0a783f6dd0f923d84579ab1d82ec290745dd69088dc733d16aca65199c89e8e9d975d4892f3e142d;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hefc3862b4685646ee6420948976f8c488579f4880f8236b920e0e78b1ddb53be0fae77ca061679732;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'heb96251b5b3bfcb858647441be85670076d7d910d195fef6bddb3c5db6f6ec39c1fdf9ed5def81fb7;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h987f80ca254d02a23f810de62d5bd0334ff9f09cb22f4f46d7f633c144580849341aa3e491fdde28f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9e56987f819ac6cf130199930b53925e67fb48c2e913ec13e0143699965b7a3b1cf4399e71fc91de4;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h44e30836fcfeebe9becd0662baa5144b6a369dc8aa9f1f3202bc2983cae193224cdf03ca289718b50;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3f243ac6b7ad6c5b82a35684183faa4b5c5abb5626e243ed8082a29c734546a47d10c346b0dd2a1fc;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h143c6b8bbd44b50a9129889ac388aa7393ab8d10227f46a14743897a03627781b2b9dd422f2fb21bf;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5ed09b79862bd2ed342bfe954d667a44d31a5513191d2d78bbbab870c88b3ad5a2b42334d3dd095fa;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h63bdf0b1025909b6cae55031c1500ac9734b81719edf11cc80910965b6a8bdfd00b82387a30b3af85;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc6ab944cda211ee3307acec5e9f78875f507c173a4cbfa60cfe6de0f4a26ba60d8d50047343a1b7ba;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4723318e46e1fbfa3bc3c60b44a7b4cc842737571d39d62b4ed74cf387b77b86efcc65d76c4a4f738;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h21c78b0573d1b76094f6e08c6657d4d4a05e0511149437001511ec950cdff8ab38209764562e49fe3;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2ac7d7087abf153f759dc3583b1f03d55f5b9b470118e11204210021cd10408a1bc46f1b8ba444216;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h84ec0a87a214e74ce005777b608adcd12c59f45c41be4b456d0ca8267e40f72e70108df20656bdefb;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'had50f2c6cff93f12c3034b782a5c347ca519306a59b189e7a91f10263b23e67b09d899077ad8f8012;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h81dd9c7bcf4e8841fcff7daccaf033c409b1885f27af32936f61bac2a9079c2234c220cead56fe8dd;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9f4db5f52c95871845339e39026c540ad8ab6b769dac641d7d487e4945fc0c729ebf3253fb376ddcb;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3cb899ae7be0a776e3e8c2d81d16b6f29d3756e6a2b6cc479f5f0141dceab99f33367a736f3d9347e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1d5f41b9336e6f58d563ce670343677da6f32e8bb72fa8d7389f4a6bc8ed1a1e0bd16236c004a9155;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3fc612f27aa1e95f7426715e769b9ece1cae634212e563a66af6519effa43184c21fb818b80dd6bfe;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha2c2db810179100e5db858178df3b864dd90f23bf6e30f5035ce58c77af2c548171e812d504825ee;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha0952429afeb58b11cc5c1ce083764797a419ba972ac24e862d8ed026f74475783039951bf6ab71d1;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'haed5f0fa89236c214e06fc7012b449c4b43e73dd9b5cc0c8460afd78674b353c8ee7de2f84bfc4007;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h87a725535704d9209a97924e7793f227062ad3a53bfc49526abf46e9a5e22c8110b68a7b133f28b8a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h601b17741f96cca1f002ad2baef7507ea130e0dd152211ddeab134278ed048630d1ded2199fdce278;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h241ab262dd466fd4adc70a1747e9fd3399505770df80ae73d4145e591f51a90eaaf69459d3d33ab7d;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h30541b3e55444ceb81e1381e37cbe68b3d6ddcf10babbc0f5155548138b4713e8e1b4fa4237d064cc;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h64fc5ebe74c903d87060763351033bd4fd489157fcb5d8376da60f96eba1bdb0d9788e4901995d153;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h51bf78ed74c1fc1149c1ce31180f57888493cdf5cba9221ecb5532e9acea81dbde4e10476857dce99;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h27b314d922e130b7f1fb1d71d1083c8095653912425df95cfb43598079bccd5859181e41184fff808;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h208da55892be3cd12643fe6991f6972f1bea92cca13151f7b662d5fcf956338b6d55f34d09129ff5d;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h41dcb6a8b63e6b586fc83c912dca5aaa8b1709deca578eb580cd242ef8d87493f4e3afe292e213bf6;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h66dbe1eb5d1a3b7fc28c1dc9cca4a1c4bb20066dd5012439142dd4b21e73a771403d8e00a11550d23;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb135b510857586c42d8fcbe6e64b43dc7fc7b0c9819dfe9f437bdfa4c550ad9d1972fbff1bdf209c4;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4dc902424b3541392e534ba64bb8390d007b1abb6a1262f0ef5ec312ae6bed4094a99e4fb1ee4e71d;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h482cc19291dc9b05f0f1355b7b432b5ba5d58de23b172b5740c613469ab880b86ccce291d10cc6321;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hea849151b62f5a8fc7ef3d6b5e39211127bddf57a6f3f3ce1d49788e4d4fdcb41c4f4118cef038210;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he373cbf13f1fec064d9440b32ed8479fc2ede7cdcbec569d3308d722bdba4b75eb4f6d152acabbcec;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7294f1167339cd45dd060cc7cca216c9a112fc0e4fb4ed0b34cef2d196ba05388cb7cdebd92efdf1b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha9b8331deeaf53bd9dec87ea4d0f320f95dd464187e8ea48c070f1a54b80bb1f1f3dec3bb818991ed;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb67573bd49454a331da50af12283b9b5390da6dc2037026036b9e95daf73707e83b30d813f64f4064;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hea02bb88e5c33808131be5f1391e26b7d109f8c8990a55e32e54d062f6835c91807112954f4eb8e62;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h17aa870dc0e670a20bbcfdd94767dfde2e2c4eabbaaf45a7c04bd13ec9aa612377e8f4e2fdb6b4131;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc55d3d9df4e147521fa59640c39eeb37ff620c7d3e02c22a6a26450abf52c58a7adcbf3b05ea0515;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha4f11fcd6ccdcc5c0278daed40fb8f86af667dbdb62f2328d373a9776c0678a197c7415dc5e458a4e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9c6793e5ba04652efb2095651081872e9fd326fda214c043003ad32b6df99e51d51d56cac6ffadcc4;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h76026df5fc9713d7de5ffb7797c33eea4f50113ae3d259d1f7aba9d9cf86ea1811fdd61f2801cfdfb;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h44e74e106b7978aefa4081fb3e98c101f66a129daeb917a77939feb5dd69a1e4edb987c25b23482f2;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9d613f88cfcc6357fef0946329f1b4119d7c7760694d0cb3971943b656904be07e2d716ed35ed0e8;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7bc81decd1590920ab3cb69e4c8b4493d2a9a670db495807bb831f6b092d42683b9dd4f5e11baf7cd;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd9f60a846236da2558bfc9f973f82c6eae4b7bd47a650bdb667f52822dc7f781752fc93faf451470f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h634dabecac349cbe247e16b0425616148a213f47591e78c4c8677b8745cef1abc41f942a7f2744ca;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hac99c84da3d7b671e3de5b6ddd823f345aebb5edd7cc6f63aa431b9cc3034fca186a9ae198c9661cb;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h84f8f43b8cf6cae6e7e55bde16f0536df0b5342d191a4b200c94188e81e7cbb9dade1a810902ffc6a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hdb0d30a2fd57c80daacc84fea7857938b82b4d347eaabdce973c5921a56fbab055687ab6f8caa185c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd19eb93c7d5e4eeeda6c4c5aaa7099bee5744d7948dcbcf124fb68000a1b4760c4024c644d14e8904;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4cb75a0567438e49da92c8f9d052c23e63427b82dc751a07d9c537e7ef825bcba983de6a31c7fcb2c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h870927c05605dd9a9be625e558daa0b225b4ff65de9b8d6051f2f881db8cf17ffd30f5e07cb099ea1;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'had90400858fbf25267c1e382c3bbff6bc2d6e6859093bc9819329f00ab19da69fc09d93df74cb0ca6;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc372f5cf2284069c444d6b104dadb0e20a0d27de46e45f56a3581fc3478a9cfee184485eed8feb8f3;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf700bb568b1b38dd62482f0633ca5a1d5454300b152b26a38871757c0cd9496302503c4dd28d963cd;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h789c3e4f9466d8b7b2e4a4780409c0b7d33ca12c9dde9321f47ac4cf44b9075beb135fd31f10d5654;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3a09039d4d0d28d7d6bb0a45b46ff9a7e1cfe6b2e7a33a615a25ed4e8a5ba01c7359978ce8e12b0a7;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'had34fc3e9aef075310937beddcbaf42657160a9e1ec82bb2ae25c22dffc46c95ae83d7bc8ac0a41a7;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1ba259fdeec83f48419914b1f019ffe73b3bafb2662a96e8017c35f0fe39ac1ddf4dd87c1f18cac3b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h926a61eeb7743cdaf41c86b9d6b8291eb98a3401fd27010e5b48314875eac30a87bda26355f699f41;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h66524715981cfd07294a3ff0fbe66400f9294badad764aa8b52c942ff536dc93cc0dee2327e4fecf2;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf80022d94cdcbd61eb2bc9b029fc28c01e54e1a9893ac42231dc85aaec4137b0ebd7a16c9bf1b6d89;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha31a6fcc4f1aaec0d1fd249ff5aa26b2d24db81cacb58fe76b58c7362abbf33c4a8d44c682895b8e7;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'haf32fc8695b312c7ecb62e6bf2402605bddd80db1b36f46c7db5de3799fca4a8dd60a9e512a65987e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3e03006b6b23eeb813d5917139db92834c8d6a534f932a3b56ccf1371756852b88d853c1e2036996c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7c6383d4a2a549c4a5a930347990475b08e4f76fbf59d9e1b87cc864c74fefc8400e1e6e1b4f0e8a6;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd685c355c73d416d55e85b8d34f3f0e38feed95d401e7504099886eb3f8154bd21d2c988afd403c9a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h34722ccdc0845df95e4845056191cf9ed6421495a018c884f89141e0e015d00aaaf2dca92643bd985;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1556aa421294b15e34f7e68bd86980692bbd437661ba85a4b97b97f8d08c9215106a652d8d515e7e6;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb13e2fa4edb0a963220c9375211372606c892397d184e759f3bad891eab1ed099a91c1480f9f4d1fc;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h52258f13e997132cc581237039e3c1abb5c107ca2685f9ae143cb6fb547f122d4b09a9b5484f0aa52;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1023ff892b852666c0e71441038ba5334bb699125d753001ba586326a52c0a3b5b63206f3fd42c7c9;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha6d0f862a9b9462866332fc3b855060563b5ba2f4aa62ddc3311389ab39190976e26eb00c541e25a9;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he2da1227be62bfcc6233c576990ce3ba35d6a4e9390755658a6f5cb3a007a244e8d45ab4233f16f3b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4cdc3437e063e3c670f7a18c71cc9be359cfb4f9a2f1968e8352f7595f296755095d0a145942479fc;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2436fd3b1484060c198171b66a527d690af5f8824545b84b23b773dcdf658d5219ae1dd775b035604;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6e4596e12f1d3057bf4b2d18738d4823b22fb86e0ef6281b2ecbf8f27521a44ef9d0f78cb2767de7c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h13178e3e630272c8c8186d38a98d611c3ab79062e94f566f394aff88c0e50ce484411560e00d0b0a5;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7ccb5a7a04b71a2a99c4d70d080ae3b0202b2ab4295c49231ff4b2b91eeb5ffc0068f9e8acea46b1a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h722397165e0856255d155f206334b49a65bc41a61eba572d0d5c908d8637e7a3494a7630a05c3f014;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h433d052f6478666289939f53f20a24a2e2a9be0fa1313e299c136f8bb246f92c8330a1fac30a3767f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1e74b5455210215e4bb0df1fe80e328603b35eba932acf57bc34ee3f640833502ebaac2de1060d133;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd0cefb5a663f5f2f1b3dc4586bd4280a47581778f8ffc945d6b7945cd1d92e267790051b365c4d8f9;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1583feb47c50f369459d5e7ae7bada027ba93d8a35514f82ac2ea097509e5d121f4f78192ba7c7acf;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h23bea65fe16a9d0a4df32c90587a6846d4b6fdc15a3f348ed6567f2234c56d1a48fcb91138146dcc;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7523801dfb9fe5198f660cd0cf23c7d478044e0d8dc384b7a45e8af44d6bc2ed956a3a2a51c9a002a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfb4ca67df79edf0bc284988eed013f1d5e82b584842e3c7ffcb7a78358a61ab7338a306427abb889b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8ff12e937c7cccf2711e38f82db5e7fe6e5f8b42c7e7e5b0f646a15ea7125446cbe3f4eab06f7c4cf;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2ed110384668bf31c24e0e6dad59f95d6a2f07afb9bc8d17a6690074be94a282b6e38999a0230653;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h77bdc5f44b76395763af1335b925dd09f9512b534981a2fe8b72cce6b7dda5f4fd85e7d58c3ecdf;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h19defe398a8a060aaae391a67621c98ef47413106963e74c7127730e29e3a87a01fad1df3a5800582;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1add59c897473ea455182564ea40f64dc9aaa046050c99bb907caa396667879af35cf4a71d38952a7;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5335657376313185547b085b65d34a5104f0120582936589f944d2575a04e11fc0e5fc2c294617e9;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'had4d1b42476ef2ee8a85845911f78b8f4b39aaa15adfa33da82c37e1f8aa076b424c492f8bdc6e649;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h14ccf46dddef896816eb38b29b41fa7e65c196a87e5833885687c8c2c20dc29a932fb4c56f3a278d2;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1a770d7c1eca04466def0518f5867796df36e527d33f0f20e713ee6046b6c5ed0f58dcbb7f4795af7;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfc2fc2a7a21f79ea4a75330be8dc38267cf8da489fc2a77c383100efd460a602fbfcbc55c3366fc93;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2ca8583f4f3df4ddbd4351ab67f55e7116ec765da521dcda08f47c2470d34406e9e4e668a2fc1f2b9;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7b7cc0c7004847f9b5ed2e80d7ca0f699bf3a3ba6b4bbe037feadc077044044f1149363b2ae529127;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha8eec1bbd34d7036114b58ade5796f9aec16156e9a0b75e21205f212b5be2265603e741bd609e980;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9c95dff0b3b2baaa08b71476818171b0bb86c587abcf7762cabc5ccd5f989f56e5fc169696b3368bc;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h87d4d6c81598054072d1ab651453bac19cf87e21ee5f61958995123b9f68e1e37cd3a23a47380d78;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2f1c7cc042b07de9aa7c24a95eaa92ed7dafe38ebe00cf4eb290d2a238829f3ff65690b58f8c348a0;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9f87cb44ac0eed23c6b7f10680860284db7cac5a896f8dcb0e183691e3d92ac8a511f7ad0bccd8ac4;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h346185dba6822051668f7a19839c82a22e97e345d81f7356394f59a357828d738c057111a1400db3e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6bf3f422c0ad492d2792fb41bbb2b3f6e9ec9056d5a8c22ecfd11e43744774da37e26cace4b6a9b67;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5b7003cdd093cd885826b50bf5a1a63b8054d43eeecd857fbb083f4e4c7db3f73f17e915ec94756d2;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h93d79243796621aee72ae472cf10169fbc1030a1fde19f43e23d0ef9e82e0ad9a56c7c86243a74110;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h90931ac90cf6b5943ef85cc366817255f41e6d1f23c36ce75bb278cc98a0dfd5fcba9e3e4ca2015ec;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h12ce154771bbb7930c21ce6f1e958d1c7410ff8e6024938f7262b5408a4d95d99db9c8a5474f597d6;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h40ac3bbdf25d6d1450c2efe6ce3e1665e2bafb8581806ce358636040c9382d77cf3a8b3e6dd9adb53;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc93fc4dcba1c90d3e128f2ea1d9be480b82fda3b42f10f30a9e24374d94878739ac9b900ee1e8141d;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he82a5b9d4f8e977f430576fde19360f51c52d73c3903999a94080fa3bc634d7901c0fca468d608934;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7cc1a9c8954e9dc1f41f4d45e516ed64df07370c7bb58fb38dcfaecaa9cc39130ee8625b9a129e798;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hda71556a94a43f0813947cfaf98ea9b724dc4fbd76a4020b91196570fbfa776068d23460fc530f6d;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb0fcacd9d3c2cb029f39b3ab6ab995fdd7f5c8ff02878105e573a58c84330117eaf0a8355907f5e0d;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'heee42009188f855ee95fdcfd573c4d06cd7d4faf8834f70a36bbc0614d362abf9fa3b708c4abccb0c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc3b94adf65b049262435b66148154fa74da026bb85ab57560071c90cca5c7d3eceb3b9ca3ebe2a434;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha7bc0653af1ab091f614a524c196007287916bf7e674880094d21e62e98d3e41a85e935a4e4361c2b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbd00914998eb2d3b28166bb1e48acba9c6b8ed8895d35f0d863bba1c9260874c57cec764fe0b88d51;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7cb6061aee69b7410822d4b03e69432dd4565863d802e48474b25c0740338dc89e9e858f4a3e12612;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hdda0833f0e89bd8ee0aa416c4b92197227be440dc87399fca4474930ed067764ddb31b6395c2889ce;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h50b77f544ec1fc21b93479c62267f7e6672595fa0f0d24c9a4808991b090f81d07d69e63a731c4466;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6deb8229c48869d45d56393a2b61f969960fefc90bda55dcacaaf41e42a9c8b2bfba5ea445d7e6725;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb190d58cec8404d1b2309c64d579bbf7673e3871155612f27d72602ab0b268a8c3db17c8a1a80bbba;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc5bca28f28338df2aeab54f67600c9a62cc403e7c3905ae8cd83dd8d81c3fdded6a04efab49fd84ac;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he19594c861b19ca4cf558220375aa334a7ebe57f4798b983a7a6a33b4c5507c57b16e84737e28a10a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf2700b9c293f530b03596cc5cd540667d2b05ec4be1557be36da6289b60665b78778e11a8fd1f6f76;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4481d8e4b634e03511e1ed872e441408928b29f269e5a8bc31cfd107f48e2089a03774910f8ecd811;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h143e8af9085d6c6429b94e25362c5200765f52058b9d08254aeb45d28c97e5a6050752fc46e752fcc;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf68aefd91981f150c49cb4abf0506925bf38532d632b29a9488eb58857b827a88e9080ac640f4d545;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h497100750e4fc21f4e05591f58a2de6c191f31053fc3f8f6b07e45e6adbecf9d996a8f3780c8c8f35;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha451208d94dc2b28b1c2a8fb74bdc88d170ed8bbb0068c8848ef2002ced79e919de9a4e65896c496e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfca1329110f0365c2f912895a9fa9aed7411b910178afd9bdf24b1ad959c6640f1972a8fd98df4ea9;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3532ee16770e5326f70fb54af9bc74a6358a36780070abcbbb3fe27cb641103bf8a283b372e0b7374;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h79221af2dbf0d229674700ce781fe3e717b4bd9d49e888744e46003fb268a97556a3f03fab67f88b3;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h165d53b5bbeb107e42e7b74dcbbb87d46897d104c05ba61676ac84ee1f0b63de304103d0169041dca;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9a61dfa7981b10e6f352ea98bb198ade06ac66c4f87e22c5e41cd02246b16e816a1ffa28164a12d2d;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf129926baec1010aec64fa5b1b08dc5112c05cb3d07a875bfc162f612cb4c3264631e2bd40776fe38;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc5ec3b98ee38e8b78fad895bf25b037e11571e2fa91d424fb8956d9c95f6ba95d3259d29e68781608;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h80991bf57120d7f87f54df3b885b2c3dc3e0d072d47cd89781c388c74f1b6c74f5d3aa49438bd0db3;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hec23901b95a80681253c7b8540af6f46a2277f931947036ba8bf22d1d1e94ce8903f2aa628d1bb0d0;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h158ae76690dceb1d19e0dbbe4431defc0b5276eacc299a213000617640cd11134593df43d03b78ac3;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5c8441b692c1b9c8e7615eb9dc9e871182689a088ea17e016511c2a8f1832c152fd246ab5b1018104;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hba2edf8c90496819815b66382b2956ce0663b740e563209690481693e51ecf118724b842edee892ee;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h16849443fab8d06218c194e31007a7f390e0f8a4374593ebbdd39f140e88f48fc9c020fa793a0023b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5ed67a0f1a03551d632ea40e8788751d890a7a775ae13c897c04f9a95db63e9856c716ef4eca9ab4c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha8027d79bdf90fe4abe09eea8e2b0995e6340b51427608adccf4060ab9b1961ff36c8a1d518b68e9e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9a9b4eae230bb1969b681e1a7adcf1cfd5d73d3a750a9cb76f9bd45ff7ca41351f49fe3d3f4542c4c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h984a4a79c914b40cb56f06556c52abbed5f4e8573addc83f51786117478f69a1e8d21c7f8a3cfe3a5;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h60e8c1fc09dd4cf47cf16298cec7f77ffb9f68c4eb49a50d018e0d7ff421b5e0f62264f918f4e7a7e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he2c6f940b69953e2e79e55c14a5149c0dfecb2d0ec1951ae5a66a935c6259721fa1e6a3824cdca6e6;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hedd4dbe3bbb01cfe8f85dbc826a9ea8be6ecff687db7dd2e2e098aea13f311bc0451096ebf4fe7dff;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h18e7913044c4f7e20b004c6814c7315d1b8a34f1a9bbbebb7549876e845cdeef6babb9eeb65e45ba;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8613b43e71a9fb4808e9c99733f484dd3c95740e9ff1ed57b6ab796ecece9949942146c06b7ef641a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfce5f8f04c25e9ececb74c69811c1fb2d769a3d1f2b5f155e1c728d9f04a9f38a6dd8bdd86f5b4898;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4949686c83189c6261fcddff34672872b3f0d8730d77d0e04454eae29793c1edc85664a55d3fde441;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h958f21431fb768ed76ac34eb633981183268a62643ff82e11914117dc48aed665dc23f78ba7f4a692;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h674985a58fb06caaaba03ee4b539a9f9a93343af829c1895c1a090d9bac47dd41add113fe65e58ee1;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7e0a21602ec3542275cf49c2be21e3cdb01e36699fd85cf1342610b8df1b95b483a31f230976fcc62;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h996a78bbedb033e7b951e05e46e3dbe59e2c80c85b6607001f83249da839747d509bb664cf2496eb7;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd4f97727dd9a9ebd273f0d393dd9b2d78f92d1e9816dea859e542b493c890a4a1411ac69911bbdb8f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd4e6a4aed02c07652c2c325d5bf87c75efc72e07c613d652cdc6a2cc8574ac086842f29bb537b5466;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h35cfc3f6e9f94aa9c2eee0c854da905fc4aba9d139cf17573edd7dc1a9a2ab7490b15a37714c6e50b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h29803d4589f187a94e56717ede6edf42e1bf3a1ded0e7a8e215f33f7ee74771b6c9c1ed11a9450a3;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4ff3f585057f5cc78ce7188c782530d62cdc83b90590418865a92dd8d130ba36339f116b7b379ec8b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hdab6ad8e2cfa16890c24edd94271d3711c501fbc24693459794d0f4d7c7703bdca99fbfb363fc9b94;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h22ad8107bc1351fcac28fbc47574d44d4d0df03d47df3a86d1195cbbddeddcc50fd3a5aa3b833cff4;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4930abf9c2c47a710f87a08309c01c00b265f9507d1b7ac9618ff9d31beb4eb171e01e75e9879bcf8;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7d5b6b3a46ae23234e1bf70f585dddbb7db26c3ee7084c1815df7280323580bbbd94185b28f6d6c72;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5256c6bf0575337fe7461c27b203503b6afde66b352f2e1a372811d6c5436231103706c0c0d4c2a84;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h241718fb37c0adea678863506f859eb876c8af577a18e7dbc550935efda5d28239f4fb922d4de4618;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7c9bae98d9d31f28e0f86f5a15f5c60dc65719759fd25242bb67ed22ec40c2f374f7ab63f1c213ac2;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h891c7e305990e0240083c2bab5a3e688ec08df6911559c357a34d1554e8d27d73158ab171ba4aa21d;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h39411caac5b44cda9ed11311a1c1cef1bc9a0c8beccc47f2f3fccc8bdccb53276a0179c39298ac235;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha31ba767136e00b86590866cff22c7398011c63a1df346d9a38a14f8d4215749ff9a16c5883ea1d3b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3d8ced61ac3e1fdd4052050e7922184e51193322753af3c34c9d7b801c4f3c6daf99aa6a8084c6265;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h30767114c9917092b45f60fc66e906f85d68122a29c0ec3e21ed28e466d31184fab36b6818e7e6d58;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc83f2b50a0bb0bc1b55d51935c72903f03bf666575e376eaca5ee45d20d945b529ab7f92c0b5d93f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8d53f9b242e02e04f6169329749cccbf07e536fc8dc0bdb02c0c29ecf0f170153e686cac75881d4c0;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha3a787fbe58c6ca5f3f7925e192964ccd8faeb64ad7fd313f354d27bbb459d26ad068e52012b46289;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3bf20acd0be455a7c32b1fe9ab41767e1dca2871068764a0889ae579515dfb48e1e298f748f26bd12;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf95529cdc89b6200530bc6964d4c450b645f5f85e5d5642d3869266b1d49f34385106fd5b2a024adf;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8492b26fbe779d5cc3843ead7f443f04719024c824ec9301648510af36f8855b13f12f87c6b3c18c6;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc8bc16e2c3203527c1f7bd2e3be269c30de561a15cc37316bbd1d1586f4bf61cc598eed621fcd5f94;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h10379cf4abd3d87e0039f0ebfb8b9a2814b4f2ebdef5a08d15acf932d8c8f42d5120ea9e5f732ee44;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc022148d356f9e66edb6f55075537aff55d22b45c2dcfbecfcdd51cdd14197dc449c11afb11be3b91;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h53e5d8bd613537c9b1e5a8cdedc4e69159146cbba257862cf518ab3ab7bd983adb1071d6c9dda4304;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6bd6c5a189593509e537bec0e7b0cc382a526e9265a255669880f0d6660f6cfa2a5355b6dd3a58048;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h95759e241a51aa8e2a146768b9b746725fb07f6e38a15916800f960e6a48c9085f7a7a78bdf743c2d;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h82f3716a4935523e6b3eff9e552cf71fb73c2606ce98d9e81192248fdc84c2daa17a1663a9ff7df1c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb2236dd09b548a526e04f932f2f73cd5d909b7886edfa8d65f2060edd7118b7e79762625ff305ba4d;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd861894f87b30b159cf643704e4b66756aec35bdbb95637a06616227e3eff110d8fac0df6bd64945e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf203fc8ca10fc45281fd7c8cd9fae51c9049835dcdbdc23469241858a9075abb0f4e05579eaaefc72;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2839b1cf76d972b954186690c44b8e18e68f80b3e4fbbbfe9e00ee65b4c80cc234f5c8203faa68531;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbec896080898166a68fa3ff263d7d1ff2b120fbacb0a352e423d1d3aea41f10690722cdd4803948c4;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h63bc58c5fd8343a9f3c20a920a459d0dd9763142ed9c822cb15003e483e41d210596478bc63ac422d;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9724e804accb66ea7f52715c31f33ddb85dd4195f4ab291a83f8255c7c4c7749865222a37c7be1b6c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'haaac51523d1734f0ac948f9beb24184ade5e756b8de64bbc3f2ccf0e179483816288df38ca0484885;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf7aeb7ff9ac0e31e04103f9bc5342ecee671a81a1b13d574a27867ddb92a1b3ed2056f1862735dd94;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3e2b432bd0f46bbddc725ec6c8605f797f9fbc2590beb1e957e181ec89e05c7a19c497afde2ff1a55;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2ad865793aec8b3cc0b676a30bad296daffbb54d71a9093c8313432ac68ad7dd2f661b8dc22161041;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3bfc34ad02d86a6530171ab7ceaf3427cd9d1e8f9c2f878a3734965dd152b4471f756572e75d2c7c1;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5ef2b02eada2cfbd20af18ac5495c0853988914c47ff093ad8081fb1adbe5599654999f60c0e0ae9a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd46ced912fd5a86765655f40d86879dff6766ee402bf47bc869eb1fce588c90eff5549a1daf22ab0f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd2ad59095e37a15590db22a6b02043750e85f983b83de74f42aecd490ea40c0cf97d1fd9b55868f10;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h167fc24505344fd5fa52ece562e463daa5b578649a5e33f868b9c9a25e393c08546c2fc333b63b3b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he550c8850684b67e93a78ab5c736921f7d281f02d0b75f0c116ce4c2eab85ccaae9524ad64c1dc4e5;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf446d2822ed99f16a0331bb90b8df4b09cdd1d691420359e271b245efd2b1cebbb9d8aa3684cb1e14;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h923fb00da44a9e6ed329f377eadcff057c18a54eb1ecf4b17568c9c5169395d1be732989612bbfbf5;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha7d2956502354e6afdd424c5bbbdb015fd66e31a0aa24a8857a1353d5d426bc6bc4ffc190d3f9581f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1d0a59a0aedbbee0485fb9441e0b262464557cc1357f0e43510a43d85407ead652961b2f580e12094;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9e140c4155bcd3216d14e4df4f2c1383e8341f3642cba72e7652c267a61b62cc41436fbedbe6d16c8;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3039faaf22cf50b4dcc7d36d3bb2039ce0f24110dac59c42a930f242820dcef5ad0105704aa8df9f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hab87c089d117a6f0ba518d011b41eba645b50b2b1d5060dad3d9dceafa8e552a13baf3710bb1a62a5;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4c7b1af12262f74b949ac4e21cf409718b26dd9d1a14847ce5687d07af5bfbe87fa6e4a2167daa508;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hba52e5ff5f353603ee8a6c2276c03f79348e28d1ac01881f82483aedd3407ab815102646ee4803056;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hea33c6c6d9ee139ff8510ed6249b1c5baf58b37af3a0aaeedd0a8d9c3f701fb4dec638dbe79a4fdb4;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc4a473e9b6335c9afb93987eadeaed1eaeaf2edcebff14133fedc875472c53f7c646c512857d0aad1;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf60f824009f3476e29aa2bd6626d15f2cd1f519a6cbed82fcf933bdc5f1fbf9b4ac2572e2110c5810;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h18336f7d20c5a145109d6af3fcd0ef4989733f976dff8c5bcd2a5637b214f056b900a894f7a90432c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfaa4c94eb4372449aae4c2fd9a76077d7a2374ba40ded493aa7dea6b20dbc41966f7f4e44f4ab7257;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h36b4f293fac8c42a7392a79caa552cafc961923cc1ce1eef4c8ae66078044a22cec7457307f6eff48;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he59600dddf45174bc50d2de2072b47c5ccb2b6dcb408880036fa6054a70bd75d42cf025cea1ad4a73;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h650b8a1d1d78835e0331ddd1101795b35b46e140fadf34933dc5c9157d0c164e10d4f175cb640da3f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h46e5394f17b58a32f93320976187fa530ed57f1b14c3202002794d0c9eaf95bba6f0824c54f62d53;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcc246357ce1ea779515ff3847c1a830624ecc3c08a1085f9991dcb8a9c7ef7b60e9d9db66617c6e36;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hae03549e654880552924ecd271f08acca8759e59aa5c433a8ad7eca62b0f441159361cd72abdfb41d;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h895ee1f3036314bb904f56eff774afea841481044119d66e46d1b98435306c9936a6f2c6f2eb917ea;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hdb7430139f5e6c92988c22993b0ad55edce297cc727c2580e8497a00aeec9b2e1fd76bd7e68bcc531;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4819cfe46919d50b7cc64b79a163bea1b211b5129841a5a710fb8b449a68a5bf8e70b5ea10bfb2eff;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h11630aadcc0ef3f74e508961d4808e74c739811d3a363ce254f4b9d937c1ea7960999576321242dd1;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4fbfa8d54236c8316d03252f62f58fde307b84f7c1e31f44ba192dd19207cffd49c85b32af78ccd1d;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf46aa419f7c4503624db5b3da8ee4d5da56b79aafb5de07758980af2252ad44ed7f58b8a3f701eef;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8caa166b2a493a8d72da680272df6a690cc50c1ee7feaa4a0e6291fdc7465df7686eefa200fd0344e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he1f11cab3f05b28a75235925a53cd82a0d9187e813e88539529352337fafc1f0e809fb03dc14297d8;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h409ab577cda2156fa5b23d44c8c8847f391f0549389d675745c1fb39271570896627f2cd46ddc73f9;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2cee4555778526395b1f213cd88e516802564d18d8a631d9cec1bcbea5862cc20c2b332b3770fb0ce;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7e5d1aea79982eae7c0ab011a55994557ebf970bf7dbc2493553015e4e1781ee0ddc9f58f5390d673;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h89b5bffb984d6f61277525e02a30a2a708596b93b35fa2448755b98301013b5efede2bdc85b71b3c0;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he9244e8dbf14d9a2f49fcaa6f3e310dea7df68e5135987504d297d885494cf8730590d5898861bd90;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h894af65003b4fa82e547a6430d892a56d6c9bb6ed8a7c2eed7bf5e84e82ce766ca5bdbcc51cd89b41;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h67fd9e57ca052a085c4a72b9449114d6d63bc391f9cb8e1cb73642f05402f1f62ad4bcd1ea26dae01;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h70c0fe6dc9214f7fea07be5c0067dd6ed14d04062afd6ade54f4b3ff9e491c3aff1ef0df53d8ca855;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h40cc4e1c7b6e4dd9fed0321a9b92b55dc76e63438313cd9f98266337097497020301dc64f52495eb8;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc48b5bcff633dd589c27db193cf883b1d54084a3ae0d074bf3e8213f2e6b0328f8658f51f4837f7e8;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hdcbc6c434d897f0bdf71b71e6285c3c597bf4101caf8f7cee87020fd9d08585b2c88b7df4554eb952;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hdba679ad931b63d883c59f855656c4ec1e3c2b27eb49d26ffb447554f3e8220530f013240abb5c152;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfbb6bfb986c635920cb9fdd2bd07132772a53c1ee8999951e12bc848043c7de0ff7121bb1e572e10f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hdd444419433501f48222399d723a500856a38565b2376be39f5aa0a7f5bca71ee62ae90376caf9c3f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hee26716a56fe2b65f8185ac9864a40cd732482c76a56ffd27fda012ed6b13c0c292740de5b37bbc4e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h26a856fea5eae39f6be6673ba11dce5afce665038640f425de52de7945a18a64d59e6917e011a2d6b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8d5fdff73f0649796aa0d9abb9db6d46ad0af373caeb063bba3839e22b7f6653ab9978f33781f525c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hda1981a7bc4d229c8eaa7093f99dbb53a244d998287d5c64242181b5812c88a7143529adca5d6e637;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h49b14f10fa872848f02c3492449e6d816f4428b1856c784bdeb71406bb17f5f4eb3a3c2d8005373e8;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc59fddb0271ad42e679535c1eb206303a15dde0be5b68e67d215f5a9c694261fa5256649e660c4cd2;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2fc2e8e1602e4c43389543c343f6380e8f9a01e45af3b98bfb1047fd1a85422ee1c0003251328276c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h35160d4cb7f8b88188b7d830b50fc2e0378b25377515832a6127291fc2f6842732fc584cfe19da54a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb530c1dd0040e625befcc6e93971f621a9bd56a1904346bfb74d6f85e83aa8f04e9bc6023b72b9793;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd6b4f18efcbe5d3b495115d16a17612fd0a9cbfe0a1732a2f125fbd2631fb2e9f7473dcef8d2b48cb;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2b8afd49ebae0dab9783d67935b7aee34d47e9e0b688855fc1a0ec26df90f2ebf327a6fa8b7ac145;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h871175c5aac6b8e8f04c57007378c0288affd0989cce9c10e2ad45df4747e278c72c30d87380bb565;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc19a147a55937e741fa3d36c6fcb9bf30052660d60cc11f7fc0b47eea63ab571641610a2ec8fe2161;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h568afb528b10955c855ecd69b419ad3b7755b97a54806373143ac65a7d0a35f053cd302469ab960a0;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h706c12a207dc5bcad8e91edc4fa33853fe44f18f2b61cb2c5ef0de9380c1571e28a915ffc58f607b5;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5151252ab9662eb63793a092922f23b940b4f5d736a50e0ae2a6ad696dc10e109f484d30afa0b2648;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hef601ed523ad3c26f4bc887aa7a08e5f421e3d983f96c548d15783bfdb608e2f337842dc4365107f3;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6d17e9714b441a8acd33e3fbc4d83d273c5533f099b75962f0441e559a20c27829196ae8bcecdfed3;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he2046acf235e431c7ba11f8b54824e07c2c73803523e9c011619ef6e181d5d57598bd9ef7f9ac133a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he28e317491be5795d7a2aa105cd3ca6a11dfa4a813db98049c44e0832961436bcffda42e4c8bc6c63;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h52a4cc2799c134b384d4bd3d610bfc9167eff9658f1f00c786f1045c29ccc2bd2a97044a85bd0eb31;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha54f85e1332ad394f47d7ec3533de986be32b7982c9942721139faf21a1dca3d933ef606b182c4149;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h48526fe970b969e6428d183e5ecd2198d2a7dbb1125ffb5b0edc2fa6548830ba5b95226c7d6898897;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h21b10e56a8faa48ea9fc2add7bef9fa53ed0d4a3c7d9e92360b1eecf06d1c8cea7da41c285f5e7110;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h43b514ac9d46f41f87226a7fff80350a6cebdfbcef56373491fbf41003e8e4d5b73f4b012ad9e808b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc489d0c96613261786ef05dea4f845187089ea42fc14117432c41da3ed007edb93f0986d89b6bb03e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd265b90027a382c49ae51a1138529d4d9084d9794eda167d6bd81fdee501195e9810b1c99c9331524;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2be1bb275c5bef05bee9f7f9a58a645284c2095019764ab1f49670e228e95a2b32d451e18476cfd07;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h64ee6b6576fcfd3dc55ae3849762f852b9b4059a0830676b69cee027e4b77e223bf74fbd177d85d3e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1be0e7f1bd50232c40868df16f92b97f9f1ae958ac3847e5692bad52f71f4fefeea9300bfc66b7c7f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h111495cc0fe8d0939803da3b06c04b17aeaed4283e2fa46fa658a592eab43db421b16b6957e4096a3;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4ebe56052ca82c88e25941d9a8c24cda2e3047b88ff509000497d903bd52d83f9be3ca6fe9dea943f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5388d3cef83593813bae2b80951ef4927837020e78ed6f8dc25bc01d143f0607a7243e70748f41969;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h57d666263ff1b2cec37df31666f285e893c13ebc29b14cae40b216c283e5c377afdf9b79cfa92823;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb3d68a039a67f2d0b41a0e440453b9310b2dffac07bcd3455c4d3d8e45aa8465a1cda659d0a8c220;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h224dec906f4b5516ce0950ab26d7658274d811dfebda0ed6c5143e884f7e62b0e71391c7e29a22d42;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1eb8f045e4d4b102f177c40cb3fa27aa03a56713af14e38b9e216a7519b7e638f4883fc997c2605f5;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc81e08a62bf66fdea56be4130c0ddbd188338bb5a4a7344d5c62ac039153389fd1ec8332ea13fa625;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcf68ddcb95c413606c8873f7704ee4fd94c42886f11d53bd891366e97e3f15a705c9195794fe81247;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd85952399cafba1d4054240fe342f4a0d19046e8ceaf6aa5f1869f79a5c4098d15d816df834dd31b2;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h670e3bad43abb1b8d596d8e8bd43af6533e68b5c69cbd8a74cf24c3a8e1bc589760f27ba5b2b320b0;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h137de38aa8bfa24b51bcf5ae080b97931610918528112224dd589a7d77432a8cd895de4004bc06c0b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h27df5deb48f8ae9e4c7f0171968fcd606c9aa6da35ba79c3e512634cf64d6cb7c579563e6700622b0;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h64861ecf869af8fbb16ce50b0f36dce17df9341c9ffbaf5910a37dcbd2defa5f38577b69b3dcb81c4;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd18891a39e0610f4b0a9f0d78649720ae529c42b57448a2545443475ddda2f5460e3f0e7e2ed2eafc;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3150e64b12e90803ff3a34fdbc313d61e9d7c905e614a757863589c800453fe80a9eac8e6ed28f3eb;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3499b1dfcbe7fb4e6dce4c04de106a0d63906b67bb67c3188a259f72763b5f6a1d2f01d088c27de79;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'haf5f0ede647384f4d1d7dff6a57ed35412732f20aa53e0ad16098708be3710a1fefb48ddcd779200f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he1455097c73f787301233db7e973b06c29c97543fc3a66963ae7863b97556d0d145d95b32918a8d4;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbb3346b39a7381ce113811493ea45b131623e30d948c56d6190f21dcfd49f774f9592bdfc79c4f730;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'habe749827e41a020876e26b563b5f9815de726c06c6e74d1bd9c374770a0f27fa58fda80e6f1d14c2;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5e3a93f39669bc0b8f60f17551b25c250b7728b0bb834428b4b098a6ea62390c8890a4671f884d5fd;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h948109dd1edc2e51e0b7fbaa5320ed2a3cde8cc4efc7b6a64638ef8c707a8a33953cb5b35388e1e91;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb0cf76db6b1840fdd32241043f61272ae4c642903b681f71aa4744e5a0e66976e7b505a44b216d314;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb781805ba6edc5016147d59eefe58fcfeec8e3e9e030ce03ce301b981ceeaf6eeae5c7e8f7d2a4f6a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h360ab2d7e37339e6d8f45809b1e8ed9dde54c2ebbe56f1e9f172e7b7495e16ee3a47b41cff3636c83;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd5d0a968a1bb2155b11ae9960ad0464b01d89d700912d12916cedb9217b7ce1c8390e915341a57819;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9cedec7faee96ab7b32728aca3b4da802ba0eace69324a2c8c2da2a6e1cbaa3f01c50eca5ccd8aff3;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfb45adca2249d31eaf031be93e7ac89a7a8c6782b21daf98b6eb760c6d672c4f6c16e387dc2920291;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h435f6870e8f17d061d3fa612bfdc16b681d5b4e100f7b7dc93f0bfa06558f91da7912abdf354d32aa;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcdaca9436348a42d4f61820ba62f9be83b707f3380b5477e2ef0030d5804545c01382f5d13fe8efe3;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd32d9612b9e1af0e5cdae8de7dbfe3b815786da427aec571384492c9393b75de34d16ad4c71154f2;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6ad24972f50164308c8e8a0feb00451ea5b76576c53ba8be81915066375c47c7c824dbb1994d093f0;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc0618c641de8e377f406b046dd84fd84cef0212cf20abe761eb446b830b40a96b95cb8a5777c4f63d;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h753893d55b1bbffe1956d2ea745c7eb261c4a0d766ab8ba377927f86547295e75bde939e63cfd0833;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h168aa6098b39ac4cd839d902e0ba6ea73a8cdf01be24415cf74b97f1b1dc0efec535a6a7acf704234;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1c59534b2ceda03976659a252dab201aabc2b79f40433180e079035d476ea61e1d1227e282056089;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf3581002a51a05060fca3b09bb89c3bf036f4bd1b26e5bbc27aa1c17a74fd47cd9bcaab0184c24748;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h783ec1e16278df6b61cc206abfbb91772aaef765033e4bba64041fe221619ac4a8c5e50bd3353d6de;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3e6d83c429f5d84f50466cbc15ec1127c03aab587eabc31189def4c8e35a76629be0effd80aedf20c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5e3273312e1db18a3acfcb5e4bdb35ea0073d1cf4eda5ec97f501047b74d35d106c5b254e96fbdae;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h192adb7b21bf42a2a2300a83b74a2c593776058610e673b16c022b4f543a66a1d4a8fa58f441b366d;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h75aa71468b526ccf38317fcd44a1cbd8f252241ba3190748a6e2f2b968fd6446fba1cb850e474ee47;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9d51ba8a42c571cf014c2466e2860d408a0b51494d677f1fded06cf682150990ebe11e61fea421435;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha43d1b1efdc084ecc445ad967e92b06b2b10ddbe59a97c2c92687477b9b11f6d02b2fc805313676c4;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h32b521dc46778f1d6934cc210f9f130612b62a2f104ab321331dd47802e5c2c879f828ae71b2d1d8d;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h15c92e966fbf46a7da99fedb0e4720329ec3e88df289d42e4de329e981334f341ec1d2e57d3aa9a35;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he3fca009105d1e430942986f422d4c16d0e0fbef4c2f5cdcd268b554bf299de1dc492d042c5486bce;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'had7074d3e36a83a3aa76f70316016ccfa174c0bce904452b3519ece9dd7499fa4378d61423a7f6b2b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h90dcc0cb68aa706f0fa03abbeced48f059a35f95cfcbea26a9870cce0dcbccc837305e3f0aa870f4;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h25720f387852e06afba4a4dc1a5f270119dc2e13ca2b27eed273673f594991df614f4e1670854b1ed;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h97e91d476af56839de073f59caab3fad300ac6399aa9ee0fa654cdc4edba4cacfba9812fd2cb05a59;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbba64080f6d2fd9d3fbb575f891f4796289ebc52780e4bcbf774f4fbf4269ee6def685bac4c74e807;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h212b77102803a82465b9f0ceb37408ea837e69b414f74d79d8ed1dde2d5b1f60396edb158258d131f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hdf171ff9c90d0fb54e644cf53bf6cccaf78b504a705950b41076f9262f8accac9cd6c986a2c2be44c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha4ff61c4c48df2949c434911338c87e249c8d3f895dae9da25e0bd6c95d0db76138279f52ca1be1a1;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h92da7899b4cb9df431e93de2495dfadc71e626b9559a7bb6da21954f7488f68494c93d66db9782bd;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h646d9d6a8826a923983d4162a7492b6e2d8a37ce3537a7f7dfb32dd7923ee30e7435ebf8c860ef220;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4f8e5922dfcf58e797d2bbcc111c0e37661d14d7b15abb6af2ece39a4b0ec1f2ec840288e6c7daee5;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4d7a8ec49e4154cc3e520bade8cd07794bc85b2738d9450eeca42453f203d720147f8ef52b4392108;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8bb0f0e1da84edefc61c3e9543c60860c08c48b92a769f6e306445e4a432d50636e3763d504d1e27e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6267c7d050ebcb7a684cd34fe5a8b0d2d30e6a1109427aa4b0701e17103c74bfdb7eb468d1487e569;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h42bf203a68eec127339fbbe18be46ce8d3e89afb90612c5b9169bff03c398a7b1dc95d10da1417577;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7f4e3840775e6e7b93a6d0c13d6cf78c95d1f467db4cd6ddc0a218c28f88b6e2a9e2d84d0b734fca3;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h70bf4d60d89089458097fa1c8f7d54b0aa2a3153a41bacb3778d409d02f9f6c5747df7c1a3b19036a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hdbd64ec164e8534167ef44f0fd5824d14d7bd6f75bdb5425ad86ea58da84503c9976c0a15f9c8a7ee;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf6c6b6cbf2a630a3fd5177acacccf9f9d019ed3416b8a1c2aa44360f162d4c056bc42dcf215ade9e0;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb8446926dfca22352b314ba01edce94e648ca17b2a6f8e21aa62f7ebea296b0e0c1a0d38a270300af;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb8823e5852b1f344b752ab6f174d965b2d380e357b95420cce0a491e257774216d45e53df510971a8;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf600e32689b2fc8adc542482ff264b15aa933bdb0125a041e5b6496460577617ebb8c8467c4b3cc8a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5e2d4ec4612177929f0fe840c108147e3e35f1c5318978bf0e365c33d4834d6536e340699e93bc78a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc822d94dd40406cba34ab1ec344b025369f58269c733b6b9ac71a025c65edf5e4112fdb158fe41645;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'haccca0994ff4ac7887e47b2ab67832771104e4a22708ede3dad163e3a63a519111337904254eceef7;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3dd5ad9a7066aee36c6527bf6d16c66c3733776cb632105611f14ca6c7e472eb405faa9a269646370;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h81a1716dd51218cf373372f9cc212bb86a1c44106d6cb64ee7d2a36cec5718c8db04dd5f2faf1f133;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2c377ff21a173bb1c935e73e4845ce9213e800cf3f194964347d55f463619d69761b03c4dbac83bab;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h952562d294b7c968a11df36ccc9105fadc6bfb73a7996431d0d1bc255e646a17bc848d603bc16e6a0;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h18dad6ab262582021f4ab55295a9017b828857799682be59ec5f0fd2a30914bc66da515c21120630a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h12d6e0188e7dd5194d13f10b2b161909ad073232480c67e40300004d7dff4c095f44d64c36ff534;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4957538a298987859c6ccb99e14c71ad32d804bd866dcf50c1f3d0703c19de4921bbf72a0c0eb955c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd67049ec6ee728176ddc28fdc37aedfbefa27cae8daa90b69476482c19e5c0b736e3e1032a72f721;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf0426a22ab0c466de6b28727c1453d96e953fddbac19337e1b68aa811c9984b20aded44ae3d310cac;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2af95de743fe92680eb332e61976e77380734bda749a8ce0389a73dbf005bae9f3b8ad5a8ba10ff62;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4ec8cc496778b7d10b99f9947832f1c72fea3f8b8b522d53a0fb3cbe34b2a02b3c16451ff277c039a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf58b54ddd7439fd1bd7efc1e5b0b9b222dd7f0124562913cf210e9d8062860d643ddec94285dd1e72;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he7ffa5e7207315e7add90619798a9bbc46ae197b1f863237a54aa1e77e2e69f0d64b0793fbdfbc12;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8e3cd557c5eca59de46f6b47c39e212833f8990d193dbad95e81885d58244a83021d642194d881580;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9d4e9965e6f08085bcbdbb590265e1f52bced9b7559c4590cc684c1f7ccbb06a75f55ff5d348c16ab;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5f5a111109e9ad20fbedcc251b07a89d64b3e0cd39434bacae3edc25de36fcf0b59b639b028880c3f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf1f11cb9b24bf0a2283cd3298b12ad4e16fd2032ff0b4a8fde809a3fc764fb7b4a4d3c5eabcb87d80;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hdafd34066d8b57601d9f0c8bb4b153f988c8e092ba10f4460be395d46907a8acd470daccc13d9aec6;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc2a11574d336e6454310e60665f41eb4c9e244fcbd9228d811c328096513cb1225a9013506a41266;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb21d11011522f5c408cb267e9ec79cb1123a4068ddf530381d331a9e8fbd115063725300e5f978800;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6f3b484faee5b2022946aa3f28111484af84fa317c755a327dc893bbc0df509688ebc4c37ce8943fd;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2bbea6888ee3de8f2aabc8767954b558706cad303cec83f6f92617a3ccfbc349834e982ad61e9363b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbb731658951b734e81f3e6289df20f4ef04490f7ec48eed99867dc5265b1a7630da10d08a8519d347;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h76e7bdb189a78f23fd316a1f08c0a436f095949d40db61a42cf2f7d9342b7ab9f832af9022d4d2a3f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7a76f323e63daf31a07f705496120b0c5df3effb020392f29aac9264cdc7b8826365e22dcd475402d;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h91c9903504e2202806f4dfb9549139fd671691db8633cb510b51f66753b8e502d77708f8986486de3;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd8bfd748508b7184e943daf71711582e5f29d492e33b8d3aa1ed0b9ddb48fb46aeb23fc5705a60334;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1eba7d43037fc8b92dda20b477eafd7a06fcb13dbdf0a6bd2f0aba34ea01295bd65b19b5fc0fccd7c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6b3594792093c09937233d6445121e8b9f64a3921bf5ffaee9bb4bca4f884dd486e2fe3747aae44a1;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha95a172792221b4a4bb0f8ffb9f6e25937ca0e674252431be5029ae162d25351aa9897db94784a2a0;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfbb33c33d08a081556e90bf06d4ccd6bc51c568f48e967557e77322f39afec0873c7a777369b4f6f7;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfe14aa47661eba2fd20320e473806d1c05d634c05d78b83bc72964590f3c4ac9bc3d48eec1758975d;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha875863b47827f4645e94928b1f02833106aaff14a26e3164f215398380bc635eb4ab54f97f6bfce0;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf055672f8530905a7d83101bc94e8f7f82802ef7db87fa4af7df8e1b586623192506567f9d3c3a2fe;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h83c052a9d665a8b5f7bb874997e6e1fde22c3954292182ea935f51f54cf5c1e57072b4e125cc71f09;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hacdb563d5753ed1b81c4a15f1060ec60faa28afcf1cb40fb118f7345ca91396dc1be6aa655b80b339;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8ac371a83a980280251087dd65a579f0435f54c82ee7ba7cfbfd7a307bb931f2b157acc9fa08baa53;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb9059152ae3d2a8f5e26210386b4a468582d59bbca138a8d581f4989e9fb9d71bc83fff20f54cc726;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb49a07cf26093993ebfa4263148fe591bcc88a38c8c681cbb24534d628c73d95a2222d6d54a40c20f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h608ddd9b91d658be1975f089f20294a182d8ffae8e8671ccde43c05df0062fe2dbda3f78b256414ef;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h10aa1b3004b0d5f9ac744340690341ca7e1776ec344f967b5eda66230fdb899cd56d0a5a724233cb0;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h98be90d42abded096bc009e7788e83ec8396d5b2dc4e7baa872d13cb2984db3274733abac25479bf2;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3c5977e287ec0417098df96a27e7d06cb67675ed1e2f60a4dcb60dbb8835226d28bd3df21c53d7294;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he9296b5d3d7b7c3d7f922da5e3c1db5ce934acbfd6163af456a84ec24ac54562e39b6a85c300b7439;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h382c0e958840e83093b1761fb6118bf9c3f9505c8243bd1390a1865c99a17d875a4673b74d3aa3fac;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf9d5e6f4f0878be5c205f6a3c8010c168107735b95aee08ecc089e58f02032ab9abff3ae94503f832;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb60d66c86a139946aa411024af9f4493d458205461ea5596b304cfc838b09b719358cb4420bcf77a2;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb604fcfb36cc7cf9e8d80af54847e0c5aabe70235aecba9733315d51f247489ee74aff81e74a38462;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hea2d830e36f43c4b7c3296725b48744a42adb620d78c9f85a6bd812ee937232fbf7140d5bc6af138a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1a45344d733b7c53ae64acc143c895f1f7dd0fd1527d93e1bcab6eacc368725ec4ef24aeef1a20b18;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3cf5d483ddb078ffbf59cc16575172e352806bd2d306140743a6c514d4af6958e3fb546d6b0f9dce9;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3334f52e04096fd5dbebfbc8b63317f383dc5dee29377086809ac349e2f61eab5c031ade93fc5d610;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4c1a631ab164364d85e642bdff02befa33800c47010bd82199d99bd5837ea3223ccb39f0c3e919607;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8c0f26567512c2fd152f399591000caa8516d109b9419be730a496a5ef490fda08f1fd3f3adaf3409;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h40e0f3aa66c5c31eaa921fa26f85daa2261a3ebea1b36450686c4c851d48d68ba863434267f1b4330;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8b2f6da39a3a80c0a9711347a9f3b0de9ca1acd0b07c9d98e991d7eae49a57176e2754bad26bf2ed9;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7fb50b2fe666294bd9190db30e812b7cca7e98540f5d1f1d855cca23c9109f25f5321febce5eda1f0;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9f255031b97a54cf7b0530b88a9143eb9d73e0447ef21be1e1c79808966faabdf81f6b346df5fbb99;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf731dc971bbe5305c35c9406871d8dfb41d64f32127507792477b85e38898d4e9672408010e12cff;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2e165610497c627c50b1acacaaf3b91919d3fd0bf633c4a5c34ae04a26ba9b8680ce7c666fe79a5fa;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha010365f17ac4741b9c43d4f3b378f2bc6b8ec49fdbab85da6d7ad383dcd37ede0ecdce7e00b5fc7;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h29b6e6fde396bede0c21c60e569ad87a4b0ef84d1ac2faa4ffb0d918426f04c7a8715f8caa41aa29d;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he65943c09c003752001167d0ce592419036962731be03856a84921c1436b1e1b4692de278864b38c6;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h577a1c7774a16ed93f65fd4e6a944877ee24814804aafe98c33fe2ca43494c8b01008a094d82b0fc4;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbdc9290f13ecfbc1f65df432d18ca3e294dda0c19ac150be303471e1ee2c023092151e842f3822fb0;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h32d3b5c15500a086edb492fafd5720b6b42e1a68713f6af2081df6cdf55e45d4207c554f549c73691;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'heb9941759332cac13f2d881073b30bba9b9e31121b0f42d633447c39429e1d026d7f16cf9eef9fae5;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hec797832672f66c5fe75bd6e18d28be9b5142e47d5000ff55a669859da4660bad8dcb28d50bc9bd86;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h63f38c8d091f6519a1cc4f75a328a38ee345d0b1e504c9e369d6e693df6a2c7325e4c8deead9a74d9;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h14d0e716fd8fa13230d14d2c45d894fd3d0a77d7a1f658f2c0250be0cb98bf850d3b9415e44660670;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h55e455b4d5e37eb0a0ecf8f9eb7ef9c99f0881af072a28407219b036e3d7a4c4c2955b3a0695aaede;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1082e7c7261c2f011ea1dc80b3d8eb799e93f625a06fb279243d1d33a25bca1ffe93d49b070383a80;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he7e2c7ee2bd71d2f3120b0a1efe4b81cfdb3512c862ea9dc8d8aff22216f98f0e630d77830f672756;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd0e460c5898a589fb0f80b3058ec5de27136942c1b78f2949cc34ce7de2cd342e9bf5f6506148a220;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1b65cf836bed86e1dbb48a0e4257f9b712ccb63f94a422ea0bb1184438e1500ffd610bbaea2ac3485;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h22c7a11d7a95f4d50c7b806770c3b67de7860a0c2bdfbf122eb043530ef5e1496d4ab6fdcdc38602d;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9bb1162e6bb9c0461e812d8929d815899d3e146803d2356cbfe2c575a3df5eba8289210c29c9e0481;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd8eca24cedae50d7dc157b8bae7cc0dd7a934cf9e7892cececcfd812fa5faae1b5a9e398abcd95b4e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2b24515f070a8c5ff7788cfabe1ac8df744b32d6d8f1a7f960bee4cc8d78322053321f7fbf85e0618;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h49c81beb0a04597b4124209801b7731c5fe531076b52ea684ef3fa94310ea6b69983ffc9a76cc5f16;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9fb5557bc817bfcd86769fccf1325e8ddf08e693bac473e7de78cd7688d820019652ec5e21d4275ee;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7bde38010f38f7314b048edbae6ed2b22e7c20cb2a5ba7cba7aacb0e3c6b41db5f6226a17a90a34f2;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h83308161078a7c85a1ee2b0887d3fa85327c34866e956e0ebc89ae4ee4cf7d73a6e8c04222916f260;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd53a880c141ce6219ec5b04c768f15ac76c48321fa0101e26ce6a7b3022b4ed3805b76d0ec8e38f79;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he8f908dbaf986be956541edc4ad4ca72954a4c978311828c9105ca3dc247cd1e92d5bb327ae519743;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'haa60c0510760ca847fa7b1e40d14f51891869dfb7c7f5dd8cf40a5712e08e3195c2938177753928b4;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h48afcc95c3eed67f86a6d8c419e39e76238dfbedad2034e0b536df15161866b9b7f839cb0da8b6cdb;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h620959f8c318507b785088e7888e5052ea7f5ca9c7453ec7d12c489b2a6155f7d21d72fd4eb0b9238;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7716d26fdacb129c9824486293a92070c4ac001aac807d26d0470c385dd52b45d5ad8bcb79d40167f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9264852fffa57c23044aaed4f39cc0ab797119c71d110a105618ec5d7838a968be748213651b0776e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8aedc1bd8d9e76fc8a4b0fc44570a5770e674a5c29a4c6516dbad3854fd1ae8557cf5b058de42deee;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha1d8db4454f0f403976258043fbd8a62d9491340ceaa8a810d9bf0ec276f8880865413600da795dcd;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h411b8891c4e74b6cbcece97fed17d5433cc96b10472bbaac076857a8a5624355a2e0e63ebec3aa20a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he2099a281c7f3da687781e1b06c51586292ce92e3ae3ea730581657d5c599d3ff44f627f941a31506;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2ed7ebecefa75d183c720e2d9e94206533466af09f2ded7af7125fdfeaaec1e190601995d13c97b76;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb6980df96fc91627a20de83668afd7023b0b10793c492cff6a022fb38e5d3dd56713217abf912ebf6;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4118fa3c4333acabbedd388f4a24e2b15fb8f854fc64578e024a7eb69a37080a05dbb6f16fab4ef2;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1ed2ee3f444a6a1124e208f7ca2b9458544af0ff86ac175af3a6a2cd8f861b5adb6c7df80283372ef;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h789364cebdd4f5b36e748080e4ad3f3a98696485352925912a7ac7d35b7ff25feb4dd6a9c5f853216;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf0cede3be589fa2dbac87ee8811f331d50469b53ebfd99d1cd6e4714c311c03d54bbe6020c9396d01;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4f320834f64c31d08808f792daf2f0186201dc5eb7d78c1676067ce3686f5ea77f0e12f91d489f6b2;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1ecd53d85f53cfed136f942ca3457ba80e3c665d65d4cb11c4bdad48d122350c25a311dbfaedb26cb;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h75370cebb8472200bb4b392b4fffa0e78310c989678598cf90698a39347f45617c5e55b52d4308b3a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h167a412c162441c26cc33c367111e0bad7e75993c5686ff2b5a6be4ca013de71db526c1f2c93377b8;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h61c9c34dc3ad7ff4a7ca7d6567db1a068c94db92f10ea6d26e197595159d77bf7f5ccee4c7596b2df;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6cacfc29f5f337d27d4237c3ea8ab53cb652ec507217dfca247ec59631da1d102d9f99e191f12fed3;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he31d06de3e38a3a7920614ccfb7fb2a44643109c32c971964d37432de46784ed5928ac08843bd6df1;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc0c03e2df85f00cdc7c14891fe9f7b787ca10cf873df747802040b5722deb060ede360610db96c5c6;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he3d8c0624c958a88806ae1e239ec8d362889a014810cdf67bfdd1ff32751e77fc8e7fae0e2fd59033;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h815293caedc603a2465207ff2d5ff8ef84257746ca4d875f6d3a2749739c5c5e94d3359c970d868a6;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha8107e22bee260df93a13fea24bf504ca85a1df6bd6c93cce3140432a5f32b8d97b2e8472f5166d2d;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc7b518ce3a2cc624d936f3715d5f4bf8e93838a98cd1d664b88562fe93ff7b2ad818a477d86874680;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4dc2979671451cdcf839bd5f1b605e88251cbe318a130b4805f1b3f19af1dd799187ce7998ee17d8b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4f572a47f916df7a34d36191e04321539a69c563fb29c693eb9076fa3e76e187f1e984482239a76b8;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbbc3f47ce869b4b7daae12c0f5c823681e62b1ca10e255bb812bd19b4d623f03baabe70ef7f7a58f9;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h13f9d7e7a97e8cbf6d8f17a7a61de609ea1e3fe73bf2ad9ad31ea8305606076561291b4e4b0d72de5;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfcb147860b188ae656b12de122ca1cfeb8157191126a491507126c5c955cd1ec0c94267ac5e04f0d7;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6323764e46ab7aeb7c5e8d7763a93989b5c12fde76522f786a31a096465e7722e123714b751becaf3;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h95b6caa2c0202b50da6d767dfee8ac4916b2d328bd3c5df21af0172bd22d633295223df17295823e8;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha8361f1035e3e5ec0fa7174044a82d1ae61e04d3bcb2b2159872c2447f830a57fd50a329abc1a69f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8e0dea23c0024a4beb06a5f1b430ec666e3584ca49db872a04e4de09158a7944983f180250f5e4169;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h480c52963bdb6e48941f195785d81e21522c26945bb4e1ce6e1e56aa142250ef3db62c76abf504328;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5772c1c21cd7b59f5df83865b156cc12debb17d5b32b081f453fade88d2efd8ca7597706e1f7f05c5;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h365e81706a37de28187408c9e7acc25aac4a6c79d47a5b50b25b4564536593dbdc1f80f97752de502;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3a29416a53519dc700a430916bf699d4c3a6383a13c279da0fee631b0d6086be492941de9b9697df8;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h60bc39cd9204f5656db31a93869c9ebf10780b4bf2d1ac41eb4685b01c700ba22625abc072d7d0048;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h914d765a7253b67ffdf247022ec9c97a3b79b09e55e0970cce2d530c441932b533c887fbc47b91708;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h45e402467ac924f94fad6ce2d47562d18b758ac3928fad36ce411c59cf8ad5e8efc5a99a462a91646;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1b726fc3bda79cffdc6d3c19f9f6b095733b183645c5ecf15edb6e04884bbaed478ffcad7ec2c94d4;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf9334b878fbf95ab51bfb25f31bffb5359bb7e0f28f0f136003b76de316786dae34d4ad5bdd1547a1;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h88f0f5216c0e9a859bd3074b95ad7011dd21444a560c280d2481b9fd0abc45d0a3997ab8fd850daa3;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd3dbfd3902249b5f3f603ace3361042b897dc76b132f833fc3033f0df82177912e2ec34a25f985fe0;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha74dbdcbbb4debde0f97abcce412797e3d17d4f40f3115b3c71addee163ac6d9ae52287cbf16ca4d4;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h56b82afd8f2d73a854ef73f1b4a3101e6d276a03ac2af3e56212c5529e9bfe7af31171461a2ea6b93;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb10502f8e8d5770246ddaa1b5f80ae6c4c9887ddd46aca75286b6673953c7fd512b6470c392cc1789;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hef8c6a2f0036a16dd48772b445e1560fd5746f0957bd936754684920d2b4bd21029b5f1c8428ea47c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbc4958c15ee797b230a379d66efeaa63ac0295025435782f574456ab6cd9455b2547d995daafed376;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h498f77169b03ad7f11ba18458878dff06295522122ae6f4e2032b01726dc49327ae037bc90d3502f1;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'had8ebd36939da4ea7d85848128ba97644cb102bb6db0c1ceb0d79cbad8725162b12d4a074a9da1b3f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb9078ba90cdb685e29a09bedd518917161f6b1758f95f5d00cc4fb401fd258860048a2bb2a2e252e4;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h81e318ded8887e729ff18da4730a61a9d1f4be4ad2eb8b8664bc689409830848b89ffc7e7aaa2906f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h10f4c0b3e0440bfbfdd130ce2e53520ab7707a06d9618d6abe2be1879e3027456105beff229b65342;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4f07793c8b8394d6306bdcf2d479bd3412be7ab29c49ea80835163e7846f0a20da6d3b7d86f87d005;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc47fb88b7370a37045b25544f2aa47cc2627d03e35c368c9520be1b7a693ba03f11503df9121e5b3c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcc92b397fb88981cb15d050f4fae881f496f8a650e21be5f76c7e1cc9cb5938437214585db9f7ead6;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc6caf28e444a6579f7a87a3f8b157f42d71e7518119063454f7844fdbda2c086eddb88d126f483699;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7fd748d75def3fe0e97436aaddbaa871fbcdd4513b34c4f61808fcffbe77d09e67ebbc747408422c8;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd69006f051ce489da42c208797c83ce3b637a528c925e8c1e319c334a258145f1066745c15a926da9;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h40313c9b85343196e4ce69d1e600fb315513fcb3539e203f9d0c6b2ddd0b6500c5e4da3be5ea26b8a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hece3762eb966864b69c7f2a7ca9fec4ed828c3714159841d8dd4c2aacfa2f641a2b36f4017bb8ae12;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5ed23b30ba6c8abc922b645b25cb79e7487fdce27ed659f3daf14f0b5a19b9491a63af239f7c44d84;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h404ea468d3ea6d3827efbd3c08d7ec2e0fb8d44c459cf6de9d5400239835a91275d76a28da97dadc8;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3fc302a5a7a6d52ad40616d59130eaa647d5aa60c18a061d49e0a2b7839cb1fe221ec89c6b9874f15;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1922b074d78ccb3af23d70101f0110ce2a267da66346f1a95100e698fb041626e582dfc37f7db6362;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h86726f12cbbbaaf1e4acfd9d4f1bf84ccfc531847ce7add7aac633a3fedf142249ba550f1aa6eea3a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2b6e15d0f18195fd3b984c531396a2c6bfb55cfa0ec952634633f6efa7626a5f50b70fcdd3fceeb2f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h536e8d52a8a78389b0df26ab4f7f1e9939b82ca4db22f0349b78ff8c01ed7a978766b7a25ae27dbb4;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h76553cf210f74f5dbfd22c20ce41cd7490c08690b98fad043967305bdeea98b457b2b9e5a73b2013f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9749805c8ce89b59d2849142ebc2c52356c0062c3421c31eacf39ad22c2705e00e000090e150da032;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hff75d39f7c2adbdbc16c4f2402e5aeb9c8d5a2b72fe91674e448420c4835333499c09a5571a6d8fb1;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h436f29867f86bc75ef1e70282cd5d264813e593625a2e5ac7db4910f13842acf8f955f5d846fdaac4;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h70c1868dded652db68752ecfc360893262fb76561857c41ce6bf0ef99cd9ddd5acc029123946903a3;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5bee4098e86821d112f72be236c21278735b4695d3a0fa6f8da1176cd4afd494822164cafe89c4f6c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'heeff47448d2e80693fc49797b4103ce4114056735d0f78c4753ba747197521df4861e38296785436a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hed20793da67fe817feab134b2bc8a2e7c8d630b962370298fb22045cd52cd2d409ec99e5c41c586a4;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd0b34a3485517d71d5d1951ef57e4759ed9457e8fcf449a66d2e9d5da91269303306b57bade5795ec;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1d3476f4b945b125bda14144ebbec59e4773169d53940b6796256bd331a533ee8c7fe2e487f4f783e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'habcce2a5c905c5310228a84f2ee7cf0378206ce673e81146e339141df8a4953bf60779c4f92e7ee70;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb7f6427a1cb8e669db227e31d79a2a104083ef2ce4ebde3453458b9a8ebb76a0b013d5ece25954ff4;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h601cb803aed4657a5325ad32279b42eeb5d070bb2255c4393c800b1c58094cd19ed9eceb114cbbcaa;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9173b4e8dbfbbaf3e779e694820a3858e337c65b8f06635ef827dc60ea08c9b6271b83c69a4140b5f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbcbf9a21244f4644cc565595eb7ffb390c7e2ba9632fdc0ca5d371085958c5e3a9cd4273b9e31f380;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h242b293e0977fb1669310ed126672cea5e554d43bfb7b8ba7aa77fe11194f9077577da69863db68cd;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h917a935f612c139f038b31eb261488a6169fb7d0688185c01ad7209f1ee6c4e7fb012353cd9b6fd79;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h13c7a2f9af1a38da12e6da8e55a8c5cba04d30014359d3d6224fe9b0faa2a394a85bd5dba0f2fadff;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9ba0b42494c663905b004d83de68799b0aa82990e97639c8734a40b84e9d5fd2902170105695894d2;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc5bbb263bc3c8a82e4569f74f7a0601155cf0ed2e36405dc0542bf1ba2dbef3a1c0ae3f1f5ab2457f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbc2bf49e4599369bb5ba1e81e5efed28184495e941837ab70d496003dbadbe67624c232d619e069c0;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h931465037f52aa24e3e917bbe3f57f2173e67c65c8d40ad4aab691b8d92dfaf293ff923584f4f3c4;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3b86236ac4577fd147c1e90ed921d5ba98c0bbcfe947a0d3ca7514dbbbbe437d01512fa7310bd9ea9;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h55ffde6763ecd6531501252259970b787b8f77a7e277654170bb7076c301cece091a6dcf56d956206;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2d29472f64593c59d659e027e3c224ebd3c56792b518d79930e7f0bedbe149704d89e65e485b4b7b9;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h164b5a5359ee4b59a291c78a3baaefb4011264d5610d13d9bc3fffabe9b7f6afd22912d9c6f037d46;
        #1
        $finish();
    end
endmodule
