module testbench();
    reg [17:0] src0;
    reg [17:0] src1;
    reg [17:0] src2;
    reg [17:0] src3;
    reg [17:0] src4;
    reg [17:0] src5;
    reg [17:0] src6;
    reg [17:0] src7;
    reg [17:0] src8;
    reg [17:0] src9;
    reg [17:0] src10;
    reg [17:0] src11;
    reg [17:0] src12;
    reg [17:0] src13;
    reg [17:0] src14;
    reg [17:0] src15;
    reg [17:0] src16;
    reg [17:0] src17;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [22:0] srcsum;
    wire [22:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13] + src0[14] + src0[15] + src0[16] + src0[17])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13] + src1[14] + src1[15] + src1[16] + src1[17])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13] + src2[14] + src2[15] + src2[16] + src2[17])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13] + src3[14] + src3[15] + src3[16] + src3[17])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13] + src4[14] + src4[15] + src4[16] + src4[17])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13] + src5[14] + src5[15] + src5[16] + src5[17])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13] + src6[14] + src6[15] + src6[16] + src6[17])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13] + src7[14] + src7[15] + src7[16] + src7[17])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13] + src8[14] + src8[15] + src8[16] + src8[17])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13] + src9[14] + src9[15] + src9[16] + src9[17])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13] + src10[14] + src10[15] + src10[16] + src10[17])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13] + src11[14] + src11[15] + src11[16] + src11[17])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12] + src12[13] + src12[14] + src12[15] + src12[16] + src12[17])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13] + src13[14] + src13[15] + src13[16] + src13[17])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14] + src14[15] + src14[16] + src14[17])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15] + src15[16] + src15[17])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16] + src16[17])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17])<<17);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h0;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1b09f18a53ac605371051c2dbb3d5e5317c7cf75e8ab85a8b8173bdbeab2520ad9bc5390fd81b3ac1;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h838c991bff243175fd1f268672a5cdafac32c44982d3962d98258c9964ef662fd790babdd148497a8;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf91adea4ca9a5b5a6161535ae1f81d6535ec6df1dcceee73300ec89ac2c42448fd77bca7516069153;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1748b0926bb3b61590e2803dd38806f743720e8a08191b015a30b39c6ce0942cbf067b62d7e888868;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h448c350f3127a9c3f480626feee81c6097580a4d412bd01d9f3493b0de8adcaef4cc767817933d574;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1431ad844b17df4648a176f76851c54d63774b85981bb30644295ac46fc2b97ac0512150dddc2ba65;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h21101accba0f901e4954196d6ec495474cacfb5fa68d99b15f6aff7e08cb7d3c12fffff904dc3fc71;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hab72315660d2a44a506365281f49d23c01ecdc7a4da7c6d8e0603ed717b8bf8e5ba6be304d1716449;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1a8b667740be128b2b1f7e853c10029577991b960d600f5a458dbfc799ba46a28e1e6bbc112a6941;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h242ae39a864b836779c1108447a72fa374143338aac71d024ed00e03608d29e4735e882d3b9f43540;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc2fa9da2a58c41bed5dcee4f8aeb5dcaa77e9b1b0a94d9c3b08c83accaf233c5abb79bcfc7d669ce;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha7155cb40e9da3a593d1d96f08370d3439920bbfeeca8863e5216f99300776d84b4b893325e1253e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha0ad9b3a9e3b6c9885fdbbe143ab89d26ed0c33a2f7d66cbb0952611303e610a079af3a76488c11f3;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf3661bda5af7e73d881db1c129dd7102f62129dabec7359c4eca38a5871fdb9c55d7e1fa975ccd2cd;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he7293857d7ae61d1529675b43089d13f010436bc9fa34d81e5c000e9f43587fd3fa371fca9bccb10f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb9a2b482321398375180f5f7c10a8050a5d22a9221e626f8247b97fc9ccd7cb98e1e9e5d456b08b1b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h48e2a17a58fbf7ef19b8878e660c7a277f3e4115de1755563279d6b22aae1afea594e541b2e45abd;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he08bc5c5b5a5cdcfb7893f06a35cf68fe292f6c23478ef86655e34d5fc85e4158d43aed0f53e2cd52;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3a01f73c9f6fd0b8fa626f65a73bfa412953d93bdea10298296f12839f3fbfe176bd20b35a3a72fd0;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he46c1cc347e4ce65e9d7e80c953141e387d4d59762b386aac41b5c7fa6d12446b19df099e55d09032;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7dd54c215471f06fc59c2589700e172cad2687489b88575519d3a59db36d94c97a8af0951c566be38;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he0b86b3dbb6aa52dea9dd10573b5bd64ce9f94378cd3eb354fff50567cff3373f9578ff12dcb70a2f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hecd5361e41d6a36dc4fb2a8b36e4df00e8e092c2848e3a4d259f31621d9cab87e597ad1a7a4cd0c79;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc60207ee18521e0d29d6b93670a5eeab394f0d588d86ffb14921248ffa495866899300e383b388c66;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h57467e4b29d4d48f2729dd0fc2d0eed4666afb50514da100724097c607ec4c9d111d8da2d927d2483;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he94b07b3e66712dddf4425394362113edf5ce6c9e3e579f18ba9a5a659ae5e56c68824fbcc1d8397f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7c80724b238e4b0d98a3dc2b22ffd045a992160b98e0bef2297760fd409e6f94d1a86ecd981e744eb;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h152225c73e339c1f4f9f9b16d454d9e420b6fd16d9fcdde4adb8ea09126159934ba4b21e7cab9bc42;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd010f52e92583499caae62949c21a2d86587bad828378fbade7078dac3b721e9f2b6f49e3093a0133;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h23e7915ee7ac53e698873d064f3edd80a66f900076b5a4cefd0f4088e0b6b095e14ee208053195093;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbb9f1a431a902282eb4518b1c1837e11401a2115fd1c06e3ab0890fcff59f066ad8e105ed3956489e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h831a11c1fdbecd66bce5d4ba082bc99a157244aff5ac9bfea7144375f20fc2157365e6b934c1912a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h443a03d77ea59bb4f7e3fb398a0c7df5c6362f73b856b8c09310a7d40e3b86489f197a9f2415bbf0f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1a36031b6b9ec3c2d203cdb21f0722d16882c39332c59409370b123834e6e84d06ddc38b64c9359d0;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf81397a99409368276971ff7f0909a6489e89c1697ffd56b2b9edeca571334f98d2484c95b8fa0059;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h36a281c6ded083e17e226aa980fbcb1f9d6b60f576cc66b6046ac789093ec594370117c339c4468a7;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h57d88b20468e5760abf021947a70aa119fc7f762829a4c6771d083012163264ae90b0447edbd9671e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h192bee42db86f067e336497ca3877606742c41d8dc0dc040a991a63d47c8cacfa04342b0124ca1620;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1ecaad0b5912578886bbde7aca2ee5849dafaac72398d6d1f08dbb087cc2e7474e2c21e2048da8e00;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hded727cade4da9af2e7e4aaa6a22745030991eb0877c4cc34c13d5af915209022ebd9faeeec0796e5;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcbbb1661fd17695c9cfd6d741fab583e3e023a1cb846cd712bf81a874bcd42b94978c5cb65266afa9;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7224843105a9151571c86afb053d6061e8b4a6676c9a45f9c27d80f291ecf54921b92dfa35f6fe6cb;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h158335f18f481685bc8641364af38474b8547811750d3888181d3cfe501812f0e061a679c641153e9;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha3e561b554f890409a96856503e28deaf07add92ac7ba68bde9591173247fe4168b0d333e24f62102;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h80ac3a4726a683083fa7287298af1b8411e877ee09f9ee4f57cbc66017dbe5eae9709e5a103730537;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h59a6e2f7cb0597e0f64e7753c0ac2f1394579215a36294317d010e4a2ff061ed62407df90b8533ff7;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf261a0cc860bf42e1c812db93904d8bc9ee97ce80c6b690cd746f8e7b1246355ebeee87547c664aed;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7fc3d452a5257bc81a39cb1bd93c7421cf842a419f6523857d4069859f6459e9c7d6b983445100dc8;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2e0892d05f2240f3b41d6f60946d5b7571ef1a9b8d32fc6bb1db2ef00fd351f80cd883a67ca4f885c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h336f884367512a72d120af272d5da29219245ea4b78d52085dfa8b7145defb51eb83c85feac05a501;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'heac8fa7c9e07eb365c89fab957bdefeb2b6fb7b91d9dcb0c2d24596337175f553f081b5ce0a84352d;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc01db009a7cb25b415ed1379bdc329c6591b36f5a5d1558088d67ecece6f6d5c1aef5d6a7696e69d5;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbf86f27eda9b3c42829c4b22596ddedf281f7ffdb2bd7da0e7620041dd98c4f67d087815a5d7a4652;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h845ea869029e7896774916755859db7e79c78f21938f19bb8a9cf1140cbab2745a8bfd07121312afe;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha7d56e3c4f59d8f54b3e9d56bfa417d41cf517f180c767fe8bc092b6cc54efab9c49e2b3bc5c47129;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc8171ef5906a3368e6eae0337cc0fc580a566b9ed19b7b8a5c54d0aa856f68a4f88b4ff5e7583504b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc368c7597b5641c4b224496780f0beb8790a40ae8c66d5f3ef626b3c0e32dfebe21c0b17f64d5f999;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbf74c961566c47acadb3443770bc48ae8792f17d0348c330b317eef037c37a7f2fcd2802cedd7609e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbce1f359a57781b107b26cc330dba7933078ce5898e91050cc8da5e975e3ed95d9e590ae992bf1ab0;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h262866426967b42552f0853cb2d8bd1b885deade6d92231cfe2211194defd583948974bbbe3fc7625;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5266ce959e7be0d43645dc319df249196cd522dc157d10e6c0202d6dc9beae9e6cb65874c8cabe11e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc9337b0a0f4f1e48fbfaa8c9065ffd3e331c1ea6ed65fc9cf973ed4690a76e40554f1fa8cbbd0ed9e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he2aaa024570d09e9ba0bbe239c5a766cda0ebf2ac3a19057b1bb93c422dee25f637dc5ad3a427d082;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7c3e928f9dd390c5f449a789ddc5d9a8cef11596e52a03054c8a8a313316822b09c47c2f3c3cae2cc;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hef6940a52475c2fa83167b01583d3ad304f2d8a335a8d31c385ce708251bd443b702649c7f570348;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3a235b1666efd194afe7020a1c87687b46b753ee65348037f61750988014f91d321e2386ee0faa586;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hee61bd971c932ee81cc9741e72d084554d42c761beb2a9f64e74eeca67e6ca116546cc13a7e2b238;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7bd5aea0b8186b962a5208906bd56a74500b0b41efb8cabd457fe22689aa6a60d9d2041f1d21bdc6b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h876ed7206e5e7d73566c38e0f070a1ee6595669c72e68b7b93888863214da71796e6711a9b117e0e2;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9ad50e30b95a197c8bd197bd153b96f3008ff350f58803165b07e4b464988c0d5c8904c5186a4674b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h14d4ca4f862c8034e0f72b085606ce33d835201608d53c9d32f6f11d9a9ed1c6cc1fcf0a5f89e4ee7;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h43560c0bf645d464f3cd0e337139838a649528b34c40d5389e8446707347022523c048c9216b0e804;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2e5687de8f09b1bbd9d022e398b8cfb7832c0bd857515e37793a7fa937885eea0079cdf397cf768e8;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h995071e13cc30f7995a1332abdc9cd5c4c4a197ad7c328cd068e59e465b748868273e954cf06b458e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2f901d67fa2617f41cdedd6c2acf597a70fd5192683567678f7c1dc8ec5664cbdf0a4200d545de9ae;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha8f12796e730418903eae6abc947b176b8fd34b5add140fcc9d28d51a719068bf637ea5277bd7e090;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he74e9247edb4b036cbf165db603e2f5b3beab1b7a3bbdf298d63e07f0b6f34b0ea84b9884b347dff7;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1f1a0ae6b5bfd89e617afbae2cdd282a4dfecf51c889b17ff3db40a968e6e80df5243d21222548b49;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hdea5e423f03d03cf6d3e3a4c5e6d028b23d160fbb0768834d98ac0a33281e80379f75c76322062f14;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb6c0a7bc93c35214ec33e366550ec049b8414eee78619e2e20994127e3a41b9c2625223595c93e2c5;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he0b62a8d7393ff55eb0903c01526e516140a8b011a3d51f9ec8ebff3f8dc63498888b521daa338af3;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb45a646de89d7b8b8e7f1dc2f29c1cbaf348f75ea19a7af1c9421964555d97d4b9d85a78e54eb62e0;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6a9934b22b7713e2001b6728a445c74d8ff3a08bd69d0a5acbdd9bffa77a69e56bde9cc8d89e44a54;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hdb26914092f82f0a8fe80eadcdd4ab81caa0d30161d083112c786bcce650c9e45c659366f53814cf3;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he477a9fb0b0bf8c99b5ab04191aff12a7f5db73b3e8f95d32d44607db5b61c757fb34536fd6d54cd9;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he3c57a09e1630fc3447519b5b248d3806d98ff7011c7c87c531e192849b9cdc49dbf041e677ee667e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1c3de08f7c7a945ea3cdd9521b53849c1d16ffc05581c2301ac5cda6d34d03352b234f44eff99308c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha3cb2d9dba0233ba78222ff13b369a6f8e004e824bcfcedf59860f752f4a3c9f59e27a067d6b701f7;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf8508dc74214a5498ce88e39e1763cb4afb0e4ffc95eabe2a8cc61f865e43ffaf9c422dc316e0d07a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf6ab50ebb5f9aacca0a74acccfe20b27ce3f9dbbe358930c455792c827bb69d75754ffbc205ca7577;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha38e9d3dcf858a6af6ac2ea27cac1597d8c707d696e49f3c22c2bfa65b605932722392b4dfb21c59c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc9c224493185daa20a961e601653b9e227c1fa76f17d10e7f2237b3b93b1995e9d3a22e3c37a4302e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4ad448e424a2d2245c1b4671e8ae1501ee3aab85db5165afe13b4556206f0e8e092865fbeb29a6d7a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfe3bb8f2351851b29c4e7e65b8f4193e6543cbf19e75b0bc246d82e3276db5a34d0f514fad9f6bd3e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h15c5fbbca34fa07a648a9ef5cc9ba34948b0b3d5b838cd763e13ec656678f768527310f150a3ddc14;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5336bf4d8ec17eee81f365e8f0a00261e6739f811113a5aab1ea8f669d0837f2b5ee3464fb799efbf;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h53c7af6efbae3a224177d5efca5ecbe9450e3a58396b94c742488e8f55e8f615aac96260ee0d59f2a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h409dd5e6bcd64cc2727abd4811598341fe481d28976f2d93a31e721a65f815de128237b297ddabcce;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'habd3a8830e80e48310a4b3e73d35cee276d0ca0ae7c67fc364376a3f59ddb10a873dc7c15965d7520;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hadca6d69e0d69be2e8e9c5e6b4699c108ffad3c72456f788a274537cc9175c3bf09784ebbd441d0b4;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he73dd7b29455128aa033be19d254ba809e8391d6a7d705dbad3b735f5be75c16e9594cefbba45c029;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6707d13ddecd12c6f2f25c4391b0a8046f7466f6c358909e655e43855977d83180d5b6dfe29d0581f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb572712b7c45df61c19026d0dcc6f3e2f1142ea483f8242335e98c647e5782d77d2836455456cfb84;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf50add81ee1f0bac964371234b3bed3930c38a18842ffa209532d3dccde8d2c85c0f660e3aab7b0e4;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfe685911b7454d53a48a60812ad9b98ce0474557513ee7545f53d0fec0755c67f97ade3654d0f727b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7c8b63d3b72fb7383f119526a27d35fc2b469c15c4b018064784068bee4054e26f2849596cfa7b27b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h65f06c47e7abe693e350ba78a635ea02405e517457c0b4adccdbb9b06d0b39865717b6e5a44ab4f05;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h38a5bd2920b894f5fcea6ac003ac46d217cf28676858cabbceb7d1cc708d8b00fb5978450e6059c68;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h24f2433c51f5df147f983ea2ba61f8264be46d92932503b964849f060a12f0d51fa640d32d03f7c5e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1d43d70f6ae3e5ffcb0902fabb83782a9a3361b5de85a9e82a5693e4e59f72fbc8923590d4ad21e93;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcc092d5c5bfef69eb2cc7665c50b336cee10f811de12203448fbd15d8fb4725f7596aa7db7fe29824;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2410276f71d1e512d65610da1c1f23a644af46b83d28d713a4ae158cad6d7f33c461b4f5cc9e75480;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8a0f88e12d4135f3573016a40903753b98623ada45bc30df281fff99a77d1a83a43ad6f6b0f2619e0;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hff8f8841a6baf5b317d018d7a266c1a5aa3d0297503768f010b66840368373867e50936e0c8e63f09;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h60a7f19e861c17104ca2dc3fb322d7d0aafabfaebe001cec55e4dd5823f9af18117ea8486c11274e1;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8ee8c6fe626353fa36732dcb94ce9cdf6897499945b0f1cf6b825d1afba98f54795579e8842680047;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h26f7758babe2e32b1ef3ceb4d5bc34ee5dbdb848e842d2e78419ae7310756d5c1ba4d0e9aa8cf24d7;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8f87f4f33995d881fb4c1ab1232e0d93a8f8a86e65f4ea0556e534f18af885e805e5195b33c3d0b34;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h57d9703528d4dd0303ef0b25065b2e0ec6cee65597179c421ff1da727d04b59c5300cf1cae90fcdb8;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h23c1ee2f2fe164f25c9d2c84b8e7091a8194ec7d82d7bd479619d4fb70c1bf398348d8df3d321d1e5;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9e9205896f2755a2d9ec9db212187a246193aa19583cd26ff7fecda5441e0d63c56a76bc45738ceea;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbc71352e2bec2ec5c6bc8ca5414568e14e0e72b83f5d0458c056012841ac6961f09ce6a303d0f8fdf;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc4d78109a118d538e8291ad33f1a04fdf1691a3c6f347694f40b2462bd87b2126c78c1944d7489fe9;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h88148ae928452531443411244779b6eef55269924a45f14631800160a7f759ccf04c04d2a3701f501;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he0d486e0fda3bbe062785e89b1c4d33f39717d4a792ca1f5123c22c98fe7cc612d407a8f75c2ade2c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hdb61710a30466d48fef849f6c91f106142c6754c9d80c06e06d4eafbf28f5b2030de839af9275dd7b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he3afc5fe14ddd090ebdadeae99e4bf07be3f237aed6fcb4f1c38836b84ec0d494454249fa3b5d6d9;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2dd34dbfb4540640c07fd45eec76b661d7a4cb2c40522079a44be6d7039eedf29890dcf063202a1e2;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hade3850687dfdf824bda0b846f0e11e575466416324869bde0856edd0761c70b5ba2554200db74265;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb9c144d4a9456f48ce251a4bb1acd90057d98b4035f02b3cd5db41510d143cdce3ec0185b4e0f160a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h63e73e8e8901deeca8e81d778c67d9627b080abb00d7d7c5346cada0fd8f52441d7d0ec4449809461;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8e95cbba3355878fa27ee74035ca3cfb8ee76877c3633e879a2c390c5b53f4cf21f2dd31cc96d9337;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7dcd4f595f6759aad84ba5e2b1f6d1cc30a4495cbeb2f3aba2192f80cb1357c9631005b37913a6231;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcb96403da307a2b9803915b4be3d04e031b7cdbf85cb71153eb8820e696f6843d1bcc210d818a925;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h99929996e18d505bb38e586df9e873f96a75cbc579ded376dc008f0a50f87539ca3a23ef723d8664a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4bd94b85279f627f5032039990031824ece1c99e3e90be0433584c2b37a5a4f2c7120a43b570a103a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1c9bf40b9d3d0cd4c76546581c97fc4142c4541375c23452244a882ee58c82b6965c8f9e4e0c618f5;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h96e9a17ce8ea5d8a8b7ad1c3af9793a1453fe6913797da5aef8fc2d6685b8a6d1f9315bf2eac177d0;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha786d54e1df95bf748c0d1cbf388c6a0590a0f015cba2e7e16b532160f581ff72167a38f73ea715e3;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7bf7c86fec08f874319d371921cf223c108346991c3f2f6e12ce54e5ec6c548079848d4daaa34a1b3;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hec776316e86a483448b0e81cb60c912bd9ce16a6e1d099258f2dfb126b0d772e2b999267a800b3b32;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3613b1896f7555c1397e496f7d76b8a44275f534c9d6c6df9fce5af7f5a3e17fac70d9149ec6575e7;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hacdb346b925e8ea204342785d7a617fbc7f43218d77f2cd41dbb56f5f5a440cce32c7321dcfb17046;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9f911190a51e208582b5d80a90122e76b4d5538dbf106801b689ebd6f0c1c30e7efefa9708a1b2bdb;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hafdfc8f5d1e2cd85241b49e759e567d5d4912fcc3b5cbca72e7aefb1e8fd8cfec591e8b23acc6b1b2;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcf434bd6d2dc1e95fb07bce690317b6ab4008d2a94b9551cc4cc2840520b9793b6ff81b3e019e2f67;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h382dbcb4ff21634b2754173936a7ebe9903a472be70c4e1d088dd3d08fae08eab0865835fa7e45a0b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h42fe423e98372666e7ece20a43a7013670435f98d5e34472f318593c7440f8c6625d319087da6c613;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf756a8906c2fdf192b36020cdc28cac45743ea2bb3504dcf50e249ef23e2212b6f52e81637080f7cd;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he6d4d4bc4ee226295439f63b035b0264a9c7c85390ddebcf3c36d811d508e9cd1009726a3db5ce05d;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h35c62738cfab2a0fffa9ad4fb3d59742654c069aa236369efc2bad2d45dd71c51a942c9df864979ed;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h935927c542185db88821ae5271fee106f4d15a480e9c28eb5e50b9bb9d0f5fa1abe91e7d1cccbc08b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'had38c5441bfb75ecf18e878c3f3ce87e6ca14e390e6ba041b9b3c7f4e7ef1e9e0e1b072173471cf49;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbd3b0bbbfe6c27d3130a054225205c422bc6bd7d157b56cddb441dfcd93656bcef1d883b00b359d5a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hdff569ddc201a504022ed53fc2802f767f892e9d857c61ae220d7c4f282bb4d07de6b76b191523753;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcd988f4f38a4929d856a7be89e2f82a7247008793ee8fc55c85161a1a6c9882426bdfccc63230b5c1;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'heef411c726e285d51291f3c493e0543c3999474a87c422098468ed2a9b2170de1b23bca24ba3ebf69;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha2173cbdfcde80c4ec8680aa2a5f4633258afd98634b8d35e782e6f4b9e91a475060c40514158fb6d;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hedc1db857dce82ade96ac601b3c79f7ec6d29e0c45672445b006db81ba27d93f64d71901d33ccd08c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h18207256d1c4fd58e1a2c32dd074b6672116707160e78556e526a309b2f1e157568c4d09c5f5d74ea;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'heac84d422a6b16c7aa4c63e6f08c0ec9a5e29b62ec2274a6f2143798d1eb024712780e4e456924050;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc337061ae1faf15189b13d0ac472068b9ca9c2847a753b070e528e735f0d52e5703d0e8c888bad65a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h88890ceaec1da558f7858b305c6cae3acd39bff140b0fff27348c4a798c0a7bf00f71a39b5b8aba09;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf15852017eb1f950970dc5087403426f3f5fb5c032d3f905bb917437ce45191ee9ff8e1fcefd7ff00;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h46ed08b56572e5826177b791467efcdbfb9bb343ddcbb402ca34f01ef17f3cb34398032e69d507729;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1db2a780423aaf15ad9a8761287c04573dd8af8abc7f77f333d81e3e1b3cc9d7ad554b72e1291b2ff;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf404ce6ebc8b022420c89c4fcdca49e099f7f71605b6d7ad64b14a23a9c894f42b429550c4e5f4fc1;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbf8c6d65175ba65d4c218a5676f6bf30bde79b0d4dc44efd6ad171e15f6e224d91cba6ee78cc46652;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h93dc23d96a07a4142d7c16bddde4e66352cf7ec281af09d99eb2b3aa1bc3d218d48143a3fe4437027;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf29313c292e464a9e7afabdffe97b483ba27b051ff817608b69ad10103c6fdb827beea8443eab4f24;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h171d8462220db204622fa2f5d8167413fa5f5c91c06752f3ba5ae10199994822a91fae9d337fa3afc;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7f4e6650c41e1354e0ecb2106984ea716c09d5992b7dda21489777746eb7369c177b3a55e9258642e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb30d7bf55d99f291f8eb1878ccfceca00cda883512a3c60f3c7836bbefe1cbd84b981e617514e57b2;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hebe3def379fa56a242557c8d0e8fdddb434e950407125a1b5cf316c3a1e283e4d170bc71228d6fbe4;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf5a59f68e42b5d2f6b79bdc8a264e22d6050f8c53594b256e6d4905695c8223927c1354f6c07a3ce9;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h96cc20c6df300ca5b4657f882158e1c50afad7ce041c8704bd0ad96c57faf71163722ae85725d4717;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'habeead044e630b928ae18399f71df07a231505b2c1c256ee0c98e7221ad330f4cc60b39e0a374f841;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'had9e253b462efa3b77c13ab9bdc6ffa957c9b67469e38aa163eecb255ebd1db696e2350ae5fc1000c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7935b5c062c46fed429127d1400a861460b79ebee17676ff33f19e0602f9089c0b6dd7267f5a9ff15;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf9ffc5f84c1fbd1ab2534f99f35b10ee2f4e6f07c282345ff758be4ebc8446c1b796082cca5386fe9;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5ff799745006abf44357c7cefcb890171f9daa72f570111726982b9f0fe56cd90843277acc493ec4e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h47b2d6750cb3d969e7715efcdb81e24e62c9c98d777d6d8bef7e7b2fee0e1a97e0e14ff9a97627e23;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7419369e8ff55814fe478e11e1ab07028478327f9ad7c9bf29c6575d63912dde706d62c8565388186;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfc2ed2d9015a4bd4a22f2ac0828b8c40a6465b812d3ecfa84168698f6525d74c5dfec0aed6df184ac;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd68d02bd3c50f7dcec7afcafd4657a0d934e1c00c502662abe6bc006954b404a024801c87121bf085;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc19b6260dd47380579a2b6ad5473b8e2ba52dfccc2337835eb8b498a652f656bfa56864890d752990;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2a19fd930921f49a562d5cc91e2c0bba11102d3aaa3b5730fceffbd1b257206e7168bceb9878852df;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'habd93585808ad0a414cadea9204b887b9079ad0ad505861adb4a2ab50d9e750abb9b0080b4ad3968b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha914644ff9267ce30580f442c11dd18ff84651d4b69d6044df2c75de88a66f3953ef6b9e9ae439839;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd9d3ab9b2b73dd457a8bafa07fe79dd3656caf50de592bbe2be21b6f7116a9513d8c20dd3fdd5d26f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbbed43391d3dee601e1c1c705b169e9118abfa20fc7d9ffec37c4e525691f61bbdeb7edf1c933985b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h24277d33d53cc2d8ab142d7776e2268470152e3f4b5021854b8cd90796d52bd85d34f37610f3dd2af;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he9eb47a4b6cf790e3fd108ae7070bd7a044732d1a368131047aef4afa58c10efd258840e1854ba19a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3c9a5908c951d813afe25a220ea4ae2a41c0b23914995c42b635431ff4ef11eda17b9564e4a21fe5f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h569e36d7e6eb6e79ecbeda01ddbc35d1e15a05ba5df2a7cbef7c5e25bbc9afab1bc25b8fc6da59a82;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf566c3b8cda3750e5f5b4bafac0e2eb435a315e95046b1d22d7452877ca6167ebc2ecedff205dcc44;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbad9f86cdb9b70287cb6b1b415fda3832aa64670aaee4058def1a7aa6b6cf29fa10f97289a52c67d1;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h811ba816f27bce740a8cc282ea57695b27fbcb96586d20f775b97a94cf5fe7e48bfa41295e7b44ed7;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4c6e657aaacb107591709c0937db233cab4fe218ba9929c2b91831b5e870a8c1b650515942ad49afe;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hea4fec08ef2a2724ed3baeae05ab2cee7bb1335cad6b5de8b1091e7f40f8a0a67905ea7aa97f6dcdd;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hafd7d9fbe63303e4d3049e7251eb782aed1225e34a4535f200b2bdd2746540c1f78e6ab3425961218;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8d563ef1dccc758806419e96042f988eb2d18d2c65a2cfea4792c8d44049e2a56b71fbeaef9b0fee5;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbd864a530ed841efcb1dd62115bed869040d711721e5ca52becdc276974200b3247ccfd373a8af53;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h49d8aa66f3d40d8ba6d0487ca23732a0459bf786f5a0b0a5bb3d4a2b18c6f8ba9dbff39cb5f185bfc;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8a00a82c8a22b648d028cc0e666a74a0ebb153e039d62f4e3acb49bbc178c5581ba2e5fb8ce4ad9ab;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hddca2a8e7649a8a4e75787b9e585f2cbe18f8ea0ff4d0730967d7b941e43d366590d737f4986f6822;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf1a28aacfa027b871aecb07838ad11b448dc277f1e547db327124be39e8b049a9389a7180151d5f70;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hdd0e428b1dd7e7b8572faf07d16393347cde03a67d721b8e3f06853a9103af255914cb9c1ca17f356;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf787a53e345bb86ba32cd74b937eb96e10b64132b23d117bd8dfa591ce33b7b622da087e03977604a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2f186ef152bc40726e5ba9f921b02b9c34e6e7d8876c0c36c1248e2bfab72277ea3828410d0a7dca3;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h509d71fc117414047e283114780d587f1f631ce25cdff9bca133a000c1c8271aff0d507bad3a5c202;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h569a3ecaed28bb871ff36d90ef258303671bcb082a2bd00f0418a07dc4e71d6e6e6f7cfed7077b846;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'haacd6bd7cc0a90f65e4933af080456cbb61f1a47e0c6f106deb6c578d55836c96372ef8798ee07730;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3459c329781f1245a6369991e5401597878b264b06229887be5ece8e5099af508a747c6b7795b099f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4d6e3d073bada2cc235fa9483dd9b8c6a8ce2e5dfab6858f34b00cf528615cf642cf4dccef9d83279;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbf0a386d5d786a7498dda3728bc622ce9627223aeb394fe7b731cb63eccf7762d5e7ca3b3edfb30a4;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4e1240a46bbd625fb337b3d30e3e0ebd8a6d3bd6fe8dbe4dc685ff67dca2ded6f2755e85215dafd78;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbab78aeba5741d482a2cb38e3b6439c4cd5246018dc77513d90044d74f81a3edb96d868ce72a608c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h19c6926a899119d28696a52dd3f8e9792b914d94416f25d2cc5ab38087cc34f1cfcdd0606c927c803;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc6c808deeef3b974fed4e2da5e3475c06e3d25d693eb7f3afeee3387ed09e3237799ec9e66094ce6b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3bbd1bb7100b778668e6515b00a5d8094f59bfcf916ae89846d47073fb817d5bf91f3a06f7366b863;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hafec10f0a897034f0f0c8ce235c4cf81b3f3da21c064fbda97f0e2499093e9d6f9778f25dc5d3a5c1;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h13507ba258662df39baeec48ab57397205ef46666fd94169a98fc3e6968b17612c97ec05d30172d68;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h235664fca46e9185004e34abc2f9b9f60d462708e180b68cde84f25af478993ee29ef3fee744f60d7;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h420ca194c093a8ab19c93708f42869287b6eb6f0adf6e4d69ec4d6867f8c80223d2fcc641fe9d5e05;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4c657e6b94264d264b5bd26176f854fd98f9e9a0d1544e171a492097c618d8e4415c59fb231582a6d;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h254f1b0bffec040a835c1d219db4f4d0c24714976bfa98f714592ee14aee10c9dbad9d7f7f83c1b52;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hdd4b26c58f19f0414a2ef886d5d45cf0b46a9ad125a97a19645f84ea1d2a10af05daf1d3bcd1b8e5f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3680e3318188947196c0e5578fdeb86a491635c6c968a4ef982d91db08fda2ba5a385dce5fae7c82c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9424a59cb5a35feac189144784d6b9eb37f980f5c60b1c56658f8fae4bbb0067d63717ee4b11696f4;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'haca08d08509c550506f77223bfae5408ab33ffbf772f3a124bd5fdb4d6c4c302fc42b1c9550fc2a19;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9cc50a7af7ee933bcf39d00f31a7575be5e121eb5cd436304f7b507d103ba093939b01dbe36e93e5f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h70970109bbddac334130e4d9702d82e2182620ac3d83127b4dac4026c1fb3d99f04fb9c406f2a4473;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hdb4bc30c30c0690e5902c651dfd6737b6cdbfab2faedf5666070a5c85368507a84e66eeb6472bb7b6;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h752e4e86df93588ba876664a63265e751e1e3daa3715e229d05e503a5257527a381bdb9074acb13ef;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hed73e76d72e8da23b4c2a9732f3092e0408b02518fa5a3d9a72cb01c509b60b15e01865480514c078;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6ed1d37c4fd210778c359fd726107f8fd3ef46150632d7667d95dea5e3cc2e1fb1dbcc8147b59615a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h78de14aa45016093404be4b750c1ca1be07a5d483273513ae92b26d8a04b900234f6a023857ff96be;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he1792d9265478b1192049596d2be5b9f81a94e43e42d06fcb6df1dd4d465b4f8bc565973b6103da1;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h88e0ee57299f9c2f4b1bba95a6270cea7ae8c79067e56350db83adcf02e77ce477ba512a407ef400d;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he3a001c96b070962398947f215a5894b26d11207f0b35c36b4069f5bd248633015d5168505b7e67a0;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2cc07a18d33f6947b67c770d67d69f7ed8287dd0c03d95537953c7f083c648a332475445a26fa15c9;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'heb08e07c34ce8aedbd97b0b56dadbbef0e1959d5b27ef764c158c06607d99ee984caf17ca835ec17c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h20a70414f3f810ed10ed1cb2addb3a816273525c792cf566fe838b7f852f408eb2ae41bc660539c78;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h88d95f1118f77ee208e2fbe9da1cdb5b6d33659c02d02ed9ce80c305ea65f4b88a68515f3de55cb0;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4a582d6ceecf348c64f6b6f2cb560e509fb76919c78b9e6496f64ba62a4704ba21185eddc1a1ad88b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h11e6e78b32e7cd391701e661a1b3e1fbbf2dea648a8c81b01058fffcc23f658c81ff8866f20ef9768;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6cf074c5747b1385e8a3e23de3e6bcbdb58a494def10dcaa2f24071235a616e378959875a517cea8a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h69813f5d0ca11dd2e490c8351e2385a85ec6369506ab8ae7b9c7b59eef3513da961e4d39b6d891a19;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h442f5ff8aab8ef04d321d201d565ab8481aa334b5339b1813e2fc8cf7152f4c625f6d3eb86c9ab0b9;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h108f5ed30ac5d80fa78d200cf7604dd5f9f8f1af50d8a01f50e6b6969758fd2deb6dd8b33eb85fbc5;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hff491e0929b460b366e26f7f271b20ae8eb4f8a5bfde201bab77ee49f527fcb04865519142d1ea2ca;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hba9c3b5b0cbdeda2d41432f08b9ffb13cef07976495662d1a2c8195cab5659c1b49849510491ced54;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha533f5da8b5ae12d6579090c2fe9422bd634c3cd89312489d0613b7c0d420a695535752bfb29ec3a0;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf91e865c14b3b18c5988302d477aa475980d08a025bdfe73374c7896c65e71a3987f3dba322b61a9e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hce6baa191a1ee04f8395da19d70813bf39d2d9fadbf85279743362e862f302bb21889c49ffe211362;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb023702a1eab73ca1e6eac4fe32f5ab0a08650b37abb8fbba1026e2c6f5d2c360f9eb5c7f13cfa350;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8458c51c3a67d9910d3ca7a96ee7c787a32f36622ea9707ea5ea7221f142a3d209304a1b8bfac3bc6;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7abba34f5fb5ce022d3d5be98fc31af2fc3b73f88afe3eae21dd76695f9835b32f5f01699d343448e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcfdc68263e113596cdc0a80a50f33b2554d8dee2104037c9c66f72287bfbfc17094de5faa7eef4f59;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbe1b8242a084737aa8239577f446422954d591bc43213bd3861d799714d9b12e7037828e2bf27eb2c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h941099328a3248a24c1ed5f7c60e6374638bb2cc9f14af11e335db6cfba0ffcd676ffd40da831190e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf986b33b90940d840c839707f2e2867c53fb236bd437cd4930d1243c021a434630eca754c09d59fab;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h165917462db3b2b03a57d69ad564d79c904a0e0d09ed4c2de8b5968d0934e571198d59d14ace985cc;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6544444f107bfa935284cb396589dce2c6acc07daf2b48341228ce93e6a3fde45285402ddd9767e23;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha218b4fb9a931f38c8139072b95adaefdaa16d005d209c30bb402f94753e1fa0f029c437b0ac7bc06;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'haea08f019f0ae2e5f078817a19004080dbcc1e4c72aef63691365f188f2181342156c938b073097ec;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb3b6399f5371e3c6d9cdb78f43209f76d4c770596e0225cdcc7fc285f2efff11433cfb7e8347069b9;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5cdbb7d597feb95233a508dd893ccee9274f85ba2bb7d570246e27946a9f15fe4230703443b6e1a86;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h20a122f6584e5ed439a54e140d38b07b8b23ad1a5d6a0fac59c7124db9592882c3c801756d482e183;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h645f87d4438133868a096c9be022dca439f4cf32a6750d840b2a16bc23fcf339a376f12636180e30d;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h26dfdc4039272fe38cf9fd3cfdff6f82ff582b0d4123da8b60644109de597a3ef572b7a0138b89fa;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h68e58cf51bda2ec390ed00146ef5031dd4cac65d39bc495342569a805fb768fc2d91ebccccde5e627;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd5f3a53c418aed0e9007b261244308730f9b30b5ae94fed5ec955cc678db1fb063dd046090f72d964;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5893a78a6ca5f2ce18d8ab94806b5a089e0ec9296b3176e86fd80870560dd3bdf6786b00449524e46;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h862f3ffda3085d8c06271e29511af4cc37065d219bd7e04da82d2efbf06708fb42834470f2a3e8828;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h404b3acd3ebc6f83fd288cf47bbb5793618b5124248efd56797dc8bf2728b7637ab13d33e2de20855;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he8e5a31a92339f85745b892a6d3995c81d014d6b7367073a1e0b3b2166fc0f729f8e5430614720a0;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha88711c3bcf0136d4f678ce13b433d63ba393e091d2cc02ce4c7d9c7a3cd2eab609e2c48dc92f32e1;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h82b073171a0be8c9fc849250129e64962b07d9e877f7028586c2fe7a69a3b529ccdc1b6b3f8dbb6ad;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha8ed2f90ba07d98548629aa8e74e7eb18a64cb94fe19f4e6a86f4057a28080c4e3d726ecd1bf001b2;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha0a2b3a0a0aee00a58998299be2b72be5109785ca05bf7faffdcd50ceff8a8b0fc5736f8d258e853c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3aefacdb4baccbd451c28090ccf7975c7deaeb19369935a9a95d67f6914fe7968b25d95f6a79fb1b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h21e9de593f8af7c7b6e02b18dd921ab88dca8fb362d745f9952b51d034a98cfc84ecaeb9386a6cb0e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h45668b8874c4bb71cd2b0be48140a7048104b83e32fbf1957e9fc9e67f6253156ddedd850a18f8547;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hde0852786e302ec21291e4ef5260df12cb5a15dc522377fa4b828d3a88ce4a74bfad3db8eca2f9b04;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h58780efb663cc9b877b394ee379b19ca6460caca787fe3745af5e1ed658e45a7e34d61c675fcc6bb0;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h18ddc518fbcee1857cd92c7b1c1f83540c19d97758c926e060252f013cb0076c1eb277a0f04d200ef;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he4f07ac5b5d2284c5241dde1b3251668311bd4a38d364ec952cc8b421c476f842a323d4676047a81c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h70d07cec16ffa7c90c8da5b5e177a6647085c186330dc1effd45cad10296db7b94430179cf2b22b57;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcf1af609847a8728939f5cbdf0d7a7963775168275da87ae638a7d7f4b01aff4eed44079db0345da6;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd06352976964cb1b678381af214a6e6ff712a0aee7e7ed29aa4c1537833696af49edd6befad97064a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6aabb8a618280ed27a5753f575895ed4d72955c47234fef9fa31288e118e9ea8406e4936965579fb2;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8363f7ac062991f4bae325ac828685c8fcbb32b452166d7fa4eb62fc4043199e86ea5c0fc74d4ce2;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h727227c02f71583e55e9c587f977051dd73d953f8a44211f2ce2d130825da4ea9ecaa230b9b840ec5;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfa13842e0387e423e564e57b91b72041d753bab4ac9452d62a792160050c997721a70b4d2eccdd6a5;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb5ff4801180bfa41b2a4369da813fc26b058f579cd7bca267cc7ddd172f2e3b147ffe301dcf4394d5;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7426ee781bb88cf3985845165d59c40c7c5e0d87937e2c029c53a26788ff9ebed2262b9df1de954ae;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6ec31d3fd42e7cbac8b41435c1826eeff760d4918803f8b998846c7a33edbe757206b35863a2ea51a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h79c997f37f283bc010dca5d4e8db485433f80d0e9b4bc9dcfeb19ce64a41df05fc88428dd35e55efc;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'habf617ceb3d82940c73c56a7b6c4fc33165f7e5773d20df2b4fc06c1544301e0dd52ebd5caa376eed;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf77177ae24ff6e8e8076fd6c1d644aa219256642fd817f0c64feefead0505889ae5b801ffeedacb73;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9d9acf35eea146bb578e3b8ae8ecaffc598e503f809a4b327bd35362232705bf326e012e5ee3ca82a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb130ce4b78bf55200aefab1e672795fc6cc7f3327fa245a88e8f6f11668a4a97c4094a1a8e094b2d;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h43360ecf324c4b7dc4dd7ea0f5ef4f170f4b53c50a2743c6ac809397a77e1010f9607ec4bd595de79;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2a0d2cb10133001210eb31f405089db89ae4676234a044472724fc4886ccfbaa5cabdb7bb00c2db6c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb31b35ca22bdef289c02ac7bade92b36d7c1d609ee970998802ad8371d9e211aefbe93f3154672d9d;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4b29d5bc05ce8ffb0843f08aec8df81ff8bc452b34b5b439edfe0836cccd37b2e641c2be2b30e5388;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hff8db833269f97b7a0fbf0bde22535e21e5644fa4abe3dfe741884da3348a388cf5dd6a5be750deb8;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha745f8bf060fdd68aa6d9a4e017ecba51553fd58affa20d0ed365b7dc0d5bb84ae5e4bb181b14e7db;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbcbe87196baecef9a35955e52c626f432ae5abf9a49c44427e39bfa83886f045968ab17a1ec072fcc;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7b87fd91906f747f4bb2efdf9239c55b714c8780e6e82a453b03f593b19d89ec0c51fcd5e419531d;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h26ea9f85a183425187efdde7d0101e820490ab91db4fcf841f1bf6c62186076b3548bc41caf0c3009;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h896386f13fb6a2396e2623df5391e10b25b4e94e4179a74e5e3fbc27074835ed538a4f89628a0a20d;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3420f34097135ef9dbfd5401bed73eb25606aaed4bd786f66849e490d7cb9bb77a985c9cbe9432084;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h596a8f9f1955f3fd4eecc288a9224b95a0d128513caf0790e49cd1b01a4d898657d06db7d40b6921f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf0133d9c5431b94b417e307cd8c16afc9667d959d25d5f7ff2705518fd8fd444f805fc9a4dac974d4;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8b4203d241e534d8868548634411e80ed05bcc520f230ea46128849e5e336bba8f60617338f9d6d04;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h930c0c4c288dc1cb19f1bf6a91dfbfbc6e374c12312cd4af4001b1b48c7a2c1009332a48bbe0d5f21;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3dde0b25c9d640e825159c8c00ab1bfc9b15d496bb64e7bffbecb0ac1c66c5c2de0388d10d68752d0;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h31d4ee631a89f480814a72930f8fae48a8506fd0177d3de8c37f50d26c796ee1e75e56f722088afcc;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h783c8bf64f3acd91b758bbe3dfe48125cd1f32a8a05529ebad644a575e0d773b950739e77d53836f8;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5b6042e6206ad57c200773def20bbcbe06e76ad57051ef1ef1775d87a868fde76aedf8801c9aa2799;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3d9ae743bc97d2656c3de4e70377fc18012b7b8fce19e06282e9e7f10e33163d8c30d1daf8c61d16e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hdb4baa5e8d74a8e115a108365c6341920d205a97992955c0821abc914733879379f98697b00495671;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hafbbbfd77c7edb39a27c0a91492c1cfcb2ba764b8c4fa151ba6f942c20e95ee79eac36efab86ea7b7;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9238bfcd5ee6b32e71ddd392eb241df4dbbfbcf2df9c80c5dd857c23e59ae2283596b5e11011fc5c7;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h539900079ec08548fc7f5fdadf680cc352875d95ce49cee27f118553b6187732310dd8ebdeb2382db;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h972fbe2b3c2f911c5b9e52ccfb2530fed35172743ac4e11f0b91dae3ef063beb7d9c1f5da38e49680;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h98eab616ad9ae49b9632208194e26ec66d7cc289d22d6098a0c96c989664f1abf88dff355e4e896ad;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3306b633c62303ffb394ff623dd7601cb487900b4eff3649427690270eade27d7267e2b23e4c126d9;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h429497ddcd2cc9ffad6b6e5d7a83289ea59a9f2104cd62af0a924afdd0aa483136d4b1139ea031564;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3f2646b776570771ac2695cd3d3ec7e9725175043e825b9f1752704c14862d49d37f10f8e29440517;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h79e3ebeeab68d45602d7468362ad4fe9536f097ab3887aab682c6431325ee1d3cad5c70e8f18b604;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'haedfef87368a0356a64cd53355f1173ca76e1145fca61b70f29f655062cbb18a70d73213ff1231ef2;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h97377eceaa10740dc897d15e8927e4a7a7a8acc92aa4cf59e8f2d89d66c61d8fcd2cd463d366b5f1b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1ff5b3ccd275956b46ad9f2c02cba99266a90219c0de6880f1accb3f1379f538847acc27d7ccbb0c0;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he56b041701ec5efa81e26d414a6519e922b6018694bd1fe1ad251d421ca81058a24f97ad22c5da1af;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h143acf4fc202934a5980f8a36ae9bedebed0c371a2f615d30fa8126dc02f8fdcc8aee1f4a4f7245b2;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9ed025c2dd2dab7100846fccb7cea4eacdbea208123c95c76393163481e52634ec50e14389b349b1f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he72920fedf470130e04c9a81533b12f4ac874297bf2ebd984d4a2e8adba27a47fd9731a8ad6baee41;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6cd865f8db8a7b4427ffac5a2c26c09f395e54e20f519bb24dcf0271d67a5ac589ee90fd54d39560d;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4547debe4e8df3009be5d66e2b313596a9eed6bb2228ed8b595edc490fd5d90035243ad2fd98584e7;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h57647fa435620da13e856f8800f533d5f214723695a62257c947f8103a76e026467ca3e969cb0707a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcaf986bf741e3b5218a9300d7287d420df232325227147b3d6a8cdc46fa9718bd9e1831392dfd3326;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4319476ca47b79ce40d07a18f57f17b31f9d5ae5e01fc1a3556f95e9743c41a124105e072af0582de;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'haf0bb078a2a0cd548692bb4955634af759be50bd7bf8e3e0bb2bc8d49d158a4d9aada38c15df6bbeb;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf87e4e0ba9190d098d6b79afc5497291bc65a49b019ea137c4c2c11038e4973c5eb0df3548a32376f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc0faf4e1dc9bc5fee16334dbc178f34219ac28633da519acde0dba405e80db7b7016d3564a1ca74c4;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc216e7ca300b7725a0c6367dd19296359464d68f6155234cc7b0ce2afd5b94017079bd662736afbea;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8ddb7b5fc325c8d3d534b1485736749c20a94a97bba801d08bf818d5bc599344e32f979bd1b3c091f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h152786522873e7e0450c19f87df7db06be7ce84d583e85a68005d9b122b90898758ef718719f9d58b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc0b4ade05db02bd37e1193f4e2db219e28284d0b37b7b109f549df3999a0f1244ce66a9b60f3fccab;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h657baa325c2383c140f0b8ac9b95248b7881e666c18dbe773f8902281a4b4f5e8e0a120007b20ab12;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h56802abc782814b107580c0851ee595765e768e05a320837b39aab4d28131a80fe29df34dcd9e154f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4e389b1ef01239f9728365b8d9c47c56d5ddac3245099ff957ecc1fa7bd80e5feea613ec93e79bf91;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h84c93f3bb36381f0c660715495836414c430429f75931e5304e44c36bc09ef33808535e5a583b3731;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4798eddd469010c87efadcc498adade9924295111e5d6d97d645e62b008d842aaed26e0f8082bbd0a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h175bee6ca52f9b7d8e17b632233b508205a83014725306d6b809a97da7542515fb9ecf01f8ef8d975;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9fde411b5f528769819e8b7e7db636ec57e7f8ca6bc753d83bc6c480c29e5fcaff0a12ebf6b75f769;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf7fb17c146f12d13de1b7bdc6140b4b39cb44b2055ff61a203a137717abc8d73790f3603287275862;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h16d628b325acdaad9babe3205c9bf69716f435119528964aae52fcf57092c635588b27d4f03d818b6;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hacb50d587d5775d0eea53ce5e621314d4be4eaf40dc2c3f2b2c023037ed6d464f0078262ef9748200;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h714d5c85793f8d75b32f7d608c9b1e93d285976941d863df9cb52d2bbd0295fda2dd0017f21ebcc66;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5d843022a5e41c5745c75831340eb952b54ec5ae0a437c89f282b2554199e0417139fd75071e0acc1;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2e757c320b58f547a9a42480e7433752a2d21b24955539918c492833464e014c98ea02181493a888e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h992b205e4561fafec866c999e414e8dc663d97bc892239781e1728a69b90fef627225626b2194043e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4eb251f18b0495c86799a454ec136dc0741b0091df44ae00bb82bb3deda0b154e572c832f73e9517d;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8e6009a87fee6772eb3b356bfead5989bad51c8e4b56a6049e829b4c23a00a07984b180fe55b1d66a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h17bf40ba6df2147df3e53c1a4bc93b48db3f05dfec32f340ce2ba4c0474e8887c6d12f440e6fde471;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb2484008cb579d14a525273860dc4857c9594dd9c8112f8907e4f9f5efcf65690e6c020030722bb9c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h72de96b5b4ea5d83cc851a190f91ce7a4eb9de60435dd90a5142bb1a0ec09b07ba20c6726c45cd5f1;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd2d2e486c296b1781d727ca77fdfe6aca635bb10915c9ca8e4a39bbab03dd0186e24f681612c213d3;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2e3f7e22e88d1784973509f55344ee1a32b4e183bea25c43d3c0ee8f37fcc43c294db5d935819f57a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2ddcc7b4f368ccc3a1a68b228d590bf1a9d6ef4762c31e8f40f121f941f4faef674c76c35da513c2a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h36ca99ec515a155fac6656cba0eb8a54cb6d7df225da922e81e8c722891a01c17df9cf92c47ff1b47;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h359ec1378a9d3de06c46f144e87303a06271e4239740166daebdba626bf2d0e81223fdc6f303b6e78;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1dea8ded0aa3eb19b2cefe2ad0a01bf81ab14762b3edab31e3034ac477c651d6f11d7725c9470ee94;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8a1ce721cae6c67d707edcf693b45537aafbd0530b050572efd49e954474ecc9c9aba0921db3c61dc;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'heea7d6770bf9565fc7f2fb51267cba38bcc71283737e6d22436875691cbf8fcfe41b349b84cef82d2;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2ae50fde39f2c21a832fd1b78a88e2da89554f0cfd4dc6530dca198cbf942c2b9d568897349cb04c6;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd8770d1206757360409080db72bf568fb69cf1648bf40c93f42ad7cfe5b3a35f009dd722ad7e3a922;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3b59fd9214d867e90bedbc7d34b9d046c98b6330ac9a7dbffd940d184105df5608e446f97691dd41f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h21e96f9675406f35e60123cc684f711faca1e2b4b40237e2bdfbff31556d7d56e7962d33283b16672;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8d4ebb9f7fd70fdba9ca24457f64cd4901cfd81643b38c04bcbf91a8e515a5c7db47b6d9a41a8336;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hef136245bd4dc19c7925e985bf215556429f26c21a3acb2cce446dcfef353e6375027d85196c8c4ac;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h63ae3beb14601b7fb126f8614c6af70fed479b3319415108b625f52c2208193d8554e9ce34b2679a8;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9dcaf6a9419c23794479e1c2895e92d122a1e6dcd1daf2b388fd55f59686f78e008ae98fb46c826f5;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd6292cbec99a50ee9ae342596d816e4af09cfe9c7a702624def97875c95d77f97ec6bbe78da45655b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5a1905f4054776bcf2d6fa76ce895cd464c3fcfa25e4b556306961e7d476e9cb03ba51457f5a1a403;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h88442cf6525cd024103f09a88323c141c5bdb073cdf06594066927373cf8390b30dede218da9ccc7f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hea03dc39d954291c55f3323af77baf31b555644c8a13d23286ecb24c5d0923a33e09676f3bfd1c704;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc537739325b92156af0940287331d9791d65ae269a9741d69ce6c54449ea6f596a26e61a8ac5272b5;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h91bc7f7411b1800a904cdf04c34b8c633d13e8487f469ed2f2b53918408add6a7ac1c5b38965c5524;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2f620d2f14e5da8335747721320449b2d30c90b5b5a7c2a07a3bd084d183c4c83d735853653e051a1;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb78ceb660cf7576ad85e051d72f435c507af5f8ca95866f4b6201b65798349d17a4a9458c40772d90;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hdfd77ff127019c4950ecafc3e2644621cf2fa23c1863658dd70b76a04f60d1303858ec6de372f4eb5;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4f739058d32716a51bbc764d67fe0bb0920f72a0ca556a199c672306155157fd8a5360253a5d4ef16;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfeb80635c56593fbbd565511f0c1d34fd05d30fec78c68b2f132cb941e22edba07bfad2bb24d99551;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1120e1fdb95ad5fc09a2e1f9d717bd922715a8ed5420741699c39d454e8fcc6bc400da163e1cece43;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h857eeb92d0cb02cd2e2452730148080d22070dbdbf3024477bfe0bd46d385fa1d908ec69e45668afb;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2467ce2961ac011f417f3ccb75ca592004b16b5099da392269c0e0f0a8b30764066ddfcc6c0f944f3;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h566ce5e51baa83e47b1ce628ffdb8db7d1e611ec0d28124319afdd36b4df261d5518a63c25e516dbd;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h75d34bb9f043b94aa9c5ae3cee19da71887865dc261a6bd23c6191508311112df93c3d81230e1eed4;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h60fdbed53a586c9e579eff1be28be0265a0e79267c4a36ea1f835722cdcdd9573cedead7fc814d735;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha0d7a44e77d9aa8b60a158b04fb558e1666d9bbb8dc9bdc4599683e3c9ba630014e9254a4dc58872b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h32f8219732a814449a72dbf09ccc34f920e06a4e5a0448ceef0d62111bca8a1c1abe2bb26d9be1b11;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h728720dae1eca05d29dcd99fb510ee1e1f216c9af6c2e6513a8cbb4120d78adf6cc0cf4f894785587;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd720da397a7f848019b6ca78146320ae14c22e34419d785aa91575117e96d892f916ea9c29ee7f43f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1a4802ea4273fd76424bf4e986f2d781bff5f5f81aec2aaf3d1d2eaf2121f8489db5012e88ce00296;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7a564427916d93afb2041f1095660cc8926d9525396f64b76f11719554f5c2e3b919b5dd26618a2ef;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h269c7b2cb598818b71ae8f390466966bcd5ce743637a5e255bfef9edba707673a5531f5817c3e4d8d;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc1e8896635d93309a068fa15edd2473e8c4bf1ee40807ea74e5d84a127d02a390dc6296bace0ee21e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he5d391b6400e3174132a57aedbc4e0c331f5048bb1ae55e052d6c3af2d95092bfa7a6a1e0030eaae8;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9dc7a52c9a54f1852cf1caaccc10028c8438b6eff2d7a08ce5a51bcd8ed091f1da226c71495367fe1;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h405592fc81caabeb4fabf12a20094f6e382bbb0022dbc76c3ac7772aca5881669e08410b0bdb7679;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hddd298d314a72453b114c834ae292e9606871d82d851aad6a911263dad8f654dffb25dfcf3b899660;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h17fe0c0ee0a7e038ee206346bce406b043f542811fed38c65db3bc6ee5f1c9729d9e40908ecbf9ad5;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcbb48f78ea2d728e11ddbe6afd9b81f011c75697919ab39dc751d7486435f024e061fb3d803355354;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h75c3e1c9f303893326b4c37710229246ea922e381ec280f13c083323eaacf998ad4e8768b5c5d0be0;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7fe831f4ac4f42b22a944a70ac84b042628d24a12985e3c29c3fe5b8df73d0de83f82871d811d75d3;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2a2277258d2521150cf9f611ccdefa8b0691832a8e11f5310ffcc928dc4c584bd33e81cfefb13a5ba;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb0ce15ed68fa8f7d4eb53474e8e5181317e4f69c26281886f3a96d86c71b7f303bd92f5b3b5bacc52;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h24d4ac9afad4ce0318f92c7a28729ac0f2b799562112b75212e465d983103707256ca993cf9783bdb;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he7f8202256fbcbd28ce4e99d3b5cc60d493582082f4825bfe6065915eed815048ad6f8664a0959a49;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb7826365f0111888ef8b6339b5b8e5c0cfdf73eaa26d897e14f884cc9f7edb528c2114eb21594d0a2;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h87d284c847eb3c7717e742ca0df8ea390af42c1b88977646e878d5607c5e768bb16e60e1d7d94ae49;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6712e501660abb9cdc844a9fe7a81b070f7af16d441e97612162ed90bc3e7fae6c76218c5949f3d19;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5ed179d17c482d8bcc1631237dde9f42b478caa56acc45dfe4e7aa42bc401aa10877459684d982ef5;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha98c9f028a85bc16b320c2c49832ff9360240f51291ed3f4ce520b2482323edc0ecb63a4b525c1a43;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'heb84411618fcc0e988e9426ad67034cab711d86787632fd32e2dbe424883e09d3ba486b7a07f196b3;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3a669949118380f3cf44dc3dbcda82801a10a7f1a77b752543fc673a208f3da6f4dba31324fefe25a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc297eeaa1c5275f7f90e13a01ac4d0780236f28958e219b79a5b2b6562d4429cd1c99162653c21d6d;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf0586441271c8f9981a2d0ef27fc4cff241468cc6c7578a86caf6358666e0d77c874278d5c0e1ca2a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h61561a8ee480c82b74b0c722b8cc695fb3c2c3dbc62da00f1d23863197789785ffbbc7aabb19f52ed;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7dd413a53bbf8b3ccd89434dd4e1eddbe638582a4348c83398ce9eb7251b856533b77ced69c08eb95;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5baed930e1cf041e5507168cea85e6a7a56724e8457a5bb2b7fc748c0ea6369a1963722aed9fe096b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd8fe8f3bade53d854c6ac0947819c158095a4481f8796d85b3e3005d1ef04a6a52f94e4bb7ab25fa6;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6d78bec75880d5ee631ab9bf29e2a8f1bcf449441883464f6793ae83d13fad654365e704155d3c270;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h541d3c2e634683a4a55305a1546adcffa027eea2b68686e33289c9721396733cb3f96c55f03f313cd;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcc9275be11fdf79938d4f1e4b9e032b78a190a4494e2f54e8176173b7ed9e70eabfe28d4cf1f08c23;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3eb679ab4b2d127ed86c18c1b89dbe975d57e286567a64bfa058c5abd466dfc0beb037d6c945a3817;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h565be4b0c6361b5a1d0d66a6fa4607a4ab9c3c2f3654476eb4f2319d8c550e771129abeed9d15d990;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcb05764efa78af9bd706984c2daab53db973fa188312094f894408eba1e40517b68224df62ab3ba09;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h53de933588002886a5553d212abdbd82b00a787959fe1eebdfe12bee9cbd90e034d4cf17b7e033875;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hdac61f04372b5d07899451d941c5af6d4aff5dd474407d99ca13d8577114c8dccdae11229563d11fb;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb009db7b4299d6455218b6967cb79db53f9690630635ad369cd318318ff7d5be5bf58451eb485f185;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h701142692305fe4d20796cbbb78fba9057d6c77978dcb98e1ce49f20cdc21174b6aa5916f0aa75ac0;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc64defe049b9932e3cbecfb90508808e96d05751fd9f39ea72ddf0c87233bab3eeb3d2cb633172f7e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9a4d75f8c56580b58a4a31527d998a45417a0464b2f7c117323be0b02129bd45d1b0be80def5d2455;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc2fb653a109d4fd08f613b33e5f8bf1cfc55f7ad0f1b112e3a47be7a4996ef9d737ada61b3b4fb321;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h76974b51c688e1846a6a25f595414f1e9207bff174774ad1dc39cb85e0651d9b9fc3d05d75951fab;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3d6b028b61eb06c237c5ba6a08c76bbbb136019327d8b5c3edf05c19b5eba5e1b0e2b8bea045b9935;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'had87591fd54dd242e4c79494f972b9e8d65ca144806eb3f65307c957d633607859ec47b70d6996a81;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7e5798efeb7de6dd0fee24521b2988ef0ff7d5a1fe3ed4e7f69f8e85743d71b7f32f6e4df55936bc6;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf40e103d7488138ad1e7559f31eebe5e59c33207c4e93b3bd94872ee76ef30d819f06a66c28f8b68e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7df4ab7a3c5c10b1076fa3f0442260d3fd24e43c9267916abe6713d6c6a0fdc2266be1d49d41d5d57;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc64fd24a0430ee0f6de16d6d9a1db95d8a8dc934718afb81909205834cb0713fb1d767e00a7cb89cd;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h54b33f4ad890899ad74a6f78fd9ac46a16c2a14b36e6723a915e155e606f119800074f6c5328b6b9d;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfc3a981a2febdededb9b79f566b1476220cb9ddcf032f5e18f7beaf2a6a8efa08f0460ef21756bdcb;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h641b5bab5bc6280fae5fc0b5263e8efc0f92144b4bcfc77c041bf5359b458961c2252c5ffca94929c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h749170a20e37d8493bd23b515b6d91b2dcf20e83d0dd8f155baa49b51a1cdcdf09a82d39b3a2b5482;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h264df9a7a6a288060187a34ac1abdfe8210f022a28360c078b8cad3006051e0e4cb940b1285a80f34;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd2fce744e490d9e8a700269023c05334adcbb22624eab78b00d207ea3a19f45156ffe6050783cc155;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha82255d72206748f98b15fb681da7fba08a404bee9ca4cfc7e39b936b02032cd7a9b63cec5dcb8d2a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd5fd213c8965d102aae6d69dfb56b9857658c3984601b3092d09c827cae428293a3cad3e02f2c3d16;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd5814fd371c124889f53ae14efafbdf8aae19069ee5f551b4069f066b358153e5165cccbf8a7d2cf5;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4160a36a6837535944cfae8427952c838ebccdbb80e72559be737021d326c0b49fe27e9af38e7be33;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h44ef0701a12a6a2628ea1c69309fe0ca24e0d452fd554a8d71c14987ced1ed9f26d3d3af06173ea62;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3cb2995e05cf13a40d27e370810f6ce20fc59c823255c69876517598c0a83629ef60b9513386bd9be;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h52602957d0349c9652c7354f42c9f89194a2378dc937a4a7e3c312a2d96f567028443484119afef46;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc27e2e4bbf5e9e19358c02576e585bfc95d0a2a3b1e47e5eb055b6432b7f48eeddb780e896e03f4ed;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5300ace51741c207d2cc74d270450b09bb2b1b9b7b1b4b48fa482bf77253b1f5d2d63212faa3aaf0;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he77eed2e3dd158648af604a6795e29987f2261dd6c6ed909f0953fa480393a7c669cf587fb39d30a1;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb329e62a7950a07523221b3b97a2fd294605240cf7b68a5259e2aba892ddc730895f183182b388087;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf1eec28f45965e4343c144039a4880bb1ef2486c9439dc4a98a76a3e4d4412f018760ccbe170d6dee;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9c6078928f97a98c2a6e9bcb79a2f1ce8e87b16a40e87a46a053472b64be9a6d8bdda0b4ec91ec7c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h93b651c5c84c46b1e207d4020784d51dfdcdd902155c07c9e5bb3064e4016f950a3a7d22c3af65233;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h932fdffd04be6f73191acae69ad868d157d6f90f7fd5044587c451bfd0efeb855b3ba87fce9319509;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1c7215805243d34155aa856583653b132a44a7863debdc948d07870a555f28689026488c3e4609e00;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8e088c64e30636c3076efc50e6e1142443daeaf59c401877e41fd1d6f72b713208aa4cffaae51b85e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc937a0d23ca2034ffb20c05bdbf24e82dd78336599ef54f44c1160bbf90e0169cd176fd35d022ae06;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1fea80078427f4b4856e0b419299020ff2086b57a55bd93f714adf3fdbeddfc40d9b6dc84ad715fd7;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hdd1d7f10946a706dcd35f4eee1a52acf2eecf500c47ec2af45006d5fcbc64a3db3f39aacb33393125;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb0ad9a6829c535e2647514385f308d277f2056594a8f0eba0f15ddf8ff4cf90f489e5ac36e3da21de;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h65dc1d3a8325de4b3c84553b644c0aac0e42bc2202d661c2f7f5602ad860591e155615e9c1a4771d0;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9c38188580303bd9f7bb79bd33269b99f36c3010c8c94b87410ed10d7aa64b8f922f9317d7875e7eb;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'haa99ab2f10171f27b2a37f6c974b139e674997f4ebf7111f24bd7aea7221418bb479e2dbdf1f2e640;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h844d3e5890a5649db5378cb8b9bee7cd9a1d7970274bc56d7fbe7e03187752edf82bebf4d657666e0;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hee9186f57e9eafb02f8ba30cc81fe50d001611e1aec7f71493136c8f096da54f599dcf9070634803;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc3e37f44bcb01bfd14a8f4c661f861e1b3dc0d6959a3ee13b28e9035e375869e37743c2c81d9e49cf;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h63461a17e8ddfc5241e1a4d60ea968c831a979097fc339d47db552c439580de6f748d00d4d6ce9931;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he3824107a4bb6eb4e56bd58bea75c72dc7873d704fff0c7a4ace98350d9c754dc1cd1ce394d18e8cf;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h86e91295ba7a5fa0968ca6097cb4981ecaa8c5bc01c7125d0211df7fe2e8d7fa0d3f7c83d1f415be9;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4be12a753c5efb8edf35bd595fe478097a53fb115fe34ef8b058e8dcce94a2f8c3218420380739d3;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hac0e80336caf1564ca1f450b979bb811dfb076d10ab7ef123110a4f1155d29e09480e70564c516a6b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc3f822456a826cc7fb6fcc4de96c5ddea0ffb8e2b0abc635aa1a54d0537b2d08f843312cc73141930;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfd9681cdc7598b5fe793139115429a20f289b2eda117e4fe43da92eddd8fdcbdbe5112caca000daa4;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hff647fa983b8ba7b56643631dc9cddaa4093d26082718c6fe4663846824618b6747edcedd08d18c5c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h916e22e869b1167e68b0884f403452c3c8b7d0172597460bc49f20600c32a10c820ca9254cf16acfc;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha0bd4e7c53c76785c2c2d987cf120cff0cd7c90024c3984658e179441c2f96e2e685a1d474393f57;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8192bcdb96ea93f421745521538238ec0796a9cfc3836a8893e333d6fce140307b5d6196fdfd0d870;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8795c91e3496ab379a7451b3139ae6f5f9fbd581e5db804f0a7d382a50bc887b38c535028cd7169c2;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2806dbd608e9e3b8d231f94406d81576b720637408b5bc0b7bfefd436ce15f8784be57b5245cd5d1b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he9f684b414cda22553afea69a7e7e58faaa28a560f3f3b620ce48d12222a0fd313fce29e758f3f8ac;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbf2c6e7051c5c19b60fad7a2ef5a64daed1a3b1e09a4b6be61312637694ff417a0329b222e00819a6;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8d2d1b1bd455b477d496f46874cef8029ab62568224dc399f3e8184186a2df0c88626b425e658db74;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2cc6da947d298a712c32df618d255dbbec37ee449510a522975a56b5f66cb02fd6243d0e2ad745b9c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h42516d5cca9ec20d0c713eebfc33643bdc6259889c288a92675f8ac5beaa1bb88a684a3d5491de185;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'haefc45a0a9dcdcf88a767396585cd2002db8e401ed7980a0edb1a83312b5ff123a66fe70c2ca8f2e1;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6fa534cd7cd412836597a3ed403e1b595c82d7a9d2ff9cca2ce5974392540675e74f981cf7af97040;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbd51134cda0f4bd2209845808525bf22de25f31bdd15843a27315e0f75112b34f06ecc1095a6d37a1;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd9876d0abd23632836ec6779c4c57b03a17aa08808c096c4bcc1081339029b0c6a192886261e45674;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6a79e03f770bc407fd4f75fe05d1b9abbca116bda0f830cdc4d1e4765085c88596407015ed56754ca;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hef9afa8e5fb6f4f8e7109ffb9d4d7e14a9dc537d49e541a6e96f647f2a32bfa774eea4674149b0308;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6fb41a3024219c607a4dbf780eea85b0a5bc15a4245cc56908a5d1d3e18c85b70e8620c938d5db14;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbb59b4f2b2d8051590f9ab590fb4aa00ee9d4cda61c3db95c1558fc36547664c00f48462297fc1088;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h93ce40f53bf8e007959ac4c8d5d3fc007f042464667ba04ca1bd66a540ea741a208216b0e38702c6e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hef68950c26530af4ea1378e3b6d7e3f7056e450b0ecb09a9e380e54fe3a40db46969db7023b1bf8d0;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h79877855bdf6073f2583fafaeb6c6527c39894252c3855e47a6e1c3312db410f7f106888b06ebc4a3;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf360766106e67588c04b70fcd0f09478f1fbb8dd09e1017b38a72c055285dc7aaa392ba79d28e7de2;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h962930957a31192b7408d7e4b86e90170b2c7d39a4101cf852319181588bcce54d1d30438bf80ddaf;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1380ca1af65c6e2b4bb1b74a5ab375b81e46a1e23202f218479410536d2ee6cb69e27694db8ee24c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h96d41cbdb1e5a74718cdc1edb9ed1a88bf0fc6502fc6c89a7f7efc2f3a87dacf35362c3e4db2a3f9d;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hae0e7066c0aae5c7264c57b53d7bfd1d7ff055ff2c129901d21328bbf0143c9c63a3939b962eb79ed;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha0725898a12ebb8f5356f2835ca8a5cdd1b6d29f69cd04f364449b751d14d8cff54d5fb8933c3afa;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha087de47eeda59dbf2d313ca8b419021b258cc2548ad0c96ef41f20a199082f85c9a45fd52fcf77e0;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfa89c7e5d0617542abcdf52fffdb7cd4c090c91ea81b2233e3480725a5df19a1ab59ed6a3ac2cfc6c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6c9c4cbb57ae178904268ae688afd294b9eda5f877a685fbb1c67844669a4d085da30df7041d160ea;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h43725cd0502ecc34323e8ad497f6039e12c66c5fde45ddb9393dc7c2ee91973d93ffe17bb84b59ea5;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h58ba6e25723ea1b7959ebfc28918e817c2c849dafb1969fcc1d0832c6d8fb4c4524c57ea4bc4abe9f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h169f08e619bbb1e4378944def933dde0d7b624663f775556fae4d2cb4fc17c0560e57fa653f815707;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9c84094bec62b038cb40909020fcc0361306162fcf885ea532f051d68176a29d60358430a48c6c5f7;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3a3f7ec6bcae3eb3f4a3593361177404f81f70ee68343a3e28a2ea50e42569aff8de83277f9b49cc9;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h990319c6cef972f9a124a0bc47591976511817f1569d784dc4ff408267f0a1e2c8317e4fc8b4ec2fb;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h46d4fb17f3a31d0734967c5a516026d4d59863885f9a1c1691026c4115127eac5300b033e35644cc4;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8361392db9dd82c01cd40baa2483ef52b031aeff157834dda65b8f7dbebb0ad753ca3dd4891e50ae9;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he82006c7c93bf8142adc6e54a525481478cfd7b4a4562ecaf03fbe648498c20b19d790458c16eacda;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfa6cf1cd633b2aef0251e30b643b28c2ab04f654cfc01f8b045331a9225470fb8ccfd247ab1c8fc3c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h32747adeedb32fb3734c06bd2fbe395e486c9ea41518ada45d2a3f6c235cac5a0d74ebc76b6d93b33;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h85d1b74f1983408cf27d358f1b12cc7d70f34081ff3355dad9166d7224c155e96b1f5dcafe7bd8f9a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h81fd27e7a6136c578b101ca69c96e3b02f56dd653031ec5c0fdba0d007862c9ceaa4a3fc587574ce4;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha77a5f64067b81f0db75d2ce5c6d468ca1f1c96998cafa43ac1829f2b25d6a1905d358b327bc5c46;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7f34fb60ef4e7ce6e9e89418b3654721809b107bf11bc88c935cb66b65b617ae3bb9e1b6b220df11e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h92646ac372ad70a471e0171722e5787c2129e3b9f9f07c378b20c24236bc6d382a11fab49ef4de9f3;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc2643df637ec6a04e80b1240511ddcb863269971d0d832938b90eb3ee94b3609399f82e56b325a1ed;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3a98b06282df3a4dedb71dad94f36edf5c7cfcd608a1ee9c64ff9829fb0d7e1ed6b322493c74d0bb0;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h83a54f34301be4060d2ff8a0bd4b84ea0a32936f30594ef996ae8be558a1e35489e941753e786129f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2211184900970adff2648b1260b07bfd9ae221a107b025464636c1b46e3d357bd9ad4e6775b3179de;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h22277c18bf28ff3cbac4125b6ce4ca6719a5f1fe313fc2714f5be9f80b790cc1b0afce78b23af9fcd;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfea728664f5409740e7f61d3f84f8b1f45e5c35e42e3d9264901fac341eaafa796fb29f1d9291baef;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h55103fedcf7eb1e025386a1ece5e77523f57ca85ba724af4b1930d6db243c75f455d3d5fc83f71a43;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb351ae9366e97b3a286a26b29a8100babf83c73a1841e8097c8b28b0bab5ebfe91990e815c84fb36c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h762b651b4e8e2e2e8c8fbaf9eebe8c45abaa152d57412faaa5df4e245123920da83ac2be2c46e93c9;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc626233cb1d1a7394e26d841606aa44a9a3584600b5c71e21823761c4184c788ab2371beed6b60530;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbc32e58dd3655faf509defa1b61467d04a351cd5b631fc2e5e44a5088403c342ce1d6d1194b747a5;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd1dd7c0674c0c22770f69da7a01f75a1c09b9bcac4e76a3fb9bad735645c486db5ea7adc0125a2606;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h76fdd4c6cb8a03bd83e60dc6d4ceb4fbc0aa761abeedb40b94b6e3d5d076f808b87ee64b9d0015c39;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7727a45a27f95789034b74c638690ca84f8c13cf17f244dbb20bbd0b447aa3be21b043f9d8ad4e0d5;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h95bc22ede470e315855619d875e7cc5fd846166df35703bbac697da045ee35d784c3f0c522bdbaf7d;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb6641487d00029fe425193a504d0ebd0d644117cd60257a623d1f8dfc3bb4e8cf914a8eab9c265cb2;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc59d0561ab95278f2e6671ebbf40d90121ddfaaf632c9c4149714532cfb0a4b48a193caed5f54492a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h979b18411c5a8945ac2c382d280916d7b0539fafde5dec3fde73b9f2b3208fcf3fba5851ce1b6e132;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha1ef8e06cf04de3d5efc6a3a6e410236e7bf866d5fdaade914a931c453d6e3a9ac4afb0ae7d5846b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hff2bb244533c19602b140a7d65be2ac80ce707f596050ff5e0a7284ad8ecffeccfa56ebee58a8644;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9ef64d1225b542a46d9270b3f1323adeb43cc1192f4c6aa31283bd7adc761cf06562680f1da77df2f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5e73d610b678e49b2b6d1491664f6ebcd5894b5839bcb8a16ffc1c22bc904381742012767c29796ce;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4fd2affeaef4a5f2c0be170772580da30d4f8e9523d52a5b6e2fb7f8a458175687d57e5a49b18b59b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha30c733fa71f1719884c96c5746b9055157505debab9abf7dcdeb89f9f9130aaa0c2a0e34336bb894;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h38e6c5f243671178e8765a021de11b76ad722f4b85366407c176ff8f301d03ca98ea025b9d62b9889;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2f9a55c42ed8d5ced6082a36c9ebb16a43602a8a7e3f57869c5dfb9fb3709f62c012573e1b5ae97a9;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd44bfc58ed537bf82b34b323190b12dd9919b0b95274525b437bf53f97da8f54a7eb4cda08e2c925c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h647738221309d147b4ac2445d7b446909784bdfff5b3036f140706ddecc50daadea4e0412b2acddb7;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc1fdae2f74c02df51d4e12a505d605116d0c419ea1a4265dcfb345076de36a68c396d1db4b06178b9;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h31c98bf9cd3fd5671155d6ff1f0b4737fd98b6d99d0540fb3157074eedf65b22458571c5436fe4230;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4a34bcfdac494bac88d90df69df338d25652a6277e1cdd22c159470f7434e9b6047893ab6b5de1bcd;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3306bf49200658988a39fa6812d9a40f98c0c81f758e6035d1d9b38e9055db076414b203a5c217f2d;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbb532a3d5836f50ac07c23c4071a8b3e85c9d2c584dd1c7886ac7d84ac073986072af3aa9b178d091;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha60616b53396c298a3800caf60e5644ee36093c62b4701e218985bc1b7db6cbd88ce6e60bb0049ad9;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbdec3acfdf3d70c329bcc91c489c7bb5985f4a30f6453a6ddac579df0403b3aaea61882e903fa474;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9d9704b7c6cc8c6375fb88fa7f939be649c94581710a3b75ee83edff19fedd7cc79d889d80ef028ec;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf36e3de0e7ab0e14954a7a6c2ff118bcf657d5aec2cd4fe95b32794ab4669d4efcd432c76a36dbe6e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfbbcfa8444815d175f513415f0d631dafedb9dfec131e0b6bfe0ef5e3bcc18627b1b0b34b2e94ec46;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd527c1648ba934121911d0e213dabb7acacdc6ebe37def139dbaec8fdef332b2593359a9fb916398c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha4229c8b66237e32477096798c6b1a3300d7ca77341e36c821bab9839ade99ccec011bc673ab0bfd7;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf468397e1bd56398ab0b96e9047c630090d322afab9b6b86442f5568821593216f3d130c8d6f7afd8;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5884fd09063e150a09485e2167cc83608d9753d33f284d20b2fabf2c246375e31bfc465a30f4078fe;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9928aa0088ec4b05695b0ac321d99357808ce0210a05e7b96894b308e124dc9f958815d6dec8c1e2c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6c0e8e32ee8b01efeae8bc9c7fbc78b6ba44053af4a962b1c137d19989d14e406232c144e2548fce6;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h890675cf305812cc1eb86425d31f37078fd5e2723d027578bfae1637e8d31bff5f933fa926417440c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb4b004030dab610cf4ebe9a4a8efefe02cc5209ffff972368ad2c364952ab1dba6dc7de32b2cfb5c3;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6f88b2c626954607756b73d66081abbb31b32a35c9cf1d2e7ea3ce9fc7495f5f06616ef6ac24c912e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hab9b35c3a11704a0c679c9620d4d0fc9bfa973c0b349c5c9e6880e1450831de8283c50b298136aec9;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9976052474e5f0be21c9929decf17861639944b3bb4e31fb03209ec096346cf3524f0400ab70a6b03;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfdd6d26738396993ebcbb8dc208f052228ea152ecb5d959b18fb32653d0b6d34dcbf1a507459fe449;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf4fabdeb9367cbdce2a1bccd548c3dd9844ac22a1c43e57bc1948d26120379a1b2bfd6c024e71faee;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7cf3456fe8b6df4999cdf0f13db7061eb14f2b27cc90296a79361b0e9a7612542de575410389d89d2;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha10ad891bb64a5db7092ca63a32c8fd22f7455b6b470383c903f71e1256712b71c97a2c0ddb701f66;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3b780836901680080e35109262b3bd3be21a5c9bd951753ff38f93bef62b14ad86f4c234158b99a78;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3cc0743da38403f3763a62f21b092087b8e3b82fcc8baaf001e2f9891d1aac458945b24a0d99a3ec0;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he6c6020e340a5ec78b400b131d6310713e30d37259716d3a8d67f65ea628954b5a5d021359a251fb9;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h856fca8ad611bef3b0694170a58eb9f58cbdf51d239c590fc780f2bc5185fba688a44e391af96e195;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfb6e47d27b32f5cf0ffb9d93cd43371c1c8d0e50e15b31940f09346755a61c36978c44931b2ba4a08;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf83a5cfc8572da2a39c400f5814c1f11e4522016301caa71a162e793533e7039dfbb0d958e1e306d5;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hdd35aabca1d97836a1ab560d3aca8e2606bd1bef65ab32974099f1a58065ea73e260afb2e690e8456;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3b3c1c46a3c124a9a36fe034a873e442bab7f5fef5390f341f103962b49df91de87a0379968bdd68f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hef75df5ca771f8a65d7462f3a083cd051aefc25a837a0dea75f529be6f36da8cd2a01b176cc7ea5e6;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5c63138c6df0c80c61305aa73f3cbb7b9862832a8690a6822944f0368ba5f614f29c1c6e683d27e46;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3b8b73af59c8318e537be07613ff2a670b31a922dae32369a656ba2c9c682ea6f89fc28a334558a17;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6d60e9b0a742b94feb0931772c6da80dfade1182ec2d17bfa227c93620b65155ffe1cfb5c4396aa5d;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h805120e7f9aa143eb96bf1f8a9f06a06156c3a489f2252e6555fc7b4dbb94e75994f233837c091882;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h784a933c68f4fb1e366e627caa962bf8e9af8b9f00f6e22eb9b5f4e596efc12f3a129c7976db93098;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6a33234e1f16963001eab5e8fb3bbc208fe49613dedce142e3b94c56d8f056ad533ac7ad5696d5d91;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6a04cf5c418e7a5606a083fe252080e3964d36722933558959ff561c4743285db1a4b6dbee6a7cb5b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2e3e8bedc20d067db68a1e1ccbc2f085cbf244ae77cbf53f99eac9b4b66122170a88b403cf96239d4;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h617d6052d1468c95a0c4eb107e9f51a3f6b4e232dabc907680e83f54639eb6d0c455c98edaf80199;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h75e1c3ec0fc3af8031932c9c12c565d67f699c4f0f3e349f1ab0985dd227f3aac4bb51eae1899f101;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h50bf71d1af6deed201afc9667623e5696af815a85c0576dc495a95534ea67de14a90eb9a41c2091e1;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hef74fd841afee45442393cc539bc629c8461cc038430ed690ecd1406aec53c707f4591a50a409a53;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h96bb1ae42826035437941e91f1e94a59a94896a5e15b0b84f70bd40e2c23f3a9d42603e543db619cf;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5ff8e2f57221166b0088ec3da9a5ed0d06c0aed45b8743b6d4de07ce48424d485605fa7339b47969e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4f95ec388a7285dc28db5ec3ac91226cb4875c73322ff9c7c353ab0c503fd1008b25ee8a15f59ef73;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h54dcc9a7cf25d7a0c43e560b43ffd7bff1d7aa6ea251784612996f6f581355771f51556cf396556d;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h710c36b08dbff068108067ab91efb01b96884d5a150188edf851b75be0ec263e158b5d2a114d3ff4d;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h225cc5d2f6317089e20e952f1c28c623e045539d5275b8f71c2f92c43e59cf5b02f4a6a2128e9bccf;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he55399e3c9bdbe19af829c30b668b98ca7a775123d4edfa0a1976219dbe7c6fb9c06ae200fed67c74;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1154540fb52776ce596337c3d794a5ce29df17a916ee77a96610a7b720c2f724a2b1feb1b1aab47b0;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h72d59144a46bdec3566b48d8e8d7216a976737671f73e013753d5b9f5782d8c9da4a2b2b1264f0431;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha3ca3da9563d575219dec04d0f3839f0f0efb75282996dc3a60076cbd8f3e6975915742de294d4357;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h98188839938026df491ecba5aaf4e876368112a060c0e83a9270d9464bb959fb57195e814dbb34b53;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h143f5323c8e942fc0fcba14d0336aefad5229509e533ec2c9d5edfd49ef0032c2c1219df07ec09141;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha57815fa1ceddc3e8c5499c6ee143f0cedb9914911a09200fd1ed1356a404eb40942f63f23ec908a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2355190cccef817344a984859ea82e5067d647cdb29f7fb719f129dd0f9b7eea9cf05f88e6fba2717;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha3b6b931b7013852f4bc4ed6f522d0ba409108f81ebca31779bc50ad4a3155cf7e7e0cc32fb84f7c4;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf80b743035867b582f3587447f680f0316f2c588bc29b577bde1c54a7fa71df02ec0958856d83954f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf74322180ebe61c44a48f1d0a96abef7579f5a2b0bd30afd6c07e7f091595692a341805ab1d5a5ead;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hdd1edee268414b236d2952491377feddb29f260c0dc8c955b19d664f7c65aa92a2a38e6df97c985b9;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5c2944777c9e6e4ee2f40d67f5408cb5042f50c640102d81759c4ee320d7b9ec55fa4c77b47687cae;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8e06a7e997d52dbccd246a1c05fe2bcbbfefa2d4e0348f4702a7b99a92477f4976d3fc00f2efc516f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc223de6d643829f560ac27f957a5c7476ef3d1540550276d35a176bf334b7af12a829e51ba2a6d7c4;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb5a979008c5196b7dba294ab0b59f118b2873150af42e236b649c4d3bd448f58367e7de5ffa572a3f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb2df5ab84e60d29a557182d9eb40b231816eade32982b6564d0f3c42463abf3cbf39b8eead3f4e1bc;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h99021499e642de046995a46eface22f9a32b95b5e6657cdbb1ef53974a35eabcc12d96b4260ad3a53;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfbc9057cbd4f6317aaafef8c40d1ded15c6e5a2fbced0b0b33132ceb3d6981c2281501f640bffd2c8;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h173767f112f17043a3b323395fcbcf0e46652177358b085ae4aa36141a0fa83b4ff802111eb69e081;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf9b3eed27eafd714bc185cd549c0b5331707eaa49f59be398d0730fa6b6d740058d984081c91f7750;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h710cdac43eaec51d84baaac950639bdbf7cc6316443432ffb453c5d5dcd5700c36c678ff6618d8dd5;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2ae4341071ec0009e3b132d6e2ba6157e60c15f6efb3666f3a6b308495ad8d818ba5090955ad3265;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc357bd80329825f78e355659f6e3bd97e0bd0257a1498144bb6bf259745815fc4c1efe82468d874f5;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h26e4b07fd835bf9a4ac9d03f125c35f51a4b013511218719f18b42fbd1562a5ec64b37d41f2bf835;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7da3b7019873808fc8910710fa8d72e948aef673ce60fc48743ce84357622ceaec83923a56a342b1e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7692a147334f58214665d8b6beabcd75bb99e05d667fb999202f450404224c007442b2f9f89c03bc6;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h60836c506f06d2287a1e8954f2bcda70ce93719ad0e79108980db46a8fc8276934c567d8795390b28;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb26a804c4bac07c068ccb9ff1a7d783a52325a900a64bea0881c49392c20b353b9a2b0cdfb6eec94;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbfce580d8e80f7b2022402b4926593001677f87dc87ad175c7fe09969a16aee73324049cd8d2a7c54;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbbf47f72e874a0b037221d58cb98e2e60510c2afacc33e3448e47ba723e9a173c44283eb7a990b5d0;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4b73244145b5c633fbb4f7ff1a02b632bd3f5bcd046f8c04b94017584f958dfcc3942fe454d00a940;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hae884df9aee755f01d03c48a151b60232bfc11f84ad5830544e20fee185aff79ba43e98993d0e5dd8;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3f5dfe715c7c74d2eedee9251fe1cf5f48464f05e2070a8a2537cabd9e5b650aa4093899f69387554;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8363e09d6657aca093a5f694e92de8c71c5e29093cd97bffd489f03f23dd3dec06c72cd812624082c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfc33b0e8f6efe5b5e3763d8ffff4b2c33ff6698a3af4633c5a58d0591a90c2c1356d67a4d08eebebc;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hae2d95ecb4df23b36ff5bf5eb9f6a511cf251e57055e3798f9ebc0d18dce205216840efd7aa05b05a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h749c5a5161f88525a50b19f61ff820ea710e2e09d7963ef2a7895c37da439f2293b606570d9be2b47;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h697892d960be14197ef2764007d71eb7ba9fc3e66f630c54237f0680201255d12197939ec4d82dc2e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h24aeaa36f8e0c662d52017b265374b26e9923641c73eef976616ec6062b9d9257749bd22a6de8e77d;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7358a22a198817eb9ac55d8ed7eb105bac0278f8c90c092bd72764397638eee833535811303770d4;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6809620a0b07b8e860a9a172bb5253b41509a4d3d96d5ac7870910aa59c66a471927fcf035e98bec8;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7ab25b90c86fc4c8a4eea4fe76569e4dbb3b9cb566bee1a896f510698f2a0e9617e157da1007a3eff;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf3d65033c59045be618ce9a2161f43f1b826ca6586b0794946ca56f7ec215f7e794d793375a688421;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h23237aa99fd3422c556af1b490447d86b31e4c5f1a5883a8228d4bd072b53560a63e12a0d1c6337d9;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc4543cacf42a9b40b031869e1fc13418f2e043a895863a45ff8bc91145633d9add4aca167904d79a5;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h44f9930ca89f1889bf9084f6631167fb0997bd0270155d88c5241a348f169dde3a9057a18c8a20820;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hee26153b0c533b6e9c7580af95f0dac8bde7b189a1148cc79b9ce073fe220258751cf98842fddb5a6;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h31453d5e754889a42c0037225558b4b7411e3d03686bb48e5460f1a7e2564e6b8547be1709af7a2ae;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha96e752a14951343625be3a5365e70f6a5de5c901ca7f0ef77c7ba644cfd84ceed4481db2c3592453;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbd61803fe3513b64d4445be6fe2b1d6564c9a85eba40fafe6cd32310fb65b76cf455d4d483ceca2d6;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h98a531bec7501012d55f92775688e734c12411d3f7aa7b0ffb50c2f364df0fa213d41fcdee6739534;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8fb13c3c09cb9cadd67ad05d0b041c024b5a39dee0a3450d7c7fc456bb22599d13792ae0c725c887b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd477f5b74c46c2a82da677dbac4e9d4474dfedee4d90f020ae1359894c74f0a1e0a9c644e0be9dfdf;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h66022746fc27cae9777ad0195d4446bbdaf731b11c1ecef01f18c25f9b5aa883d87ea0b5387bbbff5;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7e54587eac93826a153078138ff85625c150805b6a30c4e9b6c273c7b039de91b29ae9514ccafa677;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he5d028abca7e9b70fda3b62131d3233308d32afb9ba3a135ac107b807d75fff41bd45a05e72503e19;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8ac1962014ccbc263d527e545e7ab42f2bf0cfa9e6943bd321741984bd7926bb4333c477e955a41ff;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd7be4489f27ab7afc2f96105e9bffd54f73b064afe85fc3f2811027a1eadcbe0e0dc420d07fee996c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf45a57540de3dd0d6bb1717e36a60778c927d45bd7e9894792e797d52355935468b962a94225e76a1;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h20194a7a036ac25dd1c7191e76af6b24a1474875b6b4240eeb9d18eba2661ebfabb525afa5bc900b2;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7996b397bdcdc886f5afbb16bda7b9db3f98b9037c918a39161a93071d137614e5a5bccc8b3254fb2;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1ab71b29e46fada2c42d4ec93fe4b2f83ce440986c1ca0efcc61fa3f4cef3f1da1a91beaa47db74e1;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3c62f03b5524ecd44ad0b68fda7330430a7836ad264ef879e3514fb7024e4cef279d93c8c77d799fa;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6cf62c82524cf3279e59041883b2d5e05b573c53c75c7599353fe2ba5656ce00e6575c67223f8ba39;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9b8cfab573a654a5b6481f85ec8e1efc23e109dccdd94b2e2180493711e88680f5ff26e4d20fedab9;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6faaf9e5d34fb5f1e5c25e35f73ace6fc6306c391fb90e868eb1723ada9867b14a8419a6838ff41b8;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hdd95b303df362f65083e8da09725a8c5c110abd650387cd250c504b5fe4022b2103d835577db9a00c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4841663778125a66088a8b0ad6d70ac9448e08ec67648762beed724ae81a89f1257b9d156dc5b9f64;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb37aef5396ad26a37296c464b1cbc60e657d3d9d2a769149387d04581e0043fd92f77327b00506328;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf43f46bae295fc12e1af119d64dfc13337f4fe6dc4f635c16f0adb6f45b74b4c5b6ea0ab0b8edc1bb;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h564f98080fd0c70e0f958b0f2bae94780f906dc400ca31f5417cb25970030cc3b0a9040a47101eeeb;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3292fd29a78231b83c5f0d033a0a908fb8cc5abbe6798ffb5e07b47efa68b018c1af9d1a1b21dbb22;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb6e90946925902984c650f69af4a0bbdf184dff1fe993273dff2fb779e2727b08ce0b8de35e3f8e86;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf48a84a6b30cb4f2b942e3cf4c5ff7f25e9fa4dde3205db645b0f1253823a0213aec4e738cbb0c455;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he64c8a238fe13de7227c2f06b2df0081c2897d68c88ce8ad199a4fbf9e72c284a1f78ac4dc7cfd1ba;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h59bd9224749c4fa881b99af33132edad92d93c77b464289d15baa0d95a3678b5179d8934bc71bd2a2;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'habc9e1ef3c57f095a6f6cc0df48d875dfa2dcc56f3b24651d789438238208813a8a65b3fa86967fc6;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb29708d3c45e1e8825bf86f06279c93abe2f09db4aa9a66095995a7a06f9cfdf23925d0be2f792113;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha76b327b391174a8552f6f7733544a35a1f84dee5b29df3e59d69c57effdbdd516abdfb779cc79380;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3d87c0161cafe881386fe23e1928f36c2bcc1576b9d8309bf75b7a99094a6262d8d39c8b40c51e251;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd9bf49145cf2f6fab6fb2b044b76975566c62ec8f8e462cb146110e388e6b04e2181860a9cc185f33;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h15215727c1e4fe97579ff653d9c5b6595310c5490026f80e8d8a7bb111c5db39883f78cca031b2dd1;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9e0f3935f17e4fb0f074268c7617629a9c94ab26c51847b858e56a26d753648a572cab9d1601b3662;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd5d5934f36ffe337ef528788741016260f8888f05620ffc8f164246124d8fb1f6775ba417f61ceaea;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd00980bfe840efa85d81237a33c542173858f5f2a76da60a81fe01765da2c192e77ab0be43410fb9e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hccdf7012d437f26c473c3e4772577bf706c5c51197c1ab361a82b0953c0a8529d81c9eaa10c71e76e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h51e9bca20ee2209e5b72da2eb1ff32ab331cb15d3e9d0639917c39cd884753a431b3f4c4a24b39649;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7c2a55af2823450eb1f03335c5af375ea3c4e2d8ce54308d649ea76563cbb5052e7615df4c24e107f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8725374b86eb1e485ac399bf31aa0560870263f2e5cdf727c5aca5105904f97610f7f19513ebac69c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5a0e7fd62cf5187c2ca9ffac05253d0befd94c028c50600d55c21c8f34f9b6b798b4a0eb262b057a8;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd13ea709aa11c8a934fdf0c23b7e10c9df314444378de0c411033ec669db658ebd23a8a012276cfd1;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb518d3839808651130ee87ef03ad4a494c68e2fbf13c3126c6535140390a97dee6c380c9fe31da557;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he0097c531f9fb19a36720d09fb60ef5c24f34e6dd71c4808645290c6963cdd12cb12434697455a07f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb88c468efb0a7dc0557e60fb7470e147fba4681fc840c2c073f879eba8d6c18867addb7e0042a9425;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbf78bcdceced397953b89b7faa88a58e264482abc83bc146cf2442722cff7148569c0043cd785817a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3a0e71058296d3a2f6cc1ef8501b1378ac90e51a1363f85aa15ffe497abcf1689d264911cb951c72c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h97818da4cbbdbe4cb3a1a44fa71c7cbf5e380e594de6139062e65001dc35d2446e83830294ecb1483;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he82d130da7144a555fe1471ec76eea89cba9013a49719193d905c16e54129daffb3bf789132d4e334;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h15324da29ba867a64ee6aee4a6cbc05a5b4f686a971ce255c0086b137d35537a6bf864d3abd498781;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd11b360bccf2ec1c4b9c1444ffd72de52b2163570eaf0b8949f91ce54f62c60d0928a8eb4b0097fcb;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcd931a05f6e701562fdffefc2825009971ec4d074277b79a8d6eac3e8b40874f230c05c2ef39a1f60;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h49d3a6a5e8a4ba7b7605d346a3078703a6084080d5968e13950e39f4950454d523976d6c03f80fb36;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5717bd1402c1f8670053c1160aa0e9890704c51d460899711bd9757be9d748d3f28cd70a501a389a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hae5f5a5089fbcf6b516a47a871e68f795d6fabe00a05c06553e2f26409b425562f8f1ba1b20bd5c51;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4c1d90dfb68b53ef6aa8e8562e84bc8fd3cfec0d03e2bc67502cac4d13123029c81388fda2a937c0d;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9fed31891b0ed72bfe3cb0901e5419e1904f2baa797427b462bb336b40389a33bae6bc720ccab79f5;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h71dd7d011eb5f3fdaf72510c786ecf07a7b012427718d03f19a4b36b7e05412ac3f55bc3347327e3b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc01377c93ab942bcb779cf2f2be866dc22e185a477a92817cd4d5209ff322ba55f6867b5a12a12ae4;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5d986e0e1a89e0ab6d9d2ef39ba186de9cc4b2f4bf0f666900d47140bec18911565ae7da3743523a1;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h538daf2e538017391ebf175f60ab49900328d00ee41eee3336a5d0d3c004d1c4df4649e1d7ad15369;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hce3137eb65cc98ba4432b635e91827f712f5437fe292e53e8f8c7c2358ee563a31712fbeae09a7c5a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h43c0597a74a87938260ea30c9f6424fa1bcc94d2602fb8baefa0fbc3177c53ed2952473f87833d357;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h11c830aafeba814e1e5f08b2b73089f32b74e460b597c647de21e3ace26229b7f3d3065a685e62444;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4a31da24c7d817a34370b9672550bdc0b3671c42e314ac36ad191173230aa53bed735b6117957aa58;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9af09f217560a8310fb375bf89b51df6d0f99ea2092944d58beab283776a40b19e0a57cd948a3641a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h72dc1724da21a7abcebc27673aa1baa1a2e707a968b5911a0d125fc6ffdb52062d6e51768c6533882;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha8957deca1a75af0e076a07e9a5b17d7ac7f3edc3204ea1aad0d143e18de0041b0314ffab437118c6;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8517893630001a45134cb8fa812cc0a3ad8227dc9e7b26a1a605e2130e35cc628e34ad52d1f9cf72a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb10d0dd4c535e4c2ab430db875bda734752428b3d8855cb5f0fc7068f8646e68a8e9e30a8e08c0da7;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbbb32e5573df560baabbf45afc910f0a675a8e4b799bc84caea5ab9b32e91373d7fabdff47f7fe48b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hab487abfa9c2f13f6276f36a65891dfc36e7baf80bf12045b91f897629b04632165cadf53c41c0992;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb79a6a14bf80ee79f8c2e295c3e956fa8ba3567fc692129c1c5f89c5d338ebc403f9beff7fc011ad6;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd225d036a9e3b7187760e32cd7b84eee9e1ad16921fbcdccd80bb63a251c288b0f5ab7db7b9bfda3a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he36d2485b172e4fceccfd115cf26fdaefb71aa79bab77746a8f89d2598598d6d57c4fa7b53a28ab1e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h74e2b2ef613312a24bebbd5d277e29b658df96b4842374c26d6643821c0f313662b817a9f587d2e2f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd7246aa8df0a44efaf83108af758d4757e855f4e9d38ecd0b366c3f2ffd3c88c19e3b5792458d2164;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf59d47fb511aa2fa7777c5134893be364934ae8cb0361b18eee76b85ee5a8410b255214deca80561a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf8a989755c31d7097c30c2f45c10eebc22356afdf9b6c2b911c457fc84c0393a798746c7d3301148b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'had19f2b94a49ac615b1067bf42a9a3a8716fd3c876d972ecb9c23f9b048876254c2b8b90b501dbc85;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd3f72fc614ab45a48b94a3dfd152c1cf23ce21cbfc3ffb4e62fdab5522ef2dd4dc7448362c14fc654;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd8ab09daeefd2cda9c72f3ebf9514920d27aee07d937f7fcf8380db45b817aa57a10255b351516767;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6eb0f6a57f4b8822da9674a67f064c4b7f04f65b46a8a248062911b9359336ddc2f3ba57f8914f66;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h78e99ed1e3345d673706b96c4b5df03f63488e8afd796daf5b10340ff4ebcbdbbd9a861061748858c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb2bb3fefffde62bebfc054e1e3ee5ebd8553a3e6627b1b53190446708c830e6454738b975c53ba15;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he4fff718b8f3b001d5d2720203e0541a6da200152721273bf6193b8a1fad1273aaed1eee1c0e0ba4d;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he6243d7e03d9384f2f3814c5b08e438593abde9d8911e6e3dd28bc1eca85022f764eff265294ef051;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1099674259d67f8fd681b3051f41af56976b1dfaf91c0bc00e5addd92913d3c01c0d4dd91b3226475;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd0df92abce69840c5f792cc549a6c83be9be5df3040bbb9328e6147e06e40aeb8017370f1efebefaf;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha15d39a3caf30fdf73374f998f0bae3adb50b53d2329446368a973faf99f7c49c899cb47244545ee4;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf1c97dcfda5ec33175ffd6a20eca8b69f6f59e228936d666846efcf3d1ee0212c672f0879742c94c6;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hdce045fc87f49ac03b58c003cf265720c7b4fd085368c8d17f96f6b9acd895012906d89f702cc9d8f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4dd70e9bb0ac165bb6b738f60a136ed2e4d3eb35ebbe819043d115bd438b141c43f1e4f9ba6725ac8;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd0ebac700d420a91d345ea0b8c9bd802180033c9d57af91021392bcc82583ddc0c7628dff95d3d582;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1600d64022db0a4300b037541cd62ba247a9b3fa549f8ebf9635e4a1c0cdd585e744646c550e357a1;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he8d56a624cde984dc178d03888f3d77f7565dc07e0f826f02315614b43a0973fcef50628998c7ab0f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h562ec8e8c9c9ca922c25e76a1e349972256b1a1d334586339cb542f3144fa7bbd407446025a4bca78;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hea1c516ff29153c55b2bab7b3cec5e55d4661a411c222aa2e9c9f4146b3dd5cb23c805f883d37711f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h931bcafa5578f4b931ca3e709a9269ab4b9c189b0108a561194eb30e5defb13b0942abec9e540b083;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h97fad30bc0ebfce91ecb49113c9b821ef184211de5991c3ff55daf6a3ab1668a123d2b1f6922d9ea9;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hceaa2d21f68d4f29cde1fc39177b2436ad399ecd8407bcbf85b3d95693407fe1de1838a0d96841f4a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hff0ddceb27586dbc2306cd3f29a9db87236bd48c871182c562260e9ae21548afefddfe36cff4e14f7;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h80fb8764e75ce8cf5c91c88c787be9efce8deb388b092556b0209c0b03659415274a0ca236ce22277;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf645a4cc21cfae9f0f86868824ea914713e61417abf37a59dd470db26307561eca3652571051f870e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7c041eadf534e3506e960c0908fe197d8caca764729218fea9bd227e24412042b91ca9c39abfd4b6;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hac88296fd048bb3d56388db29e1b06d35e8e56f3e54c118ca169a96bc7cd8056db797a67d98e5fab2;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf78158cff766e7b7fc739ceb24912ca7618cc47587523851e8a5bf8d97b7fd55387b5daeac94aaba2;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8765ff719d763269982ffbe58096243fc110d7e7bd1222f3c9af63f7ff7e84c4f2947ed1e3b04a163;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h95e9dc49da64c21d8882b9712d37fdbdb37c18832fcbedfc0e6aca7cf0006beeebf7646eef4fa7ba6;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h57788d5101605d34ef70d3bea97b261f4cd9182e779fe6c0db34902ea8e5e279d05b45375b4716fb2;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hacb5eff0633391b5a6254ab69d1188700785769f509626426478dc28b626e22be90be0d1ac513b927;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf716e2d2481a899cf252881f249f8fb023ecebabdc0b6d9a59ebf13060ad22e456d0dacce3b11a8cf;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hed957632be0dcc7ac6700010d0b9e51708e5d75ad8e218fa03492a31bd6677a7d76e12e40e53186e6;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9a156daea040d666e9af11ae5db3e42db6908f54c656585e82cccc916ea79067104ea331ec1951799;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6d5d157ecd588950100ab23c414deb8bbac21868f40060df4ea04ecfb9dc3e25ac0fd7679fd8bc6b9;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb773fb98833712bef52ca35e8dbce6e2fb43a6dcfd6490d06fb1667177f0171b1bca76331efc664c8;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6daba0584db0809990cad0dadae893704483f439fff82df08320342d145e5dabac1287837e1e0af7;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h69d5405000ada1ec4df3d4677f40947b9cb0fceba655c95d10b11b5274e7c4df752877c7bd2390a4a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6bb178591cc7b7aaa9b5b39162e4eea3f5ea8818d4f1905a761440d0cdfc4546307234097d28120be;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2fc023d95c0126f55d43f612c6c25044bd805d0f0379e49e8538e07f4f3fed24e6df878165aac20ed;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h119bc54eff99f84afe7ef07b521a5922d2ba11dfe33f67f6662a2df0467abaa4e182ac37c9ebfb9b6;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2b265a62dca65f19c783754afbd515bbb3f1adbb9719f684cf54eb3ebbb667a3d266bf40fbb69e123;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h44729ec95edf0c941b97dfe5e108e81207d0b1a7e0df52500090faf438aefa623deb9c19b058cdec8;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h260158815f5f33baaa8022c49cd32dcb201e7045ee090989aa8275153f4e951dfba596731f444c4d3;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7122cd8da421852a6084e98d3e02bef1deabc19628cf40fe37124a35ade7aab31dfe9c0c136a8c7fd;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h74e30d61b7ceed4de98d9ef288475a7118d67e53998d79d3c58c68043e10e5ddfe1213ec28203cc7a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd2cc553365997d6da524ac0b4f33c18677ddde3af1be0717cef92e38a0ec8a780052389c799a9069c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf89805b1811cf31f5a5021dd58cf4c44d0c2099b73bdc9b97abcb6514c844ccd11b9b21da566223fd;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hff7fb561772f87aab9b411ba81501e71ecff80ff5d04baefbd8889b528c9547ef387c8b4466b615fb;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbd56a3e52975da86566e29f549281c8b45360e0ff96c483d489a34a421d7679460c50055f6a3fa667;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf01ceed56b0dd9260ca24a1e06ce8d44ebe1381c3eb62199da0cd839b541f04865b29c4ed96f72088;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h335456e0a61955d12c7085e7c766eea4f6b5073cfb9b4915e3293ceba62b4b460a7a9c875291db77c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3ef897f530fb10252e8e0ed960a761ebbb8fd57eaaa61bdb446dd4a6792218f13dd24ccdddd6ec360;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf231b61e88d3a016b4f8c02b6f6fa08f435854ca1824598e240187798ac33f32ecbb3917eff780f0e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf278b95e1c0de753475fbe4d9456e15ffab75c9e678da6962fdf4d1556db07e4c85695ff44fe95395;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h591a5107ad890acedf1af3520510bfc84f10e7ca1fbf24cca627f998f6a89a9489248db96de1bb871;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'heb7962904f56137b0fe79203916365ba896f1c09f1270c50bb5e59390c99d01bbad41b545513ea3a4;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hce700f57fcc423c153ba9d2afac88595def8aa1e7a29c278928fc655184078f1b30d48b4b395c8f91;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9bea0d638b360e5b12c76f130b78b687b583d2fc5149202e84ecedde49f43361910ec8f021c067002;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbedd63a22377d443e0156154491f05b3fdb651f62df08909277aa13c87ed33f3fa4a51ba260005843;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7af307c1f101c5055857b643eb38563cdbc63749312863f839adf673adc3617fde059a59325ecca39;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h551778d345a832be2bd710473b9a375627951ee7984e7f19dfa52434d5d0159fa6cd964886c13393f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb42d0ebc0e98f8e587ab4a52605df21420bf3208bdaca030811855fb0213f36e674a0b3ef4a65ada4;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd05a7d5ae489c8e59bbeaa7a5287a53a85ca6219ecd757629fb489e1ab5f402521832abc654797db2;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h286bd72f57ce9cbedd582932553f292829e4df66edf9a8be063dbf266131df26e2d3930d1ca52234b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcc8a7831eb43cd16bd96a208dd2af1853e1e267fca8def74badbaab5fbe2dd6e6e12049a85cc9c342;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6f25876d65eb70b2ec093ae4772721ef0b6257c8b1e6411e2e0f90d30bd986895854b73eb817387f2;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h331a675e64d6f9b0088bc26f578a98f09049267f6c2521951f4aacffc6fb66118431766924b5aa86b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb2366dddbdda70cead14bbf37f786cd9561f5d4c93a10a1c649179eb633d5e4c9062edbbe1818d5bf;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha2e877d6e0c536030c41395e4a13c75a4f6b70e5af1379d012cae6dfb016ccb2911e6dfe512454212;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h874acec64c13f6e428074efe198463384e4d0c654b6acfc5f19a0d36f2e9eb486c9a8940f5048d753;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hedc7dd2528ada0243ed4c113c480d2f4bacef1054c934f9e3f02ba89b8de28188c8a3edce1e72ac87;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb2b58be0b196f5ace15f17b1850a652c41c6a4877e0c863d422eb7438668047e167439e51449c5d5c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h91dddc1cbedbfa5f93ae73fa76759ee668ce815c8171e218d80f5b8b2670a4d54a3a8a5703ff1e379;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h570f715102e41e3736e206958ad68d798a5bca3b5b92420f0f1901ae695a6e664c4aca4d1f77c4415;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6d349997a434dcb9595be873eea366f0308048b938c24187d5e74594c8776f946dd9fbef3fb4b4bc9;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6f482405981fc0b2eaa6443f447a1d007c0eac3f60a78a25253f93caec0fe7ec6ef3a2300c4331cf5;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7b29a4fe2c3609fa62361fedaca10d302ac0b20d214f73c7504c111af88c34b53c932fc946c4bfdd6;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb77ff6c92a845bcc22bf366846ff8ab7c04ee05f95522126f53461d0c8f7ef5d6cb2af898708f06a6;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf0003af40ea111b9d576bcff7f2b03126ef69d86369dde934e7b580081db97a31487399da0edfbefe;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb1d3f35edfcc14556fab4f41233c7d87117b5f4a6048c1660553d35019d676ae4fbfaaa582e0a905d;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h711e8b4edc3f6505a6beb2c8015861002e88bebff09fe725edb15b734fc6fdf512d28f2e73022c4ff;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfe105903c51be4cea1e105f3b3b64b2828bdcefa2c61f81f194ec52e65c2e7875c89d0c751f43181a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h72a5e6b422ce23f43ac06af3df13de59593ed798a9960e361c491d751e61c51e4ac0a8057be218280;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfd72c0554b22a4663e78220a6d35febe1b387550afd46dcc8791ae6e1df7bbf539d9b537ae12b71c4;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hca6260c201d3635354248c4be18e377fee49319043dca25b524af791b00b7338f8d9e9d0c7f98e711;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h51fd18e08c0f9c42bfde1864c7d04cba12c2d63af2185aee13fde3cbe32a9fc8966a1c6f0099871f3;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5d66aec426e4dfddddc9d74f0c21415bcc98a42394f511261175edaedfddd9bcf7b6e4f8c40a04be;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8dce49cb7f99eba63de8928ec17d6e6e8a6c8ce5e2deea1d96f0edc000e66d4091862119f9943930a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h716e287c88291cb1983fd51d1d1bf892307574cc7d07f47776cb3c8b376f374db4c79a1031173547b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf7b366e590f55b7c60246c01915f36368c7ff0dd83ee3f880471b6af7e6e1e9df561c463754cc7081;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc2fa8b6df88f26700ac8fb9845363ff4dba57dd7cd08faeb776d0154f5fef6af408456cb3a17efd3e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h27bf6d25c7dbca56cc8a60cc3419adc4da0712d0fdf9226083ec713d10199ccfa31bf80b4f95b62cc;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7b3e8474759915ac8dcc521fc03c6ccece2d34c651e47d966ad06255ef38763f7a5812133f9341207;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcd049a662a19c411d85ddcdef00911a9037aaeedd47fec9e976a9c864204ae620d8abb9625a8f6232;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4985db6a97ec712dd2dc3e7bd4d02e3eda21fac54bc4d67eb12a1e139fda650301a34511726478498;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7bab67f7e32a0891958c3a18cb54b846f099d402e3ac34e1e6f3da5f3d181b42bb61580406d7cefb2;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4d99d312aa3de73df02e30878a471b2251643ef67ec0a7eea6b583038ca66ab310ca01c77b9eea0ca;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1af498d3a39ccaef02158c5edb79fdd2b5f0876d93de6c4032f2556d9047a70482d05df18184b5c35;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hff9cc2deff121014e9800c5a6f671c62772a6a9daa1a3ec80db60cef1aded611b7cdcdd5f39369cb4;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h723162234ebf90f48425581a16c78faa25b125b05036c1c02c9d165e129497262ade7e1a7e7bc7ce0;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6aec0ac6f851bee5cde8f4d6a130902bb05fd596e3dba5475c773c2386ab85da93b39125dc2664597;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb935210b8312d855a6b7eae2dfabbdfe90f55f0af6a54f6c082ec29274d0042624b98d3a5db920487;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h953f4b0ec6bef37ea6b3a9819d9c1fab68a50f56c45826e54bb58f662a276d1999c35f7ef3a31e1a4;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h835d7ae1e33a9a484fb5e603940ece59c183c0d10884664827d922761f01034130d608661e7b62bbe;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4fc3569b463173c5436bc04e6a92b55a6a63c9c109b24a1e325b3e9af884281b1795bfb4be4f5f3d5;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc98209d3f5e53f9dc066ffb0995de32adb29d2fc1d4f2e4ed65e82de674ffcaf6d399fce7b66603cd;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h729c8135210058d8af2029550692a33a1ffb9c9061eafca620347519fcefae34a7487a33a527f62a1;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd5c5a3f1fae20344e37f605307e62f0c0a9b6e89abda0cdb91a3e7d76f3a853ef0200b9e02dd956a4;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h17a1739c0c9b7e45bec0936258903cc7a6828f4393525ae2ab50bd154162a211741153c114ee093eb;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'haaad144cc7de9bae7b93a0845af45b254deb28ccbdefc6f4147cd5422fac76c66dda6670e03462b6e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6c6458d10aba7673b217224f6566b82bb906609fb51f93a148ab74b011c70a6fbf3b7301cb8727c84;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h58cd38a13bed5675d28361d67761117ad7600ceb99cbf94150f496cbf7bab4a2e628f299acdcf0450;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h616e02949bc73bd05ea1594cb5165b1f41192afd802a76e5e4d693443b875e25ccf542ab47e7e8da3;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd923534a0f469446defc6a8712c829d5e078bdc4e02a36ff8435f1769b5e5c660e288ba8d6cc05070;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3b8484f8c5e4791e492d94ee5dd501854d5a29adc38cea6fa52d98623420687d571a9cd71f4ffede5;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5c4a4f9db85ac58671317938d97618e0e8c3147c160db6c74680b2997adb6cc310d7e142912f6dd3a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h20c7a7d849b776c77364285d4fff56efca2b9337db15b89473670c5c2a84475c37a9aa8acc3783a45;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h767fa75150ce80b2957d045318c60a3465c83d39fb33491055afa724e07272ff00dc55cac0ea3cde7;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc0064b9797443c35e92b8da9d077fe68fa7b02f081910734ad0934a1dbfd63b375718554a18fa7d9b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hee64111339fb9fbdec27c1a854641d0d6fe865e59740a8f50fbdea0d3da2de4e45212c242bb0a9ce2;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc822c39e31e926fd687985d153ff62e6102e8f4cf6d91be2a78ecd117c2b2198543fce799053046a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcf7e8148376fd63c0bfcdb7f955b2f171bcd01424ea0f7d5c2461d68362f82cb568e28a31febedd44;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h384ce781c547080c47b8f8e7513fd5f28cfa5930ae926d5b7a2724cfd3409e5c45e814b50ef347169;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hdaa3eba0f5ae8d678ce33c6c43ee0af1a99bff7dc49e029cc68fed55d6abfb4984b7e8cc964bad0d3;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h60b53d66ca648628de8f9996953f75a8f6b57007bc9d7e3c517d36d9b7ec48375264dd4bea50121b8;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h19cb957b810cd3e388b4b95e3420f2181ace935d324ec3f1d0b896779a246ba78ae6b86e06569db9;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfe66c9d41a0b36d0663faf555ae47d06cf9293e6fe5ac3b324b0e8f1c0906330238b339a312f2b649;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h712dad4138013b92bfc1d46a0d1229846ffde5ae6adc202657e28b16a8a46d81f9914834853807bc2;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3176322c272c15c48b757955131aa467d8b0332b0fbf2e0c45d437ef9280d143609bbd61fbafadfed;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2c3a333f8e9f2e4b20de649da94674fa492d0ed85fbf2c39997509d0f77f4a977de1c1a58e3fe29b0;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h435dd1278ff4156bc8ebf0dac940c216ebae4a967061f0c81c521fa2cd8cb42812a02963bd118b5c1;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h29daf32abdf6e890e3a2604c22e76fd2d8b1736507256296045d515d6af1ba25d6bd5c4149ee05297;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he15146b0d0501ad92b570983b5147e9e35ff397f095d543f423165371b0022e4755914e3b434fa5cc;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6643f3d10cf89f8dc3cdb4dafb2aa9656bbd69608026eeb3ca02c2a621fe28e0eb1378db7aff20e17;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2e4768af6e776363cdd3f38a5dce3716f3ce0f10bba5f2d47cbc3d682e1c3a55122feb75382d4c45e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hea65b9c9a2c5c669ac892f943d16676443f906ae97cf7a1b123f773c29526c1029ae920db7334bb23;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h23563fab5b8c0643d10100a75cc929eacc80359fa81e30a0dd3bc8b2040cb2c2ddabb5736f585a33f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb138c76170e3f4d132f1c76f9505153de1db2225047062330cce203034cd5ac1e5c8d025cfd437bc8;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6842d05c747634fb5ee12ffb777c431420d2a7f9b4a59ba9be3a2211079c95f4c9745806b142c78cd;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h42e4e97bc33c10047a8539d4d3c2860bf08bd3a1a2c6aba7d616665a6418162f2906c9586fec03464;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5ac27259c2e3fcd9f775f168d92dd5889b8a25a021db96fb3bee9b3df31208dd21431af11ab0093da;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9aaeb4bc1cd42ed76315a616c1a5d953f63942af123a52c15698b82d5d11eae56bc72c7912c481c4b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6458d408e1775b22859a21e9694f40d5c9a22130cb14a12b4efa427db9d3f0a767a6fd4214819af6;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3ed6db8d0d3d1d21c6667219ffc81becf6ce29b4bb042e55a81a620f82cb492591fcd4dee78fdbee0;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc1049b93c7fde04317fd0fb8c189bd5026a1921212ecb4c0e9bf5d854181a28c0e0056071b44cb5fd;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h256172ac6b326cb3314ced72f6b121fab27947fa1feed8f803b2e202c4cc5261a6eccd1b470d755c3;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h92062c1433813daeb19bb554c5a7c747d3c6fb746e71650f95662c026c2027859e852df70beb0da08;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h18270bc028e3f60cee789316de249b71cd80d622ea456b121f02415779b53d62d2e5107c27d94fd61;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9acd5caeddfc0f0f98c9bd43e8ce043a3bc84ab246e1b38e69ebb2f1574035e41bac639634748ef11;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha362bfbde47b36349248a5ca5935176899d9efba98de4aae9bfde8e4851b605c200fa6ba27a5fcc44;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hac273149450feba1fb2d45f94ed1d1431f6d6d9f5df2a20dce818a873e401cbdf936cae9709d04fe9;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1d3320f90f58ef50df51ff54df279a3a87f405a071a2d7565a266b4f45da42d3f6625e864632d5559;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h242a58c5bd4e1c2035df5bea67528f95560567bd054e336ea1102bcf2f145ee6eef01fa4d0ed2db47;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1f6afa315958982fbf2d2eb6e605c4350cf1dd0ccb97c4c6dac5c0b0a0ccbd614cfdbdff6c9820ad9;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h14beda3955122a75b372f7771208a1a47b1ae66865b09426fe5d6d849ef708bad5a80b15a708b309;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h268b2a689b0e000b0dcd2d49afc214212afacc8ccad3e002a03a20ef7a019a7ffbcab4d18c5666956;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4da6375c4773e2c44e628103a26f65a5e175aa246d7849b162a0cb5cd5ec176012f2a69887b0d94bd;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf681567e4f588c2fe861f869c1e10d8d63129b92212e65461e40f1304222d745fe4cc3b0581737a2e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1bff1dbf9d275876e210565dd40ecc6ad70ca934f7283d64307064ac8a1a4c3765abb9df915e503cf;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h54f2a1338c5538beb2e210297e6281d810a5baaad876b09650f7b8f096b612901cf5ca4817a917f5d;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1a38391027a87d920fe8d28bb13e8a8c65de514024807f8ad44d1d64b5bdd683107368cb89a12f250;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h67183299f3d85fea0e621dab8dd8a5291a6227d0a612228bc3b750950f87c818050e742db91abe2d1;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5504f3014211a4a4d026bf53a3ce28339d40b51c308579cdd6afea0652b9c9d986d91f2695f79ac56;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8e4a44f8c71d0ccb66e7dc263400e7f901540bdcc02c5341a33b6595944bd38b8b29647523cd8c83d;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha981edb2a8b5f4420feb1a37ff11a5b00f8fafb353e193306642c536f0172ca49da127d84a9c74e56;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc5fc5a3f0c1af653c0d6510e2520e546bbfa63dac0a426737fb1c93c2fd531e95eb10c40d17372be0;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h75cda14c17062cc319f04ead727e65c060632a649be8a2957833266f135bcb8c34629bd153a64c6e1;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8631a9fbb1dcf7fd0b264cc80aafdfdabbb43510c16d98ef8382898eb211139a549cb44183ba2fb08;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h467b88336f7e70fcfaf6f69e7fa09c8817e46417fa1fe1b9cd33b925280cba6eabc7cc7dbb1a2998e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd189b8c1a88d26dd85f17a3b6aa681824d95217cd16e7d6609b247365a6a3be10a026425b249a5a3f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hac023682d97b5cde9b5f859145221f06620a110a8c3accfda8cca630efcda6419b2b42b059fd87768;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbe24ddedb0bcbb4d64b451b87c97a80e5d5cc1b8657047b6a3ec6a3dc2d1c07e9ed1d396628c72e43;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1c4a83061f6dae21f06febf8182dec8a0c3d014377ded2e15b9164757c5557f0e4d11865ab03cfcd6;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd5d489c505c57d99235a341af1d6b056062752a8dd21361d87cc6169c0d20784f00419a8848b8f0aa;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfd24ce9dd5b5e149b4975843356a3fb077d0a9356729e96c986786890c3f72e52bd2d71edc1a48d9d;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'heeb2d18f8d68ba3cf7a9d8d3f0457d8ca6134d87d291a2df5420ea14a00a3c84ebb0fe6765b89d3a7;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3e5bc41802f539dcc2472658d7c92803b2b943cbfd7118511b814bf40a4cf1225febc1a093f1d128d;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb64328e92e5cb960f320c7ce33bc4aca288c526a6bc0b0eaacfe025c3af801071b2b54654be79a9e5;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7bbfd3cd7a74eb0f2dc8e46e0517d3ccaa2585a448f76904bed76ef63d753a5d3c2bceb4c53c3bac;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hba18bb4c6b7ad8f3623feb7f0a97c4bcf24f05bee4d7e978a0ea30654b9981fe9a9a8cb2b427afad1;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h58735eaa1e0783bafdf167b1f18446b3c807d66cbd7a3b5dd9264ccaf38992d4c2613611756603df5;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb98dce7750a980a81f846385c47fd0844d83696924c0861ea5b3738b0646dfabaf2325faf51307ac2;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h530ac0916ab18fd839e2f6b2900872a0b04900dfd45765dc68604f1f3394cefe0beaaf36c79e39d01;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9a69d42efc4eb1bc943375c9241d04f5536197cd314ae5e77326633716cc4a1b57f7e6f222acfc5d9;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf7b60cb5f604c66ffecbb84ca4d419890cc9163642cb695da4a068d886a5056655a30cb2b1a177b21;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2ada193764852b8073471873b767f6bc4b0e62228ad63a40be548d088bafeb8c304abe938e9bbe0e4;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h822a42c9caf1110c79d13f444537650d315ba31903738df1d783a692f94702c3f9c468691bbcc3d02;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9fc4f450d16077d5ef83d7b80863e62cb2ff5a8d91bffc7cd539a206de96c2eb731582c53eded8b7e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h63e520690265205001f94a6f1e91830c21b76059cbf3f91ad997bad458d036cdc5bf9f5e026e7c941;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hdd22a92200c3a42f742e8cf8a180a60339dabdf6267cd0c5a18f8815cc9057ff23a3abdba2284b33f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h11028de590172f272c46601ad497041c5d38e6ef86a3a5789b38e012344c2b7d3bbb534e73c50f9c1;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h112fe6226bdd553b2de4523722f2d5591c69faa2a06ec8fff9fd011fee6df2e8b1537ee3e95d02c74;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5c072182af16f93b166893a1495bc2f8757161f2e6b1a687822e8fedbd634220be19c19cb5a154cb;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5dec36782b08b0f87a254a49561fdeaf26c34180f70975b1fb24cec6d46c8ed6efae99d609e06eaa;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3340a3366226221df4549f473cfb07c2e0f5711f1de425cb1288a3f2a9a2b7723ee46897a5d2ed86f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5991498c756987aff882dd88e3700dcb1f1943e7bab1dc47b321b386baf76dc3e608764e470389536;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2fbd220491f3f74b2b0f08fc60ed59d1b7c08baa5872ebf33e4dd913885987076571e58637cc551c7;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h86761030cf20b31a6afac952e21cfeef58f8c779ff2b8adb21fe6c7c9924f636e0506baaf1825dc1e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6d192be55bd7537a359e67ba2cef00490bf5fc46cf365cb936f98a3c12c84b2ef3b7687ce0e782bca;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbe96e4348b686028c590388577034256fddb9294a62b167f9fc696c24890ac2b42776d7aeb93aefc3;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he041f76dec96f39e48718321ba3078edb526d9f942753fd8b6c4b257bad20ed2bb3a6fc75939c6ea;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb5e2f8939d8f6f51c449d6fec379fa7c6a2d2320fd4745a5b75510174eda0f8285ecf1a3b65e0953c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8d7bfd21201494cd58e9be829873f1a3c66c96f2dbb6f41858e20d195f87530d1dfab786e3427b44d;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h401635bce7da78d31b124c6cdd553b3c35fb42870aec67fb882812cbae5fb60df766c4687aa60ba77;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd5580659bd91eda948dc4f31a86cc7ba1a519da2e7fb2a1ada1bdb220958e3088ec252c9a20af2206;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc35e2d720bb5665b376173a658040ff6978143ab6ea00c7b4c074be6f71f1eaccfc612631e85cadd;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3098fa399387d4579b4876c75802210657ade60fbf1c8ffca8411d30f4abbc766770dbee647dc049e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h58b38ed3c4a473a9e59fe6ce36fc14ce8b25cb15e958dfffb3aec99d2dbfd0154a006a3f0105c1008;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h84eff4a51c4c5df82f3677da571521807a059d3a056fe8ab3e642db55cee2da13f03b6e114524fa49;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4068ea66e11af15b1ae62ee5b8677e66a9b4c322f28a6d9bf015922a36942feb0b72c45680323be71;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h221c72d6fd5bf27322e3bff4d27b0df9f9274e20c114e406e96c2b465937c2e939e2822dfc493a9a3;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbb9ae099e033d226635a69c993a7f591fac4f197034bd6d5bf30bf97bf36ee701b444cbf5ae836b4b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h445000c5b21dece8a4bc5ef3518319b3f68d29fb87115b493be3bab964e82b81f867393a50cb83099;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfaba9d5bd15c03427e9923111c341f89dd2680c6f8000d3caf0e52a4eaf06dc141e06e8abae125650;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3ce81a11697dd7781ba57b4816153bed76e9e69266600e2cc3e03d404ce9854aa16632e8f4ff458dc;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2099452812685a0c05bf73233bec08d9d982f0024db8f9bbc85f5494a2e69ce785edee88ecc7f764d;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h114ee295bdd0910faafe94cba999c421a67b3b82082008b3049520fea2ae095e7a6e23993c682b952;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h810754b54fa4285e5674831dac7be511fee9a23cd0bd210a537dfdf68c7d53b929108737397f220f7;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6ca610a685b16ea5d9103d015524f3b1e78a571c15a3edc1dc2168fd56dcd9ad0f9b877617bd63481;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h65836f76a3b3c85e2195808800ec5aa3076f9f2c7d1afb5c7b83c31c9494e17db8f7ab85910c9c0b0;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbe090729089ee8986a9c3682e639582fd084f101ae227dcd7d3f586574236d2c0d5718ca711421ab3;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2007749e16c64a31c1f02ea5f7c08fa85023489c94cc9aabba1037cb9c8728a9d05b03fd3ec9f11af;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfd06eb7d90184c369f5bc0906c78be1ace40d7acc1644d690179ec3c7bda08daafbd8d7291471c2d;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h70bb9287e975f39a907282f9bb7caf1e98e1e8a818a22c88ea2016ea4d76620e062e0cd2cf406e507;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha39e44256c8d3bbe3f575e5ea970bb78a24572576b871f090017a1f85f7dda6b919310cf0d9ee5d4c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4e04b84d51a4b0cab7debdd80d8b5e1561042d87c124157f694a49f106325d2eb247cf26fb8b382de;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9addb2dba3fdf7fb134afed534c0bf4043c1c587e354cd6896dc8b449abf8d258460cb713cd65da92;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb19ead5ec3ac688b762128ea62880e7a5671cced47c71a0ee5df1fda5705c3475a7768d9a4e240b0b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc71277d03968f912d8aadd71535e585baa7dd35ba8dd8680e9b818240d37f32db5919d81aa65d8c65;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4d685f2261f4a8bff945a5775f8fd6670b51f81f8bf498b3a8a882da3918e864900d228e2d73b3466;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8491d9e1ab387339f7d09f2db34236a4524020217df59279795966065991b6e38445a9c578d4f169a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he707c91ff3951da344cbc7f38abc4f298f176884669a2258a704b97b4b83afeb7ad216ed8760a2123;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hdf50ade5c577579abda16a073b2455aca22faf1185c80a45a9edfa1ec9504980ca2ae0859e8bb17da;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb69671853f62b39b45a523622b0a7a041ab0fb7c3e05dc2632d8d03b0b1265b95b6a14573a9384f2d;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h39146fc550637ade550deb18110c72e70e9bfec150ec502a6489e1fc09f5300606ef14dc10f4671bf;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5805b11e3cee6f0e1743348d453bca1eb1a88e30812377758927fea46cd7a932cd934be966daf3d97;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7aaf33683aa491390d446666abcb43ffbbbecd14fa4b8d20b396c60360fcfb91cdfd20707b69fc10b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hce780fab1b4f82813672d1a111f6d2d112e69902f05070eb890217e5eb8f163ed71ead8a98d80d366;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9d2a8b54a0c562f8d1acc34c36b82a317c6711cfe0463060c5e1deba03dcbfcf016629fe5aafd43ed;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7d94821be01f0cc7465e708ef0dbdda5046a159dee661d0ca2b770b14a49c05e1fde3c9f0f80f48e3;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf424a165aad10655f38825d48e6947cb8e71213e0f947e6ef3465fc0ae1db4493c9728db328a24dd3;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h640d70c947ac2079d96a054b3c3a7db48a6f6ebf3bfdee172195e64d069bed4c96beda9e6df1d46df;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8164c46c71e200f5c508a5cd8f8ae0442c67e16baa605e907f31c09d6f21c328a5ca3811014b01539;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6ccc3fba268506cbc75d917e193c1d624b9962bbcbf052b245544c0cd82503e8c066d78ade6aeb2f7;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb49ff676283fdb5f996332b34caa290028bb3f4d829188cbb9fadb4b4f09bcc50d568978ff6d3057b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h680b308129354ce5d29fb12de52ca0a01c07c1522261d2bf308d22332fabe95b51c44fc4766f4c0d8;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h43314e85fe2ce1177ab6922ef2226102c2e8b5b469768a25a42aaa0b5953f564889f9b867017b9a79;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4d4f29be69cf5f8074791708c016147c06953cd048989f6e98bd77aa23080d33ab5d5c300e3158fdf;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha00609dc3b47e3ea583687d70efb7ffb7bc0cf8138e405f9775b1a4dee2499730ad7392c21042bd02;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbe21d91f8301897d3228693dbfc4f29514a232739fec4d4cd09c2aaadb64b5374def4fd86abb325e7;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h15d40308f0289e53c554f539bc23e8b17a8d8ef4b41114f5becf22c934f85284541ca41124b16bacd;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2925a430b6afbeb56690f4032187c1fec9a072259070e295a581631fe1e4079274fc4992c6417d9d9;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc7e4df0bd89e9c44496d773e4488efca37e9be57f45af6d386e6370a6098d5822a44298305d786dbe;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd9f824fae2826f37505405a49ba9556f1ea6dc47dd8fbc21480bf570ca5c2f2f78523519e008774b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2db271009706d4495ab214b6dbaf861655e621094feb6dab98692729f0be88804b6f63168f6950bfc;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5970b65acaf1520defd7d66335dca196779251978c97c38e2d0e0e352bb609e38790c6cac20eb29a5;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h74e9e382798c97f65711c6107f219b3fb23041dc59af8f09cf331b827ac1005e4232b8bf5b137c749;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h863c27f635344476284ba0dc6baf7b9855def8d23b3f5ba9fe510cdd8ca3e9e3f98e981b2f96ad00a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha6666efae50725920f4f0b9b39a16b81e4eb201e91180046c7368391b5844095ebe53b16a84a12e40;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb0dc71445ac8c221e45c842eea4022b67e83a8bd6284d45e3185755ceb662e9a061319da09d8aeaa3;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha5d6950d1c723057fce1f4d9ed8beb5338c4d3160af83334b13f0477da747b68fcbef8c10027bfee0;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6ec765f2fbad490778022ef630619204579418fad93d5418cfce752d2d6acc39f228caab8a7db607d;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h80cd22ab25fa0d0fd7bf8222bf9b1d181d23a59f1149e2ea595f846c20c9c4802f074c5b9914878e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h419452ff01615d25dd5cbf4c4dae7c0ada85ccc761b08359ade547614c8a30d5f28598d807f04f420;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc8e03a8d3f99842aa7c52a77db9cdfd3b6672dd941b9091420f3cdef9226170d78600ab517f99c8f2;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h107297c03a60a19058acdd84fdacf64aa245f1c72d786005693b4e54e4d460536dd7fc1f527b33fa7;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcf625868fdc922c6964dd2aaa4e8c8c49f279dc513751838fb3acc6842587ce1bc14f6291246a4c98;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h37e097b62a170b01afa02c9c96505041b9cf07478a10464aac4102978ce25966bab5979f9d4e52476;
        #1
        $finish();
    end
endmodule
