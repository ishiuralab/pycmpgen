module testbench();
    reg [0:0] src0;
    reg [1:0] src1;
    reg [2:0] src2;
    reg [3:0] src3;
    reg [4:0] src4;
    reg [5:0] src5;
    reg [6:0] src6;
    reg [7:0] src7;
    reg [8:0] src8;
    reg [9:0] src9;
    reg [10:0] src10;
    reg [11:0] src11;
    reg [10:0] src12;
    reg [9:0] src13;
    reg [8:0] src14;
    reg [7:0] src15;
    reg [6:0] src16;
    reg [5:0] src17;
    reg [4:0] src18;
    reg [3:0] src19;
    reg [2:0] src20;
    reg [1:0] src21;
    reg [0:0] src22;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [23:0] srcsum;
    wire [23:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23));
    assign srcsum = ((src0[0])<<0) + ((src1[0] + src1[1])<<1) + ((src2[0] + src2[1] + src2[2])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3])<<19) + ((src20[0] + src20[1] + src20[2])<<20) + ((src21[0] + src21[1])<<21) + ((src22[0])<<22);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hffffffffffffffffffffffffffffffffffff;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h28e9c6bc671a46f24db5b08b34804c4df040;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h459385bd45ab1b1c9163f06fae05a19b12a9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2bc7f8072f3a7d0c7483a56968782521e9a4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd2061b6af842e9ea07be4d9cf7078fd83827;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf2c9de9c74ed79dc84e7ce8e799a8aeb5c1c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc38813d9317b25a3272cb12ea4a20ae16cda;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hfe8d49cf5ed9693f75416a0ec025aa396561;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf2cfef58dce3ad2d673a9f198ee84e2bec8e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4c02a65180bdd76276fda4992cb156d00ce6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h84585d8a00c6f9f40e9db66ddc2e86a8aad2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7b92908d4a8ebdbf06733acdf7eb80d857b5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h30f0c58fd4939305d111978e13cd826baeae;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7f8542f6f553a27eac7678591bb1e05cda66;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h43e0d90da9c3221bc9b110c5585556d5c297;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'haa92e2cb34873a24e8a87b4e46924c9418ef;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h148d16993d98b957fd066967d19e983d88c8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h11fe64c85e61d377c621d7976281f7b54fad;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hcb5f95734dcf8728a160b8eb23c4c3a0a03;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf554bcede5aba8ee74b2a291c020b35c8b4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd9f351fd2f075473a66b14357d65f7756782;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2dc6329a648f36060f7ca7f12bc7f6d2b7e9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3568a7cb99d0f9e4ba051c95176f99502d2e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h99496112fd5109907e167e0139dc82022ea9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9c89e53d308e3a256bb540a8bc68a78b1c9e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hcdee38d42f50ac787522878ef420aa91c993;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h31461d964d037d7e0bed11358daecf4d9f17;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5145b14526a2298157b1cc9968a3a92c4353;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc4332b4e31b43fe8297ba0c5068aa9ba0fd1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h60e93df86dccec55c35f0d5c33d4288789f0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h123f529e7df452d83ff2b7a3abe5e61771a3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h41ba916ba0609a95b784e5ed3fa39dbafc84;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1c1facb8cef0a9c67eb188e88111d1bc4f30;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h670f55f85de8c1f0838a09cdfce89a4a946d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc1532d1ccaad02497a0f32f6c1742361789f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hadf4250506be25fb2428a3f3498ac155cbc4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h52afd9b1b837f36cc7f625399cf94a3564cc;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7e418dca88ad9fe20bb7b01ce12041bf8914;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7af222e8dcd62a31befb1add50dc51525257;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hda612b17f5769e2e60fbfe6d308074c38da;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h34af3fe78f687b67e081e544df2cb2201976;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf96861f326bcd3e699b1b970e85077f3b738;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h918766ddd14da462f5f7c55ab4ecfe1362c5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd6ef95e48e95f417a9990d573cf63da262e1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7964e87fe1c454cce5e91ebaf114e13d77fd;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hadd0976efee0e6690f1714f2707899f15f9f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hfb2e0fd61c14353cb3e3c689302144e6333;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd8fd08b076dd2b8cb498d1638dafd149f6da;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4c12bd17c908396cd3c49a1356a08acb03f2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9093e890c355178433d89ce6c00bb88ac4a1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf3449e67c29061fc907d08dbbfb48e5182a8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h37ab053251fcb84decd97ae7caffd4589bc2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd8f49d935b3f15ae8e0a7e0f95976b4dfae7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf7ecabd7c6b05e1c4796761a60b3eb0c69c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9c4f8e33305c2b8d41f4dc586ff55df5beaf;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h31270cf6f538419d7bf0c788b4a1861a4838;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5e78d77e09affe8c55f4a915b8c95c252085;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'had5f4c8adf6d3dc77d95f59457ab2c7385c7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd0f32eb149a8407740616fe8a6d0dff65347;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb91c01b6e42b6d4dcd3f226ce1b7af93df81;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf00cc6b2bfd8a5371395b370ff80601391a8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc9281659b544290e8ccc2868451e5f090b1c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8812815ae1fae172f4f43c5bd5d753e1b68e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h42dcbde8ecb7f9329d8df2b57006cdf8c238;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h57b026a082458cf832d7da4a15e21aa7d627;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbec10f63a8e6c12da029341b035f7e198163;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hdd8fa11db265f477a53bd6150f937e5a7764;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd8f94731b210b1979f34d9a922be2a4f8f88;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9dcacb9cde3e9acda99a7b07f741b1a9e8d0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6d437649e38e9d3ec973a077c4aaf00ea960;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9c3154dfe7246f7fc719a8a575356118a0cb;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5d437bb66623fce2ee56f83b5224293a5777;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8f1f3efe3ecf1f5e179933545cd050c2ed2c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hfa3a2a9e0cdb8f8bcc5b1bdf1b599a843ee0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6fee61d7b95632e93b9d491a65b26f85fca6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h556b1c38885b345b1f96c7b8d2dffd97e1cc;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h87e8d2c517853240117b0f8865085175ee6f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6e31a9479aa9a9a3b2f9ccaf2b99326f84;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he693bb023f16dd05180958f0e3f09638caa3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd9b0786653597916ece5af3e42b3e2bf87ed;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he8614ee2e701c58b9b6e124fbc62dfa8f335;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc56205063aed0d5b5ad55027b6c03b5849f4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbc2f83b383b2e20612cdf62a1b6660552627;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h59c3a76d59a7d7a2dcdb59e3836f21272514;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd92d8f0d7a51bc94f7be4e527a183dab2468;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5435c67237011eefbf3b788a9e42ee7091af;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7bcfda6d60c44602dca54b460e4ad0f4e70e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2105ac010038ecf89a62c98c399ff27b81fb;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h67ff0ddcf4f40c34eff60ba460e60c0287df;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h98d3dc6f68598150f6242e04c1401b2c7a4f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h643adeea7ba6356c6ecfd6769946e03e6e54;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h633c043007313a6391ecc391dc9fd5119ad4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbff8d8fdb5335a7aa94ffe89cbc2472d88ad;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc01edb18ca339215da5664ceacb7f9d0256e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb38fb37749f12aad90b7bb2f23af7d02fb3c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6a4021d2e86120201fee6841c0d772bbd8d2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hcc165be62efbd47c4890d564abaf3e204701;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6b9f657b6d6b80f456e2f0eddb8daeb5b189;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h610ab1afd05a56372cd8532db9574c258098;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5118142242015584a8095f9c54cb035dd23;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he3e83a81e1720db4e287ca9cba75debfe899;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9b6d86c495dc3c61776555bb324b73079b7b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hce3598db273213f3722b9d5e84c268cda0e2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h60e6f39dd7badc10332bdd1304413fa29ea6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1920050065116eca889fdfdd34abbf976efa;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h51c5aac9896d8f061799fadc707fc2f8796c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf06463262e484562630c0479e6a3ae209c37;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd9617e86d0c3c85b26488a4b2ed6b0eddd26;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hfc35add246eba0f4fdae29d6c113c78bfead;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1e1a09ce173f98b6a24e0f55c30c0f2b0e74;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he6f4cea38b89d4ce1524d9c1db8577654ce5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h41e5523198f690590eae7263dd25c50e24aa;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbe505d2e1f454264c6fa1547f3a2460e122e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf1bc81c8317e0ea9d5cf529f8a2ab8187857;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hccee200a53dfade8b0095f0873ba599b4009;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb0ba7232960dd3a13ba0c30ed439506a3e96;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he105b3524817016a42d3622d2c30fff0ed1f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf3e2d59e25d99ab76542066fbacc7f86525e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5c267e97684df6fb8ec7e5cde19ee81c4bf9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'heb1263882aba9e42a2d80ad1e420ee848d7c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3b680b84fb87184525abbd8bd3076ebfd0a9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h943b1019e586668a19f13c9bc657bd426c4d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h489632c0e914cff96304d09f793daf150ec4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h47093ca85e751cc509cf8d447b013770751;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1473feaf2880f90668d3bcd32b941ef42c8e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h902abe87f9ce9983d97e280cee7f34d50125;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h60657f9d0d60646a393a3774b9b9dca45825;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h50a9e6a32454840048f86dab17cdcdae7b7f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2ba4aea26b81df96a521fdb559fec69f23f6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7aa2d28ad0c694698f1e4028f7635e13825f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6626e2c31923f51883338598c53f2e7662c2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h580ddf9c1cde07e97e1dce628c9d59bb831e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6a9947f4759edb68078cfee29dda9976e0f2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hcd387df1cff3836af03ac35b91f34694c79d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h864e40c8072ee4095c8b55ffd2da7bdb5f70;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha97697a9ed90f8801be73a8b2afe833846a3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1f4b30020b14e76964a523dd67811b02497e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc0ff69a52e9a500cfcdbb569459d60058ad9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hede1176229d291303322d562302e56d1ccb3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7de44d79ad50f41408d42501d873849b4b37;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5b6888a7e53c89f162ad9e82f8e5c13c2f23;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h74d780af6f911ce1944a90a3c871b863ec24;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1836f13f72333f5035c850010cf7fe37ca18;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf902bd1372b2fbc9e231b62c1113071e881e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2d9500db223fcc7824ec8c1381c54516b1a7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h72a9bba612b905c23dd2df1d115b0fdf1586;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he98f336cf0e251a934085451d9fc86e76703;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h70f01b66b29c9cf1a0f888fe4ea37031c1b7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h337e4d0c263dbaa559b362e431bbafe7c40;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h46e9dd66c2b44ceba460b55c575936380b26;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h46a3de92929b293f90c5ade1f7bd6b4799cb;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha1037eb59e82929d8a5a8a0a54199505cc20;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1ac6eb99ef8b245ff8c278b2c0eb69e83367;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h13965de756924f0b0761ace422be64359d37;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h587d2e5c5254d99bad9e1a5b0711d9db1e44;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h96cf23b9f9b6f49c01af8fd75d971c8ca107;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd3099e9b76775196bc314ed3767aad9f0be;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf098c2f325cc14d2c7f02c9649cdbe6be5f7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd18f038c54f0b314a86858eb13a5d7b63931;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he4225668c802ac6e8512f0442415ce7e83bd;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4bfda652acad596955e367feb3f495e4eb20;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1a5a073754846b58d9b0949f16d7e6a29f1e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf8abdc9473801d319bbcfa8dca5deec90458;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb6e9f45c77a15dac53c28f78c3208c39ad3d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd0511989e0ceb8f478ae0178c5fce2a10e4a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2754acd49da0c697eff70562c6f974451417;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hfb4eb9bfc85ba236193fdc443c1bc5bc6da6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h71aa9c59d27d8ab520cba0bd01ffa21d8fad;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3f34f7bb259f90c6caca0c0d346956075114;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc2fdbb8b3ed00126457f65863a459ec9c6bf;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5d0174dc649ac8773f3d52f591e343be5c2f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha00ac173617f8ac73eafc2f7b9d2789f00af;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hcc6663e147806d4fef2ba66ec1f00368da86;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc4e3b1db8109f6b2cc872a6173fe89d794ed;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h21a5bc6b24824d7f46a1a89b5501c9fe938b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd3048dbfd7b19155ecc62b6817f9c359e00a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc09e91cb4ab3e3144de7b3bec98f754eac9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb1125011729f53cf9ad296f7a883bf43c8d1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb748ed6468173eeba4c3e620cb78e5e95851;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h22a30f87898b39a222713c3acc19c3bbe2f4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha69889556c9516f59c01772ff31c8a75fb2d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hdc9e9fa95de201ae1bb15038141c1e640250;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hfce427d87d234c460616962fd83036434aa7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h131a8d607f92b16e7ddba7e92e7c27daa0b8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9a425f2413d6e6a5b09fae821e96976619e1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha461468e2f93102b68e57089c91861025c41;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h707934316093bec3e66384323e95d969415c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbe1536e97b4ce05b79439921a5b474131c87;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd34162ae5b9a5db9fb6ec5689b5892350f6e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h38329c028a195d5ec11061c671133bafa0bb;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd0600e7b90f1596d95d4be2aa9eb13947f72;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5426ca537274001051ba7b72db2315b9ca10;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8479835bbbf207b2a4d2b9beed27e53431e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3b77c048a61c54395c6e85e262e1fcf74663;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1ba43d7b5f28a4fd5ad75c674af63d376244;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h406bff6b2e91814c2137c3762f1ee9e8b153;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h20380185df79fc69f644b7f0cb332279e144;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hef352e587499546d0bdf00e9c41a32a16b6e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h273787e3226f11a82cc9592d3eebedf38557;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2d0c6a1a5d503b6349ea4dfe3a6f725680cb;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7efabce07e7bfde2ac6807c82c76d8d009bc;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf33a1d99fbbefd5de292a813125931d6fd0c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb47f847913aae7d566b1c4fcb3fa9c211af4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h759766b62eb895098962051e7daa53be6a7a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5597de69207c74867284eacaef19c9d29f9b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h697086d986714ac9bbc54ceed51d7bdb743e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h19048a4395faf6c7f479394d7e71d7d83034;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4c0e03f8cc5b8d79ea7e098da6f72a2d931b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'heb958f04bea8234386a834a0b29f2e55738;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h29cc53426c9698d86574a326eb4777b09142;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h606ec2a806815812142dff8c1a41a76858e6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha2f5e9868f0226ccfd8cad5281194e001296;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h94cf22bafc8557aaa5baad4b899fae75ed98;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h77d916b164d22c323e59faf9507f144e97d4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'haef1166f0f6ed1f9301258bd49a6e9b9ed5e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb5c0e747873b320ee8d9f624c4ece31f7800;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h20b47cb8e568d1f6bdcb5be1e9439c1a0bcd;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1bb2ee4d762ad94c8cbae16abccdd60e638a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he155a4c0ecce21b4f4a1853afa3564d7c076;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h27b1660d12ee82f44a0c54a052c0cc7a65fe;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2813d8d9490876b62b7961bfdd8e8d06472b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5662d41a36d00b433c3edf9934af4d74d3e9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5bb6aa15f07a76808b70e68612a9ad20cac2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6603becdfcc4b5d73b944b6ecc8c3a8574f8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5ee0814f39fa5cdb6ec26c02398bd0d24e0b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h650295b70c49e6310602216005d3729be5e4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2b4a219ba00698c60383e7e5f06d9085902a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h70aba6c6644bb4871360efb0a4f0596e32e4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'haef96e53a611b7305a4b1cbdb9b7250325fa;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8227ec8be95d6e4dc4f5da30a215ea8b6477;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he28fbfb72b0d90a71fa7784efb8e222ad141;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he2a7fe4a65b2faa65b23b8aaca25616e123a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hebc47fd961cffd365eda05120d87e1357d0d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he5b1f5210160253e917faf32aa991e870f85;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hed9058f54b7e1176358a34d9a307e91edcf6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1ddb9dfbcea077da62cc557661b7bb03172c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5c3651f2961d68ae3a9172758486ab7d7e28;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he80b0260affc562c5d5faaf5625263126b09;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2ac9e16aeb2d76b5039e941a320dc61f9a62;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hce8b26a4e8387e25080da292b11354ce9cd0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hcab51d14ab9c81376d1c19087ddd5e6e7fc5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5d6d1f23380ea720a7c6b1f83c6c222f53f6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha123cb33a58a8e5b4bb74b8d74be7d1f8d28;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2738cef283a697befc8dfce1e712b727716f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2b7c6d57b22115253fccf983292ecc6a00ec;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hed35ed57143960883562a40ba462f2fdad27;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6aa0a613e309a037ef83a45d259e99c99b17;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd6bfdbb84d15b509b08a2817d5ec02b5a37;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2f830e0d85063f69d637713107278744d494;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hdefbbd81d40706159ae0564b1b9705298f67;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha203349a0fde4f9fadafb15c2ea5a7e9484e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h681d9f8cfc29c0670c045dd62fffc0dd5dd4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h77c4973ded44263ef68960b481680da007af;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hca15e5b0e947a33af9f3444641ec9963fd2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1aba5cd99bad9f93410bb929807c2ab16c86;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1bd676b07ce32b1d64d625cc153d83964ce1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hfd482d44c95c497113205ad02782b891352f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc9e1c2c86e7eb77b9bfb00227bd91037b5d3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hab7135e12dfa15bbc4c2a77d0a50cb72dc38;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf81e4b5af1fe0e03690067f6fc92823567b5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h630d0d65539ab7edae8a2a398dc0cf5f2e21;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha9c6ffafb4e79127856753dff00f002ca1e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6e3ad302090ac5bd3da0d252077f148a7be9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd5f7b990e1287d8dc50c3fc8c8d03c45e63d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8953511d9268e5dc5df04a0347b1d70a93ef;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h702723c9a88cbad8b59a78157a8bfd7394d5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9bb0fbc05f228ace1812a49ab1a7ae9a58e7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb88fc32e8f1b1f67d29d12ff6703edaf19de;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2651dbc7de170fcf5201d0decee1d5b3f407;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h10f0ddc523de7dc854d5090653f5a286b4e3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9391f4acf3bc9d80d4c145e7e7709b2654e1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf960983aa86707fb79d245b3381cd12ade7c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hecd78d350030c3ecc8a7afe1309496a5920c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb2ee02efb53f97a2a62dd43c7ea0064419fa;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he742e4a805370a796919cacb5ab5b6397e75;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1d6e6406849cb76027421e8fd81452276a16;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h120162342a7458655d521e0a083f76708f42;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9b351fd72feab99ea4a7f6c263e4bd8d31e2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h689090418c2554b1d15338157238c22c060f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd4927965a5e97fc21e038ce7d5749f019a69;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h66f9c19d920fd9b4ded12043aaaa3b812e6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h606b0f105198ea11ca4af49e8c4800e8e87;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf5beaaf736dafc2643ef1167f0e2167a4e0e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf62ad1a1d1e42b291f70b836be86c6722369;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'heed33ee6d1389bb8d2264c980a2c442709f8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h573c20d6eb2bc8b17c919247f2acd1f8694f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1128ac58e55b92217db59a3e55913420939b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h60110016e8f7fe2605cd8f8174f84962546d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h589fd37bd83c3e807511fa5614f3672e81aa;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h30f01a118bfb0864cebe434e9f3d21164aa7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h57f38277014c5b2f33caf52b06435d23debd;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2d52da7f6e3b654c46cd40bcdfe6f000041c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6a721e6619d9d39c475e8d7d391268fb08f1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hdbbdf3ce647c16b821260cc089526fe11eb8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h10b7df9d3742d51eea6e2a064d39deab681b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h839d42ee82cb079ff2d99b0c75a10b956cd7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5a3d1a6ba3052464e5c6829130caa6b7e9e2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5402700dab55272a0a09bf8d4a5ccc2be90b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf45e5f2abe8bb80f80d869ac9db55a1359f1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h98b4a7456a3f628295f56efdfbb5de93da17;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2270553613f1ebc6789d710a9dfb0a11ce0f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h445eea758472491de5cebe3800f5ab979783;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd5762765f237fe91427cd324f0d6026c7868;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6aa232f6a97b6f034bee8ce4e053bb51e768;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2caf441110409a8e253cb42ff0fb7c65fdb1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h81d25500352852533b35dff01b386039e50e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h60f383b06ab24c6a5b7d8e766fc965a268b7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7fc71cb59c44c0ae4c7515bb47c34413f383;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3b334e37e4d1ad671f9fef128f8df0066c3b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf1bd0397c9a79152892361962f0773fecc81;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hca0d6a4adec5d206c2c58f0071bbbf9fa4be;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd4b420d5c0d9f09d31636e23382a8f6245ed;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2985a0bd741b4b3b2826c1db32db8e4fa8f5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha2d1eb93bb958ce04309359b2c754e869b7f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h25d6dee7106e38eb94e69980e2b775b00b15;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h548b57d31b8bb93f689d6f31b2d345fe457f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7141f1b56b3a9909e2ce4b8314cc9a99d451;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb05e7023c82bbd62dac27f9675cbcfa8caea;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb95bbdfcb785630452bd4257e9fb932ad31a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha10a0c11ee4c7c523f3374668aa160a3016;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2467999254599d669e09bb169e262d33ce90;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hce49c6386f4745777b6e310048563222e99;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h430cd983cc6d11540809d97a3e00ffe02b41;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3b31c12a4b1f8537f68483955711934a004a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1ffde7899d2340d3c4f48e4b32e1961461d7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1dae0f15b7fee7125b3e28024d2bf706872c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2b71882d89c9a8757c7653d87b22024087fc;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha59a2ce562716106b153cfde47b09bd4feab;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h408a65b5d02280d58ea603ee4a92c0a112af;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h908f82057b8752820c1703b52bfa74142e36;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5a467e90186a01eea0b4d61df62d41f2f230;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd6efdab67bb4687fbfc4fd6f344db5aef487;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hcd0008eca943a6fc83ec50c38f48dc8b4f1f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2c62a4ae366c8085eeedebd7f110990281e9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf5eeebf54bc870122a5f20b983a91441153e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h65f60c2eac74250c03a2d347d4882e359204;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd9b52fe83a101d3a1496798612be18c397e3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha292c8c9162769d52d135f12b67558598829;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf31f893089efc55be5b382115a99158b96c1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha36e126eb0521e925fca76d13b329065429c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8bb12774ad2a7f8bd309e258c52335fa5032;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc81344ef075ef817ebcba57d7b3b460d69a6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4435dd315f155744e4bbb316c4c2f4cc4103;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7f130363da8b6f5ff0ae1b07cad3dd86ba2b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h601ec451c5187d2dfd9807960bd09dbbcfce;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3e678334afeae623fcc23c7a32288e47d253;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h538f0391e3915b493efdba5b45146e9699ef;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'heabbbf61a9438796a12921abfa411f3ab787;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1be618b8bc01b5601c1e19650ee8e09cc21;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h87979f4c4a9a279be2c5f35809add7ebac8a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3f176e2819d0625bfcd76a0017ef508ada9d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9f7c63060195a3b538ab46ab397a291114c3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3d3d7224bfe56ee30308ce50b4127d6823b4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h455350e1bb9e90aca5274060528293d350a0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd6287ee094f79361f4f8a37aa919cdaa0ae1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h46a34d2df41be6306828d53d67252d37b591;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h49b9111e8a034328aee5a5a8c79e17031c5a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'heaeb4c081ffda4ffcbabfc9a2326bb625c8a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he4a748dcb702005af4b71c6fffa015c1a9dc;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h717eb9de6d7f4c929121907dcf881b9cadbf;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8009373caefa4a6509709e2beb0a8a72fdf7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h70f0dc91e818a5c671f342a984ec7a4d6f8a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3e6f98cd094c6d25c5d311d494d63179eb92;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha46edcf062239e371a0adace90225c76f1d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8fa1eea9d8511e4514a5d68c89e748b47eda;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hda4614672520ba61eeb97330eebde841b945;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h668ed29f94406c837b2444cc95280dbff3e8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h755911100de0bbdd1b5775a0e4297e66a2de;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hdf384ac09e77aa64c569fc67b7055f81cb69;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he9a4d54c9ae34fa7cd2108d7094a340fd493;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hadf4f6b23808890120ae18d5a92139e25773;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h16720cc369d94c32e374e5c78f50f0e26720;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h59eac4d718c76035e25c8e4dd10c3f4d5f1a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h632ed78c21050dd2bb430c255611fb629761;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf37c4505cc2fdd3c031015ee2b1d62ef8709;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1bcefbf315b01cf09fc6174592ab295adacd;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb445e9155c61448fa1c387bc1c1cdd4a9efd;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5ea9fe5ca2c0e22d64f01636c92d4830b281;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hecf554fe6d50224036991970ddfa212bf453;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h358e78500fa906bd868218d2fb07ffde27df;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb58efda35ad21967f7a5ed759d0bfaf2f258;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd62779924f024283091020d5aa0c8e23cf5c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hcc241176185daee913bbcc872ce1e53ba85c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha73c267c8c5a274f018ac953868bbdc69c4b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4787fe47431a92f6ac184b7c46bf1340532e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h241c910fdaa0c77ab16e0925ff58c0b33122;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h34324b566cef94464bc4ab8855770906a399;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf9d745fd2f14107447514cc61fe002bd1a25;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'had3ca2e848582aeb6926f161699801742edf;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h290abb876a383819996a32c14d896a0e8fb2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6ebbd5f99c49be3ee57d4ef8951496501df5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha4eca3c31b396ed864b86bb3a8f5e19626c6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc15bd9c4dd6c5b89f93ffe3a59866e81982;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h297761a6c2868dddbd409037fc3dc77b66cc;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7baf539558ad2e5b64188080b58886e798d9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7007d3f2d48bf625d67e6e78b9cb6cec12cd;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1fe76724a6f1c954d36445993c858db91f0b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8d60a59306f84cbc7ccaa3ea0dbe13a4f4b0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb1bf491e5b436c0e0ce5b895f9f1e20f0ed5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8d9e362ba3751dd84be2ca9c0f4e44e20f5e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'heed2da81ec2b073befb18ec2efca9b7c1300;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb7d31e143315824440123898a1630da991cc;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9cd56fb18a2ce32100652c035e075591365b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3709dcd0141c7757fe0322b6f91342976265;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hcda7bc2d439201f9e2b5ee563a537f3168d1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5aaba21e3642f96768c420bec2070f7966e5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h16bbd713fc02290264c1079965d932bde7fa;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb4c3afb9343199e8faef6701b439b61232f1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h425bb55e1dc8df25881128cbb23db017ff3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h683217bde0405830a6692e98d84fe44a328d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h26342cd7a8f05ff14b7634da39b995ff85a7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h40ef6cb42c61a2109c139f0ae2b78b14ae8b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4c36a732ecb4867d227794b130fb3edc3f43;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h602ce77e39acd57962dae9c8b7c9e01afb19;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4e8f027ab24cac76f202ab82aee9f57adcbb;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3867d2cfdd602fd9d57af92254c73294ea68;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8696e7eea82108deeccc31eda2e8f958943c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd78414ae24481f9211e4a90fb3708fd9f89f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7d83413a49980f8b1df5f92262b36375886c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3d3b438c6f25e1da05ab0744d8ba6ee90841;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he13ed7115e5d5de62881ee7566bbba3bf65d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h961c387941ef18241b06ba3fd32433809c6c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hae8a07c4698f96ccc7937bb2430c120e72e1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h18171d09fcae7bed778ea30a608fb600bfaa;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h74a72b9d15257f10356b9d60a9b88efbbdf7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9a35e795b47b8065c021265928f3ffe5da23;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha39745b1b1eb851857eb7967baf9c4f6e368;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hecb1bbe3a0de0bb442a0823eb098bce4512c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h896a2d6836f25f320992c54d9efce2fa309b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h70fe77c93405b2417407eab100b9cc43e7ed;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hed2ad0c9d4e4845a344449ba28ca8473ecfd;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'had8103101f981ba5765451ff7466455c78eb;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h11cff319ba71e1f9e0e3100ce39a3cf6bca3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc13c9cddca4ccbf47bed826c11c148ff27b8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf39dd16438a44aad0303898377bc847b6de0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf8e4a9df6a7a9683673524c167daef786012;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h570028e9eb69c592f90f6e28a8c8ec884e56;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb3fcf5ccae1f16a0af9e8efd353b054cd804;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5b7e549237aa4ea257e353a932defc3c5b49;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7e378c1fe18912713b751783d9272bd7f4e2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4b2bb1d5559c741a50c7637cd0cfc3030d2f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h26d59445858c7b77729ab30696621490fe99;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hafba094421743b6ef61c8a7d5cbef72c3f9f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h595002c32d8352dd9a22fc6ee3a039fefa52;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h18131b276f9ba05682c3fef1f1b9bea6762f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h72f9134b53e31f119e05756d5a8046f434eb;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8963af43e247fa2133d7c2b46835769c2f96;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc322bcf815e6a71176a9f22d812a6b9e1403;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb253f915daf6fa159d0b6781d115fb2d7989;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf0e0cdc0af2364d2c96014941ef9600a4a60;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6ea0ba5038f1c44dd007911b7fa7a59a47b1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he4d7d6e31577564c91ebbfe0b2259bc73894;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2a67c91083c33bccca9c616e392a1fe5d2f8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5d1e6e82fc89e423683803e73f18e6900dd0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb81607f10b1106379b72f48009fbe9f5280;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h458110320c295b5c5983fe4b24dd7079a478;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbe8a8b75f31a1994dc3021f936919f8629fa;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6f9aa528bd95d765ebdb49ab5a7a7162e8b0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h82450f9fbca921712cf2fc4be79ae5f36fa7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3c89affe3c47c2d98363dd206c80280dba7d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc65acb4d264dd3fe4d8125881a1f15b34637;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2cc93d6d5194f457b71882123de7a763e40a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8f1dd572ab7381a546a86084b9c3e5722be1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6954431e571d3ba45c66024803046c25534a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf1327252e73dd8004c669d3379a2ddd02bf2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h48721abbc7eb5b6ac083b661db4d3b6d7261;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3cc42bdcff35ed51c4b2e224de1bb429bdac;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd1063dcb86ec3c111cafa2502ec4075fcafe;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9f954e8060f0f680d9e928dad4fff1d63f20;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h682fbeb89080b686df67e591bfc9a33651c0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h69c0fed295672c684c13b499f76d28472296;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6ca47feb9b482f4d24f81d30122d5d7bc4dd;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h610718dfbd02e9fa2c58e4a439ab8cd3d71c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha60c4e05b4c18d4b4c565cbb38f5d515b91c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h90eab4fa41c8ed0f98d385c2509c7f7378be;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbe34016bc7b4331c8cbeb9c180ecfdfaae45;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb3e32a34a252b777f36896fc2e41625af75b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h559820948ccb083b137f6683090a47397824;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8d256cbfe41d8867fe736635672164ee9394;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb499991bd4e3bb14a7cb6e19ea55696561a6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd57a49cf99984eb101b8ee6530243f709ada;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha83ef0a24f307c7490a741bd0198e906bc72;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb85f4fd3b849d88d95e167193874b1c8368f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h40a0c154b28a0a44169294549be5d4342944;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h37053a861e6727107e7f1048bdb7aadb48e9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h68931831fd815298333df80313bc7af3eabd;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc4f4d72d461f2117052a76bbe655dedfbf8b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4e5ab142f8f271f171e88e8957d8d4d1b326;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h59afdc1923f2b393d79732d965d981475592;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h86fe9ffb9f1e23da67d194cae87fe3c52b70;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h621766c4c5649df3305a1f752b94f22af09a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he3a9ae6bd74f3f1bebce6b127aa19df19ad2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbaf6aac331aa9e78b073fa2280ee950675ab;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8af5d8f61c50dd7af64ad096cf880536e6f1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf2939c9136e0a1af51b4b3bc6dd4fb216314;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h716c3f7d5408748ec006490eca19d65a50bb;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3c7e5ee25fd910c4d11d26ed0401d5232a77;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5680979c98295e359fc4671eb1a6b22ed73e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hca03a88bbd497caadc8f3225fdba4c52f230;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9bf5756f1927a287e6cb464e596e2ba1068d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he7723cf5944677015955071ceb2a8fbc04e8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hdf609538b9cd419ac6347c22fc38ef58964e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h157f5c8af2db277e91dae9d58a2fd4dad51a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb955fe39c3a2b36ec7c8a1f7de3854778a1b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h42b0783b46e51a5f5cfcefd3c17e1a152784;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8cbbe3d86fce650fa3fb2c9d4f45a4ae60ca;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4a3d5fd9604752b2b19eb6bf52f86a0c7473;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he7774b32cc169a209a825e2c60d99841e834;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hec22fefc132dbedc03200eeeb637a541951e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h638edea9639d1f17a9db531fad9eebbbaf97;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he4589c94abec9e001a7c5698aaecaf5bc69f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha39c696456953eaf823234c462881838ac5a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf17e1f160bdcf7ceb7b975487e6adc7a64f0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9e2c3957f9121f548fada3431e15a2a13bbf;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h715c97558ef5b6ad574f141bde7f3e709745;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hdd3b9d4ac7f663fede4230cc0f7e9e117243;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h95b77ef1e4a66e54c270b3be4776318be337;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2797d4bf2883ef8a4212fa50ce46d20e1f41;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hab9f6d6acb963eb9b4755916bef395638ae4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h994bfe5c4dc3cc7cc1d20761c8ebba4f522d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hfe2d34fdfbe786d99e5b7030272634143c7e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h98b07974b5dcb03b5d7a4294fc77fa018bc9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h95766033ce4b1084713d0f86c063853006cd;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb03a65eacae86dc1919a70f1480278432c43;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc0b5b93b267f942b075be52e53ddbb6ccb2e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h497d9c94959b760bfe344b163921483db0ca;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbbf7c454eb0db41a3f0a4c3265de6f14dd29;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2ba67c3d941d8a4fc28e172055054c01060f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha16b92d22742aa60034a60e35d253bffa7ee;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1d5792b6efe65c10b1640f36dec041c11824;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h93b97db130490865755e39d92bfc4b5e1eea;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7c3b38348f1b275e876e3109a55df37d8912;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hafc11061c9abb3326a943c973f2727524702;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb9ffb1f417c005d31d25e69b762b0e5ec08d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbedc9ed415ca75483752a308688d54077069;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb4953d30d6f84df730631a6683704b71c3ba;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2da28f3dc280317dde56b6406191427a0556;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3a328b836ea344402f1089ce01688d6c5126;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h836d404cccbf045fc48b66784559acc2d8f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7eab946f02c99acb3955eb6bb653ad407eae;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha811ae808f0aba2b01236955cecbb0cfd5d0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2fda05408504f9e82aeaf5846d252a3752c5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5b1db7d2e67ba428e90a58f830387e6e1c7c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h270d310f0dcc31e4a684e53b042dbc43a247;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h31e789878a3b08092a9af7cfeff9491e6d35;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he97b6b64964d4eb4aa7bec70fa545278a2c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h181a66d0bf57474aba7d7df121ce97eb9c23;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h30322513787985bf731494de7602af250249;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8f0cb112a2e68c532a335b05ee3322aa20b6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hed59343f9956694cb7b13e443cb161699fa2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h21d7968fb69127e7e78ea3c53fdf870248;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf48d7aea3e75c88823ecd975329b0208458d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hfde6a7a7705d1ed653966c21966fd3525d12;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h860ce0cfde9cbcbe4a28f3828554b55b01b1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h28d1c25ad7617b5e3fec44ab483a677ad86a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7cd7f1c56756aff56b6d2f4af723c7d3dcad;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he440ca9b5ed66854e33da28b361807e337b0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h82d939d4117c9b06f48bb8559cf394bbf420;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3e5c074173cd91bc5896917f5cbc5e1f43ee;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hab9ab7098b0fc6245f21a101b349ace52c55;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h82ac4e1fa0e240583708ba27ff74aba9dbc5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb60cade79f237042e2d7f1a29137ab7f9876;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc8e14a51aab3611d3398c66398b2c801f0cd;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hda3ae24f339544ad75e7c3b48b6db1e7e17;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h58e624049667046019074a19943472e6fed3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h867aa9a85bad36f3fb8a1dee89fc86906f91;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf36bc6cec58cdeef0f8e270b6a6537311cdf;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1dfcba2031ff5e10bd41c38a70519ca6f11e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1f605cb25fa1c114752866c7be8f8f23d2c3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbd1efa7a84a7af5ac96dee8a5a81f1484f82;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2f080883ed8ae2f9654117f563f1aeff0cd7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h53d194536e3922c716a11b7b6115c908c5e5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf410db77803d7bed2ce1512f2f322234c91f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h364ee593d559432f1cf78c0db4c0f793d212;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h625e635a4220d625cfdc672f62f692cdad62;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4be6427289b090d04c9461739fab68cfd4be;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1f5413dc270d4c97759e74b65de1bf80cd6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha3b4a87ff6caa3210a6236eadbcbfb96f39b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9e04181a3081e3a9aea1dae2c8e1b2a48afe;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hade896eb2f16196fed1415ea777474c97949;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h711bd330722a32f32861ccad8822022db1c9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h251b935f2538a01a116fc4258e1e77571fe9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha4dd91e86e9baabef909bc9341e225c23d36;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3abb2d8dea09bcd8ac154b330bfccbf838c2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h113fca15eb0a8edb248569c194c940f41dca;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h39cda619dc2716a41f642930b63847ec463;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he839f5374e3242dbf1937fdc2599d579eb83;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6c1ab6161a7b73889bf4646e50320a22ea39;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h99b9ef6669843f35661df01b2310bb3d1494;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h493a70ac06a9d4051a35ec1ac59527a8e016;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6ef5a52488e713f8e839c04cd2b1391107ac;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbc63d5b42c465f32738832c9a8258b1e511;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9814ac0b4afadbb2fc738b359690337468bf;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd9681c295de88fb04b4fe35af37c8432914c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6b9baeaba811a9bf2713bb7711d7da2ec99c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7285332f06a15bcbaa447b99207a7eb273d9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hcb5ee56dd929ab803e4a67cb3f8c8bc9c1ae;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hcf69d7ece8d0f38042a2eeb3a2b2e3130641;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he79eb9cc4bb77c8eca0a16e36b734ac51c69;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5eaf430e1f536dda10a50e2763322e9b07ff;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h11869b9ed49b0ed30f8a9e545127e7df9d5a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hee0b8cf5bc89e472175917bac80bb1a1654a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7098b93a4e8eabf3c1cf71649b8764b9e775;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb33317a8d15b028d9cd5164c3b4611b19e98;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hdbafdd339377c65a79e0644c2100ed19f1d5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd7ec6fc6ae3bf83af131ebfa597cf40a6d60;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hdea549c73c7135141779789e9d8c38d03af8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h50396740191552c60e06225de760b622e4b2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h15799b0dd1a5f9ea8c2c3b8c11781c1a2eb7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h23b14ef1c86efafbfef3bc2cca735f8a7ddb;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9536e2914a2ca5962e75d28d7cee593b5c18;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb26f9653389481743e7d820e24272b87a99e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hebc8b06684baa3d94de4f0a2fd2b6fdfbf1c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd4394dc480ea5afbbe9e630df651862c13c0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1d148ab04a5c9ae63904aa0e26a8b954566a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h18cc7db4dfa1d37d3657353ecf886d356b54;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h35e70bed09670d4fac94de68ff6cc14d157d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb4732f5d70c39841a606a0319ed1301149b2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2d5c8b9aab9021e69e50e36b0d489e13d290;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd24d9da4eb97262b301db6a0af5c48ef6a7f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he31c5b9d7fe1c65fe12cfc7ec4b2a9fc2992;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h51afc9f405f7b83711ab4c0efd087092f78d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h869aa2372375c9a512f9e07a127222fa277a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'haac1193a8643f8e2efbb9cb6c22b7f8a6321;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h35da3bf6c6aae90155e7bfd42ed724249518;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2d56f65d0d8f763bc05c1ccb4f1990be3118;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7ff30b2c22e3268964797ed13d0337ced417;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hea3452fc3e2967eb214c8e0cfc357f50acd3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h69c6334dc248edae0c399c116eae2b891d70;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h855afeffd6fdc1c8d204a29f5e1386289e28;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h61d6194473818e4574d81113730dd0af768f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd12b4a3e0dc3567ea7ef43051fdd71c40fc9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h68100e092cf7a9984e4e1753ec69b177a8a8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2043852056d3e8071c3a3471109d33d4c96a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9de0bd12f60308803bef01a63dcfc628f80b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h92c64c321cc4487653e7ba8453275b70f513;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3c9c9a8f94c6d50c9fca89c2297cb4362bc3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h57c1add1b7655071851b454e38bf268efd30;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h92f55223d93e74a0a57228c64e1a4e33b6ee;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h357470f4bbc76935e79daeff7e0166de5951;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha70ddb3da23e995ff693a6ad77d45f69e8a0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha96970bc3f3daf08df4e07302fdc945d68fc;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h54087e8b08c1cf57e247f84e95d2529de721;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hed72b0638c8e148a0ae84ffe06abf7bca16e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbbe0041bb5480815ad1ab3fa24d5c39fd5e0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he8ad9e96645b76ee1fec3d4a8ef611a15d3d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7cee44ca4f6012f88159440941f9bb636f42;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2910c9633e2b376775e9b35e377d72a847fb;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3aa5c7ddcf79b85538b63c77b172a04919d3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hdaa5d42d8cfa3bff129c3a872da00acf3d78;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h37ce1c6bd95954d85f0abd5c8b1518ac6b55;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6cd0426fd9d671b22dafe2b786dda9e8f153;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha1f086df549801e8ab915f8f21c7c7e041c0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h52b687b3b73f0b35c662236724d898eada22;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha4c197e2846520d0897c60193afddb144bf2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1832acb4c8fe303fee8d757ebac4783cd8a2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1fe91ea711527942330aead3efefe1c37045;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hfc65e4bb3a93679c7f179ac783a4fdc1e573;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1f67538c6e0819b2a8b030a089a8c1b87e5c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf2b195f347db34d93321911b510220a04dd1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hccc9e4e75dd73a481230cbf3b9d91b8fb46c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h355467c0a94c2b5bd7a89d26f61ceb65014e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha81cec6238d0c5b2f8b30ea63279510ed149;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb0e270dff7503544725aefab7a2c143c2b5b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1fefcf25ec18b5b4b8bfb7996df9f2b0c3b3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7a17f0c6f29936108fd76094fa78e86ef10c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd771a87d6d226cb0621e2e24dfaae6dde59;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf3f6999f9772b77a3038840a3622ace9a6cf;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7c1dc7b9c141957bffd0616f44923d883f3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd837daed18547070a9e607ab6d4e214e0adf;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6808fd7d244dcec702248270e78f2fb433c5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha0fe0934a57e6197c489223eb42d187eb59f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb037307046fac8d195fa3dfbe125750932aa;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1624c61c6774fa8d24af1b153cd7059d627;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hcd3b3289cd02053c27fde08414ec872d9bb5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4ea6b8e6c5d838814f4c0e2ca39d622e5710;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h668190041ed7e0f005c009788362cf914348;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h26e684f1ed54e4766d43d486608cac0b1cb3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5ce07577a4ad77838a5b7425d3b9b6b689c6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he254f784806842c318274f8d2df441d867dc;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h770becfb29f198da2b735a099ac886ed10a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8f29db186f403b99c2491a7cb6ecb43bb3cd;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7ad2c33b021769bc793ae46fd8908d298c03;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd5d6fd0fd2e288ebb22169ed1b4895b8249d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h543a2fd06c7bfba8e0499a760c382a71a356;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf564555ba51f6a3b4c97527ccaa526fbae61;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he985dada6a2a20eda98c0131db68dc2bc912;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hfaf2875014d5d79ab19d5fdc7b8a9cedaca0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2100cd6e7c492ff00d8ccdeca0712c6c24a9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h91729727d7a98883c3c472b742caf29bac91;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hcb49d5d8f1078d15444f8b0be1de48672d6f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7b7d91fa9f532622f4bdf167341b07b027fd;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb52c2aa269ea4de609e1a3c8b9ddfa9053a9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb72a72faaaa3c817357aef0fcf926bc63a0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h35c85ea8a5f4fb26058ba449c803767dc0f5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h370a618a36eef1e9a8fba8dc95a999a87b2d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hce36e400b8f73ce1f3d235960ca8c6eba6a7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5affd7123a6f21a926fec1f94110457d2081;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5931dd0432641eadf6d254b10f29144c16a0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hddbf4a2ad3199901bc1206f16c8fed654ca9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb65bc2462060db85cc26b759c6c280852368;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2832daabe1e9aa613531c338db5b212657f4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1aa1ad437eea01415876b65e657da1e31b60;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7d36c025cdddabf7381552aa7221dadd2594;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha1d471428ab2988447b0d58ae248eb053287;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8ccbc698b77fc7aa1330fc19c6930e1946b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb2b300c578b36a8bf5e0285eefb021e4cf55;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc844bb6d04acf3c3c8f2699c6a059738a2d3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h13af0d5199a000925dd9cc3ef6bd5961d307;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hffed0f6e621eea5e0d376f72463f436f8043;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb4c1a5b6336a21c50881f8d7a6514547016b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4ed5222fa9d2bd4e966de13e23b1da95d67c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9240bd2a1d8e23d947575943b871664b1210;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hee76432347e34fea9f50d983d20d5a34624f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf61e335f04ea53afb502105885c154051b27;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h209dd377c8d9ffa903bc6dd74002b47b44e1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc5d0de312d455fd365e0bd7be415fee70e9d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'haae436039a7acff30e7df77e1151642be650;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf43a1bcddbda89de7a762a3520ad51779e45;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf463bf47c3608325a226d5540d60b25a431e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'heb9a05a071d6ce37e24ef92778b0976362d0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc787c5dbec54014b9ca365a446166e3e6a24;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha9e98bf5d7d2c12a8071a886fb6bae1c8acf;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1dbd25593e49bb0146f93d536acdd5d82eed;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3e329aecaf443f69c5dd4c7a38d134a64ae4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf6a4e207c4e99b940431da8418da8dccfe4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h55140a7240be648b1d62b161bc1bf64e8618;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb51bd8280d223ae430fc33af54cb3d7a78ca;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf1c67e4d1da7127549f6e97f7e0f2ad52ba8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h28d6b5263b7e9833458a027b2d4430cb63da;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9dd9de28d27eeb0cc3c86f843de4a7a84099;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6c61821b7e59bdf625abe1ca61d392359804;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc326cad5569681db2f71e1cab6871c2eac5d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h86245b21ff6689033dc23ac2e70e0878041;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4d701950085cb9b028aaf994f5ec7336d934;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5354733d04aa029e1f5dfa1619502dedd514;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hcc1e63f3fb35938f37375f71d944fa2616f2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb6a5d102c66651a4cdb64aa396ba79406e84;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf328bcaca5dc99cdd58fad07538d2abfde12;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h63cf944ab620b539d3f39a7a08163f290b57;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha5874ee5878646ad38f173c82d30fa062e66;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hdd784ad079d46a5d439b48027a922ade9be7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9a56252d00c2de0ab0cc066488959c97b48;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'haceb446f5d0ad050df14aeecc3397c0c6b36;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5768aa0f33f7ca91b89373c5770e05c26e8a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6a52a401360d07f3f954295074d3f5c7559c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd91903f81e9793f53b2df150d611b12d171e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9e82199fd46143b68beb0ed73ab517aaac7e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3be98d315f45428ce61b09e81aac87d0599b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb7ea48264eac6652f4377e985c02833e5535;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd47582001f37bc4b4c065aa0bf22e3b04187;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h17de58864560cdea1b91ac35fd9b419efefb;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'haf6b631fdebeca38c87db4fbcb7f9e4b03f3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7526c7ba0ea8fd57f6b0b7a4d71336f885b3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hec4420e8a2850695b33f793336e83011158c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h173ccbc17ce005564171580b511c647add9a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2ceafa5f17f3c19031854544e05c50bba86c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'haed79c0785759c61c3f3a966ee4618e319c9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7589cea46d6142e9fcbd2477db07db993138;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5812b7abe72038201e63d10bd04b261ebbfb;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h865ad3c9adadcad25e42f3f7e15013ec1d95;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6deb70da15e542f75082b392caaad1d4aa86;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8968d73b202fa6003df30b787def93f1c7cb;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h40db7d6e925b0fb02a7130f01aac1abf22fb;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he77f333e33e1740181f9ac0fe0513065be90;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hec13bb123562d1f6b1a0be69c09a05788b0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hcc98071048c6110fc703b87145d8bc7c20e6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2c8e0d4fc2f67a9cc295e506c89ee54017f8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4cae475f07da91ba3941b2a76d62ee94fd00;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hff3897e03c701ba9deb2668106cb62966f1b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc728da209ffdc7704ce842986c477f51f4df;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h24d02eabf1d4081bcc1f9f1718df681643b8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h172c206e4bde06abff07112af40666ecede6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9697ff30b0a5a5c65e6cf3e90a81b51ec336;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha281844b55c7c48e22d88730e35be2f543c0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha94d527ec1947d2361312d44f649ca169634;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h100f85bdf3ab668e0c1c69a2563c5b70d8b3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7004683768d29e62bb73b3283e7d4f39e2dd;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd29bcf471f5d2bb1434a9e22f11de8cd1922;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1c0b57446fd62686d02b3139344db90b903c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf1223c32516970dd6d988c6a70b27d8a019c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h88a7a62edde8d247ead4c49bfc9ef0aa6d71;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha593a34e16a7e6c5db9e7876d1b3e38c3fdd;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hfcf462c30b6df6184fb13fd1d5dbed82a1d1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1ae126150210cd35b78c86c77dea387954e0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd31d49b8ac65cb2c6c775b0fa1853a6f983f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8d06d4ee07eb8446e83e8f7cb97ac1e68253;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc6bd7eaa23f78aae24e36d4207e072100234;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he403438ac60852d99fa42754f597692b4016;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h191cf17f0d2c0f4ef7ff75398d6f68fb0a74;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h418baa1d5b0cb17c36bfd25f78a0b281e66b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7240f2747e574c9ab00253e411c1a5326c5f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h56c2176c0ead8744ab6d0ce948572ef41bca;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7653abf62df84dd4779fd73ab7e6947ebc4c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'haa4bf43eb348b4eed96f8d9631862e3446f5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4608691dc54a9b050e6d29a1136d63b76f9f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h384be165e9c8cb53d2027940752f5e405ca;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h464916ba4d0f7ffb3117394a3da68a1e8793;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7e1ce53ac7d0342bf87849df58e3814d6dac;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h712e103e12036b333ed949135b4f88c09a4c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4cd3267bbb063f6b7399274cddab1f6ccd4c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc9fb6b8f14f6428016e3e45d90859cfa8aac;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb350d3d6ec2dab8bcded202c55de80022720;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h256e6e8a6c2a9fbc167d9e672881116e039c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9571ccfecdcf50977f6333709104715f1950;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h50175a8a314b6e13c9e350ff1fd9bc2f05ba;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he2ab7ecddc45903fbe455991e7971ea8d365;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha9a75a6fc4f59c194c39c8bc77e8d1a05bf6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h328f2a9eb083391128e1699ac8fbc06692d1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hdf286bdc2a1ba562841075dae440b7414217;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h822356914b195c102f1d373a693740d17a09;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbf3814d23ce6000c0fcd342af2a2f939414e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h35e7d4d3301f89c4c0c902ccf812827e669;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf6aae5be7c29b85bd6a1d93c7b7b6dfb3b5c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h65ca3157f3c36497c041b45ca80a0ea712d0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4bbe74eb8664d37c3f73b66dbd013b1e95ac;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9cf3470a09c6c4549755afb91cae44776442;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5372ac78eef74d9ca457d6ea6795b8c81333;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h29ace6507a1b9320ad66d38fa29bb5ec0296;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd97c2a7276ff39edd85b2e9eb74039d0b1fb;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hedb2bcae24c24d475131bf5e149919faa90e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h989a9a530f9b68e56d2bbf75a60b1f4dc824;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hdf2001adb9adfd6c15ee5e10df7234b19173;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h441d6b12365f333fc681b699b0db880a7d92;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc9a3ff111e5a1bd7cd39a3b6ffc44cf407a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3dd23c508d1cd8e8e42313b4280b60e81e5b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6500a22f14854465ae383570947cc2261418;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7c1582eea4f884157ca62c347cbcbd209d07;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h94e5f06aff069b3292d64f2c447e7d097e53;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h21ff93e0ef31b90997400285ba06d730b36c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h34f29c8f5d6e2f0379e6a83e5932d0f5d4fc;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5e9733f9500ff266e4bb3dc77b7cc90cca03;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbbc813d1b13e545fced733b06724cc36dca7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf740b1970d2fdba5e3fd760c3ded50f8ef4b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h55790d3bb55da8cc4ec3f5acedac3b1f77b8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h14f188df7942714086fe33ddc30efa97213b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8c683111ca1bad5771b597551e256f88e1d0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hfa17f47c06f271454f3e897901fc9052bd14;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9fb8858f357bc58535845c0136a923ef9424;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3899067f3ed7cf0be6f937bbd5f7ccd53815;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha491671c55251285b2417d2392e0307a48fe;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he84dea48f8ec78ea935f081f78e3ab435ce0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb7db4c6e140de8fa3c7ab36872c36d47676f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he35468ae374a7136896420e2bae2ee994cf4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h33d2116771ca96709d670875ab87dd316f17;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h382e29dd584602634de7394cdeb5ddae594b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h85e19b2d9e362db46f6a91f5ea0d0b705b0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2df26251dd308597abed889bea384003da06;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9232dfc13db4cd48dcd32f100f48807a1f01;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hfec59c37e1bc9dc74b6f2ecbbc498f7f62d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3f64b75136523a8eb9d0acaa05a8dd440d8d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbdf4a1af24396cb061e9dff54b4d25572a22;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6fbd395c4fcf58c4e55b1bd2b8f9f50cbb24;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf952ca7e26a7a1ca7fe1d92df61789bc2a20;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha6c662260c0f27b32b375cd9709de6389470;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb756cc6c0b350f85426c37ea7fd95311139d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2ea4afe97b5e55ff3dc4b891c329a92a5bee;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h18562c983ce13f44bd56c87007a3dbc2df67;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd6788421952b2ffd2482c08a7d5a5c6c0b60;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hecea8f59cccf9dad0cb2fa47305c9af69319;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h27b46b12ee701fb793891d71224bbe49bd7f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he283cbc55917295c791f7f37d3b599b6b6ed;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h38d64f79c7b472b787ea2503d2cbc77c939a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h79697013e279dfee89174486ed7bde9df495;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h62d416f7252079368ee41fab415d5bd4bc21;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hec0bee9ed85f562a4d9b36233754b264efd8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1a987ffb9d57592be1f05dc2c1762e0d76fc;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hdf15e14d322c35382e2a01467266d99ebc09;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h231649b407eeea4e5b6d9b9f6724c73e3183;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2a463e5734c6ee63dbc2a41d6e405aaf54cc;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2ac339e847e15828ce15247d0c8975aedcfd;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8d0cdf02897cd91c268aa8dbcd771c44969b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf9aa56c6ec2ca0dc5cb1af35e7c06c8479a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4463471b7f4aac702f08408e5ed40c2f9d93;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf5e2639572930ccc8f5e321f6bd961c97dbf;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4ac045b7444d2db38e58764ed8d33f8bcc7a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7941ef58ceff24ebce9bfd7bf6d9c00941fc;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd1c3da6b0860c736b75046e1994e240b4e3e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hde5238ce08dd6265b1a04558d08ea578ab24;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1b4fb98645327848487bae280c52bc1ccace;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he5fc5f948df2516cc322c32b28b09c3ef906;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9daff05e4979568930382c14a4da0fc13c2f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'haf758e610726eb11f604fc7b9e8efe15ef62;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc6660b04eae86e5f0ab0867ccaf314ef55e3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h195721676d9ab101f723fdde40f2cb7ff2b0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hca1e625f87035ebc5ebdf50d86aabdaa164d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he9657b789f137a2af5734fb31213f19bcbe9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hfcd9401df75c73a23a7abc69370b792ea7b0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1b45423510564a270a425d1780f69f0b1251;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc5202df8797b6f2ddecc236786eead314c39;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8315d8dd446947afc186da0c0e2ad12891db;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hdd723e3226828d8dd9d794c79d78ce7d444a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h37feecc6b4b94c1e786fffcee18e3d83e773;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h54687aab93bbe4e63673d4cf8902845141e0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7d6122636908c07b0da5a0af449a7b4cb053;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hefa087b0f8ca86288d2a9f6515e3e3579d72;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hdd7858cf4c94b5b7110c7824cf797525671b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'haeedbb33bc14f7a48fe6447b91e214f0e539;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h88071840f457bb70ab5abd263f0b92e2fe12;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6e7a46e8663cafd881c284d3c96f165ee6e5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4fc66eda2d43f372cf90ec06948002d02103;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h220e1bd32dcb38f44dc86027423607e5a23;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h827937169d9f600b49b6a8c7567743edd55c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1704fbb6be31ee6b45a5d49b2d685930d7b6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha883c4800a309ce84eb829cd5ce7c38fed2e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hec05ca8e7467c56110dd9142140ad3e5f7e6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7b779e4def67efecf2bad234d6f874846587;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd29dec1737f86ebc5c6ea6b655c502d8632;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8b8117fb80cbd968aca30d45e318b6efa9b3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb8b3d749f8204515a748f6724f78ce99ca23;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd4591b471507d45634e0a86ea299c2d2fdcc;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9c3b44283d70220818fdfc0f68404444f70d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h55e7f305ace3aff6939dfe60ef4f351a2373;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hec8f5439892ec321d47bcfdfd577ad499227;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h982044aa7a8c173f366144af85de4e76d645;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc886c2d351e02aa83d32d41cb378b70054b6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5a9e927ee52430b4951018941a447cd3398d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd88e7314104390c40a372ace8362f7168256;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he30dc8770500ff0220ea94377abf26145eb9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7d52a22cc95d4035155ced55cf37fbe29439;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf098d45853767a0250e0a638a28087a3ee8a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h24d762285d39460c9552b1c4085ecb2e64e1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb012308305b239236a318ad083e70d19034d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6bdc0035df78e31076f99add2638fde113f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hef0004bf863b3080af72a89e7c1ae7654210;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3002199f37d9554c4254ff5d746898a034fe;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6a1d06ae8ee02d69ce191c061c30ed81f19e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb2f2b426fde1f29be9dfd88e7a8eb5cb7a78;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h50b41c13cf40ec48793026ac1ebefef422bc;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h454e17bbd04a84225fee246d9871f6de0f41;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2e2e4d005408c85631a965a8895fc0ba0ba8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h47053b379749c8c94f322bbd9c7400a35024;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h25738c4fa31e1db8850f12877777cb4a891a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf2bd17164dc49260b73cf7e76cbf12802448;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hdc4a2dd024a0cb73562d81c1bc919b3f3875;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1c47135d04b9c84ccf106b2752e30ab2c2e6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3519ae1df4eef8a6e3c37237b0d7b6f19731;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he8f3e43ea1ab7e133a1a6735410b9c145c00;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h656372a8812cd53680e0b8b6cbf9f178ae1b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hca959b5039184e326f9168e86f4f93b146b3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h10af2d3cbc869c5088981f2618fbe8e1afd1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h45d6dd5d62e2ae919dd2f9cb3429200d007c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6967fb552682d669e8904c08dde708ae6bb9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hef5d38cd24ee3d921f378b623295da052526;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf1c9790404bc754d9c100d14a1d55afe37db;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3431b532cd1d39a9f922a693711b92abb89a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h767e4844be856c858960dbc193c632af49eb;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd60639789f3ad81d77796b58352ea4537da0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3a0ac68c310a7ed7150496e060f128cee664;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf1affc2721c034c804f2234956aad2f177c5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h46bc154d300db82b31f4eb6ee52648787541;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9baa1d0bcda753f0a4575d7621a7a3275f0c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd08aa0a4d6b43cc3eade173497381a305495;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd1ef2873fb243a317f4ebe54a73e5dd63c6a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc3a7e98d451281ba0039499db29c48b01b9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4751aa3bd210952f0ab387b4dc95b2bd078f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h50d705da840e5a9455303c91f05dfc7095da;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6de6788f84ce2d629e864a5daf57dca181fd;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6ce8b6586991a37f710885fef5b930c53ae4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h65a5cd844368ebc59cbeed9692b65805749;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb38c27f039cd2fdb8ffc0fa9dff3aa1201fe;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h36a25346a1874866b4a4c4016bfbd4ddb0c1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc79ffd8ad30d8cf4608dfdf83490f28588c6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h36842fbe997c37e4f66c9b0f64ec1fcfcda4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h621c81a24dafbedd0cdb20def783da60f8fe;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9b1537f2dfd39391ccc9f21ba34512630979;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hdcc1637c943d89f2f2fb1a69e031ffe1dfe7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5f65f23303a7a917b6d8bf8f13f0bbc74485;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5fc163cc85f352fe19c9e273997dcde1f1dd;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h22678314a114fbef83cbb6d24dec9cc2b833;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h342a0b694dc6d2e741119858485fcaa12d98;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha07cb22bd8e1827b711e865661dbc97ebd6b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hcce4a1a2894c14177726b0ebde40c5705d9d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h555127ded46d78cb2c20385401e1307f175e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1daa8c24b3d4c72f8855117d097700929dfb;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h51da0d5275b1613108794c56a53132923426;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h54f39b83b32d7010d2416cd336cfbd963d48;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf9355df508c3119e5212e36dde5bd984bb15;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h99756db12347034af1029aec923afed11284;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbe0a45ab75ddfcd2b8661839d163058f9d3d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3365fae1cee46a7b3810ceeabc7f31691ced;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9eea044cb086a8133a1fc64ddc65ff5c0193;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc0365267df0525dd8176a444ec0eb823c0c4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'haf713c5e37c642cc21d7e2c0c8360e410b7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha75fb51bc4232042e2d53bfff0c9651f24df;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf2bbf6095e5a9b84d3df77a3a75359bec8e2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7ddfcb8a704ff08870c40f53f1bcfeffa3da;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8475ba68a3daf8fd11b1fea4ef36bcd8a613;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9bd07e82382e2a9beb84e56e923f84e0b3c3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hecfb2f5536406e62b39e1d82df67c1e0eacb;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3131224427bca4c907faa7fd9b554c59551e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5449f362be9dfffcf1691391083daec3c5a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he729314421b4015bca7776ab2620fad7c30d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'haa4946c087be379b72d519d5c1d8d706a54a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h67155db1e4aa6f6af19f8d942cf90b69aa3a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h62fa1e20b83fdf93620341f4a54bb492c144;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5164dc5669478d1092db39d681ba2efafafb;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hff3a93072b1a5b0a9af6ec4b17fe14807672;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha7624e6ebab66a13f5043e36da8deeeaf968;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h98306df825806f7643d6536245ddb3972572;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h87bef1f1c1efbd96b3a036e32c38b043b702;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h67fb7ec482b20865a742d0ff039858e78196;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9a497c0874e3b6635cebab6a36b5b98b04f7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'haf2591921bf12b0521ac1ec484145f7bd392;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h61b26bd6ecb67d880bff528a4a92cde2af36;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7213dbd58d2e723208c4925a346a4ed0c07c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hac4c2766bea0861a9d343ba6d064b37528f7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3648a95c0783a5163a844ce1cd9c9e0e93a6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6023a837b32e2506ee4f4a6162f802cd21f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7bd14be422c0e5379309d22369e471fe3807;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h845b6fa8294f48886c5061717404f4022550;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hcb7b042542ae106670ebbf4213b88bec86a1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4369a07c733f637be49a328e9f8070a32ce5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h14a70c2bb07daaa5b4c3448086cc1091dab1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he937390b57476af3d54aa575eac8cc0eebab;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h32557858367fba34aadf018793e7d4b0688a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc0703fa974f6542a2c6e0559109cd5a6af36;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hff35cf35a066d1dca0392a24dda337dc7faf;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7f3c8b450b3911cd1029d94498a2852ea5c7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4a37742ee6cd4849bbde7eaf21f5ccfbc9f0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5cbec02e4086b42205089de07172d4db8dc;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hfaf513972730865cdbfe4edf4c780210f498;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hdd75b29918b97f4d31edb9362258fb9d9acb;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'heffa64209a9a8f9b5e6232d97be8bc35b84e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha201d053a696ecd28bcb4fd9736145f72427;
        #1
        $finish();
    end
endmodule
