module testbench();
    reg [16:0] src0;
    reg [16:0] src1;
    reg [16:0] src2;
    reg [16:0] src3;
    reg [16:0] src4;
    reg [16:0] src5;
    reg [16:0] src6;
    reg [16:0] src7;
    reg [16:0] src8;
    reg [16:0] src9;
    reg [16:0] src10;
    reg [16:0] src11;
    reg [16:0] src12;
    reg [16:0] src13;
    reg [16:0] src14;
    reg [16:0] src15;
    reg [16:0] src16;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [21:0] srcsum;
    wire [21:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13] + src0[14] + src0[15] + src0[16])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13] + src1[14] + src1[15] + src1[16])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13] + src2[14] + src2[15] + src2[16])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13] + src3[14] + src3[15] + src3[16])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13] + src4[14] + src4[15] + src4[16])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13] + src5[14] + src5[15] + src5[16])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13] + src6[14] + src6[15] + src6[16])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13] + src7[14] + src7[15] + src7[16])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13] + src8[14] + src8[15] + src8[16])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13] + src9[14] + src9[15] + src9[16])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13] + src10[14] + src10[15] + src10[16])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13] + src11[14] + src11[15] + src11[16])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12] + src12[13] + src12[14] + src12[15] + src12[16])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13] + src13[14] + src13[15] + src13[16])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14] + src14[15] + src14[16])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15] + src15[16])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16])<<16);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h0;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1215e434fcc806d236606fea547b6d3d27aa3b6c0dfc6f39d109e44ffdc884a90673c268d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hbc3e66a7048d0704f580a5922227ba1b56809c52d63bf3a1446c83878ceba9df883863ed;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h21273b2a0798bce33511b894a51ae6e64068db383a8917a1188b0b819e3687d7f75a9bde;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h747ca6512a9c4e3efdee04f7dd913836062508c363008f90264a0f529f2a681cd02c9b96;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h10606f3cc7006390741ba8655d67c812bdca877c47fabbff04a87c12c6fb430aa3effd2df;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h50efc12656d6c5b4389d351e753699d00b6964383d76ed80754f36982bff679ef88a827c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h512928c7118381a9c2beb5c666e363e76ef02d20e6450e4b2dc7791ef1231ee6b8629dae;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h11e39dfb2cc71d2fa04c8d99020e10901f341fbca8a2a332fedc12590a47eae3a6c83fc1f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a285e7f75eddc2f78703d769761f9b3f545d22b16b64054cbb321993176b0fbc097ce783;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15794140c9fb55839d7da01658db55e46c8df323aa960c5516617ce7871f65190aef161fd;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f6fc492c0441868bc6121c1c50c635f9eaa98df34c7f6f6554d7ff5f0b50fb1738eae841;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h165eba4f17437ba20953cd610309cd510e2a5d5803d760a7f7bfdbbc3c14fdb039da74029;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h7271140a3dfa34d1fa96e60df35403362cc23d2b9d53ba51bb92f1e727fdfda35d6e5f36;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'he566a9f577253bab939c39cedaa11afab78ddecfa1da665ca943b03a6dacd55da6a6ba02;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1051e6bd71b974b1a9581963f82df38896a69f8022e6c6791fd8f0621aaba01d5d4ffd2ce;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'he8ac9e1f76048ac36ac87db0d2990a769b3eae90714433458ae5f56e7ea2b8a1f7601233;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1cdbd2b80692ce591af04cc802fb22dd0424a7216270b3820b81ad52dc5afa9ac86f78c25;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1364ab009d86498b11031ca326ff310cbbf67b1d429ee2d700857a50d2bd472360bf9b29;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h435a4a4f79dd5f458f8e73611bbd8294c1f36975a6d18861310dd82013dda97059b91c82;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hadafbfce23f1e2e50996182016d264a56924d2747e5b4104a5b2bc03b8a85b2b48b86f2c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1003962e1bd41cb94f78e579cd47ff286ffdf9eb7fd19b7dc1a0bf4d1002cb69ae12a83c9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e6b74a166d98d0a6ab28dd903d8c0e0b065d3c90cbc92a664a10a90a9b1764e10c23fe0a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h88a3af832bf533c67f0ff22bcaf8848cff372261ccf69283d5cf9ac1cf8f556a168e89f4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd0a77760be7661c748089f3deea76bcebeabc7272a53271aac80d18a51b5f50b389ca09c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1df0b13f5c2dc35c4683f13239a3b019adb9ae0a6fcb8eb224fa1f57a7f8f914dea8ecfe4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1fbd6e7f83171147c4d4d7a9989493051ef4efd8b65d4c39ab89c933af228093ae1c69c0d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h192c81dab74ac2ff48dbd06e5de1ff612c642b9ff2f6ec56577dbbc42657184f0ff186f3c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'habfb81f177f10fb4007daa5fee6519d673cb40c4357ed5259094242bc7efb1d86d5beff1;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b5583b0155c07abfb25f81045997aad3d803017b37b35518fe6b2d150664cb8152439e67;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15a4258b7952fa6c155076fe773917c858bb88001bf9fa630847be753687035656041301;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h470172ec0242e21165e3047bb534b515c46d737f5a548d25561eb2ee76f0783e9fee998c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'he4d21f5c904dd15832062428cc2f5e7dd355a9c38493df546c4ae50f9597e82a4588cbd3;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h53a338af6d88db8cf951b8cd18bc4121a84c7ed59b970d2956f0d8ba5b52563b43687404;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hcc6c36a7f67aefb4f79099b95f379dc36b6722f3f4dfa8abb2e68ad0dc159eb48f517287;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h294760f5de3df2f4fc89a17de41237a5b6b7155b9fe235b689d42b95ccb4473e57e94fdc;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h77a02d4d16b00caa06a2012dc562520406050eda3a3c0fb6d4e57a83dad94f9ac4f44b49;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h10c88825cafc8f3a4e9a88c9057974df4b3812617169a0ed4f3eb5dc304c89ad07e56e1cb;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h18d39109ef109995272316451029617f2a4ae7e33c7b1ff079a005bf4d046d669564ffe5d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hfab9f877e33da6a18348fa0abdae4457f2ad25228a39b45075e03c30ad773e1dfaaca316;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h182750bb6c9f5e1b91369bd835ffd1431ec31641b5e6e8abecaacb42f1b166e58875721b7;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'haf2d3c22ecdc0e88ba5ef4e8f11d5c08bb2cb04d5136ac90c46e9d3fe50c5f91c639f8e0;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h81de7426a84abedf8277671d71fffaaf0a43247e346a333bf589af1c84df3a209c836213;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h14b40d874b15cc3e415ede1ec2bd07fd28eb4bf939e2c2fa6802f4ccb57e1e06c5d6395bf;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15568e55757146d61716cac9be245ca08821a48e5e2b90db24122d317b4a2ea9d80149b86;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h115c0a3d702c70ace0cc2ec37d66fab9f61b9782f1cd5a796894c2f5f89a97273cf7a04c3;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h18968918dad18347740a409c50c329550be1ab40875bd2eec6e3c36d8d23ed0debf1788bd;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ecfb793d923555c6b15b197b2db43ffeaaa170018d6d07e82eba139511871eb1f5a16c32;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h14f1eed9f1e7eced418240b974943d98d22b7d1c76d977c31836befa009ec20fd34baedeb;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f3737d680d10f94e564c5e1e71169b073b09f466d715954ea30b27bc3a50b02cb5e2a0e0;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h14b9bd2e03e408f5f26f44c79b9800d6602dcfa3e64f2579a0febe2adf67bf75db1a2683b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h126be8e6e9d719bebfe9fee8764bde57a45e9d1509089d549ecdbd5c511fd946a1dfde72c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h325b2aecfd5cebd8a2881010a32a4649c19484d3a2a349aedf66439f7b851310e3b905a6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h9c9bc70cefab21206e16090f70d53d8746246dc56c7e6656e0769cf37f5779081202e4ef;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h179df8aa816944d54b40108a5a7c0da6ed139c177d3eac022376bbc1d50d20921c45265df;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1faa58ed65ce323e41555cf66ad9d57ecc0aae318a38cbda99dcb114e432dc0e119856b34;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h109bde9e5a6efbb1ee04fb361633959ca6cc98715900d040619be043d753064b864083c02;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f683f2f5951de272e9143a906e51b89b50dfb22409d0782714f3f20f5bbf6c7e7296f7ab;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf7d38d6d5aaaf88cd2041ecbfcd6f284cee2ec0f4e6140c538e805debc50ae7b33dd924d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b9df121fbfca45bc2f544002b5b0bd24f709478d1b9478908d9f0e087f1033b334517fa0;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'he27eb6e6def353a0d3d102daad713f3d92b377956bdbdfaff12e4a63b3058d39872ea454;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1bbfb78ce7a6dc341dbc28f29890e4a214546b0d9ccdbcddcc32e4de6890e400b01f510c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1450928961871442a7c703a9eb782ca86770716b1a62a7bba1fc254a578f7ad23a2cd219a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h6511b475cc52e2f5b97fbb8c112f3a40cdc3383904541736b180361bf2be9fb32d2804b8;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h5857e67ff709ca6e1912ffd0ceae9be3e236d566ef07c0cc194cbda1a85d33aa3c3f03;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d1d655896d5628151bbee535b15f1ab364811016e5ea2e1d61d1408b7f47ed2b8fd198dc;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf37814e034293bd4c3c1ffc82e257cc4a1d85358d5f80944dc0effc21dec6d1ac63ba1f3;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h64b548881844682a2db94596789d0b10e1f7f89901d83cb6d943e2a48bfc43605f8f9cb3;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h182f8ca2786fa285106408c93637e33006e047d7ab97be905b5c6577649b22e27ac4ca95f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb4f805790e6045b2e815e72f25fcc8d346f0de8f4ffd3b08f7a7927b76013267f13e5937;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h48b60232ef7a4d2c7c9b2739d85c146bbcbdb0f78f39482362ca2c8f3094a8e9f2a07641;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b0994882e8d2c0e5cee9cc25790139624ad97156f12a3bcbde2d64cbf13e4b6b0093194;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h16e487d17c25a4ca8a65f5badb7f9aeb1b1d80743aa0b38eb5b38cc7a8a54ff0c827bbcb3;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h6ce6c186df1e801e0446786dc2248d9c9b9fc96d2fea50f9e652101c7ae357a924342db1;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h483fa3b4598a012dc88174603153593605a87e78e65ebddf654a713503a2690eb59a08;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h9d9323478a80922048d913cc73366db58c39f45d2e3db95a2afcf4d5fd9126e2f2426388;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h17de175e42543ab9b1dc897d565e0768aa21dd4c9feca71118a380b41a71082e55b1e7950;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hfefd582f4e07f7cf4be0dbc9a55ca2a54bbe4ad0fe9aefd3e855b0615f083829352e6de3;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h55115a911ba2df8220c5510e34a331e254fb056ede6fc1dc87421e6e248e4dac0556d91c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hbae7c03173d06b59c623a9ba25fc41f5ef679eb3bce4b9b99e3db2254b31aec543c29978;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1decc6d87e98592a025dd6170ef5b48fa5fed2a3f3e532f2e572d811f7460069b05c7bc76;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h74b2e47a51afc71e4794eec21a3b50ac71fcfc437dfc726a865d4c678c0203aa56c528e6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d5955b8afef0b7602db166f22587de7237aa8a5c283ccfd51480dd269b795bbeecd63ba5;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ad651aa4065c879a0891a2f4b2f859ad464f6a8368c3ea75c31a1e49feff9305b2d7c7eb;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f4212b6b8c131b2417faaddc32832b178d7f99eee99676fb0418ee7a9e04939783921374;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h12ac084a51c346c470134a8a089a382d4b6af2c3b780550e3cb85ed5ef60b6ff920b124c8;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1bea78660cb68b66c38feba8f140f51346335a323249b6f77e757a00361bf962d411eb698;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1acff95585a5fcbdbd1afc87dec636d75dff5c73da60a9bcae708e6a01f0a9a456c19e2b3;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h337119fcc91d0a0e99ed5c9cd88e9f09938fa76c21b7482992427e704618e8c093d51bca;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h18163c555a10d022c32b7eb126e5fa19baffbdb115bdc0e057d5f79f247b058cdc700806e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h194273b722e5a9e4c7d5714c68d682aead7255f0da9630a01b33ceadda4f1b0b110fa318c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h16be41ed5bb70e7cc1dd1d3cdb1753b61e6b958a3cfd7f3ea3f9b98d0207a8bc7a1f6ce4f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h601cb049b5218cca78b9c4c56ce896742e990321d8231aee19a53d06381e2a5c8da57875;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h17cf7fb74a669fbfefa123db6c79873309f29a6cf8859f7a591dcc4df0ffd693c7a2cd073;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h927369d9df8250855d2ae9df88cf6a68ae6591dd4b65596dd8cc87b2029f59c41d316634;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1299445aa6bf32de96767313a2c6889ae74a0805f4692dfc8df807882f0d76245a562b91d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h7bdddd35a3ccd99de31771b381424beacbcf89ea22b2e023556c5ed4a7cf5f1c6db2d1b2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1023b9175ecb08a255cde818486eda28dd6ef1dd0db721c45cce1aee013ee30136db73c5d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1885cd41045c9d7cfb502e5e4f22e331ba6961e7e0c72663137639d7b87939ba722637e4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h18f4b91b2105b8a1df64ea6deafaa6308d4c894d0eae39d71752d5c3df28936f9346022ed;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hbc29475e988461d7b5a56999811507af7c87362d15fa17bac4117e89e4f3fc59cd866987;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h66759c362bd7ef417bf4de5559d9ab385393b913f78a4943e25b6f8c6dafe5f6a99652df;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h2b03574dca46d448577e221210daa5f4ad3e4dad5bf6d6802b4933e358f661d6dc1aa59f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h127a9860081257fb0099423e7cbbc30df4178377dc5448894e653bfc00d16938ff06acf6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h2934bf1996adba2ec3dd3ce371169e10170254500fc1de2545dc3bdebcdc13ac332239d1;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1449b06e3a7d87f966b434e6b46452b46e4f6bead7efdd74eb593d54927fd3531b44f425c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hcb2f393156af3d0809c64b9447087d8d20a500fc484acb0e4082d5951c1e3c3fb4a76617;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1282888311cd559f6701c2aef7e0d9ccd1b99f045432a8aabdbb72d0d141720abbf0dfa28;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f5bc0672300744b3aa7acde84143c904c8a16041fa2f2838f9e285b2b5b714d4081c552d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h17c2976a1bb1f751fe4f6d014fbb56a9c749c1280ea715c3dbdb84588266fa884f80b9b81;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h198ad1861dedf2bdc9ba3a0da5d2906d12914226f5c6f70b44fb79d315c7c9844bffe9ebb;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'he916c5c2895febe8fc80bf826dd2ed49a25665da0107e15e07dbb8a82993a1fb703bdacc;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hdad204cf4774001b8eee99176d21c82d833e71f3c98843adf67d57be9d2fdbe4863278ee;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h156b31a515d2bd43f8f804537bb418c55b5283c461d4442ea8ea6b331d1185b213a98019d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h6f394b95e7f7ed1a904540994e700911d8517253dddd43108f03f71f0374644eb573555f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h69176355b0bfd8028faadfdf9747b6adbcfd0fff86e2c4892dd322468a838240e913fcc9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f4ab387cf7c35ed5eaea8c3472f82bc12cdcf080c1b5ae489a02f3da89a78f7c41cd244e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'he4509dab7a84ee717e65cb48ab354b92dafe352b0fa7456c9d583948329a50907419ce27;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h7952b7a412234709b1742265acd15168adb89151bc16472cd8421f30d1b0363489d9d432;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1007d7aacc509fd608ff79fa6890eb00ba48252fc740a4f73de32866fe5e939206aea9b9e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15b07024da35e2c4f80272cb92a70e1349044315a03f2ed960432ce67a9d9ececbba02e75;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h8bdff69f2d500b164133a53fb547cb8bd5eed182a976f666702f53dafa215edf0d03cc60;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf6f06ee1c14db5e9c6e8265de300109d4b72c935099b86db37d78f49f2c0b090b8152a75;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h85d2322cf351b496c021f5353c1a761ed94cc969714882285a9abd0442d0efff6b420573;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf93ba692176d3d46523a8361755e9b0de4121742815dc89ddb94180870c62d29e8b8dda1;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d9074e0180207ff9caa6e0da7753cbd8e530db2ec7bcb684b0da30f7de5ab8f577064c86;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h6095b599353188b4c3d835d1c58f0f3b8195dd430eab00584307275959d0b68e02c3b8ff;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h11294f921bce99d90740b38048cf60429cfe4d7552fde61aee61b12d995d200e05146c69f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a58014d8a8c38406016d2a13626e37b99f49692696734431b91eaba47273eb3e595ed025;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h17ba60768b66eeccc4e2d7c0ca7e31a9926788fc15b732268a13f376d3f979c9a76e9a13e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hcdceb99dee488bcb147b4ed2bb2e9506a21f0ab11a646c7282266101042d7e2940a4b3c6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc87e1d4b58a88a7825a064f472e198d940e679d37e6cfea6c812a3ebe2a410740116f378;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha001f7d0801ee4e85294bfcf44811c78ff4858ba5c686c0b19124428d20c97006f296960;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1cff1dc01f7e93c1980c5ce5cf59d4d5fc0ffecc42e51eec98189aa601fb6b8201b9d157a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h31a0c25a799029d30e8d1ba3f154827e31ffbb9f1297efa9c97e6243aa84b2b82aa55b89;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1da12d591f3f9a7acdfe9950cf42c1a8730bdc28ebd44bb523a5f9b835ff7442fa102efce;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e190add64402ca25b0f5aff851b0acbaae5f40226c66bc3029c31f6b69f84eff2d40e927;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h11136bd26877d9c7cbd676ab3474ca3a712a8bf473188aa3b9e1be82d2a820d03029c9b0;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1dc44306994ed0f80496e4a65386e9728dec293c1c09b673ce71475468c9eaa45ee6df05c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d68974af2624deaa63a56d7a0be75f6598a92f1e3f6e51818af22c0c43c5c15a54d7f25f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd5b444da738d3ab524ff8b1eb8fb13d968c69880f759f3a00ec4b4d1fa851157b5e4663b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e81f9d1a3621f1a4ea9b81876267076f38206a873cac356c2a73edb41fda0d49418139f5;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h17f6d51d3da91b4ebba459cbc72281922e3038fbf86556786991ee4ed261b55bebfcefa0b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc06c725c38922c8bebbd45717a3f2fc403091bbb43a8a8a32e4bdba90e8835984a96fbd1;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1266f56e997b650b5a12b41b92cdaed83465871972f51d2917c0bf3a2c1fc2d75931047f0;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f961172482d30175f60abca4ceaca30566ff9daec66f58b463785bae55f3c9cf1559525e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e62adfb29e2b30bed1ddd60781dd473a637ba652e5fcf59b4d248d94a10646109b209636;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f48887a4e00862196b71b0bd49517481d9d1bce8298eca545a9a9077c1f572e854a3175a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h62690dec70065e16b0d40d27713527415abfb0c46ef95b4eb8df31165c934a59f01d3ae3;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h115de9c3326afa6a653472f8a0df866679a7a1396796d0e9c15f68deda3ba687ba670672b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hdae5aebb1f9af381cfd56661ea7264e4a784390f69586acb2abd4c3380e1989532076903;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hec4c777389e19bc8fdd7f2a1a841c58f7e7c88e02080177b7204fa3ac3dbcb378fa80d99;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d744eaed7319e41da83a1d2c992c881591be707c429d2d9eea809af017dc2125de61960;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d0cf6e0e4aa494cdb758f957c5351428e4f61cbcdc9e9df50eff93da0e948f3e06797364;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b26310fc8e33750c3149686a861d6eb5507b51cc60e69d9b1b1cb2d9136de100092aa4d8;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h5f27c3bc7c3101792dabe7e3931c4bb105c397a586836eaccf718dfb992207e5de03b4fd;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15a974977b33e4eba3c385c834507e4038c8707dc10b15bfd0ea51f8e0d72369df59aceb9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e21fdd569b9bd92b1c0d28f654f1e29c50b57647f11c0abfabeb8d1dd95fc5a23c3769cb;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hac41a8da8eb42354f3bcbfb22d6d582f4c8e89338013a486b1285ba30125844d4277e1a0;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1edbde67ef013981cfd027105660f459ae8bb6549a08b52af7716ea5b8fbb4a6e2323a210;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h84e651fb0064ac78f89371f6767eae5e4f1bd0367a421d65ecbd9ea16caaaf14bd065b2b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h14914f5f9181b2cb7ec7f26d4aeadb915e3c804271f606143ee41a00f86da97eb0b228cec;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h62a38e53a10077e1b321d43a81e60812b09b1e80fede55530fa81e787155906a7c8ed99d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1342d12a0202437a797078dcc3aaef5ef76d1f139397557a12e0a582be41da720ba564b10;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb9e0a5c3f80755665e6f8c77bf434b4ec555547b2bb007b0ac0c50c532fa24bbc426281e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ab789bb8add75807b7a776d1ce8236b1a129975677e7997a6cf1ca5d1c2178b79ed89d4f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h17756b447082741c18634ad1fe3a80dc98a3145cabc01937cae656698d8d9a4d0dcab7508;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e404c0a70be8972ad79094be14de8c105453686adb9f60bcb63a8a998e602d84b8aa44a2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h7b359c40f6ec1df7dd9fea4a256802b27d26512a8fa2188c936265e2843d0e00f314c41e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd99db7be75262f92ab06386b50b6031ed3845c7d78f1939b246b362c6371215e2d3cd89a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h8b3bdbf000ccc22904b74e09e8cdad9bf3e8eb257ae29e390142792acf19297f99d8e616;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'he62cfc15fef21ef1f781500bf127ac856621254e7755056ef7abffb8725dbcd2c1b955ee;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h51afad4e3969cdfc6aa03452933548ef40d0a89216b97f4c30a38503b4dc15aa5cb2f112;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1fbba9e2c84a7efc5933e0b6544bc87ab5831874947775ffa51cf5e2c6fa67a30696de458;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b1d7b75c8b9b5e78a47533237b1a9d397911bec82c0f3f007c00d390870513416808bad3;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h18b95d4f631f30cb48fe269bc8077f730d71d448d23243189c9593a77f9e5156e29842771;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h151f3a9dfa9d29c50fc885e85a402e084dfc00f0808f5b987e9bcfee71788e2243ba3f690;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h707a05c8e76ceb1c35f9d1c793476ccce7ca5bec0635cf27ec9ceb34425dd3097345a6b0;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'heec30312394b282824d20df1c1c5f748fc8e25408c4902d794d7cfcae1c359103611b505;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h2ddcc62375a1a30bdc02c02f2e110edf1fea36c538443d81884a042fe61d4aea78adb2fe;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h143ab9980e41bfecd29f5b1bc890e81bf660a87f433df37cb0715a919642794aafa91eb49;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h4b377abaf3c5098341f2fcf65e096d00f997c4349caaf207f730d4fb27ba1ae8bf399e78;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h621cd8166b304374e1c15cf5f740f41170b2e11d992717c2b39d360880837d98d1049474;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h9f77e510a7c508568f474f5b6f7d5eaaffcfc4a54b5876e0d621421a16ddd06e8a95d0ae;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h3b1ad86c188bce29c6354876f43af27a1ca5a19979aa560c7e0c728cfdcc582959c17fff;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf870592f677627882f15efb59cedb48143454df8ada0cafe50c04659773fbfbcb27feb1a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h19c0ae5c4d64a7f038c1ace7490bc680574f16f904043e4248ae7ca3b4686680a4bbb9097;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f0d52d760ff69035ce2c63d6f271231b782840fe90001124431581d469d0e91b65c1ee9b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h86a937e02ad9d2ecc6f8efdd7bdeadac36560d71dc5ac291f55a301d51e7e7e3fe4f46b8;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc87daac38a3aff9519e2916304d872a93426e15877e45ad65de06700105891b25fc2162a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h10cf8512b96543b7c3bbab4b7ad7f7518f361d758b9f98e7e0224d8f6521bd958876cb2c7;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb16ea6dddfd66c26bad832312829b75dc3275b5aef03639c9485ecdbf21b04dbb499bf8e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d2c9faf19d04c4656774101f51140819d6d78123196164d6ed68b9e90c0920615125518e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1023fb0933bab4933b7aa62b091b19f9ff690a2e9d7202c9be3c7c862e3fe0eab1a90e478;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h118f0a6bb7b15e0b4a8366800f054053124f280b50bd53e39f02aa19a3acb9c484b5b9974;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1cf1fec5f779c611b30d76d94eb63194bbe077437373e7c0e2735632fdb582ee7cb0307e6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d93d3a9e227848c977ef60f8d7038b2d58a9e55af978b59128537a5214123267c26d78ac;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h11c1c624295e4b0654f0d68e37cfa9c3ada825c93fa3d20b7af8d380f3a2ee1cdc77e1fe2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h5555393ac17a9cf75e7db88f1f4deb9be617479a947f044a0339a5e0cb42d605ae11f615;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a5a76ed49f2678ce618b5bbadd3dd6cb1c0368cff6f73cd068cc24882ede96983e403a69;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h505e294abd376ee35cf42028a9fc3d04876401be18538061c22e76093342db0bb7a757b0;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf3262656fad8cb820ddb2547513c3b4468d4f0cf4b8be3d46a38600818d5e221339dd9e6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc62607f967fcf34376d330f74c22e23f54d1260afb9a2410a89757e5e04991b0d88c59a5;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15e3284eee1b5c181ac7631a501e6d1ddd495f4cfa4f1783ca2f9af0a73d394f38d69d4b1;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h94942a69b14ec677b2b67f4bd6474abef1c986c38ab339a2c01eec775fce3783a66266d2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h12e2682d6662697fe7a7fe6c3b06e738180a4e122c9a415d37e3325d9fdd32a828ac29ea2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h73b17fda88b9d8674ced843476095e75952a490c36020ae2c6c097ed670233251ef8c09b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1151787e5fb06937ab903cbab9ba2f0044ba07a2d1be3e0214dcbeba54236a591f05de2c3;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h119018ed562a2e6b4e4a62abf1244405807da0d397a60dd9c53c1bb56aab99ad1dfcc086d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h17907d8a6c34b0bc22fb362fe023b342a37f141088ee30b0ac9a7e528be90d654683121a7;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h166fccb6f3b449e1afe72a3054f453da917789ea88dea3cd98c07725ee324d0c7e6a09fa6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h155a3a4e7e6472b61c1dc08251e35506f42925ca3c678ee250d1ce5dee8ad92406147b5;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h147f19220f700a65ff25d1ee224f529977a3ba1b79ff99688e8adacf3c935bb3e69988573;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h981b4dcec308d0326104b8840be2d71ad1d14823666927c686254cab6a3996cbcc231897;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h2250a69f56deca59e86ca8dd8706947033976923db439f36be0a4549e8d0b156fe75945f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h166a28f11d28f03e3f3cf68790863665cdcbe98e99a4b515bbd58568229d2b60239502d18;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h12e548810f444dc6964605fdc31003365bafe588d2d1b71464f54604e35a1464136a2ef30;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1187c9f0329130420b099700c17a64a421518513f5ffc080bd3d1cf359681d3a9142b5817;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hfda882db0a0784a39d7b28873bf4e31a8d6524052e0f53827901d9969dc011806122a80e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h39a15c58d47e24afbc364ec76cae559997a90d12ed96c0900f6cefb84495226f3e8207de;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h2160c25457da01cff3e1a6e974ae21e89581edc9b3e5b0c36d9998a723650ca1ebd7db9e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ca9e32bdfbfca33231a37bdecd09d6165cf33ca5d2260b157ae8f873f5f8c7a4e8a5f98e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc26b5118d6ccaac8c6c0302754153e27f88bfa8d3dded18bac8067fd0ce3b170812cc96f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c493240621f3247f7f949820347f9ecb3dfa9a756d3a896efeddd6a646bd52d6a30fd29c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h19d0b256ecf609825b63a4bb953a6a0d4ad9d2a2935fdeddbbb9190cc33fdcb932a5ac3b6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1397f2852d7938190f105b3ee86e9b92c28d922e5c2b9bedb4f4a658ce8c8072c66a6af9c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h176c44b25c07222329237bdc91f8b621edc4a89fcacbdae1d46f46598104a6705a4890f65;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h7d6fb2cc038d95b851e4b19cfbe793f14833395df21d9c30d5df05f465560b7c78d4b687;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ab111b1ccaa34261982a48145542723e9444cd15fafb1309234bc59b7ee447799439882;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'heabbbfe054140856f158fcc4accd255a0a4c09ebb6248a2066b668943c45115d8d562db5;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h126054c8daace299c1d9306fab29994ea2dfc53df8eb80b22e8f4560a6037ad595ae081f0;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h114cca7026466825de62325d672220b522cec35d00ed7babdb9b978da11535acdf350df82;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h12884fd3a13d08aacc8125ffa8d0f95a5c39492e42a07cc023eb847d124a2398ba655a3e7;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h47b33efd982afc743abccbd3cb5fd27ee65227ca4a849a8a64c740830c24787bf3952455;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d77a54b12820263295e2af149b4248a5a17d4dd32efa5306f5e1f9d63bedb0ea15e18590;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1acae3c36b7be22a6d49d8d4f799318dbfff8e1e3fd072b7154f8a1f5dd9a968a22053ed2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h6100a663a09b086fd65fe3dc816bf4fed18275f9f86fd14006aa2b47485b074d771abd59;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h2f04419abd1d05c6466ee7e6e2227ef609c610bd2ed0febc81bd8809620a94139e22ce0a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h180323d5ebcb4f0d53c52600dd89f864b4e5ecdeaa669fc5e8fbcfdf382d354231643a46d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc610a4dcf7fc8af845668d04176ab0af59aa4938359814408caca0659792ad73a630f237;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h14f7e25a7621bd6c39a19cb449dea4faad115fb99a59760874f9898c8a69742beee65694d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h16a8ff3d780e645fd7279b317688873c7747fde8657b8fcce1c4950605ef71cf26b2e0fb;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1bade9743fe56cb640f15984a21b1fd145434d2613b94176d7d67b2bbb1dff4cfcfac4e66;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h81b1263e530f777fdabfa4261ce81d1bff9634739dbf7316deac2914dfc39d7dda62126;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h169e29b272e5b171f34098c31a84249ad2dcbb9777f0a7edb1cf7e7fb5500f1ad50af4588;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h941377d2732991fda87aee5c02e6c41799ecd42ae50de1919cade21e05602f0b62acde6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h10b0b2919bd28f555830cb5fc33c62df64ae058e53f0b8075ff84b4698fb0ceeade88d789;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h5459b898a2b13bef0411de398d0b9705b33a0297fef29b2955225991b5745938462dfdbe;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hdb3ba82e4d1aa466ce3c3824e2dfadcc1abcd1843436de00a958893d996fd32c0d3f3152;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'he9465b594610d3a9f44f7ac779602c0ac95ab9e5a3adc78a975d71f24f24996886a824fa;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h12b1c0fee4d310b76c2ac8d567d7b9099920ad1da433f326c35a5af25638cb0dcfbc02b8c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hfe9130c0937c29e06597edee8b26548bad5b44c6da3fd0b320c70dfbea51aac67b6d6390;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b426e1b82eba88f6ca798c6a90cb58e6d3ff42a6d5529828ec19a3a712fafb0b2d2379d1;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hbf385722df263509161aeddbe996ea7a0955d07ddc2b3213f6abcc0ab096e774716a4a1e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h19890db39e27ff0175b858ab7a09c3df0e8f357cfbbb8d7fb3fe33fcf52bd11d2cc204908;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1073e120d58a7bdff08db263a71ffe0c243669d3fa83558fcefb117f89fb374b9dcde6074;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c45468462d2a155a426d6998d338ae297501e743903eab9382228765e71d0b5afb4c68aa;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h192e2517058d14cea45b821e25a06f61c07395dc546c9bc5fe80686b8df8887d66271b57b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h711f40d7f9f257ccc3e8268fce82a6772c8ce57539555e9ff72b4984ad104fdf2a15af02;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h4a792f036687c12c49a479cbae59a6f60fa7c82004e87d906837f12671190a98e2897256;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb5f4cee837c7590c66c1138b040c146a92682220d711c72f9cfe3cafd59ffa7200020c1c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h19a58637cb7397f69aa6ca49cc041268e8adc52edbc09936081986d82f97da911956c34af;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1955af7be06cd6985a7623d2c808b3a561da7be268e63774b8d7df9f1fbea9b6e8df9966e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h192bf60769bc07c58652c60f19d54261d580bbc4483edc245b5f4278ee8bc6c44484b707b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h6dd33f1423145cdc95eb270bf030783b1cfb6f8e145ea7bf5f4eebefdc1a1e2dc0819b4b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hdbc9d77d599fa8e655efc567c8a51a3b1dfcfafe89c652e42243f48a4fe3317b9f05add7;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf1664d5bf66e174ba229ae7dae2acd9ece21475a12562561cfb4d3e9a2462a49d111cc13;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h95ceb79f18a57894d8040550a328e7e3f51bae118afd42236360588122a8f850ffda557f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb220cdcad0ed39f8387a1f161e44a1da31bebed6d9312edcb0b8c1599531737477cf0b88;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h19466da98e66bf432dde8bab9989fe3ed7b4fce03df8c0807fd9b895820f3dc182d1915cc;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h184c83e132773cac9326c172bd2f7d50a0d0db521a68e853c9ca631c6b6098a97a415b29f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h10e9343200ea4d9e9bb2b6b674f28c7c8aa39b8882173ceb4dfce55faa7c79965a0af713e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hbe3a703551c5708f8bc67bd2d4170a7b89a55b01daddee46290b79d1b1e10856d4290397;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1bff0ac34f2a40b6cb200ba874426a767d35b32c4bf647853ade722da1fc0d8e758a75aa9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a68ee17c26e3553560812ddf28d6e92c804252a70f7b9a83b635ed23a835afa0a1024d91;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e4856e61717a9ead2688032a5e10d00f90cfe6c20e7c2c8df4ab9ffc11081e8294380ebf;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h86e1697c9f4093820a254fdfe985b0ac52367009de7057b72963296024a2397e88e1dc3b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f72bf5c3a3cb65b25205215f425b6c710d8f145e4298854ffe72bdef9a19d7f0025eb4ba;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h9e95930525bcadd5548d3c48b728c98c59a53bafa999aae0086b5f4e360025fee8f9fc0a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h140cc61884b1490ae99ac0ba244ecf729a7e6a3c19df1ba4e5f60ca1cd6fd77a3178f20a2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d634103fccb2a5b6a60d1642b5814d2e1a37bb6a2c6c7b45b6849c352606cd63ca37b6a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h2791217a1563a567b7c54ab3119ca0ac7f58d0d03ff3b361ee4b375e31a8e92379103f74;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hbe18ddba76bc3fa4f8fcc81c5f69ca67cbc854b02e0b39bc7c6ebc0ce43c673419ea7fc8;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h68fae4fdef957f88078e2e521e001b9b8313082a98d09c4972daf105fb094b867c9c7e27;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1be426332d3141e1278915f786a95358bbe44f7a2fe8c90a1556933c6bf501535362f8e76;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hcab2aff41844b971973864eaa94d0846548b34f03609eae85066e7f19d850ae89791be93;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h19bce6688d47441c39b59dd0a47ac1e47ab48f7d78fe4c9e583a84266e34ea3948c5a2c26;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c4971adba78511aa208f8d2abdb0eae7bf6711bfb1a7e10fa7d1af432cfb28c5a5737523;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h10867f46a41697e96428797ede0e7231b2b2d2eacdfa92f5c01057f37205d0144c733dbd4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1833c6597db3f4609a96050ee7597cd70569bc24ff0fbb9851c85ab60243446dca5f8d82d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h8195ce38faf03d733bf76ec1e8a5d94a02b48272a26ef6ce2cbf55aface70559d0e019b5;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1bcf3f3908759647a2a04e3f0516c3daeb8d2e1286ee6aaa8c4cb8cd1b228982dcd66bde4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h100e1dfcb32e35727f02b2ccc169ac89c917c24fee5bdc2e1db9bc4862cfd5a8997be8092;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h74f33430502382502e1e4e7d118b9465551dba6533f587dbd66eb4dabed38da919078b33;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc161c0ac6447994766dd99a24a7e65f3ef2bd49b144e17ab7e000acefd2011b23706a650;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c1e4ee6777c63ca26baaafcb28463b9eb1e62ec5eb9751d7ad0ede65bb8412d633e69e54;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h24265a3e42261de2d8f60d4adf78646e499dd81fced4c8c0769ac4f09c3b05a1e7ab4421;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hec37c73cf06f37faadf1576e6c107703f73b1afe8c361c56e31fd9553b52091e73c134b5;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha0eb77e8d2494f8f6bfb8e3563008b4f51c40740d2e47b2575f1db28752a7367aa6e3f04;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h568de4e77220cbdf6dfaf53a55282199bce4e20e6b65fbe27d90c37eac5d65e699f9e697;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1beac250684c34077c0be27acb9cfd65747bc40777bb0f147c9d468ca43d42b256ef64fe9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1bb673ec70bfb4d7d702505525d0b40d09a6fc7289e9ca659559400277b67647831ed7de1;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b52d3a95646544ed069ce6178a47300b74fa42edff482b4c913b71279f82f7312966437c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf202767d6645a7ebb4d75ed15356d87c3e604d480cfe1f5316ec8aa0c9536e018f12653c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e10a3f2af053bd4289144416f06bc2808a519721f989a6f462f593368e4450aaafc1bcc2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h14aa71eefde07a5a8a8caab7788425bb3373a8f2170ad4d6fd3bc11f1f8a1cd400fae39f3;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h5db9f98a82b31c468ebfe03a265c8f381ac47d58b91a83ec277a5822bfdcc37ccfa8afc9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1af7d47309b009314987fefba802fd7df29bbdf3794ba8ee8a3ec4862a9a527735d67f98d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h132b766d3024ca292bfedd1c8a4a89395a30aa69fa086b6908e0bbc9c718d4cc6f091b096;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd292d64d17265e2a6a46dfb99efaa186a42b8cd542b6cdd6b6b5f946b2b0842349b7f969;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e92a511b5620c729b5f62b7994a38d901e2a9d725b964722b39435fad24ed2f65539a4fa;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h12b93160388bf59fd47dd1fc3b85237e20cb8a5b4fe8cfff89e705a7f3c940622bb35a0bd;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h9eb95d19173e4d20cf23faaf2471f06f9214502f57435dcf82fb70854c2868916d9224b9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h47f7d68c8bef84e9b5478c60d00d58bc6fc3f8fb5a22b8284fc927731d4e821b488d146c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h16907cf7b9599c75436385b9294752ac60af2462a961387631dcaa84d6c4c322d649d1c0d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf72dbce4a217086f4191bc173100def5b3ff630332448ab8bf9415d737622ccbcf738e4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h5ed55a3e81f400992d01f8be067fb460b42230670b429c94dc2818c11baa2f9fbae3892a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hfc510a2e08ff3bb1fcfffe76e2e6bf8e19158fe14b6fff1fa9837239ea5f3c8531aeedd0;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h3c29ee3fb361e55217eb73aa7310f08bc119c1d45cd9a31b0cdaf4ae65b32b84bca62a26;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h153cdb5db24886d7cac7892f0adef28a2f43da3b7b9b311f3ca8424da904693d1b43b3ba3;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h13dc28aa78ff626f7ff70746a273367c7e85e210602460a5f6874831099bc8ed50738cc12;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ed8210a94d162dd7dbfdba48076ce4788eb75f02ac45f995a94876481358d58c78ec0fb0;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h30910bc2266dfa1223dc72f159394c0b9afef5170bd2e5de11766699abd5135515848060;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h2e57892ac7bfc1e9317f37591477b04837873b5f797b7f7cc5ab5d320687a1cb41844475;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h416e59dc058b19c2169d6a6858347e6c6fe867ba7981b502ff1e58e08011e8b056601471;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf5b12ebd9ca9127bda30a21830a8c74de8626429e133ab2974a8158b8592829f1731ea76;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e131d55b6ff4c9495c107129367493bf304ec6df4d589e48875742778927a1e892a74622;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1fe79188bbf0fdd94b15ce1b3c9be0f345876f084f6dc9caf5d0f87f80829b337f174ec5a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c80c055f4550668a0059982161f994b677c825073f85733c7b4e9364f0e6550f25edc4fc;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e04055ab4e77037d5e8067e89d76e666f03cf176a0f33b9e86695cd41c6e180dfd197140;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1059e60e900dd3129dc899f7c5cc15663e41b3f9022804f343f98c6a00c1a917528dadcec;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h11fe705baf2e4c68671e713f16760c03be8d12538f5b3779a7d361f6359104219a528362c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h360b283e18b62057b35900cbebe46259dd9265ff8acab26d27c1c5714619b9d8e98d15e6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1261b3e0c8b543d76fec616f28c837ac7ecf515886c3857ae33099c00aed4c97fd2d82c36;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1aa04e9ff45981dd746d72f6e55e32f0fd6407ba7ae1f968034747ffd54dd8274e2ead8d1;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h16df2c02e1be798054712a566fa8f2fedfb3607d1def3c2433d3150fa21cef73f148bb8ec;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h20cde6ecc42dec56f0169634cf58b5410f89d66bb4cbe2cec7d469fe7984f4ac73d397a1;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h69dac60f8457a1775dd75fe3a5031c76ed6a604234178d37cda2787207f16cef2a2440aa;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h8075263617e26de9e08c68bfdf0deb91c2d605e0503aff120054c2e46db34aacf44a5a65;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hac7727b257324cae5df98ee00bea388a45484315b34cb6c01373c2b8a669785559d9aea7;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h6f00fe9c680de151feea2aea12e9a3e572d77cd862cf577c21f7b2be269531fe84ed2afa;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h191bc62cec52d8328692010c29fa9f07c0a6a6ffccbd305c31c90e128143b578d17a1da80;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h54db7be4772922785fd6eaa7ea98907eaa0ff8fc4cf8dd48d718c54d5c53c1a1d6625818;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h68540c42f56501dd0ae72e5078779cb39863e16048b07d7ba51a6d5f5f4a5f2f9b53c5d0;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1de1f703f1430e7e5f15eca8fcce25c20714e7c743cb6692a991b13c9ba24ed68b085e404;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc8966288c9855ceaa9eaa9dc9efc5201add1ccbe677e81623997d1fbbbfcb5fa5c2206f4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d184bf6f3face966f30e5fd6754de21525263caa0661ddc6f06fbe39e0de5253aaf8bd35;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d36628be66fc59ff4795338e50330b07290aa71cd279205a1a8ceffc9a3af8ae5c791206;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d11f41e5e37f904c0f481f65abcee7bdb220c55e67c8b8dcdf15286fa6afee96ef38fab3;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ce9c964741a956a8920e104683900e8c1d205084e0b2701beefee5be07695075c1b30c91;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd8716ba32f379d3c122b0097ba46278ed61b7e8b8a2bc8ad2ba61592e809fc915088695d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h33b21bb0cadb8dfc1ff7cea2d6d190220b630e862207bbe6ebe13604f3988f13bafed9ca;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha6ad55cbf951afdeea1338bf6cd537aec671b48a1b3536916c3ddbfdb2d0bc61d9db4bef;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1af86061453c30254b39f438e909f1550ed14ce87a27d6dbfa1a8b6b28f0f944ed65daaad;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h72209e717a068fa5b775a201cffada6012863e0e7c57a67ccdf83b303c0edc5e73a7bdf9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd57c652ce68ab427b02a939c40852768b71429e2c4acb824b273c23a50955ae49479f267;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h10c0a87a8d3bb4e538033ea8707fe37203bf3152e36dc2ba30eb507cbd8e4c1b1c5b50c33;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h2d9daecb67becd2522017dfc46d0ee875c4c8208698cd75f74dc196e5bd4bd8eb39bc11e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h19e1e2dce441e679dbd39aa0cec2b437bb7b2efbe0f24b9c15745f2e0074b569b5e7552f9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e5b1be8e7eacfc980ece9e6cfa83576ff427dd785c2989b7741484c1fbb317bc92c53833;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15d045a7641f6e25385247a4eee54a14389c84f9179ba614dd3fa2a11a66030a7c2bdc6d7;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ec999ab50dcb68205ccc7a540257bbfe2939426088e6f483909df9fb8dc50ce02e47b594;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h182edcf936588c72d90fd3384f7eac62345bbeaf2b39f235a9c73b49972655b7548f9545;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h924c5546bbe6881ecdc2744dee5c639d2055e1635d89f2dc117c3a5528a6446aed16e7a2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h87c85cf72a0e321d63f385df092f29afe27c2e13dee66296e0411b7eb44f349a19b6200;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb55e2806e7a930bec62357300563ff08f9c71b45bb581dab9f22a0e4a372916f9ee50838;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h3e839fea5eedf5da377073dbf4c59ee5b8f65e19a274ba52dd8bbe808a4a2ef1d02d4f97;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h20845a803e05cfd92fc7c9992a77aa455a0ddea20c4aa0ecdad2699e321bc06d1a8664b6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1585788d20233c98f3d9a4b9e5d4b863695a15582921030ff39c4459f1b53a92d378a4c3b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha307f769945e515b88a1a1929970d23b20f0503ba32558def3327ec1dad5eacb6ac9112c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e05bd0ddacde234181c937f321b1517eef7608f6d168fee4e393987c497494386a6d7c01;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h7ba36b4de934e8f0431fc88b3e48f3a0d2d90842e5917279a46ebc4882fed11654222e95;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h121af997b11ad998509c9886f2697594c9f44c2902dee27f87cd13ef04a849937bea63ca5;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha3ec21e5e859dc40abfa06435cad44e51a3d748e0a60d335a425c7b845f23190bcc4853e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h515108c233348407dc4ab7791d278c0d085a278f9d9a9d9ffcc29509a3b55232753e2298;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h55e893804e8c71781d40413dbc8be2d726ce2a1ec09c3b67ac610531174acb2577c08522;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'he4daf5b1644858c584fa082c0cf8a89389a7a54794ef0ac2aefa8c92e1bad1ecaf5f28fa;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h61cef69d18501c532da95b7271c612e42a7987994db9098a649c484e699e22b3b094aa88;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb2af977b990356ded607956a04557a9a6b8f295991143cfc912950258ce955f181f528de;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h32a8829c1a7b07d07b28a8530fdd5921f8413681e84139900c869e1110efd67ebe025d2c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h67d157070503589c57bfbaa4db92a193edc97a126bc9a48610ff327a2e1a6a0d09bf8997;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1947505133c6c6de328a4ca95f5053fb3e1eaae9e7ccdd7da8be75288b10bbe9c436c31b1;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hfa3bf18a3266c99eb8eeb4e65c36f45cf639579162d998cbcfd71f6b4f6a7dcd0dc2c85c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b5017d30343e322356863223b3b8c2f87f4ed6aaba15e8af6dd57ebcb12b04471fc89e24;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h18fced7c5d42848da9447d6b583d5878977ae7c31b2822c412ff3d052760e475e361b4452;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha261880cbde9f0dca9ae56be3b34886fe9b5957d9187d919f9aa4dd22ef17e669bc3bf4c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h89d601aad5fe113240f5c742724716b0accc17efe9285d1d8bf900df8d128c87b343e959;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h5972ca357afec6b8a414cfdfa94a19638135fc21ec59009dd13929e8dacb63611191ba98;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h153ced1f41f02add622c36d4e3c461e947b4523707e4c5e4f7a9130699673de197de8b1b3;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h10aa049edd92bf37ea9d8c52b68539ee449dcca0915886263d38d15d309233d853042bc13;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h18d9855c9117792aa124cad088fa8864a18fbd312381a91a4ad62ead866c6602367787ed8;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b992223334c7fe20ddd9f3f37123c5622c24db98ce7c66d6bfcf54d7ace0fb0c4617db75;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d4ebb8d0696381d5ca865edf2e895d383b3263c4cf2f5f0f8489e63af114f6565e3f8d77;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha2a45e1bfa48d3a8ff40c812ab234fb1b574b1baa3277533ad70c338ce7642825ab497fd;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h4e3f5f2f84b3068e45534f2fbc5b889f10fecca7ff83faa4337c7658fa8b853d97df8359;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h49d842119157f1c5e3326240626b669685bf8a6599ea9f7ef07090e990ca80bda823011e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h113f83aeb0676559b14d10bc8dae79a38489b96f31f825ccd62845e539fd65c4c89892427;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h43ae489c1d7732f2cc1c44a837fcd4bba60298b95088ac5d212ed4cfa31007a5ac57d885;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h10452bb175234d327a5e3348a6ce2e48a26bec02d7edcb2314546a2bb8c27209bb6806a72;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b9bc60086be8853a867d76c1cdae429db3789b1291ac517582871ff5ff99f98b49ede978;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf81863a2d118e9c31e37208f69f6403c7ed751d06a54cc5f7dab0f7b8f46f942dd6eff26;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h14c3b47034b0278fc6cd6f8750e1bf89ea5c9286a2055d5b6129102398cea0346f453e975;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1075f786680b705174e8e91c349e93c67f78ca632c614b77f0f9e97382be2fb944b08194e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h7e06f35077ebb006b8e39b67e884ec0e35e2d6e6c937ba057aad257a16805fa6833e0d7c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h901617b7fba93a31a6e6fd849051162ab1bf3aa335f8443c9d83904e8ed31780c2dc7c45;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1883098d6d37a4412a2958076c23f686c9f08e38ec6ce67ff15746b21d9fc2fec9e5da85e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c66ae11019748de819e5201a5277f4282e8951e633b4cdf4ef51943aa0ff633bcb260eb1;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hea589a465f8aa89951af017af5fc92e9575a978f6851644597eed15ba11bf8a0bbb9d2c9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d49b206cccd8b8aca9fb34f07b6d24a1c12d9f60ef13cce8bc2d245971444a600005112c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a1c4dd2c03b8bfd0ee673350580e4f9c140428bd10bc892cd0ec8d71a933d164f8b840ae;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc186dcb78cab06dde1016da29746dee5d232a9bb3dda8f8da42781e833fcde46fb2e6595;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h119542b3eb48facb924ae223c59d6cb7d1b3d70da43fcbd789755af1b5a364e73ccfb01c0;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f54d2ead2fcd9ea5a4a80b71d6b8c66198523d51dd4936e06f2f58d349275919caada7c1;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1721f3a136ac2f2d99ed1a5b05cfe0fe60273e1b080e5fbf624ea7ec0468fb78895f116f8;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h117a96ea99f4f33d3e9bcb775118e9284305965d5e614d86b2eab1f35116f3c891afba27;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h2ff46623cf5d67bed738331f862cacff59e465b42bf68aeb9e318e67d804eed4fdfaa730;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1eed38d7b5b9b3e70cc257c1be1e5ec32b57e15133a92746d1977314c9d1a072eac327418;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hcbe9004c7d5a4097ff590c7ad2f96c59aae7013f1d3dc533ab2d72ce42572f40f3e3405d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h12da1ac63be3ee6873bd338644ae5b08f0aefb1644a636c929333e23006137d01eeaba4fb;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h103bc00ee22084182faddceb285efa2b140b6b864d4c1d9522d5ec07eabfaaa32ddac6574;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h180cc76b521a58d8f41453b8decdca1f728462da1b2c452affbb90e131fa12bfeac1844a0;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1228bae2465625a190025d13b474c219dc4060f1967d034d7434fe39edc3ca97b032b05f3;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h87062763e0543e11faec452c4d851e279c2ba89f4bd7439f74bcf38f0450f6d25f6bd6ca;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h59572119eca9d5bb48f57c8ef74bafa62cee537b19e965e1e582648e17beb0b7cca18583;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h8010279f5ebc819d69973eb09fc396d391d223fefe074f54a22e6721900065b9445cdd59;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hecd99d35777ab5c44d9df3f3b8dc5d4bed9c9715620ba40cece419910e46ea874e67ebf8;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1dfea0443566b692298ea45a6d4881f9e94d98f8867f3c8ef34014a34204b8a117fcb7dbc;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h3bb5cc6efd01e05db1b30ddffe26cec46435d5546865f57406e49e30fc077ffdf488eaff;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h121dcef71ad26f93582c1f479eb18577dca638a0ccb91635f4d0ac787a0428a3c7744ed13;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f145fec304710d44417c28e594f886577a1867718dc3e85f4e03a01ef4c42d4577f42e30;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h98379b635b8ea5694f1caf9d146cbf107cf5a7e40fbdfc02f28a36c3db0b1b4ce63d6f17;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c92b71d2e434cee7422e6717a6dd6b6ffccba12af83b16cdeb54f216a8356e63a1999d40;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a042662240a303f0f979c526b8e60eb1ca0da9b536ac0ee9e063cad7be9e35adaf9dcf9a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1cd02118618006dadf5fe3ce5e857485aa777aa913bed9a7a2255f584c64f570a715d13d5;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h4f1011cb9d7ed3b99b8640e57cc81d1c8e7d37405eb32f3707109cad6becf5daba1433a9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15bda5e46f5f6087f39b9c2b9f025922daafa79134f6cf8a128b7e1bf9dafbe9da1f836f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h4cb230bdbaa8613d2a3972a2b77aeb3d42a7c8ecef3f2ee3c5737f0891058c70a35ee4c7;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h41abbc5844c15923b90670d578c0f513bf9a9d4773bfd76658adf4d28de641c8333ca970;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h4855a405e891bc05bf01623c8c3e0bae4a108f316c069b3ec9be8df3ecfdb453139e3a31;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h150f03cc5c9b115a341dd5ea25470ccd375d424017e6e0c0c3b4b139bd40738111f0296f6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h10636c3a99ea0ef80b79cb7f0f826e82b83dddb8c3416c974530c1b4f27e7e8cc926c4d5c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf040ef3a764a331a147f823640f83862657612e6daa1e1c15fb81ca6c1447f98c0f65764;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h2f3588b1642f8ef748b1a87ee16b84cce6ba9ce2d645bb91413cc2638efe14287cf2f41d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h11abca51f6383440821f064574084ec390d9c4572b48427f2a2f84f0f908e9623bc591871;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h133421ca5b2e5574f2fd1ef867f37791f39342b26123615dcfc3af50fceb0e6793bc0016b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hbc8ccab9c6723450711b6ae8f8a980f59d21e1a77b4bca418c33f040c975bebf3770b896;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd05672425332d9a7e6522469ce12aa98e89aca5de89245536d80467f8a96fe12ff2fe76;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc92cd5291a934867b9ff98fa8b8c6e05cf02bb35f7b7e75438dfcd0066f8bf6a722b367;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hce2278b820f77fa977e9bb85633820907290d54de934f3c221edad04035040fc00e4a836;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h14d0dd9db4eabc9cdb7aeb82f604bbebdc0a0397d1556232a4cc431e0b0aee893fc6ae71f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h17bab376aae4c9e7d2b7e069a3db924e56a163e44cb1b4b1f43161efcee9d83c5e6a39c1b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h17a20b1853f4e5ca91116f2da3657b6617f116f561e1e2e4a306621640ce0c67a931cf48c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hfa621bda3eccbdc3166772332a0ef12ee8a8739450dfabd2d076a6312fbd59c79d6bb9b0;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ad7cd06e7f83e4eab39a3249d677d4fa05ea89f740118e6d4de4f32a2eaf88c98987ebd4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h2df7ce82353562e6d400a23a56f3d91816267d7f112bc8ba0c0669dfde0373e661e51403;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15e2ad7b7dc8a8d9ef8bd0d4d34668887d1df407c045ece78959d2d3674b9a1581a248561;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hcc12b56476cd69625f16e5c5c80ad87cdb9629668971b44c84102ca3008354e23b785cf5;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hfa586edb9e4c40b5784d706639748b6aa9467367fa56936032f5a4f288514052674b0b5f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h14bd0b8b35327cf1ab733a1df16909b1c7365944addf90931eae74dbb01ab270431e45224;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h8cadf9b39c925846600b30c4ba638a67fadc49576598348236880a5ef28189ae54235f5f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h2dea90ac4bc695a5b2f850a316899ffb2cb799f7d0e87ec105ba35639f2961e98fe01bed;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hcaad6a70394adadd0688bbe677e1a53b51a034dd5c315d33acd883ae0f9f6d16f4f3b89b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h4b6480011de46ece756fe9e4925b79b7e00f365a55db8a20746a38e85f87c6ef03e44279;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc1683e61f5961711296b408dc905af168daedb881d556309b35206623848a78304c665e3;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf0687ddec36c23acaa0347863857df764baf305a5e760192ea4f73d50c6118ec636ab1ca;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hcfb9aa5656215314af82c31486ceec7698c817a1f504b1313fe4979ec90d4f6458b5219b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h13bd526e302e06fa690e0d723cb09edf6499b909e47a2627b27970e9106027b8545ac4dc;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h11793254f2b264beca8396a25083f6286cd035c630c6693ed2fcf1f8b66c8b231b2320dc;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h13c5986808a14a1ba7918d285577ef7b89af0b9c2ed5c372a6dc8cc414a9030a4451661a8;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc052c3021d5940050b600202159544c61175e473487155ef254d07b82b7072ecba2956ee;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b84bd8423d019cc1d65973f8b6b7e5059284a81e25c6cf903f7c56b6f58327d0f0888563;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h166aca9d84518fdc123d47d3eaf8b3cad9a3e2cbea12ed97d7f9aa62f533b53135e2d6f15;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h8207afe7ebddf9485d5003382845261c1ea2fc544496f0346e64926b61bb36c088bb4929;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h12b13426e86b8fdb1730376772b0e4a46e66fbd8dbdbb258da5e026a5a7962dfd5d3cb600;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hdc973df3575be7e6262c51e7d52962dae18f50fe3978fc0de6d0170e21e3ecdad27e3738;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d02b9605bfad501e0e3baa0a8f7a65f8b6ae5d58295c11b4e603101bf553e0a8ce0ef68c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h275b952ba998b507265a2a820f314d041cfb2851bed865c3d40a4e92dcff5e5df1c8a6c6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1289334ad657a4a0a5797410da3334e6ea79689d222bab6e939e332e7dadb549a341789d9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h672774bf26cb372dcdef36c2f66493dd138448922dbc4117c1d325d3f199d8e4320ce49f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha8e3f8fd1002fce7850918e0e38861152e5813bcbc117bcce5973f6172e83f15048ad395;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h74ebf2134fdcb33cafc9923c427596bd5468e9da8b33ff8b78fc2dbe5312002abd064bc5;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h788de63f937506370e07348f6752bf0ed507043f3a3e3ef2c8e9dfa0edaa3e8063d6328a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h12f4c86b85942f2192fff02871a335a3251c31912a66c724f2647f9c0b90c18907c70aca4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h61111fc96314f2ca5f3b84e389c4178d54876815a9ed2e1086db22dd5335430ecf70564c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf238a7f20511c64e4620c3f371dae9fd9405e6f9149915b16f46fb8ee0ddded0221ea58a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h13471296dd7408fee4ae192ab622f5c9545201e28d348ff8dec30b9535adfd9842ca39097;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h19ab3e1713559cc815a57af81acee33c2b4bedb25c225caf7534f1048898e7d8b8015f9ce;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15fa18ca80007ac794845dcb45680675248d3d3cdc22aff9d96efe30d19abe0493bdcf6fa;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h16687d9b62a18875adadd86863b7bbdd2d5692b5a43c7f97295d525e6423541dc26b4d3e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h16d8f318f12a8d09a816cbf141d511c01ae551c19d60bb65740f32487a4f4cc90a0dcddc1;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h472216bf809ff7cf05fc7794e9902c61c7b0e2afc3da01e5c3e06d3a91af7b4092772d3a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h19a01ea189b8c8a94c87030d98d4ef4ecaa3515dcf2cb2acb697845578dbc37b3ef0d9031;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd282a7d247b1e70e1404f9b16b6096e1d529338273fcffe73b38025b782abdd17218e69f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h5f9460c09e88cc4d1862556ad25a1947478722fbc24f1af9ffb671959bcaef121a10dab4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1eb2604fe652a7c4574d875d04693e099eecbbd7784db39656030b7f33d4331b1d11c455e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h3ff0332a8ecafe2cf44be621a2d8966ec517807265220610bbb03e5b6e4b5a3e415826c9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1fee8e409d0e5876ac4d6fee0f8e46d57a00f9f54a38898fd0424fabdb00352547b5bdfea;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h301902340780d533d12fc048e550d5752128e11642db8369f344f30f5bc2ecade68dd474;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h13cf28e7de4f1da4ee7e36519518a0e9fad70267c113be60b28f8f7bdfa98161d64c2014e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h272f558e26c31ef31ad8bf470cb0ef5707c34e112923f52bc51acd869a082672181dfd54;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc57f3c4e93415913ddb91e1aac8566d2846e85be566c9e41f2ad165ad51e37010939656c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd7458d38d99b2ddaa6ffb9e26f563b1eb3b9a53110d3e29341970e21a59d9f44ae72e8d5;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h13901a8c43ade123dc1a9a38e5c34b3176e1f9af7e52619511faa3cf14b599417a0f44916;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h5182a24b6f8f27e12dda5d9f45723bc9033882e2017eff6d1c0257fea2d7417c3036c928;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h176f1b43991256e6e6bdc143e531b4d7c9a2846b59723dba5d4cd54c7be2d754f67ba0a45;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hbbe37497def7349c83f49909456f3bd7c2d9eaa00eed7ccf80ab5d45716be720c795875e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf0f19c5ced104461784b7874604fc9bf87fea711d58c453c2c00a14e71a7278d652abb14;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h562fcfadfa35fb24f2734c940d60f186fa34c6eb04a1af21258d2531975f318fefccada4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd3e873c6b53bdd197fc37249f1d9da827e65659071a80f0c752051983f6f45ef421ed3be;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h8df166289ba6337505a8dc2a128db1c7e02bb256884ee0c4c244c9f740ce92fcd14b9617;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f91f7dc82e838d6e141b90b4db19c7667d7a5956c8b888f9b15c7900deb4b8236cbb5dba;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f9cfd704fc3faec45d7be035fb1201bd8bf3eda6bff93b8a16ce0fd80c31b4f2e92675f6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15c2b91533412816fa6dd73b1743955f008e14001a3053673d8f6b2e71fa3b9f227dbdd27;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h12bb155894a4dbe5fe1f4b40bbc8fd84441c82d72292fa941073381ea7a11add509c13eea;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h64932373bd7d11b62884e83e1986af63e1cdd09237ea3608899a98ddbb4fae0313ee7026;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h4999e905649163120dafcab82a10d6d414c374b342c1ef38b7fac73e5d202ca8ac8a9cfe;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h4689b97bbcd79f96e9a77a5a2524edec344de203ad1f11b575016c367fb6171b38b17a45;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h976dc28ff9ab8c2141081cbcbc5093504679cd027ad04f57f2548d12fc1a88b1ac25f283;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h758941ed8420e825a4df5d764048e9550b4d3ea06626ad23a9d90cfa89a21463106fd322;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a25aaddd584f504521fd24082e4b6ccc3f8f4b5cc586b7a7bc1cf00d70d8f58aa8c83cb4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h2d1c6da5833b77cc8ce1aeb7a4967f1ca06f75dcb13610eb2728a477052441f0f5e368cc;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h16a06e3778f1cffb6abf8275d2f0e295adc17a2add250e23f568ba6359d40734019c1ce61;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h117d1b29d45b9b7f29d3e6d78f917f495d1919679212753c40272d6ca68d02a80e0de14f5;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h17dae836c90c0f700de23d1ff735913502e16db9ee0af48ec69081edf2d6a981473a5b1bd;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h251bd116d2f10d2a5c559fc0a9298e3f9ddc44f3d7e1090a7df6da2a2ca17393ee4dd8ec;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h4d106b34118a19ce3fd9b2fce11d3f4536c755c3b9d26e4edd4ced4fcc56e97622f60a71;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hba3120353887eb2a0fd3664fecbb486be705a847dbfa647a6d05c3d23479c8d165d70133;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h128caa857953a77a52e7f78650ad44274fc0107ace726bf8e9eab0161e01b914b1905756;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1384ddbef3dfa1c5ce04b9a8c081416312ae89aa3be33cbfa50f122ec30db83178dfc02f1;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ffff1f76fb495c29c7de3c12608381ce0cf026feddaa8d145a3653b1aacdef422ef6138c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a716bab05d02bb5bead65e017f78e850caaaff8265876d4814321ad3445615ae6a1f3df8;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h33cd6e56f6f4dfdc2156b81509fb99d793f170f6c951307727e476c0c5672c333b20170b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h622ef72bdf23cf223ed8effecb0d1c9b75048e8aa1125b0e2ba49aeb46a67c8e1dad43bd;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1fcb5035badc7c4cc76b838482c0c33bb82ffe370f98d497c4ed91a26eae632c698ad8a3a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1bfa9c0ab35b7164965af948f04e7b2622e34af0e5925b28adc9016e603bcd3b9070fd51a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1edf8157e7cc480c31d8acd3474f4991cb3bf05dae4914ae04236627692c0d8563a58c905;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h5820eefbdfa69d4bae55950c7ff727f813c2f456c608874eb28e1f3f9a1e0ef5029025b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1900fb74179749aa3ca4dc8be281b0b3bc0b12be941ebf5253a942ef1dc67ab5fe1a8988e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h72785ce376959d12c744fcf3b3c1fd8546be3022d00adf28a172a5a71903b0cdf9f09774;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h9f93ab5d58483c0da4af210050371077cd1b88b527d570beee8b9451e9f44dbf3bd7c8c8;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hac6b6f3d61d87ab02583b98114b9413c759aeab6973bc3ff5ad0b57d054dd0f4a2d02512;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h17245f0b01c0c969a59287d357a15b93c11ddc42d3061c0ece369ab1c9d9ce847a85c01c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h226d9a00fe386797e435f08bf253f4fc1f728c45dcb29f364a3d0f99aa47f72eae0f4b04;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1222cb7ce99d3d50541ba2e8881a1813f11f071c617bc16ba86024415d71fc8fd411799e6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h6dbd970228edd264ed06281f6712638e354db7ac64aa9d93c8314553f8db73bf9cd70f9f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hcfb17e522461ba73ad04c566143531d6d24bc267aa124ebb29066949934a399dd17580ca;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c2d16dbac5547d81d012a7466316939eadc199b21f388a4088908d4869e7c38130c2ad73;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h91ae335d278405315590c8f57c1a0eb4cfae58084a016ec80b1880a5fd2dd6320394ca11;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h4b339c4a42d947120626cfa7c44e0feceddeffe4cc34bcfa14316bef9907ee5120674dfe;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h78620125477a5908938cf55b3c59c15f326e21a6a5458760bbd0b58f125dc4e5b8966dc1;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h2e482f3792393f84ea1d9a19d9b7265ae6fd71396317e4606ae822350759af39c423e34;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h74b75219500e6105c645bda4154742d6c582942a83ff3938d4d4c3bdaa5982dd981164be;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c4a0bc5f36d7d5bcff99bc7a07fd93fbf9dd3a42d9856799dcd9e1f52d1f9cac8ae489c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h142b730b8b904a7ab185ac6b207f307024f1d72b1927a0f4b7f5f6e4565aa31071dec8c66;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h153ef4f0cb55f36030748feda078db9a80c183d1924d06131b6774fe05f08cf68226f1123;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h11abf4484fea500d61f9f835b5511c42a74bb9ce6abd0a2790e663b32b827113a0727c9c5;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h9125526cdce02c8f3e5dd9f4dc52b62a90ce733c4458814c3b149c390a5245a6f234d50b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h4f5d886b63e76eaff087d9f2d10058723461532c9dbf95a71fc9edefb2dcc96d3541d71e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c5da958d14bc3cf9fd2fd717126ee5f5b62eb92a798842f53b51275333771dac3570853a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha9bda0598bf6a0ab0dbf51aaccbfbf640df605e0af0e4532e1e313b3e559000c3bc858e2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h156ae3c55cec25977620e681c85795402cc9b4497de37fd51828eabba332bab411ee1acd9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h11304e341bf07d5802d8d47b23377b783fca54ec5bfcc8515de81e43f242ffd3754241451;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hfa2ad0e985d487cddbcdee3fd74bc1d2b3a5d8ee4e1d051a5d51ac6882cf831f8a7f8e7d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha7d8ae72a5ceda9bc6ae90ac88205aa0f7695afbaee203389f1ab397eb85c6fc5cabff3a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h11bfad4a90b1fbcfd00a4d338e89e8da1e82b39e44eb53b8714f47e0c6a2e1b70e6c8ede3;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h182ada36083fec9d3d77adab75998ca264a13bbec606a8c55b2ebaa328826626f1917e104;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h19e962e03f4ba2448e054a4b60c7a79ab0235993d46256ff40ef87e19581fac9de8a4e71b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h143c623fea3711de19635ec60ee7f6cb6b8599eccd18663a6e4f5873c3fa699fda7120cda;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha98f5fa42c3d4036fe662636e210adb9c3af852a91491ada683c853b12b59006b3331133;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h102a1f806fc0523ddb0dc26f2217c6bf1972c56e1bd3965684b36396d7d385f412ef37dd6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h6c5e1ada1e245872cbeb88eedf959634a464cf6ca37d7cb83de1a12ffa9b3949369d5ae5;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h87f949c528d5cca1fae8016d5c2a57b58f64e6d4d65551893b23e33ec11a4b89fe136f6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f2af6b07fd10ad21506620148604cc4af50d679c80102ba8e6c60244b4cd7a59c47f9264;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h59eded00e19d2d03e5da6fe1b9c1f94f5bf9456d697ac32f595b09ed09911da50e8d1b05;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h10331fd3aa653a7e285189ea901d67c0057f5ac3c9720c9c9453a28d2425387eca1086d86;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h197020bb5cd93b83f3ffd4dec898b818ca3871a06061d2596dcc6d34b437dd9d919ad61c7;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h718d46f7fa7d0c2e59466aecc8dd08b98abcf04dd7495704d7f5cd456a72900c07de47e1;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hbfbd93bd3020eac59c64a4cf8de478dd6a5585a286eecea025aa34029c58bb668212b247;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h17cec20f6dc8efe26f344b6daaf19df87ef10b5bcbfa499d8ab7c6dac23feb9538d70bf5f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h71d9a8081f9a9be5fcce75f81ea78b7afc2418e1ff221396c14a0c45d596c9641dc00a23;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e7079cdc1a3bfac3bbdb1db1d898d80f28702168e2cdf080b3da6dc9c7bc7e43b4087663;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d59605a77ceab95941cc11e9822f12a081eadcb7192a239cc5d58158c4d86901ac5ce6b1;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h136478a57868450b14bc69a57ff9674e8927c2eb404781d09b10596b586da6897cae06a8f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h638366dd7f43cc41e9ee06a471b699cbecdc0c62ff54bd131c6672f48a1aa80e25c0ccbd;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h75a23a2803bf6f6fc0fb6ee3c1cccb67f4a827b359a37a1f14dadbcf0f8379c24fa62fc3;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h87eff7f5698776c006e3c54ab754df77525bb5bccd7da5c3045f3b3047a36e556ec3ac69;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1dd48cefbc9be6e4dec8342d1212c33201bf187bbec377f883337ddd2090377fc789bb3b9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1978181a920cb8784f4202f13d3c444ef781c16b27a087076df52f030d0566af62c74b8cc;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h54b05a6fcd814b5d5c6a410fb20146cf20c0eb84e33087c516d6e59114fa8812ce1214ae;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h13641e79de537ebc1658749798b0f41fc5fa05253d544394d333662760eda54cdc608d6f4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b8691d8f2b9e6f3b5b9471fdc017274b80780db8579e5563536d478361ba9ae15b62870c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h582ad2165a3203500382dc59c0a12875eb5e596f6befce14a69bf74c77f6bb6eb5863a23;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf230695350e5e98cb64b092c0a048ee0ef528f1ac98749fd019de9251c57527dd35d27fc;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h8c2d6e4d3f7dad94eb4730a5a3c6e5ccbd8a21285cdac2b94c1ee3292f50d017aa06fa1;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h57ffd651d79b4a9e3daf3789e1b5b6a8861b331043571ac2067f5fa0ad451b5e6139b344;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hcb27dd8a6cf7f1ae2d046ee209676c537859d4a42b70f0450de19c423282fddcf116d4b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h18983a9b3913981184717cdaa3bbaf5ce201fe33f61a0870f1fe4033b18ca302940b88238;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1869ac237f21c3e408e9d341e60918bcf646f4c9a963eccb5f25bcafcad9c47ca724c22bb;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1edebde932aff15bd0d4211ac71025fce21ed6bd3d3d364d6609d98e39e11cd257a50433b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h859ae70c7da4f0f1a5342c0585742ea4c3286e8bcca1c840092bb783dba8cb96137c27a2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf6be3007f41ba41be5619ff4a869c7d32c8e6f05e3825bec00fa15e1e1c15ce1216fc01b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h355fdc73e31fe7f1dd3e300d485dbaab8d128d93336d488b67ad24ea9d201a826cb8e06a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1cc9a166ae3dff62cfcc69bd6a110e8d3a4611e54fc3d62094e250d9851bb28ea87021a0d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h9abb9e89076a07c18daa99b3421a29f9c9bb4a0d69ebe6f34605372f427b236df38cbff3;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h54763a3be4001c7f9fae6560723897236899c5d425e9d255b78d04156cf79439d8ccd94d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h4e80d82082256cbcea72470f561a38aaa7fa08c6728683634d98cad1dd4e6b631fb30839;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h175bcddf562fa1de52a01ff1a27be0c542dc82cab5a7aaa328b82c6e26438b60671f45546;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h30adaa7fe7adc20aa4368d7d6694e292e51e36e32d407d6b94ea9a8f057c34aa387aa739;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a968498be9e29c6b71c736e76282a443dbed8cb346a2a7c87822a4a428ae656c0b3ef11d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1988442571bdf9ba8441f58e186f6d2869d63b375b65c784943f394d9017f2297b8e94d1b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h189311ac60ed3d7931599bfbb80f351529dc5ef0bd0ded67c216638c84b596bb0d002d3a6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c7acfb6ad4c23e7ea184e6ba7eaa63c9eaeac3a276dc116986b3637e32df2b314cffa7f3;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h61c2295571f7120e318dd96a9fe6c9c905dff5fbffad5febf1bd1e98e46eb60a1d0cbf3c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hdb9d8c312a87290a026778745fda7db3ac96f327a41677db7f1671671db72ba1c6c96b76;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h131bf5ae9820d12f00008f374fd8f61a24f0d5b28f6e65ce435c9bf6c2b9167ac373603b8;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h7dcc84bacc2df568b120090079cbfc308232c5d96bf8e30aabf8a6ff9d0d6bb4e571360d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h11533078d853a91814fd935d7958efde0db2caa0fa8f3984e7247ac38a61e25d1d2e5deb3;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h6a565cf9d9c17e35fa5d05e46185a4c79374e88d699f66f68350b8a1edd22ca7cc39c548;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc68adc94c588fc6aa6cd36106ed4933361cff1e4a3d875d8480ac6f406362e6a96549995;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d0abd1097a2e0f234a482438bbd359490d8f52c18a5e765f9acef3e0fa20b93c6a5a0876;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1322080f27263dd65ecc79455711386251a83c69e23580570fc3c38600b37d4eeded06e09;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h13efbdcae1717db19acdd885cb74c8f29e4dd69f7c786423065050ebfd9419dc047119749;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h16eccc40152e10056817f8e2ebe858496fda9505ba2625db9a4ddca2a1732383515c5c7a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d016d4de6ff9a4db5fab7deeed1543c9923108e120ceb88d7a6d15fd9c54026655381e96;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b2ff2799596f3cc48b6dcc858c759e9923df01e322a3824ba88bb37ed4cd396aad0b014a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'he372b686d644068b899f814fa373e4bdc408708dc6feef370b0076455ed2890a93b3e0c3;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h4b3eac1d2b448918f0399c222e1c7b177ca3bd32d8791a79a039b9a396ecad8b016efbe1;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha3639e4d82f318e23c67cb0254f8743ac42728f6a9e08820c96301e7ad595880e8c1d011;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1212a45b345556cb20500297f215ca1f377af658cbf0d71be8b6dd8603fabdc069a00962c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha6f50bc83d05d7642aada0a165acec6d73c5de6af1c13e231397e8487ae0c94cfe02af66;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd737b0d0ae66f5e810b37f28f9bdefb09a1c663bd2dbbe8242d255d42cebd460e045564e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ee885328a701405d57874698bf5576f60007fc3c1d9b815e402663fad94468123264e1b3;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h27f8fffa4887cd01fa0187e70b247ae11852e5f1262ea10c48c626808a7bbcb3ca928534;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h18ad9bd1751d7f3592e002d6c9dd6c07d56047436d856ffbce52ebca4732a91536333fe46;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h334587324cbb3457e23afce5c5b7d119df60bc23ff19084819f9190efdc8868748a6ef03;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h5ba7b728c15ecbf6be65e79c85854033b7ec2be96a0a6453035a8dd0b508d28281dc4282;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd677e498a5c1811a324cd280960028d973cb9356e7eefaa293d153a1546d67b13ec6afc7;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h230a96ef716d4301bba95c62474762d08829f81fad520a483d3526586e1cb27c97d1bb5a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15a0933d9ac0a1d6e69389968ba3d425ca9750410a223cffe51c7a66b4e21d444651e3c32;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h173458d00674f3e4b05e68efeccfa03da99e7a04ece73ad111b3707e3cd9a94fc163108da;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hcfa3a371d51c94e10e669e1c87ab74286323e02bb1d9796c7ff4fd83d2bf2b03e42cd823;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hfa1130e520b2f3b5ed284d1086898559e8cb6753e6886ba71a9a4cc7d6bf5533744b09e6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15a38a984d6f93c3d4d1cc80f0c5ebca033f2a063e410e2089a7e0d82cf0b6e259a767c05;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1040260a77df0f52c4e709211f56622dcf192c56a727fa713f11dfdb759f146d15ca2af26;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h10d01266049bc5a30a4a35cc641c3aae3d4bea28acb1b10dd3e8d7d631851d12110846e52;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15f053c78e4cac845622130a390b78336181e21905151bb4c9321e4a065b573f79aa85537;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1084b833d02a819ad1829625a5ea8c22259eb734ff29c2b4253a6ed5eaea62e2ee8b1e364;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h4e89e9c3ea82374453dde32fce69edbe0b624d6c7b29be0f5dae37674bba4976475490d5;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c5354ff2a4dd60e30cf1fe6c46cfaf6e181f485a5482fe25a78f28a33591e8523bbf94f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb15f16ead18b864591c4ecefa3006f048b40baf6d1eb41a3f2c66583f5ce9ddfbaa11b66;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc426a9da833e300c6133e71d54baeb93f57b96256c2f724ff2615a3e1349513b0d80143a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h16dc0aa666ac9fad9a21f76fdc181b02402f7a474803463f5db501b83d334c29678b0d7d2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h113698947df2555dec8d0d96f3a2bf070e963c951582356881e7873ac599a968d46f82eb8;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h5468df7d7d7f8a6981d7bd89116f8f706b6b341c176a34d973b63a605ad1859245c33bea;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c7a0c6941c07bd90f74a29df48d287f41d11f0f312d4532def7e84825ab9e858cc7f77fc;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h112bb1366cbb38fb7738c5bd1ced67f1f6a62d54758c4fa585f37aca0930be41c17870bdc;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd9fe7b6032e45c27cfd4b6a489e00ae3fcf1435378e1c7f926cc46ad6e56e6c26f07724e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h7f4c867fe91f57c4a1587cabfd2501d50ba943714ef20ce0f1a4c49f709b8bbc86cee67f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h9cc01c1c2b9097cdeffac120bc129152f10aa5b7587ae23ef0da03a42db825175426231;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h27978be433bcfa810dcbee1286de4967d590ed9dc6dfb58fcfa67953433eb73d84568500;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e10106c4f998d7ea0acdb412e7c2381623b7ef603b6e824a207dbe1e9ca2af4a038848c9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hee1243e6baee24dcc0a50b8c876e9f0dbd5656ceda96b09f76b82264fcdb0205182320fc;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h20d1c3ace59a6f13544cd51ca733640136314f5ab0b7c0d49a6728ed6c5b1490846a3be2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h5636517cd624f18d684d112672b8432a8df45bf2e384ce6a42add235153ff55d1b427b26;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ff458b489bbee1675df2a5c6357d045303e6ced620a667d585a48374c5daca9eb077742;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h4583ceb871d91bc76d04810e08d07f2332e8129d8999d8b98cb701d56c4c94359ceb7a57;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15acd61488d1ec933205ad0714650673b0cb09944e92852502d7f6609d456069feec0a93c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hcde69883bdb5e459daedc718fe610bf192bd275a640245cbc62e24b9b1d38882dc980246;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1694d4362012cf05679fd94a92d47999f37fad20ac486d039539ffb63f71a73fa06928dca;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h100412a6f8d24c499c25747e2b0934dd2fe4139c4ed7b125f2b909c3c318c292afe6a8ee2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd6105cad5ed3b1621d4ba1aa7b821a517d3f297db7bb4f30a755ba32ba1a8bc36bbcf439;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf7e485f543f59fcdb3847bec5404d5e772e5ada8b77660202abf45c3b52e29dfbb4366b7;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b4f0c9cfcf10dd7a474098d06dbc0c12cc3fb76cc174b1bcb8354c87ad5cb49a1f375493;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h104e971e94f69a5e40cd0fc8ec5dc9fd47ddc4444e3d7e7844c5cc72c3b3345673600f93d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1bf27be19229f9dd7f21cfe8aed93d79905fc1a237c491dc5b3906f3eed8d4dfd7ec0e8e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h107e31cf5b57eb01798ec907c2b37ee286b061c7a5ede64f2b2c7a22186866d9bf69f3773;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hda7b673013449fa042695f2ae6d509f3a65d36ba07437525ffeb88a57aa23bb0eb70be03;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h64993b20269974f23a364fa980503094027a84dca3d02aecd940827dc81327bc0c98263f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ea1e40f770e81ab87744a15c46fa8709e868c2eafc94d9f70182c5298d27339ea07b8220;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h59a47e4737d7ed799d3da068fb4697a82bf006658bbe7f36c9fd73f520ee4679feea8562;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1213791beaef0ef1105a37501e6e84583c1e3b8c4824b24a70963c869e43e0b53e1c65ced;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b610aebbaf8826169b8ca95fc9a53b592ca5d4a94df58bab5165943474790f50718a95b2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h689cf4d321a66fcca72c9ee949077f548716606975fb5a82342dc2abeecd7f7c9fad85c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h17e364744a1fdebca8a29f9b1d13cbdbcbf7e83e20118cdbe628af92348f10939ea754fb4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h13067dc6a1765513b3154620d1752d65d3605081d4db4de79706b548bbfd222e9d21c3d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h96fd76d4b2a766d8640da600f91ead44fe64d112d2ef9502ad6c6c1fb6e96bdaa60ccaf4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a902bd355b3d5e10a38aea99ee85a05c11afedaeaa5bc9219920408126f5f7c34c04fa43;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e9b1f6a60bb48f2946a7b9008dc39a8bcba9af0496b839b7ee1c1e0dbbe30efd72cc63b7;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1942b5f2035f949a1e64da161a083d9d712e102f6be9277021216202dd49196a6be1a9dd9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h12f921656056aadddda99e13c4f598c09f99885946c35ecba4c339dfe907f63e1026bcca;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'haecf68b54acb8bad650fc767e06d2f92f5bfda9809e5c86a3f6f55fe7724177147a2c9ca;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1abb6851bac30ea18a9427797e3672505e4a29ccd57fc45d5a9f8b11e7cf3607475f83d17;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h12a0be62b881b414bad2f758109b2e02ffffd70c173def1eab13a621e84253b98e0653345;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15bc19b0e06931d35fd93e225128203eb8efbe422bb06d2d5fcd0436e6d3de94d2b16cb1e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hfb925129b6547875301fac68699488dc3eebfec71f551e5b7f500c9bf454b6105d2a4caf;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h19a12d9de46c5a13a5b2a59863a4dd32abce3ed09dafe896378ba7e7169518ca1a62342aa;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h10fb16737e74505deb45c46e0674920ec15748d02a24ce66da1cea11ffefe01650956ffaa;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f79439d71c8f5499e5af98b3d824d6c6ffaf155723f1c38f3fc397bb01f0cf678cc2623c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b2278d3756e976b0d0dfd836b358a86daac42c200b48303acc091a89bd41712e858e3753;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h10b241838094a9afa58c185c1be76f6b21fdba4e1a3a6883d86eeced3ed501d0e555f4c7b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1745569e87f57fc3f2ae5cf953aa59f059b85863f6290be2e28ef52e6eff146f57f820bab;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h69ef9d90456bc911c8303ee0637fd83108085bbd834bd7d4a292af58ce10ba1bb8c59e95;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h17f09d65a69e8b65e86b042c8f74f466013163aa4cf17c52ab8f2982deba3cb471da9c886;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc96163edba66c0fad585dded84e6891cf3be41045e69b57fdd00fe98c9832bf90f8bdd3d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c3fdf99b0614feb73555298c59d83f6677a07054e402ee7154a3e3972bdfc4f3e04132b2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h19550def486ec036b2f39555c5b1c8f302a1c028e0c6c68cde535c4381674be4c9ab89aa4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1de6446ad00739730c0cf55aba40db1156b0adc60616b970c3132332f8d70c0aa385cc15a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f9ae6b0a0964d4cddae2db082ad3586ecb4ff10817a4de746ca78f6f8e95257d54374098;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h6ec8d14aedacc9ab09195446be2f043d01005ba8c6a761d0f9ff65ec7157e8ccb74d818;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h11e0452d20d577957b9a98737a6a770527dbf20306bc0b439793fa922c2d2bab117199d81;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h145693dc0e944ab28038b810b7d85f90e2764f852e8d9b3525071e8a91e6b3a880d5abe6d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1cd20d55efd896d8075981b67a78ab3002645a1a1dd7241b6d6e93d96f8c6972c5c3ec2ee;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h19db3fd9347d5d9a53ee353f26c3bd0821fadc35a999536f2c2b9ef76327953342ab7a05;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h18506ed47bc7cfa36ef81e2db468a1c838e2ae92b064ec1f9564751d883c7166c25df0af0;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1745b8958089d3d4380f0dd59d41c57c0000fd4cf2c8a2bb3a328289e195f0abd00133a39;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c8a810273bdce97e8286caca79e95b5552090f654507b698ce3cc762bc90e9d73b1c9829;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h759c5abef8d8f5b9c36fdf4544c57fbeefe7aab2eba1c7031fadae102383e7ddb1a631f2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h19e7bcc9b3f993ca5efd72c2cff8fbd46bf772f363ba0b18f5e8094736fa93efbff1dd477;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h160f568a794af0dd2215169224a4fe0fec80455d74b9f81d5e473ccadd9907a527c4e8b29;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h5bea5fc7dd2eba66cebfb70488c0a6335fd6fe440516ea988aefdb63ad915e46e9ee5050;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h187ae49ede16a52cc156a2266a4f6f8338c4e251a2f0a0f97e4e9054212bb224c62061f02;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h3dc7eddb5a9571ff6d30adbbe64354eb67d2bb616304b04cef7842f4669a8a3020f37fc9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c2e69d6321a87a7d51b46e3f1c13c1ca75b5b0b2e5874ee80076f9807afda3db01219d59;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ef7d9c2fbdfafeb2dcf5b37036c942baf9cf5ee2cc6d00733dcf863523d0e8b74d1422ff;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1262cdfd073812bcd41b17836afde239fc4f8f05d8c09f9d84e8e27435a418ce8e3dc04fc;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h49810b32da02b630a207539876b41dda55221bebbeadf90447a9bf603110e10d22398c1a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h99c9b6c3572f9082be7a3410e7ed2af95f93bee028b91fc7c8113c0f42faefa8608a7484;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ee24de3c95682c588e05b6ad30a2e001781bd0e93b49524c95d29aafaf5a3a43eecc639b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b43d8b6bc0aa6587011a2abae49f9c813de386c136ab3681b5c925d9cd25a9aa630c1e65;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hbb8a82f1e9bd1bf89926eddf437601605da0a80846b4ef628cb487d6941bed04f53b8861;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hba4dfa801dd14b1482e222cbf0ead17cac77132defa23fdaf40518b8f4bec4729112fde3;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h18be3631634b87c0c00343236d09d9223d7ba92c3046b3e3e5859fa96c8e391180bb69ae5;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f9c71a017fa53cfaf90fdab859c21ac3ec04101628a3771371ecb6318e9ba617a49c8235;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h16f4f341911e978f0fc02229bd2749c082557f5cc78b50df3b58483a2b288c45457adb97;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h156b69a6aba4862be353bc346e62eff9852cff793ddcc041cbcf2a81be96df82353aaa1a2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h14d42877b228155fc0c870df97b4ad572e91b83d6d440ec7d85d7ec43d451981d434de691;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h8aa61b1d17f88012c9f2935d10ad42468e7885cfc0cfbb33b2300628cae3cbb6db1bc55e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h5d187c276ac501ca5c0e8138abb8f25661fa78a5fa2a24312c8429bc1b672834dca50ded;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h10790b61088c45b217a2e8903641ea0fef31283cfe7f1085f2a4c31011b7a4771e1debdbf;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e0a56f244038cfd4a2fc3fdc4d071affb4fab04b158a519d49dff8332a35d58ab556e61f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h183c733b3dfa6775b54b78543bd27e62217417268800a8d09c9d01122b6b978a88f280b63;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h145c29f876e9b695aef95b7a1359419c09bae5ab1754b9f92f6b1242bae4f3c335d7bee4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h469d9a5a27a3c6501b8eb699c377a6f53a4d822d2cf689d95410a01febfb86aff7ead170;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f91ca776520733049205a54b8ee0f4d28b5edbcd3dcb0c9d406e34fb24d5a902e4d2f98e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1286c778ff5d71cc0015ce3b7d3a8344d6ae6311d863ebf45017d0ad8354c80e11335e0b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h2394d148ad0ad6f5816f79b214d38435994310b00619bf007903fd22c1f43b272c5ed0ae;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h812467113865ad7596ea4836af4fc661206c7855ddb6706c396a488f46260bd252032e97;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h19d51432fedd53bd7f5bb3d6c576eb6dff7968707a98c339fee7985ec03bd070478fd8a64;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h7803d473cbc4d80b4abb3364b8d3322e501734597037a5b64564e7be6335a37d696fca0f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h4b379041f84b5b0c7cc537839ec8b0ad9d95e0c368062ed1d48fd274d7e63ff69ea12cd1;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h34f92c0a6160888d1adcdaab4fee6e7b73dc15e2b7a6bfe03f81c73e8505928de886ce5f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h136dc5257e3ef45aacc693ccac9b26a960dee5156f2a27f9f4857fe222a290d85c491488a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hef7ee416d6d10134e9b4f0c8d9103a5683874785706c3cc5fd9e37f8b36c22e54dcdd91e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha0a01fee25d206f0b50bf31dbe06639226dfc62b577f1936a4ef6ef897e9d8ad615746cf;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hbf75db4e6dce01ff6eb25eb5581e3d61c58949ed73d44c32b7f5d4134c42d85b3dd50b43;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hfba72af4b6c9706a5c7d206ab32eb2387f110654b0fcc55449213e1f20d94fdde3db82b7;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h332f788ae874889690a8069bafad9c9c53817b5a82da56b7af7274fef899090d3fc391ae;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1964de14620f63e35cea5499a2d5de792555eaaf8b26897dba95cdf33b53b4a85e5a3301;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1eb42cca1c0205ad6c3c8d144f4739178abd13c5da40508cf6940b65c24ce475b8fb732d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb37350bc8db296f3607321d826acbb2831acd92c259713a66454038cc024629cf98c52d3;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h32d2e75b9bedca99f0412d67218dc4b38f97955770ec34bd4443189c5c27113476e6b52d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h126e20532b8393b21b707f754c9116e54f5b3519ceb00e2282372a37354c425eac1ec428f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e1826d9d518f1d5f892928b8db0843def8cf07a07212e49d13374ed7b92b4abb2f306b6a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h7ddad04bbdb833e5f871ab0b36224fb55d1bda7aa5f8fdc641a7ccf13db6465debc68bea;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h932e2403d29e3f7def8acf67a95b2fa0e8f5a5f640d0941efa8e6278e2ced161790466b3;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1da446685acdbbb610b059ac5ba98d2198520dcf29e2b2dd02eb32088590857e6fe2a44c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h10633bc877ac9b1ccf7d386502719c20198c19c8615dd63b07f5191973c6319a692893f8a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h8df0d486cd89d7007c400875a16fb39d2309bb18ef74d7666d3fedf53d598d3a63dc302a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha13fa5146e3b18799ae8852d346c375bf7d26b1a886401a1bf4acd1b3d456851fd8674cb;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc528c18322589d161a637e8be5b967f08df3d8b72ef69aad21b2286b4b17bd0ca6d7efc2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a0f130461b162d101ca9f5194ca63b2402205d8ff8f9dbbb40b12e750a9b65a0f239b833;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h5183c46409c22399cb7dd37d0806e0ee867fb5623ddcdcad0cbdbd32eecbd0b8885b9c11;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf95ea41f06627ed0a368fa40624a4b17bf54c40ee66678ad501caa7ff983501afbc35765;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h3c68c6fdf159f88658bc4d6b9bc902d73917798edde6a1e4a0842b8c4b23a812e44cc805;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h2786ff999eb100edcf843c2235bfeaf196055b53666efe3ed78f898067ac845dbf063a54;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b6af5f074fde4dc7a1b844b8786a0f3b4c753c6b74f0cdf56c0bed5627c4c1da9853f292;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h124bad808ce41566d2fb787cb96c102da53563d925ea6666222a9ec9466a4b41cc5e095d9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1867a88fa407435b836f2bfdb74a9c1f3521acb7e3c85d86ed859b2b2a25cb37e864a9307;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h81d5defa09f3c4051da6efc9d2a604961104a59299637e2c38af1966521ccf836c2f45fc;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h131eae1f79308ea46e491f6efd242a17eef04689cac8b58b0dbb8bed106fcc63a866e226c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hcfc3aa9fcfb0e8c4f0893d2ae37794446b3fe6cd5b6e08b8a349b9fd97a114623f3deb83;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h191bd7666713b943c31d780564b3cea27909ead8d92bb7f97f7aea375ba44fb782a2294e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'he1dd8954ffb1b6671df19fdafa43d9adb950a13b924e7d18d9dd2e9056d6b5cc096e123c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a11440962228b49049080e5aa3eef39399a46c09db0685b1db593f9b25e2ffa4db29916e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h138c6c41c45c20dd11fd4350a71635f36a8e77f0339ba53528ef7a0898be0b495136bc69a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f9e2b12bb4ef468b0b06c6b77b684736470f9791aa034a70077301e562b02a5ef785b68;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd823e09e1d77767b21c6977c42e6f4383627ef071271d10fb04c3ee2820d1fadf52b46ce;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ca8d4fb402c1ebeba124db48b9a6a2b71dd45b11dbed5556802b471f9c063e68693c0a85;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h3c29fe0cad87261c2728445f77ceb413dba196d7fbfa9bf52169436ce8c96bca3c7aa511;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c12474933b66c0489a889cf1e9792ed4ed5622df5b007f32879a2e69659e9caa58d7280a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h12faf8ba2a40f5e320ffb4fa62999ed5abd99bf7f853be62568da5f2c66794ee91df20cfa;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h12b8138d9516af70d430ee0fc513d2a8bdc2542aefdf977459aec46ed1fd42cf8ed0a613d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1df27313278ea25140c664184a24f525bffa42b2815bf7152255b844a12e558ebaeb3663a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1fa9274b8c61db8040d15d183c6cd3b4a717db0ffef12b5a1a8c74af954e88d9c959c3169;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h13fbb06cf3c5c4dec6fc36b9c54ba21155b3f8fd77ff04c852ccfd1b18a275329a7a9ff3c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h656e39e2509936daa4a40f06915248c031e627c3de46e820b4adb74ade1ec0abb02e4103;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h4ee3ad0835eeebf2c47d6fbbb333296e6ca23644421f4ee838129f4da0af2d94267fbd16;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a1e10b479cf3e7500ac315045a70c5fbe4519bdf58ce15213f983fff839ace88c3c481af;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1141ef7dbadb27ff6377aedb726a293c6b671b0eb57f4128cd8de2fdc881ca6b709a33697;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h84df76ae440668f2b1e703af525258f538e778fe9b2352f9f2c46d21de64d160fcca0b67;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h60aa28130451aa2169727f88cad12b97bbe0b85fd33d906ecd252cb8541daf0aa370e12d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h153d3bc1fe1e9c6ad5b0c854df1f027cb67636d66156446c6e9671542527bcb5ccbc7402e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h3f3886fd05d527f4494299acd35b57e669ad973c189bf54d4e77ec62bde961c314b125e1;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h19657a34fb27b88ba41d011ec5506ec250d28f6b71a01cb4405854d3f2a2cc377f70f98c3;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h80da56d380208e3f74381353ad25d7ecafc93fdb98ffa69469441450e9455a750af50318;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd0c2f6c4ee8f2ab3ae6aa95c9f7c3e20e4203b2409a5fc6d13c00edd1ddea9f34c64cf5e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h4e6ea77dd5b08c90a3c800b30077f621f7fdb4c1929dd4c1d78930bd94a93de4f4346e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h13da7330b9036be9bda938b7b2bf8b70e3c33772de74b45765c3cfce0aab2079dc57b1655;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h147123449375e0ea3a160a440b2f195cf44ef0593c5f0eeb581340cdeaef003c05865934b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha6eede576388c18df85713f36b84f5093bcd806dd242e1ae7ceb3123586c8b258521edd;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd3a6879dd6aa0747ff5a3ad4cb09eee8d71aeaf6b94bbacf46ef925326fd4dbfaba45ebd;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hbb1e41cd3e3fe93326fd4c129ff1d2cb1f422946f0763ea42bcfe9bd3a8e469c39508621;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1917296e255f25601317a82431556e06efd3d03702a3c9fc422ced779f2d867193be9744b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h8aacc5d5b06d8e7ead40bb611beac06776a9804247e6da12d141b047b4760beba230dd61;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc7a44ae4fceef78f5e0dcbc3fafbb6fa269db91e701ee0128b84d10da351edde39c2fd16;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf82e9ec60ba0852e55bdd9aa9e16f88c2abadcfcfc421ae1e3c54abd8cb75c6e2933779b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hbe7115e1da255168fe93e47b2c37ed5bd24fc990f40a1a1237a837e7e4e664bde47d5b54;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h12a51c799a595b3ae181fc5569e13a03a7f59fd1a5edcfcdb5fc7168ee2802524b1013cf0;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h107fdd03af7e35342296ac7984d42b2c764c52ddb0b7a34d8c8da00c80382e40ebd5ed29b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1db6f6603297fb22b17bde54fb10e24d5947aff4445ebe4808123406ac56a778d187cace4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1603e2343eb89e1bbe6d1fb6cca44e6e89d7e693560c2046190f74144e7329aa6beda0736;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h13423db329be63c522dff16e1455a9da504e333671289f945e4b39c6e27386ddf1d28f0ff;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1bbf7e95f8d3ccbbc1988fe11ea94a4580bb7fb9db86684b21853148955391a4eee031513;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf2c8030a47c54b54c3091eac23c77b79d6897315d9d15ae9415970b31c4c1d12516ed092;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd1073b476f962825ad1f78d7615156f1d43b56809c17b174c46ff2731adf740da4e1fa5a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a50ecf6a8cfad74358e7862e7176b329f60477c17829ffd9809b81dd96c343246446eb2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h11a90c43775d24cdc57b722553fd5e09b2d8f5d456c72553687772d74ac359a26b2c87a1c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h9defc78ea9aa739361ac149850f5c59e6e8a0bfb7d214e28aa47d9a092d7b371e08e23fe;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb2afd6b9578f7c7a3cd4426ec78a3b3156df78cdcc68ac6607588643702d48b60600b35c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h12dbf3f6cacaf4ba67521aad0b022bacb6880652021a0355c47577b1770e58a918aee78e3;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hcc7fe2a8ae539d2f703f4c0f1c7abe3aced6ad9e9f9885eeefa1939f1d3e9cb2517d3ca3;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h8409abee7284791658b948e72a79af272dc814570ab3d4efebbcec85bfdc77c60560b5d2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha7d1240338fe0a63123017d59436f6757184c07e518b17db7457f8793c29a0d3c59a80e9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'he7f50fd6cf1e231e40cb3405f2b2975d907efc60ddc1c4aa5a95d54096fc3b2ce183ff73;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hefeeb05448859d10812e01572109d8a8ce2832bf4de019747a5548226f4be6a849046c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'he8535af5f68c32ef71977018338f5fc32705d0d26e60e4e274111045d23dc3a776c9b09d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1fda709f4c448a6f754f7a51923f6885e78d3a73fbdb33656164bc5a97c986dda81cee68a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h7052a2600560775f711e05f59cf005f42ed8a5330db21ab721243394f454cba88dd90da3;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h146f353ce6e10f3788b109b879826618420f54a369c9e5f2ccf670bbcae178d7d4f9889a1;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h147ce59ac3a80297833a36743aa33fea59a78fd2f92b4b895973bf329ec709ad7937964af;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1af1d6905f1ed47d168f0a6101fb7d9bcbdc827603c00358076c683b65e186f40d4919a8e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h903b52e806f4113505f57728c7c8230eac861e83b9683e72460d8d71a12d57cb99ec8db8;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc37b4c67f19affc372be18564e2233e606f7d6d13d57cf06e6ee7db9f83274974c9922b5;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h129fe5ad91b8d6dc0f4451ddd61656baa4c6fd5a7ca7fe6fca4beebdeb5edbd69c42e6572;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h305d9748c82b170ae693838d8edcde4c9f7628150769c8b5e7ae2d5aaf51a0896c69002b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h171fb5150415b7d4ceee43fb0c55591ff1f9eaac82b34b1b382d25b8bd102bba749477923;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c3b4033b4df7392ac0855bdfe772e0d347a0ea464ac43a088bc2a13e009f2f9507e4bc0;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h2480549ba3f961de9f5c767a648c306813379d7c79407711f0e6bb23b3d9c7c3a81f4312;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc1ba58ba88bba4855c603018eb61949e9a55d200d770422c80a68f939ca06a41011dec21;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15b54d221526d4f6593f9c9e9b4ff1d5b07b9d75a3001a7a3e0538421334aecc57a52edc7;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h9d0dc2e43f0f2eb8167f9c02e5d22cfb7c0c19904a97d2ebdff06f34ad73f6f59694dae9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d213dc64fe18a28cb98cff2aef9dc7568b57d12790352531df5263122011134312b61680;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hce80e488cf4a6a3945689b1e13acc498f7a22feec76c510e4875669d3cdc7faa3c906710;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h154d1bb3b1cd038ec64b9eabac1f60cc2e5d087052a24b100291e8ebe3e9103fcafe88b47;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hfb7a4274ba55803a67dafb85c3f47a5d38b3842f3583fad0044faf0e304673d09be1127a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h42f3a39c9bdf1085bbdd9e185ee8846b1bfd6c44287c479bcf7f787cdf8626cfdc8f4fa3;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h14ac9986bbe8bbcc42e64c026b21f1c8e56fb3bf23ebada654ca3b8b7aaf22f56a8e4b0d1;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h959305b69e5ba993cfcaacedd7ed08e6c09f52c2d9e5e56c57272c9e1a9a7da625018448;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hfe0ce6180e22574f042e55209eabb13e56703976e0ca5b25f9c61e9902f2d016f2e9961f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e24fe7ef1231c4f90870ecd9634ad7ddf45c930c8c6d1188528352f6f49509e5a0de0aa5;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h14e5e7c639017e79cfca6c1e4a2ea975fcdf15f660b6c60078e60c85dd254d6675e5ef313;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h8b3c76636fc3f1f184b3aa1ecbc1b0ebf81d81d8ed9f9e7fc2456edc2a145bdd5468ce3b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hfb3602baee00b92a8927de578eba53e18091a789c5d0ee8bd2ec0d309cf190b83b61bd81;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h7e0d34bf4955d0a86f63f4699f430e4b4709563c930025b7cee5e9cf1d61b428f57954a2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h9c60635fdce764b0a16eddfcb3b56c7e2329e18c2ce932e299bb6b08263f4dfc9e13d8be;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb88f3b566596dc87b9c8e4ec81858b9ca307069d3ffa8160eaf776b285d1c1dc3db1dc37;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h48af975465a360f3793554500b9b044fe060ba1911efbf9bbe3d07b27d5182cd4391d903;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'heb753f4c0990367d068c8c67ca7fb2edfb57cfff2dcff93e0afd1275a3ca83618b15ccec;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h186b6127304525bf0820d4a4a47e90e35e91fc3eb9219a6a8e2353e07f1505cf89f74c2ed;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb3b686862ecfb09e6519f929b123ac68d6c3f8b0e855f1b55e6d40482927dd66da90dac2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb3fbf5d729ec3b4af8e45af81259c9aa80e02a51d5453c3c13c8ae54068f8f3c424e89b8;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hbe2489354a602a5eaa76d6b2806eee9552b449c7e79bc0d95eacac04a2e8ebbf38d3d1d7;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'he32f9fa8457dbba678e05fdf19e0e0da26501e901abef33f922cb1830296dcb2c257660e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e875fd89d903e8e211d6fc654137fe4fa39ece02927d7241e9ee6e9b8c6cddb5c414a38f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h9b6e52d82aa93bce65e4a344ed8a9718bdcffe3aac431201d4f9c34a84ac79fef10d9d80;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1477e8c915cf4c405a290a67fba9353b9cd383eb295a2bb4c289742284ee9c1560b141227;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hafaff143de11cef349268b0a41a3b649147fd7ccea73bf41558234a7156d4c8b19e7db83;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h13bc008ee3a16da440f0318b448e3b3a6b41728f25cfdd8f4fc852eb0b5b801f5db3eb722;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h12494df7c1d1003fe651fa23dfdf8b86bc23546d91a82ea3602c0a1ecd6981c5b8c125e5c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h9b5b60d0fb57e2baa8e132fc48b74f12d9ea1e810bd14fb2a275b418b2cb6aeeec09c8ae;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h5c5eeb2d206039b231b829a764792bcd22ffc1ae8f853857345a24c947f160deddbab8d2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1bd811da15cfa171eebb302b10060ba13fa10a96c8d760deeda5cd3800af4357467d1df19;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h194bf48d25099e00a18d333a578a535d7eb67e3e696f0ea1e04289b1a0b7a5e7beb6c4542;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hbfb7d890396ec9bcf9cf701cdaf6b5f5366ce6dbfba7c4043598a9aa9daae101c8c900e2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha338292c12dbb2d07edf5c70ba14d17b27c0c66d841522bcabb1e881fe383aff2548f6cd;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h13f3d8e2328f08350fa89d6ec8b188619ef03c331b741c4d7ab64d5b943bf064764e19238;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e3f994e3a831a890cc5f61ce27aec184438f2ff43ffa2922d681ced88c52fb9490ebdb70;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h101ceec290456e2c4f6ff8a125be54b0bfdca3f77cfadb02091ebb6d169b6f99d5b14da14;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h111c0e20c5ccf946cbcef44e19e1c9033fd8918c00b4576aa3963a6d331eb3fa61dff4746;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h6a5cda1a03ed14dadf8704381e397ce0c643a110ece816cb6fa7ee91fa0ab2e954a74743;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h164f66e207c53a9428180991d18ac74f7fea0f147a8faf10e3c1fc427be9d711a5ef132f7;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hdd5fe2fc01c2ffa6d9d944a790ca484ec91ba599e3894672ed81e339152d40d8182a2f48;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h14ebe735d59c151d2f9f5c6367dcebce825c5d48ea686642770f607d52bb47f384e629a4e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h55854ede08c9d60dc17c4aa8438ce54a656132c718329f83cb769de55d049f2f7bd67e7c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hda998a7b47d1b659db713a9a736d3626634c86f3d39896b7aacaeac8668ae8bb4ed7ff20;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd14ad4049a803670ee8f6c86488bf55c3da25163791158ea4f656d72ffa7d16dad0c8497;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h197ed852ff095375aacb365a5abae22274328518cdf5bfd49204798a63c61b83a8bf37d6a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h5fcb329bbca95868d89acc1d9bc4808b32e8e425fbf5b86e201bcb99e8fbd1e6b65cdf10;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'had1bc76a603854eb12309012e8113154c83240eeab6580105295965345153fd649fe1e6c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h153949e151221c0eb1f8470f091d38180963878da0391806f2c07c095637c380843130650;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h58b6bed40ebfa45bdafad9a60fa166859fb112244f4d1622af51a08f71c4581123032f69;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h55df1746a2935bc4b0512f2cf618b322d5135d2ad09846dd89b1bb8efefb02617a6581;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h147443b06167c92f411765f57504dcaea30bc0866e711a68b04d290defeae45de45a6a8f5;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd0832d6a13b4546d67683d535ed5206c62a6ee29e8f4ee73431f86dd39108f4321495ad6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d79fb0802c1f2ddf83770b367578e57f5d6a05aa44d065799ab21206b033ea480fc32d0a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd092d3d9b9d92c28e6ac9e6b5d60594f0a1df3b420528d4e37a3fc6b1f9b2b697fa49873;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h86702b6c6d9ac9b4580d300fc27ddd8f42658575aebd9716a22952af37f824d4e1ab95fa;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h17dda2f640fae0c2b7427198ea57935da64a5bd5809ad73f1b3b770acd207fd6034805ca9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f0e0dfb0a908346b29d24d6d6bf4073b4c71be0a4ca396e1265381cf47b5be33e56379ad;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h109aa8fed0e2d774ecc9e544b4b72294ec197863cdfe9b3280675eee53e7306b8d7c6a488;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h11fd39b3a4b97264b35d1aa9d53a443f4b71d4f285b9e39fd3fe1b1d6d23dd3b8ec66d33;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h38f80b4afa09b28d2d72a9a212365c50341938de7ff97b084d72c41b3c18a7294a1b2b3;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h7d3313649b13ba54a23d3dcc77836cb387249abb92ce21023874dcd99c9abf108b556a2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hcf67671c64ebe196083ff36ef71754e8ef08378de2e8f5d16af799fd31a229775da5768d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h104eb7930a451b206b413489854e074e22c02c42b115ae162aa9b449a8c234ca2558fa8bf;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h845df76f533f90dc37f897ef4b0df2a1c91e6c7e638b6cd41686f96093f6700566e26d94;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h19639253ac90a7b251053de8210cc48c77ee1abb9fb3390a7d87ce5a0bf7311074b5a51df;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h17a56304bfcde8f14e5c8d0e4e512f909b021584ba5fe0b3f887100b0c8c0eeb1958b0658;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h9afb08a4cddfbfa503b4114a2a55ecf61ced2f47a48638a67ce237863426d92c2f9d67b8;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d83b4bae049c934651ccb973e9a1deff34e6ee17b854a6ceae7c9185df50a3e9061b04bb;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hac0e0a1c874e7dc8589ab88dc0ff5ed5c450f16b5dc89812f2a8698dcf6524770e31fb3e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f364bcf05c38e40f4b8cfe86c15e501b9b2ba494a175da2ea9ef5f6bd672df8e39e5636c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h18163c4baac9376a4bc91241708ee541032c5e999c8144626ccd64e87c6ebd76f32c70c6e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'he9293bea1206189b7331243b9a0e1d6706e2f998389ad857aaf386f1e06d4da94943f370;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h130f7d22e5e9bb267f7f2955404db117b8073fdf78b64e986608fa037c1f6a61a8877a0f0;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h66f5ed5a56198b0b89b80e9791bfb274515be86d535296f53b2d440b5fb3780545695ed9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a94d43fd978544565a92600bb1f3b84412c7967ecaa1f7dc1ed5a6ac7853ed6cc4b83400;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h12b3aff9050acd878b660536fbebfdf651a87aaa8f0d7609e7d464e15a5e3c05d37f538e9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h184da690401717e87fdb50157315181475f5fd90ebf22f04716760955b67f0840bf5621c0;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h162ddcae88a2e25d02a83ddd48d28e2b24ac34c429cc65991d6072c04c4806f3c2646c1aa;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd7c2ca2300848668c46c74bfd05f45ea1cad2cff7ef24f5558f241adb79ad6eb968c9ff9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h996ed0c340c0c71c2a7a12944e77713388e1376ff97bb0b0103d7544b8776e9f3a47b460;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h372c360c4887b9ff02c7b59ba58e9031d7b05ed859748d92915cd94b0b3e1b29d6c4c8c9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc9083728301ca995e7f8258df14b600276827be2a5d77935093738a6c532ab1a15bb820d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h16e9821985e4dbf753f864232c2ddd9c4c0e396e3645677874ec2dec0485530ae22d5096;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h88a5da43b4b8125cd6585416a425cd041155182de1ad0f9a070c0dcca619aeeb4d38925e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b3c6e49e2ba9149b3604ed8af857c114c2bf56f6720c03ff39fbc528718f643e02490f02;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb2ecc6d187b300bfd3660908833f29f08c73e7c371b8dfe9b384b543063a44cf59fc317b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b3e7b1f724a4cba0b04278fe5f804fa5577990b31496c0351b64fdfce591ddd6ccf5dcb7;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h2fcd59c000fd2f9b58db1690c49ae21425fa013b977a5a27e8c0c60de7bba8f9b2731b58;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h49f7cc739b1481e679bc9f1a2eb76a6edb8adcb4aa102279ec5e30242b2377df9904bae4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b23df6174cc53605080d9583dae109e2aea592af6ed6051875a95edc34a97c90c19c6dc3;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h6261776a7e29400f249444c4dafeab10779c5b32c682ab2481219679047251f231db08e2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb3f3e285ea120e94f514d3163938d1df81483409e1dd6de03b94ba14d5cff31463804216;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ecab5bc2c279d63d356b7710c4e51f546e205cd3cf89b54c9aeb3af17ef02f4215079fd7;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h19ac2aa365b3b54f2f37ac79b3d6d3e3b3be42de084530f46a3c8afed2b8513968261d5c8;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ca4e98eae64f77e4383941b2f18c762e0f02cd9873d5c5851435f50992c05e408be29e63;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a6ed703abbf455b458e849469eb1c3ad2012c05fc8ad55879eec5249e1caeb2a3d401d99;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h16b2365f812c3f25b7a739bbe34e521262d5e3c4b42a75488bff28075ef88ff834837fcfd;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c29726795166aa97db0549fc27abbcb732fe7f07644f9549f8c1f31607198d41597e59eb;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h30f002203c6cd4d7f84a93b34d2a009f3e19e2368d104c42e823d3ddeb754752c943c77d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d19b17ed0baf9ebd0bece629059f4e52f026906f70628a3705cca9d6317233ebd862a4d7;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h6635f6d1b3cdcf9ea4b7c67640a0beab8a28a1dfa40a0868307087afc96a5e649fd5f59f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h11aa667bb8096c52cdf677ec89b678a4353ab8b58f2dd11da3ab5307f376e2fa9f1baa050;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1156f0958fdfcd3a9ce0a3a0a503192fe69f10db14018dc8fdec693e8c979fdad8ac27e97;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1491dd747cb53f2ccb5a5684ab6dcb536234802b8ed8577af0b49b1c80ca962bd79029185;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'he7ab8197c2c8ef0e6eb77bbd731c2bf06da527bfd0bba7c51a3bfea2275663f4038233f2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h166eba3f15cedc3a1104e5d7485ee13e3ae391ab6ff3d3d5551ddb385a719012cb90f220f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h11afd983514f2806a91f4a6d8778a6d89085b2cc27f46ef3480a0a8467b16344efe780693;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf724d0d14611307ba8fcec8fa622f0ac731cb8af3f3897dcdbf7a632dfb59ce870d9e4be;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hfa3654b345a3b594e9ce0a660e31a5b61b453a55cc1471c6291e60b9f131cf8d458717d5;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h12c539a81190b93f334f759e0cd9070d37000b7f6bcdfcaaf22d3eab8cb5f85fe33cce173;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h22275dfb438b7ff06cf275a71a3aa78e01c1dce65ebfc3e23226cd07a41378fa38cc0133;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d462d93d6d57764482ee341ceaaf3dd6e9157071c4e1a0edfafb4e4c921893ad26138f44;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h71257d94fbd97f205925524890523003b921991d3cb80ba28376f7b7ebcda3f047328f39;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc15b6a80bdebfc82641bd34fc78f5558c71d5d6e970d56b163d651a0d69232897f927adf;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ef11d8bd1ce4cd4c9f3e4cbf796cbb5fef9ecbc2dda89773b40490c51e607600c0883718;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf1cc44d0f9adec648abcedb784a44039387c3455cc7cd0a32143a2a257d6b444ed0fec5a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h715765f3b262e6f345a4a1b0e76941949e1baf803bd613a453129908d943516c6541d4c4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h160ca5570bf545f32d7df3a2277f1d72302b34eecee44f9a9bef516db7413479e0bbf3330;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h9fac2460307449b36e876ea96acbb398b632768cc475b2981a5e9800ed50e1525e739134;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h5ecb6b6bc3731c83d8f75177bdfbaa270edb3e4a66c5b9832f7c0e09705f8b007515c856;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h72aa684dcb3ddde4e6b97996ac833ca276b4f01e4b7face0016362fedcbb74f461316631;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1bbce7bf50be6cfa23d270fde63e3f4d0c5f4d809c8cfbf1c6e36a2c96313fe15b1eb183b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b01b99d18aa753d5a77765c83e3215f7383510495201257dbf6663b5530819484daf388b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h134ac6d1eeba6a790e4860a7ccfde0d2d9c6b1df025a30a1dbb9d8ce7b472ab630f0bafcc;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1faec1e862e6c6f98f36b301851c64fd40b6503f461af1772d07168402b5fef200e79d43c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h14db0eaea84e4d5f34b5f3963c5d0069a3f3a64e2dcdbf05d381d1903d41e7d2b715ec341;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf1fbc01c9a07d00944d2dbbc592620d49c79db6bb690f5b4172f88e99584d731b501947c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a83187d83c4749a334d0b16c96808dc2c690acfa6822f9d620d53eb56db29d736a35c270;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ef3be0d9f8f3f69ae2b50d84c1c328127c6539937dec8c378270cf42c06c2f85ee85fefe;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b927d414eec86f8f892fdb231f9b535e688b3d10cbbc2fde88a2ef30cb2c2cc57e8f206b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc656a86ae69c92f6c2f2d8792f01f3b3e740a607ab9ddcf9106687e4dcb7620ae1101313;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h12d3ed19c34a3ef8bea0da02b74bfd7caea8c2930f052b521edf2f6e233bf1aab32e7e5af;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h67c6014fa7a311933665f5677710ac66c3ffed5143d95e85797754c0c8cbc8e157cb2795;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'haa656a6b94adda5e55621f7917b15c7c14a6fb2b3eb7896fcae9800a18a714e51e3acc3b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc0240154fd59d6e56f2f82359a0e07fce3fada2a1b98d37435969141c238e7b22c78325c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h11939d7d81086e541fbe8e7a42842ba403d7c0b53d377960f5b425d6dac24b3c6bbba2d3c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1de891284fe74d89fcd3cca6295832a450f0ac0a93639af868c539011c3501f71cb7fc49f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb72ad7b14cb077ac6c331546b95cc357408c3c7f8c6384c4acf37af5dd243b44923ad42c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e96fa975fe23f6f0e44ebca217cea3855a7a9c760f20d11ac1c13eeba4cb076c0fa2cc11;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h10a07941e8505e73e45f4c1e2a40c26390d8b2ed49bddfa3c39f3f6dbabf3ec0197425638;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f2fe85d7aff9f87d33bf65f4cd6c2cc46dff8034e9a8553308fc243a678a7c1f18aef412;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d831421cfd59444e2455f240a46116a8c56692525ef38892b0a110d4a2c2eb943865483e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1621fb814eaa46e3c04ab94fe2cb7deaf88f87ebdcdd4d1432165035d92f47431c04c8d48;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h17793b677b2f17aa0682975903b6e954abc20fe6381a0537186ba1ee903763cf74af62e5e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hcab7e222641674084f9eeb39c6708b19edc86827626a93e465465737566a8bf2f087f669;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c66df23df84b7a3e1800a44c31aaef81fe260c4679fddfc8e53fd5e79f2a3750b4109e15;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h4b0a18a8dc2effc99699a37e43de335b04316c546f77da4ae43040103da9e9bd17b4bdab;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h18e1a6f6e8500b1587a5c3cd3f9ce4780ec1e3ff1504d745c88f5570b97db480cac675247;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h6cd8e52b403ebdaf7b2204c1a5b358a1083fc030792d5e87a721df0820c835247f841f24;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ced78005196b48d30206233912d99fabe155b5b6534126da8b6539b6b5cc18cf2ea1912f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h137e3bd29ee378f06966e21584b965d616bbf2cc5d5d53324c85f6781f2bcbec11c6aee45;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1142d2b400e6bc54cf7f3d5328a792f78537268583ca2d477f7a5e23b075b859adb8f1b36;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h16705de976d7430afe1b1a64838876a0d9ce8e96bcf1abc7b39de00233227028cc3297354;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h301dc1f9e2a1036c3c34b93d46a9ceec6e377ff5c91f2e5a23e7c1f6eb02e218d97bd03;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h68c2f249daa09182c68682a5b67723acda1abbac97099ecb2935c0dd9e75001475133c28;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e9215a34724aff606adfb8881cb4745541e4a14d2044cdebafd7c356942458e4e1ac9b48;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a069b4defa032df817e00b515a9a6df42e16a83400af5fb8b177c364275a59d07309cf94;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb2407bc1e04ab58fc3bad6fdc3c6a262cc5056ddf6ca1d099de345ae8af0601d477464e4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h84093a942dda2c4faccbb39515850d9152d0e9bbc294376ab0957460f5c61008e390a967;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb23ad842860ed63a4b9a369029cff5e4477387e1c38d837bc6c79de1b8f426ac91777420;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1fa782e6369cd8463ae4cb276ebceeaf6cf42907749070e3f080dcf3c03f35e3ffa2a7c3b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h146d94ca69da8bbeddc73017ff9a5315924934e52f86058abec7bc0372b756a27d8961b78;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h3cb8ba002a2d1e3dd8c3a75b92c20ea48792ff6366ef3d4fc57a6c7d1d4324a7d7b97bd;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e6eb254c4fbdc0801ffd4ca134ce6766cd318ddb61e46e1ccfa965a61da6067dcde65c7a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h2948bb4cf7d3e1cd3100e8aa7419c47c2d841f11249ea85d1f1a1c5c8ca4b9db2a25eaf7;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hfd4982a7fe5d477df23ba98f356b763a213230bb3194fac4d4944e714431e0c154a98c6e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h54b06e0a8f4d03384632a646d864139137a9a9ff179d2cfdd43f22e8c2f8de74b600b92;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c59714b298dec0a51424e84c044194349e37a95038ca51deb1a392ccbe576388eeca5e16;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h8e009d54b3f333967cdcd4871d693dddaa9425a738c644a0b7c087c834e06b6496872c0c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hdc4e55416ec1c0c0c8af377764d4c60bae8564c6bf7b9ab944cce6b686daf8044aaacae4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h319d5171150f36aa160f3197148ed924a9c1437b0d9e85c1b9100f601281878fe018e39a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h160beb9793bfbdb9723c0a52bfbc5af936aaef09e5dfc5fa201bd2b4d2abb5dbeae6c0a38;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c6c0e8ee0f835601020a5ce91c46354343003dd7fef39071ad7cc8ebba250371c35a0427;
        #1
        $finish();
    end
endmodule
