module testbench();
    reg [0:0] src0;
    reg [1:0] src1;
    reg [2:0] src2;
    reg [3:0] src3;
    reg [4:0] src4;
    reg [5:0] src5;
    reg [6:0] src6;
    reg [7:0] src7;
    reg [8:0] src8;
    reg [9:0] src9;
    reg [10:0] src10;
    reg [9:0] src11;
    reg [8:0] src12;
    reg [7:0] src13;
    reg [6:0] src14;
    reg [5:0] src15;
    reg [4:0] src16;
    reg [3:0] src17;
    reg [2:0] src18;
    reg [1:0] src19;
    reg [0:0] src20;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [21:0] srcsum;
    wire [21:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22));
    assign srcsum = ((src0[0])<<0) + ((src1[0] + src1[1])<<1) + ((src2[0] + src2[1] + src2[2])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3])<<17) + ((src18[0] + src18[1] + src18[2])<<18) + ((src19[0] + src19[1])<<19) + ((src20[0])<<20);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1ffffffffffffffffffffffffffffff;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h33e497d94fa3fffc49b9b723d8feab;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hdafad417cd26fba17656a5c62e3664;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h199d2ee21a3e990a3ad8e751bed4de5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h18b7ef9a40e1cf0fa8ffdba78bfb96e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h10147c0bb0869819df38e6dcbb629ef;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1c8cf8e346e9b10cef101939eefa0ee;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hff2893f46fc4035db296beea444268;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1b70265ec405be3e939109767a58f82;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h906cdbadfedf6f533a17a1ac27875e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h11a37cdc524cd8a75732d8142904130;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h18fd370f9158ba06d62c0b38f009f3b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h724d74c03d334319281b3a7319d71a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h12750d3e311c8ae42052471f3be432f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hec962580b02756b23f47fdafe2f4cf;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1527d073c3ec8e1c259d9fd957f7385;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1cd3fa16f959cdc075d40aaa2c7121d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h5de1100c903722d6a9c028fb233c30;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hea7dfbdfccbbeca8ef6d583ef064f2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h141956d5cea2ab7ba2fc839fe0ffef1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1c3ea57b945aad5e2a9d91d0b0b7c32;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h196c0cdc47d5d8c94f3772aac125215;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h9323c54ccbe60399c940dc3ee134e8;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h13f45591c8e938f30d1c40703d7385b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h5212f177a382667fa6bddab219a362;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h90d283c9989480cdd616de680f9b3d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1d6ff3795611b889a5e3b89e9eb6f8b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1d6d743d62ac8ab6e0d89023acf5adf;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h839df7f0c78306a6651e45997e091a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h186783cec665968a798e5c263b55ed2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h170d3dcf1c0a802de398ff63d33c2df;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1e599dde7c16ba06c7e4b943d82c1f9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hddadf53b0b8acaa4a55adccd9363d9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h12a2a73469c5b417cfe222d6fe2ad73;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h10dd68ec82b0d31e5360a2d32b0f50d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h7bcb15c5535b1a23a9e851f0be82be;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h12a181115096a2c7c608912bc818338;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd25ded79ee9da04409218f4d93ac79;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h3dc536fa27a805a253c84cc08d8b97;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h6128cf4ad6c0d5f8ff94d0ca294478;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1b47c65b423aaa7be1b8b3333d08051;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd1faa5a0bd63a2bb0a19134e6475fe;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h19a424c8869b21cb2ca501b9e611aef;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h47181989e04edbbea01c36c7d884f2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1ffe9b15f3299bf106de615747f1348;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h7e19d20648c3d1fb9e07a033fbbb50;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1f9cc57d6ac8a63e116a650d7e7e210;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h19a4e9e4d4e5a7a0ac9729250f57134;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h9694469819db3c9fe2bc8b552c95a0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h7a36d5f9605f8aca8aba7c06b1af93;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1bd1c17137296c5163a3472dbff629f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1c96312d872286c0444f4fe96538d7b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h147710a8189f43da4b171edc73803e7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1c0d4b4481565d1387f8c3a2f35f2df;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h14a853b928aeec1187d9171c7ef5b81;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h80fb6ad9c80239bdddd96fb26f148f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h183d2564e3309551d04b2f701770536;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h886dfa15f0f52af21fbd37391a3d34;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h4a5a93a18730a285293f19c3af4980;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h105ac4e5377c01faf0faf9ccadd6fb;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hfce582d162c7151b86e192aea9c8b0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1a7beb8ce64c3babd2e311c0b5abcc;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1951fdd50643b6908b2697a3081bc9b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h10b2fb365c876ab3b0b1f30cc5f94bc;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hf31101478920b7744a904b66b666bc;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h178fbfa1b211d450c5ddf1555a1a067;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hac7bd4f6c6bc452c1f132ce7a882dd;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1ca674633516c372a90cf56cb631273;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h93e2d0474f7168f33c52c632713ad9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1fdef8139766a5a3ef457d21376522a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hfb9967aeee151201c28d920095922b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hc2d53f9d9012afb67ab719d0d989e7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h12ee8628c8d08a2317c4c93d6a6527c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h11da43746323cd1c10804c1b2f8a9be;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hafe3c58abc6e86a253df343df04233;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h57e5e46971971390654c5e48259fa8;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hb33dd8ac1e22b24fb76464640b5e98;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h19132e791690f4b99fbe8d0e1ff7924;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h9686874fc4cecbe77530a70c911791;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h5bea6cb0a4e401a81eef47351bf620;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h848fb51ccc0746fab099e15ad0d617;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h19fd34ffde9b38eb69f804b93bb64f8;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h10a1e0f1f1f56d123404861b2c69f08;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h77234d32477922dd3638f4e3e33861;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h17600c1928a102d281685b22773b308;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h7af74bb3a37a48ca0a7fea37f0f833;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h5aed63f2bd1fb60d37b6619e35efea;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1589c7d958d257b6684e45d17cd82e4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1ef1d4624baada2dec10821d295a95;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hff31324e8e18d478e007211cd48935;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd5f84203cc95c9775fcbb253270a4a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h15e37fce89e1a72719ff7a86e41a411;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1ebde317ecb5e726223fdf5717d9ca9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1774caff23cb11dc4187e8b96d2f8ff;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h4f358e0e602df5cf7c5f470f59ec0b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1f2e9db730ac74368b873a985c222f6;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1f342c5bd69aee437b4a97f38f499e9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1eeecf5f1866ff2b966d223f65857c8;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h16b1c580e34903a6b9795b1681c85e5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h6ae9a45181886edd0f40d7755721d3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h16bc4da0c542004cde70308e172feb7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h19b009307cdef735f6e07f50aeee8d7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h132343ad2f07957308bb47edf3da0a6;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h403c96f877ba7f4107be9286f5f34f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1221734ec8ee42dfd5c6929d8795c63;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1bfea19be0d218215493f984b9ec22c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1565295d8fad84c6079dab1a2e1ba36;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1e0e6ab871409d207b57c6aa85865a4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1911a2f8a775d98ad5d824432bc8b08;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h17b160001948447738f79843dad9398;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h13f8b8c8f70f41d7f86e72dcde26f52;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hecc49f63d64a29234aae8bfa867cd1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hdedcf666767a3f4af4cd6d21407687;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hddd3470080ed39f3a80476d7d2ada0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h18eb85bcaef282ca8d4fe5bae7e3772;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd4033ad40671579f70229c873fe1d0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'he8c7bdda0f08165dcc87221b66afe1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hf62137e0e95a75bf13d29580768a1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h10371c804cb6f00d6d3c0b666c80826;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h2f5dec9cf19b952792ee4a70c133ba;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h14b8292eb9d50b91fc9ff8437686b08;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'he16956197ff86ab5b8769813f02aea;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h11f0cb9e703c8eb4da83999926aa63c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h15550f04e474cd47b6df940f626ee5a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'he2f165cded3c5e2a6c16aaaeeb89b9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h583a49a5c879c9dbd973e902df5685;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h4b83ac508ad5158352b22ab53e5e12;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hdc8364c76de610ce0c422087a741a4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h138f26117d7f51e7c6402f8bb9267b0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h89c718a0a49716a30c5d1abbfe215d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd783f85699b770858fe51d1906828b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1c3b0fd1017ba343e2e24de9b9bd023;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1c28f550f7db3862ad0391a8cb187ce;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'he2dfe96d720a5c6b66bc0c8ec9ff4c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hcc8ed4aedcd0155f3b3abd792e90c7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h10cc679282e6af7c9cf2f55ea3779c1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h12c944d01df3f17c340fefdd7f0087d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h18a9fd7936d28108bd68bae2c311d01;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hc79c87c35a7d4e15ccce893dc15162;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h9fc2511a1392c194ac5c2bfb3b39b6;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hb51d15409c1446f833540fed3f7ba6;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd6c17994e13d10cdd5dc87a7efe072;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1a8686a5d177a24564b212f244c1562;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1ade5640906264d169a4db3ac32f37a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h118dc595c5d1378bc2d75d8d2120c7a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h106c0f0248e934810918a0bed73475f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1fae13a49046db60b9b8deacf7f672b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hf26ddfaac5a753fba859856f4f048d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h12059e1929587aba2f9d18e84122b6d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1a99a53b56ebd61156ce06adea4f376;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h67486d9e46d69c754ca74a0bc61ddd;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h143a430ae395d25f2fa1dcb51377732;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h174a7e94be00ed5054d0c8f2a37e50e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1fddda8b35a4555903d6f8c30b88c30;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1fc723dcd7a3268eb23a6d3c3563b89;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'he79bc0fa3bfabf3d3462b5c4c3e047;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hcb61eb06d654d1ae8f703df828e633;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h16d92181c4e0e93c130a20a4aece04e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hfe0e2446fe66015743c726b690e878;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'had36d6a5112f7e0405d7fd51bf67b2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h132a99a291ce56c7c64af409d8d15a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h87fab0ffafc29b556c0917402d82c2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'he349bd5ace69e0de0ebaa04c2ed70a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hdcdfac2ff499807cfbd0c8fa766d31;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h17a23ab8f73305fa75a6719e3138a14;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1fa9d1a79407a58b98dfc08f843096c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h2b2601acf897a7ab4760abf6f1c1ce;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h280d138cf71adb0a9d615441de88d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1b7622e7ea463f7bf3c176263ef649f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1c0f76208e2b344a0a2e3cdc79d53af;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1f466997ca5b8613f1cd29659765b4e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1cc3d3a5294eb93c9dec51ce07bd482;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1ed784405160f8abe9ca9a16f49c441;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h136cae26e3c5694ff74d8df618c99d1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1aaa57c75bd4f18707f46a6c333c202;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1478aa8cd816f09add8f7a8b641717c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hb779d009d48c8d9444d899ee1c0b0d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h81415639a6a69238c607f554fc0f6c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h15f8ccf8429863713d0df0008e380cd;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1c052cdd3d0b81f94164d888e92b359;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h98d62555699600779996cdf41f225d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'he8ddaab8c30454b3cbec1de13b0d2a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'he722260e56e0cdde71901c7ee8d440;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h17b576ae944125725707514305f3a29;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h26a684555e6c292d4383b2ababf2d4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h86f29c3caf6aebd85b0e34c389f339;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1dc842ca99f897de299029228be48fb;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h52c4a3d2e860149ee9dc89d5e72dfe;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h15811bea47cd4ba02faf9d48b9ac59b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h14ed0764358e82f942cb3c24a9e3335;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd58447fd59f10dab90b323f59d2be5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hdaa3aec34f9f72accb57a680b3a2bc;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h16227e2024b1b88b9db9ad6da4c1577;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h153d0ea89989c4a91e3ade8b5793bf7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'had69745393d3c4d750b30e9811f06d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hb58d7b232f58e0f7ce2d4bce07b274;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h13f816c93c7009014a79bb7b492e5f8;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1054a2c2dc66a74442d869fb4436bbc;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h2f2e943c2037eacd6a716c21d5df0b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1e1a55373383dbc6f0fbd6f6f43a4dd;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1feb4af75db0d759195ae5f8bc64463;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h81cc5a18e46a4d7d7f062a62f51893;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1b0bc944b386f70bc41f173e98105df;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h120f6b2c3d5ccafe8addabf5c3a9a97;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h174eb86fa1c5e679c0aba05aad675c1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1650268b2ec92e64a43d31581b179a5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h43d023aba63699fbe688271dd3a430;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h17e80bb967568cb1fdd79f29acc19ea;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1e26be1ad9465a7b521baaa25aace20;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1ad220dc9ea3315945c0e5f7c8d1251;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'ha0794f62865e34470665f87c8b42e0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h14073816fb2e73d2a630ca0d81cc2d1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h14bdc1de99496c8d06a3cc20a9d6907;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h188a4c04b58873efaffd6a1e93bac7f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1b07e9fb6ffd9fdc00aec8aecbe4ddd;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h82c916a70904d93e7bfcfb50d9d930;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h11e4698eb302169fc651862de66ec98;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h660cfac8ee0e090ead61a21ab9bce2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'heaa19d18ed7f81a32b628587a3e61f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hb8dc1ba107b8ca9a6177374cb49a6;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1a7b3bcfa29658b7126909c238dda5f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1691641694e657ebe2183e06022ff67;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h15bde0e355e89f60bcc86f3e955527e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h3966c72b9ce8a60152091d8e6b741d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h19c82eb42305007bdcffd4d4e4cba78;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1e47afe81f83b3f9b91bd24cecdd409;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1bf54f3bfc47d73aee8d45263f70c20;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hfa9ba0b33c0d8266219271cd1299fb;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1594f111dcb53f3985cdbcf6a955eab;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h140490c77d6d9b38ba3b51cdb47c5b5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h9a2ef2fde5a702214a49b0b55066f6;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h2cbe35a1ffe15a375cc72a186c628a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1b59e35e1aa7e01d0fce21a7e1140b5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h3d29590b1d0ce7590a14bb9b2f6446;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h5788cd8fb45745116f5128bbf4b819;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1a9e63f2dec8adc9b34ae9c20fa68c9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hae72440c8dcaecdf5dec9208e11414;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1e5797ddb8da2b1928406a41d3df0b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hfc28a922f0dc5aa58e1fdc6d6652a5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h17477f76f8db7b04d577e08800c8af7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h2655ad38a9ec6264cb0bbc5ade0e8;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1689d7ffd4227373a057ea9e6b6c650;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h126f5599fd91e421b9613907420d9a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h19a0ffe1685067dfc14499ba7e91d94;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1547b1f5b673d6aaf49c6c4bba8b1fb;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h33c7646e6ca77b559247aec4ca0977;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h182873bce73d1a5733977564fa8f4a3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h18395bf786bd421469ff031c5d29658;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hf76e38d5085bb020e85559b425bae7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h2ba801e1237d6d6a8db4ed9c774228;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h8a24a13f94894c5d62443bd0c659d7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hb4d101aee5b9d5da93122e86d6455a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h159b9b7bc355fc1e2d485bf922bd33f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h122724bc69d859b605bc0b35086821c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1800f03f08aac2a2a91ad0b291833a8;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h189e7fd8a372143276b1e86b4bbb8c8;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h11cc8e493b2b3e28cf3f4ba25df2296;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'he3b7d30fd8836864c08800406c3c37;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'he2a23271e38894344a338d57a0189c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'ha4b3c17344a6b16a41d3e5161358f7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hc98be32336e123a06087c947d343b3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd1c507bd525a11f920b3d46e7e7f07;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h44363d436e99e601fe9cdf5fcf904c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hb15008c6e3711ade208ec4002a49ec;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1d93f52a231eddc5981b6281d7ff172;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hfeba0d66cef4cb38ec26f5fb584390;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd840cb7203aa823151f4928d824b64;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1bbd3903a77eff779413778e3f865e0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h19a4bada33a47bbb91849a6881e50bd;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h12270373a28fd5c255f8d62adef3b93;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h9d6aab9133119aa8ed91c1bab8d762;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1bdd39665034a4ab48885404bf9478e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1071614ca550f0df1d0bc7d463e5ced;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hcfdd4bb3b16dfd3c13ddc10854ee88;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h77f3c02a656ac8cb26496e516c4cb7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h4151238d083bb14e79f875c2b2e5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h194ce21bfe3086a59825aef9d7f01;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'ha52b0a46f3ab01508ceedaf221b6e1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h195014539a6f709bce46135951949f6;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1995816f1da0442016af429d7ac3faf;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hdafa068d14ed15f4071ae5de4e13d9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1bd46c48cb858dc812ce6114c00b2a3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1e759dba58a9287ec182dfca07ca47f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'he4ec47da89dad12ef131c4b51d6027;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h17a8f773e7ff0d5f55d6f5bc8ff5ee0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h3905d9588431f53ca0ed286e68fdab;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1482b3e196171312889bb41520b7aed;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h10564a15b02f016fe85fed5f25df8f9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1bb2b02feeb4894162e8aa1d49ab98c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'he7dea46422937e80a00bd82de15bfe;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hb7bc921c2a5cfc51818a5cc393bf9f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1988b34af9cc33370b14256d7454582;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h196c428baf8c2d98909410840ec270;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1185e24e05dd7ca1cbb8da2df283285;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1d54256b320c7bda1d9e7628b72ed3c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h15e360902ea8ea75a4ae6d87cd2c630;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hec40842e3eabdaf01d5aaf9db85d37;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hc08984bedae086e9b22e3dbe9eedd3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1cd16fc708dc1e15071a6fd0493615;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h103f6da9f3aa8f97cb79bdb81d9293f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hb1ec57803ab3fbcbbb4e98f04cb5df;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h832f298b380a8bea40880d28ce510d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1c79e1dffcda6664c5c160c1541a5f6;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h516679e28754f23fc966d48a91a0a6;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1a9dca80a2d7db4447d1bca48ace6c8;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1f4427f40d871e06a9dd75c778f7fe1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h314a52757d6ba7d0ef2c38ecc1bbef;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hdd5b38649e7f1dd6da2b331b208914;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h121d1da290ad8fee3431d34f8dd5387;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h7bfcca5e9db864cd37bdf8d8671bbf;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h4bae41cf883e0689ab8e7703ce552d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h22f0877f59d84e65756046d58bb1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h5bcbe1edb97404da0dc35f4a5b786;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h16e8b8819208a6b120c4e1aab227303;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h107f454610b4513a564f3a71d100d39;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h129214a260a9d62e67a14ae9fa08bb7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h4f2190993596d8b89142782733a783;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hb235fdd2aeb88e7a167a61b42a970c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h174f063c247a5bc6a4ed96900cc6931;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1ec5e178ae8c380ba9501d16eb3b5cc;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h128cadff47c61591612e4b17f97c602;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1d0f1de5f30f7655475cf20a271703a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h5706148359f698b7a12496e2352b0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h114a42784a729d0d8243c340f0a4b1f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd5efffbc9f85374d6f76439f2df3d6;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h404775eb018bae79b0110bd9a90cf2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hbc23da9e05d1cef0d9af244421f6f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1f8ab2c2147f9977a7e9cde6cd19897;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1a263d3c5ab5824db7ea57c08a2c6dc;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1b2981b8e66851829d8927a8a1addc8;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd5bab104e19786948bcf0a1682da70;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1473d4bc7ebd8427546165b1bb34348;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hed7d9b491847f6108d740c2b7ec8d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1346cae622d618324f56549158e907;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h12576ff8110cf6814ef62bc36ee1cb8;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h19fbb233369f3a59f0a609eee827b03;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1890d215da883486a229f1f39cc8f16;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h18d8067403e6abe73c40fc66e34d25f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1c35cf340846ecbd5f6a0314218148c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h21e6e8a4ce29ccd1026cf05b9b8ca1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1c8c16ed2aa2c570fd9f153918ae3fe;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h6580750bad50dbef6d152576214969;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h82b0609616208c6bf8c6ae3d8b0e9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h18f962919277614d377b415b905c61d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h135d211f8574a14241ee8f49acc3da1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1e5f82a319b945999e67c82219c436;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h99f3309c0df7dfd05ad81c40676382;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h11f5115c7e18ad13da5411cfe3017d0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1c768bfb3a7d9302189b656b13a1a6e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1d9556264ab8fe689fb76384e60cc55;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hadc20ad2bbe8e5c254024e53936aed;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h19462f1ffd6500e6d2cc8a4e03e03f9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1f5257ba4ece0bf1b635e3982dde1c2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1354d78f927c73160c28ec105aab269;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h18976947828433a9319a84cc67c3ceb;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h18b03c2e8cdc9ae47942ebc9fc14292;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1876d6fd49c266771eceac7493fec48;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h891bb912b9de6bb779587009892179;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h13abd971bb5ff1f6cf21db92e32fd70;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1eb248fb3a804b5959171f8491cbb76;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h194b22ddf36ae67aa354938d80cff19;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h11c555e8a66d7fdab1cf9a652795001;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h28483a314bd27fa667713b3e69e69e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h103636e273db1f8c340ce5a361611bb;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hc67b2a3a0ec7a6c87a394dea825ca7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'he66ba613b9c609a33b618323ca50ce;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hf41472691ccc20feba34c751401149;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hf6ac0df9998377dec73e55fe5c6beb;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h10353387ff68bd0b314f70ee729571c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h11d8939904ab70bf84819932c4aff85;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h4fe90ff841bc24092111a2550fed38;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h2740a24201e0f1e9868324fb6758d6;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h534655df0cf674c2eeee83b8211c03;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h6b5687c7ace639c7a49290b061530;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h73e9c62835d68f2c57095e3b15376c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h11845ef603ec66d2e2ccb1803236ff1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h8af43a44279addb966f8f63cd80a83;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h162f5b366f3318e56ab86b96873d742;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1f01ca0989038dc7ed4b4eab1a4a824;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1f2b8c20db4152bbc9b8a3d852932c9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h111626441c39839810c69a7bb3e70c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1d54c2b144959fc046ab9dd287a5735;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1edf7e35cfdde45dbcde9717c908ba2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1e7688e68b7cd4e84c96d9750f9ff19;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1cb6891fee292e9ff1c7a9ea0bd012;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h10d5370c7b40c04bc1ea49d56550dce;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'ha5ea6a2f95df62dba5e930a1a659f0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h138337b46b0c86bf3511b8586f51621;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hdedc4fe04a9bbbaae022225968f3de;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hbbf3241dd707ea4b6041851c00c249;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h2abaaddc03f85259a33c638b925008;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1ae0f84e6fbde051d3aa86dd3a319fc;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1bab9423d8574aef3a59adec4f35c8b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h118fb4a7f4e4a6c21f96c0df80c0690;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1345140873b23ba92d8a8f3aaec6d4a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h15a2e0690cc0fde8a3e519ee1bc4d2d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'ha772310e2f632e225282f96aaa2992;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h151b8f0392a28cbefcc7941e9c92fac;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1c359b5a9ad76af40ab460ad6a69e8;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h96d97f93b3349f24396b7549fb9eaa;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h3aeb8b25b1dca030fd42fa847e7f62;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hb71bc2341174d40d306a8f2e333723;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1cb0065e04aa043881c0d26552e07e8;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h446a00879b0b30e164a9ad2597924a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h9f9e81f8bde94560633e08ba611056;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h325661ab32b19bd490a1bd5feb1fab;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1d8fb4d5d4632f8f6e624716c407dca;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h128cab923a760897d266145be979ade;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h10a524b55476ba25f6519284ef0bbf2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h479f49878b0d722fa7daceb4a70cf0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h2b4c70df0eb3cc378cacded50fe08d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h16c76964bf1a96f1c93560e000601a2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h123338db271e83cd12a73d0d2159aa6;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h12583d118e96ce75ec3dfbab799e5ee;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h673c0a2b263220fc4b1fd7a6588e3b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hb34718d42e79ec4a61b48c562d3c6b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h16c43c7a3ed3b09a70edd5c98f8580a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h9f4418f8eb775b674f229bf4a6b569;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h2bdcffeb528ca72d06f52d7fcb15a2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h62a2715958b42eb009b0f94bddc2a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h3ad00e4ba0febaae15f8146ed8d6d8;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h2dc0e95d32dce0e64699e33d5cc470;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hfe1044aa87484d8ab6e9f34203394d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hc99bea289b8b26b5a1309a5ea281c0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1551997305bf577eca03ccbb7378f55;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hbf0c2e56d126222696cf9a819c6b53;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h8030bb6d4f790e3c848a8eddfa5b1b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hce75766dab0e395816a77684d05a45;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1cf45a1413147f8e79d85a1bf2e649b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1c8e1df62ed8704dc6b22910e390c7d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1e787d3f12821a33fb0e15b0a15652f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hba050ae80bd7eca5308a2e01581ddb;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h173048367232ff94bdef640988bd5e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hdf00025c4f736b08b7780f403711a7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hb1a8cdf05960e44c7c4ba7896989e6;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h79090f259e991e1665c1592f09bcfe;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1b659840de37b1c60fd1339db1fba47;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h15cf844b4e6c6bdba739c73f2e4b426;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1b642aa904c4565aef952931d2a0cc5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hf9085244c1dc92fcdf095f87ab535a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'he06c29b0df917464ace5e0d9e5335d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h3f9b77afda3bb9e46d02f114dc8356;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hb670cac75bbffa6cb947346f4ab802;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h16fd4ee277f58d29b686970fd65baf;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h11031c49716257f70810cb5b01d52cc;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h73b671b1765aad2c1a3d0967051d8;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1109ceec2a5914033db92b826493f8a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h84be1a2075bbf0a8fa7b7260a812bc;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hfb6fc4200563ad884d2a1f582471fc;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h18bfd04278b7e4db9c88152ea71e0cc;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h3d40fdab2f7e214eaacdf8dd2b58aa;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h12765a0f880ff44872dcff3c2df834;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h19bd228e4b2d55abec360717f52b3c3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h3881eb6c79f745208765b51b142124;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h16c9f129c7f22f99170a45e7b9ae656;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h14f9500b4a25f9397870aae5998ac0b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h83b84f966525a0995c2e7ee90c844;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h15975d69e4400eb7127b9f06ee31d15;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'haa9ad4952704c98b0b83c1a39c0957;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h491b9f6d14077188487611d4a1327a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd803ee62d9767dad0b7e91420be9e8;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1b5ce9c6608ea3c1c7d3d3e8f5963cb;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h668dc08cd148ee1f51ade84a4de737;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h9eb2408b1b31e346721272f1c76976;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'ha73e5258805b6e67fb18819146e7bd;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h10092b09bf4c40cbf6abff78012994a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h9bf5b7a5ba21acf0e833c2a05586ef;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h16fa8c6d3f9e6ed944982564ad1a11f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hcbef8cb90b6419a85a53b63b5739fb;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h8303700ff238c1655c1b061cbca1a1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1e552a6a715c9495a0e8a031c49b5ac;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h5fd86ed00cb9cb63da867213af0b5c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h61fae42f6e15c9f65a124f16cd1a52;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h53a5bbc6ffdfeef626da6bf7e81cc3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1b40eee62c2bbea43b8b7490aac68e2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hb25634b5b90653e74b1cd1ce088dac;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h14c3b3ca296ca23bd45aaaf5a572c49;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h58fa3c75af3e24728fc62d55d4c585;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h3b55cc1ed71bec52050b7feb5453e2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1bbc673663c2f83bc9c54b2396e3de1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h3e42634be342672901ed9fde88abb1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h9a9fd5acafce74d3330c0017f609;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1af122070b049a2a4ed11191b6d134e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1f821b2ab6bd5cf5dada7093ae9ce3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h7d9c273c4307df076a8ce84d96bdce;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hc004856c4f00188129c5bef80a525b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h19df127e1df88453233b1307594221d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h8dad79916bf6167fdfb20171a5ade;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1ab2415c7bc6535a40291373aa9705a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h17c0ca223c09e1059702afafa5bb2e2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hacb7f3f6c67f5312f3bc9d47de94d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h13115dfe228d214a7ef4a354252aa00;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hb54d249f33509fcee5d13e6a76648f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h9671bee37447d961bd420bbecbc151;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hab7910ce8a726f42e13fad061bfca;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h3edb8ca1ed1710b6acfadd1a7ab80b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'he09c0e7e98615d9e01db82771b87ae;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hc7cdf473bbf9c5de16121ab1ae4d14;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hecd36d35c4f8b79397318667a818ac;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1924282d6230f3fd66e0972992312e5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'he66b68a988ffdb5e59918133420569;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h641219199c60753c8c9df2326227cf;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1a797c4db32d1f0eb7bcbadd0a812b7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h600006ac4aa26d812f947dc3b9189d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h8a74632dd701250e60f3ffecae77c0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h15e0b262de889873caeac64ae73c7b8;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hc7b37e740e4da7f82c85856b475ceb;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h17124897e63e9c0c495e3fbcbf3cd6b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h47f06977af15950d8c02e0ad21b952;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h666d29c4ec570743124af10c931ac4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1321d605e550489b33473961cd2338c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hce25a0fafc42f80f4e1cb59934ecca;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'ha3119301435744e28782525b34d660;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hf4dd584070d649d92bed8855ceb4b6;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h781c29a17e18039ce96d0c8a5d9b37;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hb1ecb946e720167af78233805cbec7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1126035863a1fcf03509aedd0e11c2a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h11cd46e847c45dbbdd32efaf766fd59;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h16ca7e71cce8e6e474f9ef750e0c861;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h11c42973172b59c4215a8b6999e192b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h199fa76c689286a3d2f8909172652e9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h18526a6f2cc0f1f0f34ca6f0c16564b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1889ed524d95575bad31e5bc8d97e51;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h12a80ff56dff5d69b608f1e1e5e2242;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h13b57f954cadd0151d10e9a56f5ccec;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hbed92c3ba8fc4d20318c845ba2fa8c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'ha8e791d32f1504ffc81e46c96bfc7c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hfec7958112c49a4223d49050e35686;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1316cd7d1b81c077b0b07b5baacae24;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h776d053849cb294454fdafc17f0154;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'had15eb2a5ed290817ae4cb3d1be4bd;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hb4a8e41182e5eff84d90401ccb8e60;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h7084ea3f082d9bcd09f804a0d3b84a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h102b8d4f665c8358211ab79c4b0b35b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h4771a092ab5e3b0b1873c77f634093;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h418cc721fb0bfe094a4f3a696b4b1e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h17869c9725f292799238c5885acdd97;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h158375ffa3e5fec8ef48f874753f9d6;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h14bf55c6c252e641ea40048f3c9e836;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1624f0fbe9205481f495d931de68c01;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1ff1eed9e7ea0646de051db85af8506;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'ha2af2f8cd12cb5de57d5846c00d4a8;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h50712686bb8d78e2e6f1f2b01c2dff;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h130cacb1e729885e81e31e62ba6f918;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1130a3e1b23a226228c1d9664655b61;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hfc5779a061747580cb97db9a699df;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h148377b81b8f78f5095651ff98f0cb9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h47b7f2f6c8658c610e24b5d66cd32;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'ha041c515520442cb5612889c6e2428;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hffb6e0380988e4660829a8d270df91;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h183f3cf1cbfae944e171cb12ad1f5cd;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h907208155caf7e3675a3953b758771;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h11ba6a9dfc9a51a360265549edb2a17;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h125234cfc2c0a8b6a834a3cb40fcba0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h4643b7d6741362ef8c12ad748add52;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h17a99a96dd8788b1734e5c61974987b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hb2404175e83f6b643c27159221347f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h9f41a018cbc483897e86c0adbd5ab7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hbd6b04623b2178d59a249d912f6d83;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'he544f2a0f4f063201f5afdca93c9f4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h140956e227beacba50d993457645ec8;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1bb9fd0ab883278ad4b61596729638d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h164b40bc912f591f744ee8ad0764893;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h2908108007bd6e3874759548ce1ba7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h4e04aa84d04051120a1b86c4684f28;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h7fec8e810a734a7c04e4f6f494ff0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1805803df557eabc20322860c218c48;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1a60fef3982b23190060fd9e5cd877f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1599c1136c35caa891b37e75eebd061;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1f74aacba5170a0d325074e78dbc406;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h4c9b9aecb088a5fd45ce3b09cfc4e9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h124b5ba16558fd12dd50682b796d35c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h16c8c90aca774ca775cfeb150137e1c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1feb0795848e6c1c966c6900b79f479;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1ce57b4b8fc85ee47164be7480bf081;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1fc6812699d7fa39d9431a3ad799c6c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h12a121befce9a0769eda269bb13aaff;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hf9aa4b41f997f9b3ad164e428098e6;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h170d84b99c08ba03f8f858b53ddbbe5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h12a741b88f6c1ab353f39adc6df1306;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hc958971e013db3e10547711edc08e4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h43b833581096adc24b5a81b8476677;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hc3e93f42523659017e3fd7de0f93a7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h82ab8515af574df34c4a5e7a4276c8;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd257f91482c886910fa754b789ea05;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h14c2f207de0f8f42eba9d3997603ce8;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h14ad98b1d4c791c9ce3d4a864d59cb7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h160e38b31fad9b29510605ee344a2c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1dc0e61f9015fa531ceef8f0216b9da;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h14cac3748fc3c65e27097254ef6b5d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'haf242670c7119edca2426841930435;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h8d3414bd79fc1663782f2abdad3bf7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h94ebcee9868b03108562d8870518ee;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1f35011f55e25e961d920899c69c15e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hfe7948f51a9b60bb82e0af8706984f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h5617efc8b3f70acc7fe291b3705d73;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h7e0c5f5b8353d41743864e17c1b91f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1984b5a79ba5eccd9e80ae79fa4a57c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h17f1b29173e1a536f86c327050badf7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1cbba4cb68a5a61e2f478088179d827;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h160d317ad6c646817721f6eeb047b9e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'he142c55ecfc5762851367daccdf151;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h17c10f1e23d618c6b860203df70dc27;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h15dc8db406b1ec4eb84ca74cca74242;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1f6e5c2fd7e5bfec8e30fcae7d5cf9f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h144947ebc956e35d6bc67b26481c904;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h9a54d06a88e1b8a8ceda5d76610ea2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hf404f23dc49376eaa363b53fcec637;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1aef819d86506a8917b0b2d3f5035bc;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h6061d492bda682a0ae0a50d145d508;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1a10339107f4402755abfef8fbaee9d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd4c5c33060bdb1b2411fa8635be85c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hbbc3293df441e09efdacf8b3b27515;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h982ee2eb388cafd69cf45734dc364d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1aefa9acea42b691422206aefed141b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h18187a0681c310393bcb84a8eec6f5e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1f177ec76fc6a5b01571c3173454a1d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h598df01d8ab23c3894d5b8b24f688b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h145404c1f36c9799454cee8970058c9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hc160b282e9e10c0fa77aee6f8adbe1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1ed1657caafdb9fae3af9440453147a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1b03ab00e5fba48b568867e63b2841f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h18219ac3848f96f002a062eb971821e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h34a62177a7cfc51b8f13f9f558560d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hcf3fd7945b2d59cea298eb15b6746e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1c24abb2ffa490b0cf8dd969c56598;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1c54d8db8d50cd118a941dae5e75316;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h6249268d83762698a168275118ec23;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h18a478afd2d0d55535bb760de70302c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h141a52ac15ec59b63cd1782bf84d300;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h13a23f372d32b02249e63f18c770185;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hac61cd8a784482b003cd753e47c7e5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hb14ed185382f3cd271da8744a85669;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h9a4e3cd042bf24f33ef689a51f0100;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1720b1247cc8f1a20cec17298b81ba2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h105d8deb7a64a79fbfa74ef78257d0b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hc5c80145168cb16ae8d264292f4e46;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h19f8e5c22de012284636ed8b93ec7b8;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hdef696b54e96d4147dc9a3cefbd948;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hb064e562a6ad0a8a7c28f17468ec1e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1c6f2042b323d25521cb0e2858cd698;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hf2cf585b7e79ea2f39f224583f313a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1239bebef62eecb8b59341e48a7f4df;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h3900d4db43f570dd59a466d88229ed;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h5c31f34b0a7f6e7a846e2c6af10a03;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h14bf4a52c2ea42ad737e6f0c7bffcab;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h7670f25fd268efa600342e407a91d6;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1f7477cd7aaf403357566ccffabf4d5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h164b587e44086872bd416f96b7acbca;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h44b90cd9b8e186fde3c3d4ea8d7af5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h8dca4064cee1e93a1a3094a5bd038e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1d67a9240881e033cd5061a23dee8e0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h31dd07a56c2694a6fc7cb5b09e49db;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1fe16caf5510d7d926c2bf28a8ab6b6;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hfca12ad7d0aa71f5467b2820fe37cc;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h222e218068e2cbb6258ae814804e83;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1676dea471c952e9904a520974cf44;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h12918a350667432dd03268b6ee7c586;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1c455b93c2b1d53e3ab45a9c5938da2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h132dd2c15f4d344cd9edb8334096768;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h78eb32dd381b5b28af0535763182f5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h123125582169928b7cce2c6bc55b0a3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h18fdc0bb8c43a20050f6417aa31c861;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h198f63425f1442823bac8f9cc6451b2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1eeec1af19eb9a398a5f5b91f9bbc5c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd7d465e65ff27f3af987e5eda774d6;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h12e7e6c3a5a81fed9db7ff0f3545f19;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h4a6182c94b2bb36df57c60ceee68b8;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h3aad41294efb391c183a6171e83beb;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h82153d0b9529ac8f5c2511578e2b21;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1b62c90a56484b824d849ce57196ae3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1df8afa47bf2084cdca946acb8d95e5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1534e6d7d2c8c8c35db31d7a533337a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1ece2dd206534fff1259b74024f053d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1eb32e57526ea1208acf9be6f5cc2a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hc4b7d9948fabfe1137e103fa435e62;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h7d69aa654e36e1bf920c345efc43b7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hf193709457c7ea92821c94638c8a83;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h7dc1f85abcf8857888d7bef167e47d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h85d1bce0ae836365b906957a36e27f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1b03906f783e655d93a7db3777b2b19;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h11c98b8be81e2894535c8509161a229;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1c9fc194d46a8c9dc6b2793d879219b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1a984894cc9c713392a9bb7a308c7ae;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1ff482f3b93e3bc5b1ecaf882f00ffe;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'he3ab113e8f9373fb3690f420b4f3d4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h169f60d9f923d2c58c15a123c050e1d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h6e32569f67d0b3fd77e1458e926a16;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h41dc3e5d19b8cd9e1c8bab8f4ce275;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h197f26302137c7659a31b6c4ac75e74;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h11073ac23299047e99757753647fdcb;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h16891a0f902c62440a8d36691bf1c41;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h168f1b94b87f62b8969da0fed0eeae9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hf399df75341ed928ea524dc5265ff;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1e0cf0fbf32c4825f15e2be93b620da;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hc7b5d541f50d277e7e798742abe2fd;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h11c5bbcae70ac68389c541d720964dc;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h16b01c0fea843fec08e0bcca2672eae;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1ef9606c802d4e09f84278a75654dad;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h15971297aa0a3cec864db82b7e94554;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h5302746940b0a83902c06a16ca50fb;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h16902510bf67dee6325a869a8881f61;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h791d1317a6db644ed69e16a42e83be;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h195adbe38b3ee9c9db94069244e0dc3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hae23bb3671a81289451198f6e76743;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h94b20f6b298ed2c4285bee6525627a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h12d16ae01e76836fcb0c88eb63a4d4c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h160bd5634eeb8e8298aef17e17c6149;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h19b0d355d03bd92c9fce25a712ef28f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1cfb949bd27e1719eff53f29b1f82a9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h44692184c84cf900ac55e5a0e87b28;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1b0944ec35111ccf5de334bd78b3273;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h15311631b506e73b4d996b1c8f7666;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1581285781f4c748190c34f6585fae9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'ha29ef330eaafa133c8f791342b61ca;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h143c1cc862ef17e59616c227e03bf1e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hb2de4e1efe099b5c5717e81a34dfd7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h139de26c6d78850b95561a1c50b874d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h171ff6da28f02021b87de55210f3cc2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hb146bfe970090a488ede5960359e7f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h12b3ad329c8169f04a0a085887dee5e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h17e83548e62da29ff3594ba3e3be638;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1fbe70fbc06414bcf66d7bea70ef498;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h187b76f30ba0dff871cd71cd114d0a7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1353606c4b9565422ccba738c977f2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h953a914c5a3850dfe23fa5eed0898a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'he235e8a2839dc42d1c07b2a1d52523;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'he56b7bc8fadad04466024a78d0272c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hab79ccccb2b901729c1bdf4b7908f7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1fa09a1ffbc742e1edc933dda610051;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h18bd4eee2336ae188d3de042d2c7ea3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1681c9a55ee14daf50a4c03bf84cc54;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h15382cdb3b07c3bf2afe59bf8256ff5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hf1386442a2ab7b19bbf3ff7c4d668f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h18c94756672af14ab0ba900cd8b1147;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h15d5ac143628c40c1104f3b765bef2b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1565ac56d4343970250e4ece2b68095;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h12767b9b85d6e609a878834b56e5fd0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h745c18cab55db8a7cdf7ecf024a4c6;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h27593fd714b5cefc5dba959a5acead;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h194f74929ea597d5d05b03f9536751b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h16daefe4086d201be998694be4b98cb;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hcd379eed6b63d6e1cbba23a84d3967;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h45a2f9842d162cae873e571f4b3c75;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hc4341da5d7ddaf1eab6505bf5a760f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd3ac86855163bb442783b8620d75c7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h30f4c97061b94dc03120261a37a364;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h72655f67e6d65570760e31aa1eb1b0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h263aedc29964ce47e76a7b8ac7891d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1266f281e78f0b51d427cbb571bbc98;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h12f92a76d906ea38e19775f521aa4d2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1d55d24421c9a9a04c94025e07741c0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h141d1fda11d410be2cff0ee1c5f7074;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1ce245d71c4ce4165928f3fe73d7e21;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h17eed842c27aae9ae1d638789261d98;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h79c7b629e0ecba8f22172522ca3cac;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd81025fd0c7c6f116a3d21f4e4c224;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hf7b54ab7cc564e18fb6f41e4053f2a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h118032a6409cb866bbf014317243ce2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hc8548ad397f34a33ccc458d1e4a096;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h56bcb785be2ca11c96a2bde96aa1eb;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h198eba2192e806c2289b5fd54749de5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1fefdd9d28d6996cfaf666d57f9e931;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h7c68f126121e8a522d5b23225e5a8b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h10aba5e72ab3f57354bdd37a4384b8d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h6bdb5b57447d10fb1fbd57b2c7afe3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h140cdfe9e3b1dbf2055d0f5cac00d79;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h768e75cd0f24fbe114188218ff15d7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1ce417dcea9d3ab289601faafbd5a90;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h96a813ccecefd88557191d4ab4c0c3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h112e4e28e5faf20bc34b9ef7d287747;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h11b363641f9ac5867637099a850a234;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h19478ca8dedcf00d0a96d46f643a8b7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'he39a0765bd92bc911b27f0ea8406ee;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1bfe32cd90d6d62f76522e39fbfa348;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hf4fef2eb3ae704a8bf627d14e0189;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h168d299fa4693f639f86787742cc76f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1d6ec614f06a2cc1cf2323e46d8ed75;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h172c73a141b13b4b9319aabf74e8810;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h41141fe23d49aef3c1abdf4ffc4adc;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h10aab08c737723d48bb29fa79d0c5d0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hfcbafd8eda4e8ea9d2667d5e9f6c40;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1af0dff8535f58974c4087c13da5401;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'ha10604c6f40646a60634541af9f462;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hf122a059a1e469a719cfd0133571da;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1bb9a802065a37bf3529647c167a55d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h6cfbdabafd5d7e0f6df3b0897707cb;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hdde25aaca112365ecacf742664dc7a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hdbb18adb522aeccd855398a0789e97;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1ef07ad4f895e2b30e0ace50404b2cd;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hdf28065d191fc5622de17138324dc1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1788ff270a372de8cb1caba52054b83;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hcb14ac354b367368982457b76537f5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1f49169c7ba33b2e930da4ef0210f79;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h2a55561c511116b4098649bc5efd1e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h19858117efae2ba9ab13764d472a046;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h12470b85725e063a463b1f79e239076;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h17a4ade97b6cda4ee781b37b0631b5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h10e6d6256efd6fc24accc8a9c43c18e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1deefa9c06ac63a7f968b5f0a1bfb94;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h863217e94b090cb03539d87d1a2650;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1c6260ccd1971b56ba0bf02e4d38361;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h42167e22948758fdfea5ed63b8df3e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h544c9cc9f1bb300c224e25eadd381d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1df5f0146dee3338544fe2a94c1492b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'haedd8791eb046c5ba3aa14b4954820;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1f476d4303546f8e49a0444d16cadb7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'he4adaf54d23c4e46144208b2e66a46;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1d8dd9b5ba32dfa962579d1c9c09d9c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'ha11159baac05d8df77674e5aa42f71;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1bfb608df2e2f0917dcb6a5f5870228;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h2913a7a8216916400fdef1e79b4699;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hadf1d2c50a0cfb27ca1aa359ae463c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1bcb0def677b522692d5a8b28c27df5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h7fd2c8860a073143c64c9a4a674a5f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'ha402a36892b99d82b8729f662d6aaa;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1287c410a59cce8c6a8b6bee9f557e0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hbf845067e4c41eca692547aa3ed99b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1b380aa8601fdd034f757d3ffe9aea7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1086a5a7a1caff4d2a64f8ee8aaabf3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h188041479f373a04fde7bdc689e6b73;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hbaea9963df515cba866fe2eaba5454;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h339db950a56346d5f277fb0027e6cb;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h6144a95d5f6291659a24472c110778;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h134dace887154756b1dd05b5d69b86d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h18a838d246a3bb14cb82a338988c5eb;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h183fafb52b4146a7e5d3695f3f01ffa;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h8b0d3b524500eb534feefb04c5c14d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd231add4927f840a2944d10d189fbd;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h84e200bae162344421c06973e8c005;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1def83df34930f931aff71dd39a479d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd35446d39bb749f19888e204123610;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1a9dc64c63c30176b95098303d0f03a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h179ee5f2739cf0ecc0688256c462bc1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h180711732cf18e4dbb1fcf7cfa7eb65;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h192cb8c82fa95500264ae4be943e404;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h9d5c73fdb40238fe30a623532e16b5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hfe0cc3bf481337872df315b9f3e2d5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h612c10923f37bc84af5980aa08c72a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hca7210c092c140013ba24e4582bd55;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h6c3815fb8216bfc1e913c096f5fcb0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1842e05dac0548658d0dfa3d5ff336a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1c15c1d8f0d662f8b5560c3d9e31b24;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h279d7816e502269445ed99096425ef;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h17acea696e9688357146d4953184a0e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h111cf46fa8433aa395b822db27aaec0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h16a55443231afc344f28b99abf060f8;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1749e73f327d91ae0b629e116be72a7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h168bdd1282412d925cbb9e2b2a4746e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h7d81e8fbcf29aa6ef282f5abb49884;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h189089aff8b0c98489e71dae15cd093;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1bf9e4a51eab9d6fcf84ccee78c5128;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1eb178985b10faaed3da9fceb6e9d3a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hb57d16142972d6114ca45383e079c0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h135c535096eebef015820dbdee6c6b7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h5277c17b479d7770fb716368289e86;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h79b616e2ff8dced7cb3df6af7343f9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hf7cf323bc19320dcb9f693324e8c7b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h11d9e179596d6102490f219b37dd29a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h25503cbefa2434530b62431e62fd09;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h4235e4ad92bf3931552e200a77819c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1a40e7f167dc50c80a3980e4f07552e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1474a04d91ba116a2dca4f184f4bdb4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h18bdeb1b45351c2b6c5ed11fe8199a9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1aa7cd52d257ccd7899f87f3d549709;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h145218f8c4a2a018728b4be919eed07;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h10e4cbbd2472d29586a44acd428f5e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1d3132f71deb778aac76736a9f844d4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hdaa7d97be91746e285b2eef2a06e78;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hc4fc9ae2e89cf51ac11ac5e48cc02b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hc23ea385ee4e8ec8f6ec3b5407273d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1bd5715565f415c349519e9bcba111e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h11c4478f21f117446135a5d95df8391;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h4a32c226a0ca88e1b7aaeb83364651;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h89d3f0e0c0396a2760afa1c048e0bd;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hb3169e6d3f84859c9576602fa750cb;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h22f8e4ebee7b6a4fa68521cd161f57;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h6a716b341766daded53b853a3b572f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h16db863e4f3a6295d585f460ee49d60;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h116d9fed886a40aa9362d4481ccbe6f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'ha3e03edd89d02ecba20c057ae8fed1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h167a757609291a235c635399d401477;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h6ddc71f71f072166736d7d30cc6b3e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1c1bf246325b60c1c83c91cebea3327;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h11959ebe7c531e8fe60f8d8e98a837a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h6934168989064bfa1b74689e9b7aef;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1e40f3737687623256ce90b789372e1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1e8a2714bb9f8fc687282cb3d5fe75d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h18d2a472109300e5bbedd6f494923a5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h12138218b2d86f6def2c561276430f5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1c5c5dc3469c66167add6ab8bf97e4f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h2bedbd8c254e4a482aad4d72e6a984;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h66fd2427fd99b584592ee17c821118;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h75a0fe21bd4dd882ddd019e3d0e17a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h13b05482e0926c81db7e8e839c2a308;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h9594357f240a9bdd48b250ea2634ec;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h12f56380e159da32db26823a07b2b02;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h187edca62e00d0855e3e4530a39b7e4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'he38566fc60a95deb96e7610f442369;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h18982d6e13ed12507e02f7512ed9a2a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h17f2b595baaa92cb53c52a7875a1583;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h159efd30e6036d50eb596e74f8fcb6f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1341484addc6f18193725ddc44e770f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1dd8cfdd24736f899c5f6f56f5b948e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd5d5a74152e434d8b929388d7d9717;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd2358116ce5130284677deefa64a49;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h2e253289c148ac66b536987fab0844;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h11c9f60e5d78d88a3d2d75e3b6efd9f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hf6c82932663c922315f0a681cb2ad6;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h15ed4e4827fe15f97224754c48f759;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'ha8629cc88fdfd7618560527e4fa624;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h21732d28279099ffc469066575679a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h13b21cab2f782d371d500fde14c21e9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h524797a169f9428e60f11ac082c625;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h106eefc3dfa89844502a5cfc274da12;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h112a0d972719c5056794d54da119e6f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hcb0121ea9bb2c046e48f4a788b6a3a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hc05c3f2f3e7f56af3592aed1ebe818;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hb8e8baa5560e994d44ecec5d5f4e06;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h167a8667729f8b0a1b1506fd75f19f2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h16f8dc0cf48408c2ff2eca6e025f4b5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h2a7dd7aadcbcd31c5dac522965913e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h42850cf3d2e294337f9aec0a2d0a36;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1561d1f8ebfff81a37799d89733aad;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h9a13876c7c7ed86fdc2f17537540df;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hcaf55c734ebf418c42c58b726c97c1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1027bed7afef9ad2ba4ffb9be0f6f1f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1952d771daa11907ecc641dddce7926;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1cf49db6a1008c7b40909e0c258e7f8;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h624bdca93520f19067cda9d8e01e26;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h720326c7d2acd21dd88def55ce0a78;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h79bf5e38f6268cfd920d6f530a767b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h13bd60e39ea7612be5478bcf8880cbf;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1a778f6707db66b57189de51ccfa88;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h56690c1530ac1a6b329b8582fd6732;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h117b21c707c8ec32ea0db86046ad539;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h19d854f3b75854dd5d139edde71371d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h51c9c5c6755f88b515e2a2904935dc;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1946d80961694f8522e3daabb805877;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h19198b49ba73935aa5a6af1ade29d62;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h19d923d3f56597976eb542bf75b600b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h7fb96da24c5b54128ef1aa6fe6e800;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h3f2a06a22c16a3f6b21b98ee1fe64f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h7e25a37cc5ad4c79e920d0432f09cc;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1d4596282838eb52d62528dae8ba58f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1b69fe2c42b9106e27ce3d7c9c03265;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h3fe08e16cbf8afa8e9ac1ad41c8561;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h125b20f2a15841e62468f51ac796fa3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1ea352259af97ae57dcc14d56946d7c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h8ab27afaa67dcb9dcf4b426568fd08;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1e09370af04750cbaaa7a5c985e5081;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hb5be44b1cf3c310e513cfa12e77589;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1bec40b5c0074787e3fdda7c879df37;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h14f3d18c64c144c16aa778a82416c84;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1d2711eb1301e9b2248cbc1de2532a4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h959bfcaa942f2d06d542c06422a652;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h2eba05f37e6c37087617275d392cd0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h17f3bc32c311d4fec11ac9a78400ac2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h38ebb1d57c75ed6155b573bbdd06be;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h125da9a8e9557c713e1bf8593b36371;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h98e8728e6aec7dbf95323286fe99ac;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h133e44a1bf20ef098bd9857f22be6c0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h5e215051d669a302bbc0ca017051f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd8162d962bc63c7c912349e77e8817;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h48ba2bf136de919d08116d37b6aaba;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hcb54e666c60a1d21dad0d54becd277;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1cd6e087fc9a782094c8505ce402cbd;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h18e3b5f506c900f72c4733afded2571;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h2309bac3a7bedd6e0bd1592f741ff;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd0770964f3bfc49ba8580b605e368a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h15641efa7f6cc8683ed1bf8c3cd5113;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hec917c12c5f0e39f784dd7a90dbd61;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h18286374544a0656c8124d3e5fdae9f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h163b6784c24dec05363b2c98569841b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h3643744da0d2d64470ee5dde0406bd;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1a481c89bb71f42f12291a88f3722be;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hcdba95a1e6818ce1cca5847e99ebad;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1b45177cc17f9d5cb51868a9b154aad;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h157ff8686a921c74b71cd30358f0e91;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1d57aa646800df285e20d60e21b5d72;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1be008b7d23ff28d535d0c7e0fd8f54;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h10370a8761098a2c183ce01878b1763;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'ha9aaddd51985dc744f2b87c1a96d57;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'he98769b4b7ea5f5c7d57909fff1453;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1665eb1acc82952c5e48ab5682d3234;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hf22282e030b9448a3dcbb181820908;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1901661f291b579921be89331c7eac3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h15c6ec6d162764fdd278bb5d936bc7a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h4daf675a9d8cb94c57a28046cf6911;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h120bfba5e2641393768bfdeba640f4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1a06587dfc2c3ca33b967c4c55b1201;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h13c9f20bda0fad3806c460e40556974;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1b5c117cc91ac2b61118e630b067e1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h8ecbc8a8273774eb0431e938045b1f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h12c32db96bd2d938d74fc202b1940e9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hce36e3eec1096c225c12065b0356b4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h18348b32fa96e537ef61aad892b500;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1b833e4c342aa983ef518488f5adb07;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h136e50d3f52ad4fa960577981d80e5c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1daff815102951c931f940f7a1eb738;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h731bd1fd95eeb2d1630c7e57d03d45;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h4b086e38389b05445b521f8e75de84;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h895a2d1abb52dfba4918111284da81;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h36033a5ac1af6b141d84deae577d88;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1be8c97fc9e7d4b9f165ab686b8999e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h500be5515648390afa56cf8552fd61;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'ha629de1592b0ed3d79b9597fafe277;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h82b6b97d0173de9a594abdbc4345ee;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1dd9ed9bdcb9bdafb056c1b54a90d16;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1b720e5de55a05a52a1a432e846cb1e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h85f9e6c894d25f351a626a525f1989;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h908269ada220d105ece63585177fe1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1d9ae5f378fe89df63abbd5c0df9805;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hc2899ba842b5b7eeeb60235718360f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h15571d140c3619953c125f5d157fae2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h179f25102976142586536a8d90c865e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h18261f3ca647c8f0073035058cdfb14;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd99cf980a3369299d52d71b0689f7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'he27375d78c386cfb8d649d214a6800;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h12a3ff8f348d248aecd5b0e2b59fb58;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h11d2c56283ac567f2a45ec5ba01f32b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h9b01bbc28ac117a70644fb3dfe93da;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h16ed9342a28ae0c9a5b9fff9d3b6bf5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1a47a5416476a93700993b42d24de55;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h475d89c7c08b85bfa073d4c29e96ab;
        #1
        $finish();
    end
endmodule
