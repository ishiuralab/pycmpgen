module testbench();
    reg [0:0] src0;
    reg [1:0] src1;
    reg [2:0] src2;
    reg [3:0] src3;
    reg [4:0] src4;
    reg [5:0] src5;
    reg [6:0] src6;
    reg [7:0] src7;
    reg [8:0] src8;
    reg [9:0] src9;
    reg [10:0] src10;
    reg [11:0] src11;
    reg [12:0] src12;
    reg [13:0] src13;
    reg [14:0] src14;
    reg [15:0] src15;
    reg [16:0] src16;
    reg [17:0] src17;
    reg [18:0] src18;
    reg [19:0] src19;
    reg [20:0] src20;
    reg [21:0] src21;
    reg [22:0] src22;
    reg [23:0] src23;
    reg [24:0] src24;
    reg [25:0] src25;
    reg [26:0] src26;
    reg [27:0] src27;
    reg [28:0] src28;
    reg [27:0] src29;
    reg [26:0] src30;
    reg [25:0] src31;
    reg [24:0] src32;
    reg [23:0] src33;
    reg [22:0] src34;
    reg [21:0] src35;
    reg [20:0] src36;
    reg [19:0] src37;
    reg [18:0] src38;
    reg [17:0] src39;
    reg [16:0] src40;
    reg [15:0] src41;
    reg [14:0] src42;
    reg [13:0] src43;
    reg [12:0] src44;
    reg [11:0] src45;
    reg [10:0] src46;
    reg [9:0] src47;
    reg [8:0] src48;
    reg [7:0] src49;
    reg [6:0] src50;
    reg [5:0] src51;
    reg [4:0] src52;
    reg [3:0] src53;
    reg [2:0] src54;
    reg [1:0] src55;
    reg [0:0] src56;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [0:0] dst26;
    wire [0:0] dst27;
    wire [0:0] dst28;
    wire [0:0] dst29;
    wire [0:0] dst30;
    wire [0:0] dst31;
    wire [0:0] dst32;
    wire [0:0] dst33;
    wire [0:0] dst34;
    wire [0:0] dst35;
    wire [0:0] dst36;
    wire [0:0] dst37;
    wire [0:0] dst38;
    wire [0:0] dst39;
    wire [0:0] dst40;
    wire [0:0] dst41;
    wire [0:0] dst42;
    wire [0:0] dst43;
    wire [0:0] dst44;
    wire [0:0] dst45;
    wire [0:0] dst46;
    wire [0:0] dst47;
    wire [0:0] dst48;
    wire [0:0] dst49;
    wire [0:0] dst50;
    wire [0:0] dst51;
    wire [0:0] dst52;
    wire [0:0] dst53;
    wire [0:0] dst54;
    wire [0:0] dst55;
    wire [0:0] dst56;
    wire [0:0] dst57;
    wire [57:0] srcsum;
    wire [57:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .src31(src31),
        .src32(src32),
        .src33(src33),
        .src34(src34),
        .src35(src35),
        .src36(src36),
        .src37(src37),
        .src38(src38),
        .src39(src39),
        .src40(src40),
        .src41(src41),
        .src42(src42),
        .src43(src43),
        .src44(src44),
        .src45(src45),
        .src46(src46),
        .src47(src47),
        .src48(src48),
        .src49(src49),
        .src50(src50),
        .src51(src51),
        .src52(src52),
        .src53(src53),
        .src54(src54),
        .src55(src55),
        .src56(src56),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25),
        .dst26(dst26),
        .dst27(dst27),
        .dst28(dst28),
        .dst29(dst29),
        .dst30(dst30),
        .dst31(dst31),
        .dst32(dst32),
        .dst33(dst33),
        .dst34(dst34),
        .dst35(dst35),
        .dst36(dst36),
        .dst37(dst37),
        .dst38(dst38),
        .dst39(dst39),
        .dst40(dst40),
        .dst41(dst41),
        .dst42(dst42),
        .dst43(dst43),
        .dst44(dst44),
        .dst45(dst45),
        .dst46(dst46),
        .dst47(dst47),
        .dst48(dst48),
        .dst49(dst49),
        .dst50(dst50),
        .dst51(dst51),
        .dst52(dst52),
        .dst53(dst53),
        .dst54(dst54),
        .dst55(dst55),
        .dst56(dst56),
        .dst57(dst57));
    assign srcsum = ((src0[0])<<0) + ((src1[0] + src1[1])<<1) + ((src2[0] + src2[1] + src2[2])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15] + src18[16] + src18[17] + src18[18])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13] + src19[14] + src19[15] + src19[16] + src19[17] + src19[18] + src19[19])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6] + src20[7] + src20[8] + src20[9] + src20[10] + src20[11] + src20[12] + src20[13] + src20[14] + src20[15] + src20[16] + src20[17] + src20[18] + src20[19] + src20[20])<<20) + ((src21[0] + src21[1] + src21[2] + src21[3] + src21[4] + src21[5] + src21[6] + src21[7] + src21[8] + src21[9] + src21[10] + src21[11] + src21[12] + src21[13] + src21[14] + src21[15] + src21[16] + src21[17] + src21[18] + src21[19] + src21[20] + src21[21])<<21) + ((src22[0] + src22[1] + src22[2] + src22[3] + src22[4] + src22[5] + src22[6] + src22[7] + src22[8] + src22[9] + src22[10] + src22[11] + src22[12] + src22[13] + src22[14] + src22[15] + src22[16] + src22[17] + src22[18] + src22[19] + src22[20] + src22[21] + src22[22])<<22) + ((src23[0] + src23[1] + src23[2] + src23[3] + src23[4] + src23[5] + src23[6] + src23[7] + src23[8] + src23[9] + src23[10] + src23[11] + src23[12] + src23[13] + src23[14] + src23[15] + src23[16] + src23[17] + src23[18] + src23[19] + src23[20] + src23[21] + src23[22] + src23[23])<<23) + ((src24[0] + src24[1] + src24[2] + src24[3] + src24[4] + src24[5] + src24[6] + src24[7] + src24[8] + src24[9] + src24[10] + src24[11] + src24[12] + src24[13] + src24[14] + src24[15] + src24[16] + src24[17] + src24[18] + src24[19] + src24[20] + src24[21] + src24[22] + src24[23] + src24[24])<<24) + ((src25[0] + src25[1] + src25[2] + src25[3] + src25[4] + src25[5] + src25[6] + src25[7] + src25[8] + src25[9] + src25[10] + src25[11] + src25[12] + src25[13] + src25[14] + src25[15] + src25[16] + src25[17] + src25[18] + src25[19] + src25[20] + src25[21] + src25[22] + src25[23] + src25[24] + src25[25])<<25) + ((src26[0] + src26[1] + src26[2] + src26[3] + src26[4] + src26[5] + src26[6] + src26[7] + src26[8] + src26[9] + src26[10] + src26[11] + src26[12] + src26[13] + src26[14] + src26[15] + src26[16] + src26[17] + src26[18] + src26[19] + src26[20] + src26[21] + src26[22] + src26[23] + src26[24] + src26[25] + src26[26])<<26) + ((src27[0] + src27[1] + src27[2] + src27[3] + src27[4] + src27[5] + src27[6] + src27[7] + src27[8] + src27[9] + src27[10] + src27[11] + src27[12] + src27[13] + src27[14] + src27[15] + src27[16] + src27[17] + src27[18] + src27[19] + src27[20] + src27[21] + src27[22] + src27[23] + src27[24] + src27[25] + src27[26] + src27[27])<<27) + ((src28[0] + src28[1] + src28[2] + src28[3] + src28[4] + src28[5] + src28[6] + src28[7] + src28[8] + src28[9] + src28[10] + src28[11] + src28[12] + src28[13] + src28[14] + src28[15] + src28[16] + src28[17] + src28[18] + src28[19] + src28[20] + src28[21] + src28[22] + src28[23] + src28[24] + src28[25] + src28[26] + src28[27] + src28[28])<<28) + ((src29[0] + src29[1] + src29[2] + src29[3] + src29[4] + src29[5] + src29[6] + src29[7] + src29[8] + src29[9] + src29[10] + src29[11] + src29[12] + src29[13] + src29[14] + src29[15] + src29[16] + src29[17] + src29[18] + src29[19] + src29[20] + src29[21] + src29[22] + src29[23] + src29[24] + src29[25] + src29[26] + src29[27])<<29) + ((src30[0] + src30[1] + src30[2] + src30[3] + src30[4] + src30[5] + src30[6] + src30[7] + src30[8] + src30[9] + src30[10] + src30[11] + src30[12] + src30[13] + src30[14] + src30[15] + src30[16] + src30[17] + src30[18] + src30[19] + src30[20] + src30[21] + src30[22] + src30[23] + src30[24] + src30[25] + src30[26])<<30) + ((src31[0] + src31[1] + src31[2] + src31[3] + src31[4] + src31[5] + src31[6] + src31[7] + src31[8] + src31[9] + src31[10] + src31[11] + src31[12] + src31[13] + src31[14] + src31[15] + src31[16] + src31[17] + src31[18] + src31[19] + src31[20] + src31[21] + src31[22] + src31[23] + src31[24] + src31[25])<<31) + ((src32[0] + src32[1] + src32[2] + src32[3] + src32[4] + src32[5] + src32[6] + src32[7] + src32[8] + src32[9] + src32[10] + src32[11] + src32[12] + src32[13] + src32[14] + src32[15] + src32[16] + src32[17] + src32[18] + src32[19] + src32[20] + src32[21] + src32[22] + src32[23] + src32[24])<<32) + ((src33[0] + src33[1] + src33[2] + src33[3] + src33[4] + src33[5] + src33[6] + src33[7] + src33[8] + src33[9] + src33[10] + src33[11] + src33[12] + src33[13] + src33[14] + src33[15] + src33[16] + src33[17] + src33[18] + src33[19] + src33[20] + src33[21] + src33[22] + src33[23])<<33) + ((src34[0] + src34[1] + src34[2] + src34[3] + src34[4] + src34[5] + src34[6] + src34[7] + src34[8] + src34[9] + src34[10] + src34[11] + src34[12] + src34[13] + src34[14] + src34[15] + src34[16] + src34[17] + src34[18] + src34[19] + src34[20] + src34[21] + src34[22])<<34) + ((src35[0] + src35[1] + src35[2] + src35[3] + src35[4] + src35[5] + src35[6] + src35[7] + src35[8] + src35[9] + src35[10] + src35[11] + src35[12] + src35[13] + src35[14] + src35[15] + src35[16] + src35[17] + src35[18] + src35[19] + src35[20] + src35[21])<<35) + ((src36[0] + src36[1] + src36[2] + src36[3] + src36[4] + src36[5] + src36[6] + src36[7] + src36[8] + src36[9] + src36[10] + src36[11] + src36[12] + src36[13] + src36[14] + src36[15] + src36[16] + src36[17] + src36[18] + src36[19] + src36[20])<<36) + ((src37[0] + src37[1] + src37[2] + src37[3] + src37[4] + src37[5] + src37[6] + src37[7] + src37[8] + src37[9] + src37[10] + src37[11] + src37[12] + src37[13] + src37[14] + src37[15] + src37[16] + src37[17] + src37[18] + src37[19])<<37) + ((src38[0] + src38[1] + src38[2] + src38[3] + src38[4] + src38[5] + src38[6] + src38[7] + src38[8] + src38[9] + src38[10] + src38[11] + src38[12] + src38[13] + src38[14] + src38[15] + src38[16] + src38[17] + src38[18])<<38) + ((src39[0] + src39[1] + src39[2] + src39[3] + src39[4] + src39[5] + src39[6] + src39[7] + src39[8] + src39[9] + src39[10] + src39[11] + src39[12] + src39[13] + src39[14] + src39[15] + src39[16] + src39[17])<<39) + ((src40[0] + src40[1] + src40[2] + src40[3] + src40[4] + src40[5] + src40[6] + src40[7] + src40[8] + src40[9] + src40[10] + src40[11] + src40[12] + src40[13] + src40[14] + src40[15] + src40[16])<<40) + ((src41[0] + src41[1] + src41[2] + src41[3] + src41[4] + src41[5] + src41[6] + src41[7] + src41[8] + src41[9] + src41[10] + src41[11] + src41[12] + src41[13] + src41[14] + src41[15])<<41) + ((src42[0] + src42[1] + src42[2] + src42[3] + src42[4] + src42[5] + src42[6] + src42[7] + src42[8] + src42[9] + src42[10] + src42[11] + src42[12] + src42[13] + src42[14])<<42) + ((src43[0] + src43[1] + src43[2] + src43[3] + src43[4] + src43[5] + src43[6] + src43[7] + src43[8] + src43[9] + src43[10] + src43[11] + src43[12] + src43[13])<<43) + ((src44[0] + src44[1] + src44[2] + src44[3] + src44[4] + src44[5] + src44[6] + src44[7] + src44[8] + src44[9] + src44[10] + src44[11] + src44[12])<<44) + ((src45[0] + src45[1] + src45[2] + src45[3] + src45[4] + src45[5] + src45[6] + src45[7] + src45[8] + src45[9] + src45[10] + src45[11])<<45) + ((src46[0] + src46[1] + src46[2] + src46[3] + src46[4] + src46[5] + src46[6] + src46[7] + src46[8] + src46[9] + src46[10])<<46) + ((src47[0] + src47[1] + src47[2] + src47[3] + src47[4] + src47[5] + src47[6] + src47[7] + src47[8] + src47[9])<<47) + ((src48[0] + src48[1] + src48[2] + src48[3] + src48[4] + src48[5] + src48[6] + src48[7] + src48[8])<<48) + ((src49[0] + src49[1] + src49[2] + src49[3] + src49[4] + src49[5] + src49[6] + src49[7])<<49) + ((src50[0] + src50[1] + src50[2] + src50[3] + src50[4] + src50[5] + src50[6])<<50) + ((src51[0] + src51[1] + src51[2] + src51[3] + src51[4] + src51[5])<<51) + ((src52[0] + src52[1] + src52[2] + src52[3] + src52[4])<<52) + ((src53[0] + src53[1] + src53[2] + src53[3])<<53) + ((src54[0] + src54[1] + src54[2])<<54) + ((src55[0] + src55[1])<<55) + ((src56[0])<<56);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25) + ((dst26[0])<<26) + ((dst27[0])<<27) + ((dst28[0])<<28) + ((dst29[0])<<29) + ((dst30[0])<<30) + ((dst31[0])<<31) + ((dst32[0])<<32) + ((dst33[0])<<33) + ((dst34[0])<<34) + ((dst35[0])<<35) + ((dst36[0])<<36) + ((dst37[0])<<37) + ((dst38[0])<<38) + ((dst39[0])<<39) + ((dst40[0])<<40) + ((dst41[0])<<41) + ((dst42[0])<<42) + ((dst43[0])<<43) + ((dst44[0])<<44) + ((dst45[0])<<45) + ((dst46[0])<<46) + ((dst47[0])<<47) + ((dst48[0])<<48) + ((dst49[0])<<49) + ((dst50[0])<<50) + ((dst51[0])<<51) + ((dst52[0])<<52) + ((dst53[0])<<53) + ((dst54[0])<<54) + ((dst55[0])<<55) + ((dst56[0])<<56) + ((dst57[0])<<57);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h0;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h733c9254faa86d4e0b4e58a678e753711d3bbb05c183b58133612ce4ed68045916ad962200f99d7b2ad839f452a1ff48792181f5c7da6942d58e50bde9b16b817840763d07e1b15d76cd5c4917160a451255a36dadab1b3d0b233587bb24e8af99be41edea8be68784;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hee099d4a77c1ddd56671dd222bce2ce1b949b82ea68c32f8fda45509a47ad4234743b1a9206773b7cc3b7428e12cd960962e6ce04b2466b0b0469c29ae9b3436346c77a422b17d99d933b4436bdfe5b56b79ca19924caffbf0d91e54134c5d7e953ca2a1f0d2f9982;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1bcc60a3c0e3d76a165defddd1577798e1eeb9f2000176fd57192b885b84c261d91e6de35454f95b3ac9e752498ad8be0192ef637b882dbe34f315f60107d8086dfcfc3eab45e1a9ea5e735a8a8c13e9afdca3bf426c0e67134ce0ce405bdca44a87b3197dc76656f3;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h39dac6c4adfb2bfe7c9aeda9868b139b90754c0a58401f9d884ceeb3a5211af94023c2fd5bc08d8b8d279161af53ed6a93cf1ae9f42ddf8daa9978abc12a211096cd5ab5d71481422347e2d2d8018dc044539116daad9772c6e5f27436d31362818d3e17ce8fc2144;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1989f6b5bf674817fc12fa736da353f070093579369fcf9f91d7b9ae1082b83aac00a47aef9534849288b25c1619c7a5771e83ade257334c58b51765a0005e0e9c6145852e2514f68876611c43eb95f2bf3528a373ec2975e446dbbce89ca17f95c74827163c5b3bbd5;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1830eef03227b9d42e5661ae952ff8ac479318cb6d32c14a6510ffb85df321859f4587cf7c17c98f67f4f7b2bf884dcf252efc5c0bad01eac5b4d3e8701fe2e382b3ff5961e9e0e93a1a6ddfbe57b3370bb46308dc370daf09f0e887d2f1d2aa7e574a5c27869c04082;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h163d452850a5366549128682896333a6771a8afd6f2e9af3cbabe5db573679596e2604bfbabb77b0a9a08ebead89c7fbe762020d1c40cb2fb052085b70b4724375bb05ad5248ec77d7cb4cc678c79751f01f0e22a5845ba81ea638fdf2cadb95246a3ed98921f4cb628;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h4b80786f013321c30f139dd6981694ba65ef6094ed5fdf2c0441b276d5cec02877e73a987e8b86d578e4dac7c229b810ba5adbc63b33a27884c994dc885382a7ddd0b480204d86af75617bb7c10cdb2aeb2da2a5ce36175b0ed1c536b95924001d443ab0621d2c6fe7;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c63d17075eca2fcb258616304e70de27e19432aa0d010822e61771735956e98a896febe14a851785ba942ac06dd756c866ad897ae700b01305cd0c3265feab034263d03393785812b67805c616006b59b025a20fbdfa3974a2c95f4c0216c88812e3126f0785bd4b29;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he5d53518f5fb2ca170496851efded5863c1b0fa9d5f7773bad4fccf96b06bc3b4e4fa8dbeb8257464b20ea3b9b304c80b2577bf4ac78883439ddc516a0fc26434055087c812a8c084917ed26446a0c962b26605673ef9bdc619c761581f7affc0e671c82ef187fe7d4;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h159ae1564ac709bc13040fe924bf913b01f1f98c4a79b372fd1da54729fe73ab5db012fe07fa57db5cc01bad05a030e5236e024b6eebedac00c83623476921c144630f0a527ec4bf441bb330108c99babae14685718877c46f06d096c66a2736ccfda359b91be661477;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h18e71d5dce45dccd326d1ebaa8f19e388c356eb6533f9529f71eb8673cd627e9a13a58b43cf76734e714d39700f4a06f27bb4c32c3af09ca92383b07a8450c52db02943eb69f50d18fa4c7b96f03afd47a675a61a202617ddb7eae6301331a5fcacb1d7f3ce757210f6;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h948b90fcfcad0699076435330463d21d6532336109f76ec46d6a2a670404d267debe4e850c89d8106ec55bc0498eb896feac855d12698cb1e62159131ffa2d85005ba333d33b11266b11eb6dda1cf2e64cd350f4a721a3a4143fba519f67a7a92402a06093c9dfac6e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h13f2cd23a65d90e03bb2c89c8c8d3cbcd4f877ccd9b2fb12eeef043a89e5a32f7274d012faa78344d956534b39206a42b0a75e018b19aedff03c4aac59c96eb039cae6c5dab351c1c4381ac7ef91fdf6e36a3127122d606128297c1fd70ac4778fa19059f7d5f14242c;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he7ba038e2cb56017589de47e1d7d76c022cd1205f26f916aef7aca1fd5546ebdeb989ef37219945590501efcb49077bb53ffd8bc82ba1d0f0d886f4f0f79f6ffebc07b9ffb423264e5230feaf1c7b3fa1cc3032ce5037562482447e5680a7c242b1270d9d3f883152e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h14a3f1fa91beb0e3aa957970a6c3d708ca275c35f9e4cff7cd47e2db0db2e6fe414f2f6b09d858f245793b451ea13f4ced01f253812a49e5e891ec7a06692a80df9c89855ef58cd41dea995d7f6d9ecc6342a7822908c6373931820d9ea7623552dc5159974e05b1393;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h14f95e301d42be16109be3b2ae6ba109b0477c5386257c94e9e40e27483f2a4a3178cba2115dc5e64923a1b78accabf6423fe016ef9118739fcb1ab9f9d39a90012838c712de3b4cd9f355f81eff01d95a2987a6ff32f96f9e2f0e6e2fb5df1c9b335be742599b00bb7;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h840946054ef5be13a1c806ae4bd4d34e3f6bdace6b89c76a544959457c802b0978d4a3c7cb102c989fe32f8f014be73f753f283b56e6267d2e4a5dfe5a2b4be9680ae77b45e76f161bfe63355e06f287713fa6f66ca00f676843695d28549fa6ed96494b3e3f4d51f7;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc03753f6cef6a0410b1dae808db0f3ac4268390deec3bf3156daa9a0a36cb9176c7b7a85c61a147ab83467a290c22da5f410063fbd1b9a4d62d7e4a414e9c627b7795d1bae0f10af43df2786bf3e7341ff728f77fd38c5a5ba3f861b2bc5bb3cf1d7fd24e345f8a9a9;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f359cb3eb4fcebf81e31493c45681c738d9db70d3261200379e150c36b4e9df2d590174aa9ce19f630a6a9536d0a4a2fafbc70a7483dd427f7eccf15eed1ba5cdc724bc0988d3f5284457847ce4e4f5052dedd74cef721834e3e030967d4f0cdb197bac6add1bd73;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a80ef7126ee8a2bc15a453a0aadd2ab8a6be485706dfaadb353276ae45097c7d0db012d8cc6702a4f65d470c36382308deafa4623610669a014483193d32110d7f28cde9e333c64384c71c81031c943bec4afc0696662958ad9d1fb7bd1c26dc4ea3b4929054ce324;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h16a1fc03be5105099bd6f86fcf3a65e1d1b5fa89c9d564daba9379d2a679965aa0a383c7d59409737e637a17176f2302dfb47c9e8a99eb265765fcd59d91ca81b1d8bac90fbe15779d52f69401de2af7e3fded09b542f8b08c7b94100cff6f81a193bc3587f32ce85dd;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h116ec47e30fddcb9fd7474e1352a767cff039347869ee58240083afc48014bd96f0de2e2e529ae4db405e318e481502dbd2279cc3082db995ed71406f5391546c895b710b246ef7dbfaed55407b1f04dde864acfc5958428140e603e94e28e6b7454ccd1ab18db0a58d;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d218829b09c328df96eb3b69e46da7ebfacedf48efe70dd00be1dc000fed0628083889dca1a1dfd79d11fbcafce98b36a607eb70e390f01fd77bd6d7962f2d3d1823b63424bf961f89859d6f168c0e8db640601418333beaccba6e5fb6f902caabddda01580a615258;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h7dac9805b72183d4f599d1f3d988b0b0649398582ddc8236f7a5d3921b29e7733eb03cc6f466a0bc534f73a948358e8e46386ee50c01090461d8bfbbfe61a5538419c25202a0891b5e88b452d41e96de032eae6bb8c2320b5e27c40af1cd9bd844f1abc7be73425821;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha68a074bbae79094043be176a28d01f8fe069ba6cf3559c96ae780c7d718b9bff428fdbaf93e527efd90b13bd3ce2c03117f390c9d16c3fe26747ef5076bc7940cea4d5685419f6f88f95f2c6de2f180b79a7900d572f3352165e2bcade645279e5ef075133f4bf93e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h7eb3eb87da0c5f0ece6f5266c543576eda54e82495494fb29a678a13060eaa0c3e07427629937c5f8aa71c7764ffe2ca3a80466ee70bfb1e3708060a52cc2e9deba040f92561a4f7e0a07f838b6f54a10a44ab97dc9cb5ccf7e62a1b6326fc3f680f57ee944c565ab3;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h18c27852111a70a68b68d37b23c04b85d05f19549a87bd9d06877900063816eda1219677b2f4bf97967f7a57561216cc8a5a8311e3c9cc87d5d4aba8d5ba94bd695ae449ccf3154ed1708391508cc31a8e9d866574cac6d4cd6ad1b37750f3b4493ef585f8de2e3e95e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb74ea616eebeafbe3a037683ac5fbab2a88489e6c01957b1665864a1c986496fb1b077255d83bc8d2b5319025e17bf04ffae990a4ac1ec8e97437db16ba99da7e8c0ab63ce18b8a162a889dcf16986ac71cd9131ee1f0b79e2cd897432125f3c15d347695c4ee35852;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h64c1eaad5e0f7a72a4f955c1cec3f18f3aa01a392636de8f9f2d2c7bf4d67d649aed284cc79493d0cef4b03fcfae1b84ebb3e64340c8027fdf80087f1785a1516da2155f944ef244ad5bebc281a6d20dd2ede4a715ef98b928aba408d5487b6fa1808185f453a18d4d;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1acc01a8bc45708bd0c9e6d0eb86720635dc34115b06e525c52a0164f7d7a8681509e4e91a52deaa98e26a088d895cc6bb2cbfa6c06c280eafb7b42361b3b3a061242e5c703d256c6a1ca6cd3178391e37a9fe9a7bb025639dea8d852c8697689d9b40bfd8751ff0889;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h187ce87100bdbedcf7b7f2761ebb7aa7167798df2838119e3229d2c37b3285682ba639f3a50bf3323705491d4b79882eef3b7de152270264afee4dbe2b569f22fca168cc75c942adda55094dd8ecebed4c83f118567e1b77473177b77c53b70ef7d10008a5234feffa2;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc701304e193a08859437e53234456685222e3ec4e413042c3ae610aee7bcd8c765b14bc29f96837d42a8f864dc3f7a817476eaf888a3f8654ca9ea9e03aeb0cc3bab49cdfe55a46ebf8ad3a85555e63e911c44980463d22d1ee314e883b6f106e59352cdbf054489d9;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b2ea129344d8e2f64088ddf5809362703469228705eb10aec882a10db3615ed9ce16433ba9bff491574fd429ce69ef89b5ceb160b0e1d77243c4e668c5a69a36f73a704b1abf9e7cce77d6a2628b44ca5afac79b986ff47a7e4c38ee90f98548dde2355d0d9ad7ee39;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h11b5f7c32b79ecdd5e96221001e2d1f9bca5a2506e33e1fead5f9e19a7c7471481a9802cf4b5b05c5a7bb1081091348f74d0d387475f506fff4d5fd466854d65c9345203c4afd2594a3dfad58e869e0ed374fb2d18b7ecd853b596af88abc111e2c8a6d4b694e07d50d;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h170b5c985f56e190148303c889158692a8549a0246b6f666287c7860cff408fe3293925a98d4aefea3a25cb82295d947403f96c520dd1923e4a8ee11783d5c87f8a7e6b1f119c5a0c4b098208521de83dbb501540ebd9f3b4315110ebcc661090ff297ce6016f8b8cd;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h23bf6c3efda55803c49ca3be3bdc26d31f4239b97417cc3744ab89bbc8efda55d768402141463d2f725e9950b473938bbc3e8f720d119cd2a308cd9deb6bc39ba72568fcb1c09be91f96e80113066a6979cfcfcd63230e282ce1b84395845421c5b6aaef491e364cf6;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h3a59c624296781059f975a71bcc873c7e6c095f0e57c36031b09d9b6d8d62f623775f2f91f61026096fa672e158f401f0e3e1f7760486cb7e6249c25e6f048fcf73cc91236487d4495329ab36bcd7a7b86ea1554ab63cf0aecc70e9ea3011c3f768baab732366a21dc;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h7f5affd04a95c32e328becf45c479357fd04486326a7227d4486938418d0fdeabe7ef5a40877a17b8a2421aa38e719ca5d86042b0b56559250020900b832a7d47e4505730c9dd3e31de2db4faa0d84ba55c201c2c0f39eacaacdba34f0b848aac7f96313337a5860ec;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h180ee81deb1c1c93a4a52fea565d44a39c53e1f61e8b2df711b5e49f84f35c2bcda9ffde2777f2e4779a1b38ced32738e9a57c324adc3437caf667532e1546edb3440d559bebb210310471c434f6085e6a26a0bb1953ad2468f3a5117e9c26f72efb1fa441afe3f16d9;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h12e52e823d8bcb20f68d2e5a4bf7b0141ec4ca48991b6513e0e8f0f8e964813de3ee8a62436628404238e79d5622a2d0f8ebb84863a41f2ddfcdcb115a65d8b270cfdeee065ee654ce1e75277be6fbae1d1e4530f9877c544113c95fda312b53cac6d8736166a1c2ed;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ffdd4d47f603f8c166d35245c87ae59c5cdbc3d4a49d34fc9ea833c42633e0e8f98174c82299e048b298b7d2c1cfce24b0a192af569483f3aa84a92283dc00ca01faee2eb32ef4de05a435a89c9599c6d1599f684d3fe0a86b4a59c58976b193f6d8a295a6616820e5;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a158a89ce0cba89e8d5b36baf8bcb608493589ba6d85b41e886522736e86d1399cfbc8a728971d5d49b23a0539b119b56e1031034611637e1d9937d9fb3814ab2eb5b6d9ba1dd35c4ac73a70741c24b2f2408baafba5f55c1304dd07e82f5ddccf7185a44f9ee6ecc4;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ff27d17d171e5eb649dd21057d619d558e276c46e98e94e68eb9530c25ca1e0bd5bc9f45b9663116a95d67b43bd69dd38b78f12a03815c4e0bf2f3057b43601aaabf821f679cb71edb261166fb6447554abdd9e20886f5efdac693fcd89c9107290daf70a1df1468f6;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1867bd2e203e9c7ce8913bc2970ce6236818ab4433f3e01d3af1cb1ea7fd0164d8f1ddcdb7bffe66246d9e9e9d3e571e3e11f5b3fbf76c12f113192f0d10ea5ef7a1a3c578414590aed66c1f84819cf31bf160d1e75105003b41f0779b6920dc88cdf42060e5eaba6af;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f9a43a7442247a15f015ae2c9e74f38200b11ee2c4fd8ee62cbc12834d4ae756c7b290090c7ea5cca28832f60942b661ea716f736bae60de219abfa1d616f6d6967a70a7c6d3cfadd77d0429a035e24a5b06af17002da3237bf9298168bdb5a287be829bd63f8cbd21;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b2f8365752e8772d8bb146fb1bdec781e7b73f8c397b997691be7fbb60d797c6423470d5932c6d120712b1bb4daaab61684e96fbb012e3b8a0c2ebc144fcae68b8e0637d8f9d67a78f18c8a40679d830a59fbc2494ccaa38a776af0e3cb40c6c56f7fd9294ed36fbce;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1499bcbceacd2f0d6546a287694286d81c035c8581188c66c02f2a771d4644ade01e75e77ebb153002cc6fedf4cfdd1969ff5b816f414f82f01f7c4362d47d7c43adb632beb86aaadcfc4b29db9858dcf62e058ee1a65fa4e3e382777fa08aa6c7105d7d73b64c9ce72;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h16d31ce5f9a723805c86abd4c3e1c6a6e79c431a88cc905971bcfbe5b98fda2d66eb207d2262ba56115e80c5da35f6b23c9a12f156144f4c0946309200ae9afd1a056086eec2e6d5c41b91ef52ae7f561c3606d13e97d4499e7a2fc89723f0f94369025eb574f79df10;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h9126cc1c963ee07b80a2990273e0844e446d0e655e36a3353e49ed8dd81630341b73c40204f416ec19ffed5d2e33768268fe8b97ef9a680adac9bf41cf4f4a12f81962cce05eb099d943b5e29f8ea6a90efc88c14c618d74d0d1219ff915ef578a6fb482f2b24aa95e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10350fd454ff68b4c05d0748e8af077f6851c4a9b508d03929a5a15bb5220c2bbcfb2d8b697e01d11421a29e26f96384c7fe2c1614eecef41185446ca2f8d03044279cc7e61897f6a1645828f73ad80254ce93da997c812ca2822b41fe73b61b5121bc500441ef73a07;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hbe0547370ab73df6397359723e5beff1de14419d13dbc10690efd1e3b75adcc607e53ddd2f2a40966b539f7cb2fa6485154e9680470a7ba614361227baff0e52588df405894262e28b8291d5cf502fc45c7d4483e5b3d0ebd2b83661c56fe9f7169786483a19e0fc50;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a95cffb3dffc655031c638d3b9ce1ea7e9d5cab0171516bb3f5a232f3064607bdec10d6c8ae31106e0d49b030688837a13bbc961eac3129b94a52e56a4ae8c73ac343f9a301a764b3d7630e5d0bd54bc0f8fbf4ae5fde81610be3556b39060134c3b34bf4d6332ea26;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h7d165af0794759f3291742469e01d9e02d9c97cfd5ce087d2e37956eb445587ee396c3234578b9b19dc4dd8ea16084eabbf7bbfd4423517ed76d44f13673793ec0cf28f9378e6e3ce062e9524ed0566b0830add64d0208df1dc088588be5e91dcba5e572ab7125e674;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h9e6b7ddec59bb95bdd8f2adf2fa70bf80bcbcb1f471abde349d9f8fc831f1dea0ba291d9c5f0800af3e54c81788ff966ef34ad6c23c9ecfcffceb113e875672121e5db1f7258b0c91ed61ea543fbedd145a6f478dd5907c18f015bb2c5141fc2186d879ff38210847d;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc7b44210da9e3bd2a05ed2323eb979c3b70630ee7e0e1579344dbf8e7a8a95b4d1cec14473d9eb4ad01078b205f5e136e946285b352815503e5a2971ae11f5a1dcbfba2ee1f557ee09a265597d8af62ab9ca577a7cbba56a225a3651ee1fcb3473894de3e808041ae0;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h135a68b69dea5f0fb73af3fa2e3c8c606ecd435ea21b4e4478a654d69e9d4d2fd2a9e287ce3cddc559ee042f46ee1f7df11f073ddb25e36ab157da5b3aecf03ad6d5b7a3e0706cafff6e26c23a3c6d2764969bc4c73ce122d514e75f6790bbe5359c7565fb949a13c77;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h193617738911a29b14c4d813bdf080589019cfcbaefc33c027f49e8e1c2d15ecb243c8d5cb7f4355f8cddba0232617a94d35053e3be22e1386626c605553a7862a913b36ce992ff55b26a01a6d3d4409ab147a2237e7a57606270f1e33e214f9a0cf36b91435860a14e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc86a432b0e93c6445047d2ed4fc9c4f11a13d1b9fb2f0832f23dfd0bdd1c3f0b12c2d0104d56fbef01f3c369336d657e41718d7c78caa93ed7f367e780dc350394f2559aefb0f026604f8676ac9157c45817d768d4b486fe15bbe83f8aec0bf451d3c982b7cda41b05;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd20735aab0f4b447c79b399078a03a81b1d80a088c67c18fe7d4d38781332f55817928a30dd843b211e4e3bfbcd0845cbe84af634b742cf690fa4ba8295e2cef467a84621dbed3cee24c57f86febb84b7a542531f2939ceae8c38e298eb21323b0b55ed2d228a80f76;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h43b44b1361eca12edbb07462f8a9348a99cc2324cb1050d67f4771277fbf4297595cfcd93e365aa1105a8d58d653aa98ed0fcbefc35694b51c24385d8c7b2e59b7adfed84232921a3778cbbfbb5f11570bbfc045966866fedd7e1499a07dcf5ecb78c9f1e19af8c0ab;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hdd5318374301336ede37e391e6e420b3c18b684716ae06a3ce3db85db91afc7212f7f11cc4b6c3a1effb9d434c980c2cdc84f91f05def9ea4bbba828c2640e7cd881af74e1d15d47c74be0b7e4f73967c85ddd1cb4ad7b041eacb73cf197baef5e44302152d69338b0;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h749799159dae599cb623a91ed971c97ee05e81a4288120db39473509ab0538498d0503902e0aeb25810d70350ee5d62e25dde3fcb27b3335d5af0c9fba829837de93d9e183312622559f21bc89082ae6da37f5dcfceae8687b1b4ddc24e7e2f56d148697f5ecf5fd41;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1bc3bb2081b0d9e6b177936bcf0dbbadc0e8fb15ec081e8e86922d4b592db270ddecc262ce9e6b586315a3a2c83dc75e0d0697184aea5cd13875fe51dcb9494577acddeec0bf160acf80c5ca028ad3a087965f8b444e0c2014469c2b0842e3fc313919350ff19b5409b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b1ec44af3598d72014cc0fc6d468312a21b16263b7a5f1f4cd6665f7de1beb9d4dd8a2f4804f33332e4e3ba21687c7ed0b6174b276182b6fe4a47ff73938814ee69b90bab4d277ccab2354bb1f4d143ef96a77a1d5c15598229cb50ccb513c12b03969d027c888e367;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h18269eb8792bc655feacef193cc0cad10c7f21d380889a48fe9219d786f34df3177abbf53c0e653e57982b28ef6eb5ccaadd825b9b96adc029518774de72139669b02813b8396a402f0adb1db506c55fac2a7ea250a27e06db00f9413cc53b1ac33759b970742d009db;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc8dbd832c668b66cb82c9a7b778b301f5bd93f962c47ed3b80d25e78b7959b665f327425b5f46595fbe15d49a98135a441e6e0ef74b139449eaaf5008b1890191a0c50af76128d072b88594179d4bfccfe66d27b477cc7d508a1f14903cce7caf6d101ffeadd7792a6;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10da3c40c93ee6436fe96fe77ea69cd3b2d0cc941f42d2a7bc59c377ccf3abb30be2182dd70eabbb922368feeaed1db218622991a6c7cb3dcced6bb76a499d1115efa9c4acfe20ba95f286fcea635f0026ea509eb32833fa96d985f68739fd884bd3ca463c5bd056672;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h5f9f1a0b9f37706cb1d57cb9fe03123c0463c61041351ca6a9ca0eb55b0ed2de0481c01b1db79349f6b34f17b4379b1cc8d1733422185ec729cb10abecafae097ef55371a81e4d0cc21303c304292594db023b2a731ac8b5f6ca3aabeccb3bfe86baa99d63d8bca066;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h159c69c2fb5ec83992f643314b998b0533eec8a51f50bf7fa26a011cd527d2c78d790c1c23b4bbbbeb0255dfb6bf32d8d97b614d765d0e63d7b5ad6199d066839fd759b7659edcd0b07f47ead28a11e4057263e47de63c86650e1d0d6287264930c55f30ebe986b81d6;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd4e891d54cb5394b33acd57c1c03e23015e2f27929014ab56e8b90f5b11fc5567bbbfce10137dd52795a9a07e17562d2fa134210fba9f34c6e7eeddda0c01d4fc13ae415ba790d99e70b806f3cd686c9491e95758a0c53a3286e49407fdff5b542064f399cde48342a;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h491c4f60ce7692b190247e643c40b22c34afa5449a9d1c61a2213231677674483000e62d302bc32d158e2f6af86be24d5086a48b4fbc3225d2440f368edb5dd88f5e31ac4a0177e1715fd9dea0582d49835133e0b201a3dfabb550616cba6ce3f2dc77c68529968279;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc9ce02fcd17e154ece6eeb7e5fa67e37507e3f9cb8c4b46bff605840ac7a36b36222c9b2dea3a1280831cf5a4fa3c27839dcb88c0953cdd0851124d11079d963e49856bc21d8eff72457af4f31af6c7c5458b5164547204109f6e30b7c564b2c20f31f139813182f4f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hfd71923378ac6b9b4700a71a368e58eb4b7ee97bf7a07838e6488e8b7bb96a4b149a642271681d5739281cb6527d7cda21a7d03a34fda3f21fe6e6bb2ecaf9a0fdceb652028c959fe58e455d77cc7751210e6dfe46e161840b1505fdaaffea57a0c0f0b3e591719adf;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b8b83b54dd2699732b267b433a84265bc6d2c1307c584b9b72d1a60dc80f77b54c4d3d58030dc888c5037d18e973bb41082ab08e2d43006d2f26cbf1f2445f0396bb58c048e328206dd1f06dfc2625f2e977b73efa7d4ffde56d539123fc83f4535c91cdba06ff131d;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he5fefb3e3853482d0ad5f9e08019fcce5593817ff3fa28c11bb09dfbe82b2bfec6bd5187b940fa76aa8135c5a3311f32e71de315ec3d921964f3b17fe17a199c12d589b9887e9e1a98932dd4271cbcf5c3ee129df6794fe8e127002e600b10a6d132cdb03c1ec527a5;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h5e69db23d2dc8a590185ab47df89e2d872bd8e99ab89d54706018ccb3e6d180edfc0037e315f926560748986b11b203f64cfc623fb717620515cf9d142b068e41a92bd42d5a8967e6af64953c7a00b03b231714e28cfff056c61aebcfa7e540d0346c07162a4c1713f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he083b39215070dc70cb7fde19f4a7b13bd080bcbca2318df9c9251401b10cae0f7305e0d9effc48acd9c122a1e07696d468bd1349c81e23618cd2cf1c47d885e2a22f53deb844142dd4ec8af090a126f07e50f8560053e59a16dcde1b3c1014ecaeec52e9bdc6dbbb5;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h760117a116e907ecf37a6bf644f0cb4c44889d00947df0b2f3269ad6d8e004d32228137fcc019b4e84a74d315e6e750f6682c7baa69ea67f80c27f46669f95ea0de9583f10a6828f166deeadf26dedabbff61336e332ebd037af41d0ff711ff08dce9dcfe7d2b8159e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b653ad151302e7c94846544ea59dc64ab113d1f46f3a1c1852fd8150375fbdf4a187abe6cc99036ab83836ca0b051dfe034737532778011d3889af027703d38dfa8dc930312abc13e0cc35330f8dbeaa08f508e43c72e8cd0c09bb25bb424a3e6e4eb697f5db81e91d;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h13e14386aaee45a445932ee7c3cfe6aed8e19b2723ebcdf5744d19934215468fded0e4e1d4f0e7074ebb79d202856c3a18592dd6850b1c04128590c250df1909512e41b316eda89e261072a5c2f8de428f0b1744f635838809eda9e89d8b4747c2271f64b8a0cf49631;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h19a54028ecce0b4328cddabca2289e10f91b72ec94a3ee13035c7c703b8e0353b937252ca35b8dfdffc590937281b0c830879439e95105ce760cdbf43450a80cd129a646ce6bf8845cc0ff30842b7984cae64bd1469b8134269a743d110436db3ffe36f6a0555e37d57;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hdb78d439e45b1321efd2f5a13a4f79661332cf3623db6434139082f448b89f29fd65947d6de55f2ed1a543743ac02413380052a8359df9ec92f2dfe9f22f078471fb033239e9d79b76dfa28a8e222e2f8115150e62086b47337e8ae6f21b5953a4b525c13e8a0f18f1;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha44046b838d21a53e2fe653f0cf160d32fd74cce36ca9f88816ea91924127da6021bfff98cd5447da2196a2f807a64d726c3f7b7099dbd2834d244a280b23917dd16912f432d80ce05cc68dce41c75409c6d98d5fbb062d8285170bad90dc694a817f5e563c43aba38;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd9d50a4d648fcbea112145439a10dbee620e60a578332a6a32e5f697204bbca021e5fe14dc6d4ae99499b14568978627858d09e113eb91262089291d2ba16c130db819792279252ddb295b7b25db4a9930ef90593b19265d24486e3baba7e758ba94479754e5521d35;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h31fe98b7a58350a1fc83874a85d90f813043d39026e1a9e1e7727bf582b86cd8afda42139c89f4c7eab4665d5c00f1eee50df51518c0335ccfc469d8d5c5fd11a94147693194f6043b00d499b5bb6eac33241d45752d2750b656f6ff097d8fc8431905c3f12b894429;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h11b866aa8bfc02f81e4371fcf4ca63fe687304ae8c3e991aaf2256fe87ebd00bac7546b575be0d64db0f2d7f3c57beaab3038d336621de638e999bcd674e361bcf75623c8a2338447a84c8d4a6ad231ca3b70e769c30480f518a9dad331250c09d22dc3353b73b08d93;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h451048096db1fb26021f845215e8c104d6888efc1efffbe8b69230d28163a23bbb833da4b21298331267b3d403adb348a52a369a29beb3cfbdd0fea0b4455202fe0e0a53323a78248c26da508bfdb752d6462b230eb46db011b3319a0314fd21aad5eea852ffe50887;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hbbb60c5a264dfce90e297dbb2973e244904bd8394b973141a75807583c979f0712abe03139183bbd453bd62709b2409d13d21888284cf397a2db381245de1a8375adda3a4aac37866f43352a0a9ca4df1460a14a3159b9b89f16a2a4593155446b9e6b93390ad534a8;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h51c442cd44dce41d3905168965e7d939ba8ba27f70987ac7517d3db910520ba7264d1a2be0ce94177dbf5932c6aa88c56b4728000e959be787fbf200ff24b4effb2f64f16d8476e531c610c7c0bc1cd5874b3ff10320752dfe971430178387b8e21fbea4e8348d654b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e61794ff9acbd254639f19d69c96d2db7c10d8c3964f2f77fa1dc039db4dfb150fade32496e3d43773062c67f64c27fde93293a9f139cd5537dffbff5f837c44fa55e2e31338242e88b59f9adf193d031dcb3cd5314c67b304281d9f33c8e4dc6ff14bcfe93f17383f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1fa374d82bd3e31753e4810b1973b32debc1892597eec38327732254a552f6656467fed17ef8a679ed152644543866d28d84e179f862ceb9e239fadc173ba472a7e2750c95707e91deb01ca8cec4fe835dbfb9102b26cb330e8fd347f66a3a9c45b476e969dd414a1b2;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha89f1ae9e19a09d060cde97eea2ce725a4961208cf6adbf69a24a2f4385aa5328cdff5017f432977158e37d3de0699f49a990396444dc52663895a7e9f06a023647afab37b556af2b71e7f9d50dbbbee915a2428edd48adf45442d37ef263bb7ce7359f6b84aed40f8;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h75d91f0bc44224bec253fd98ef7134b923d0a357b6d02e469f94a23d3ef5848e1f83c4bb7ff1baa67b95691149bb51d1a44433ae7b36fb3b4fe055401e8be17e0072c747ee7bf0fc16dbc618298382253cc62e28bb76feae596b92303a025ec1e07f87c22ff44c7470;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hbd1b2cffca803e0c4fd382c51c83e9c6b26aa1ab9c1b0180a7d44864384d4dd4bac69a4187ad462fe1a76fd77607bb954e64c872fceee0e39c0f0de3db41a2ad3f1c95294ff7fc8d2aef1ab24db58007cae1c2d9187642b25281640f45deea94e57d444755ea8625a5;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1640022253d24a5a0bb479eac4580329406c59b3e876b80b9c2806de8ac34bd96e6745abbf0a63966c542adcbfde9944bf450b32c39de818013a07931cdcec57511bd53fe4b5236e0e94006e530f677bf4389cae1bfd7cd49c86ead94afb843cc9ff957c82a95235122;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc55ab7be48a935c3d93ecd729a5e4d8ecc0f6dbaf970138264293c00aefbdd5f14cad5444d7a1ee4db27455ded15ebe1bf346a50dcbb6e02c950d61f6a3fcda07b398eb7876e275503efd38e571c2041b4e1b9fb59f25ddb44029d24af2a8ff8eea9e0c8de3553ee61;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h54c928d6e58d12d77e3da41c3310dac02b99d71235f73234519242a805043df0a647b717878ef2d0d8609a8c3cdbb4865ea57cd6ccd04568f242cdc55780cf8e95fa88bfdc7dc64ed76dd76f556ca1744555c8809cb28697cee972751d133d420add7d19954b71b126;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f9c7e624a8b9f02195e40e7fa085568082f9de1595e59363d67ef9286df7750eb72cf101bdc39c66b1cef6a99ccb4a121db1140877d8936527f070bf1eae4be9d3972f1b2a7cf8c0c626cc7de7b19a543ba13f6c84862d53487c7607cb1129f498f115c36984225618;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h9b85c413712af0869505ad1fd62a17b18cac690ab3131a35984cfa68af2631de3f8b3427dea6a15de288932d5056185bc6811df94e1a244916f6474f7a63b76965c586cc8cf6d053fe88a93782b27764c15444abf36b773fe67e3216e03e50ccf25b30313596efad5c;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h2fa17a6af16c3c85d82a00f37254910c5d2fa294b46e8f2332b6dc9fe01f1ceefcec94c05dbfbcc46a5af62548026bd51f1721d534ddac4c836c17cebc050d5d3210d15f69a8c8089c83c552de22b774984265c1dcf9fb691fbb02dfb05365388bd35c33356f01597b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h193e9043804b67f48b212f98eb071c0271c8f0527b5f16e3c160dc840b05f135ecea174b2efdece685639467a5d36fdb975a9bfe4cdb959d60bd908920f830c10c80a6942c4500db63772370bfe0a5464ddbe7850f5c8be1895469eae6701f7dec80bfa4a8907d99811;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e10b4575f38d20bda068482dab03c9f538194aeaa6540710aa80af858297571de1c17485206eaa04e9f3ba7ebec96baa6b9065b52913b522c80350ce563c464229029a8b960d3f467ffeda6cf83f4a7872d4b46934da5df9d9b844c173d927147e2f9f6841eb552e81;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha3c037162dc630c93395ee0d85d6a75570a2a826ce6768543e6b4813d35a7daba2a49acb90b43181aab9532d7662637c87aa89571b885c8ba68ad63a58fe2635688cca2a3ee5f09656752303050da83c3550d64c3156cbe2f57b7c4a2e4ddd48fd4c139c24c1a8c1cd;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ee350b6fbe51aaf628e31791321eff2b727d3ad2b0fa4536241a9c2f04385b41ea4d6a3d0227e0e960a75457a221b1414ed211a4a52c688d0a0a2d80a58283693d57bef8b23829c2a5370b30e4b4c2779f5386d2547237d2a5405556ade91746ff1139b28e5340b9d1;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h7d403d27b3ddba38d356bd3d58ffc555f479e899162a8404106ad84e5ed4462b350703c7d06cfebda77bc6f51e67533bd940e8c709698a8b7117b9afd83bd1709c122bd15d0d6b18e1e23eb0d133fca2640417c975080fa39f3a920de4859d0501d4df64b271d76f3f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1128f0d108bd030f47149dfb61b249e5ce563e56b90f98690743da913407123a8a05af12610de5f8dfa236f73582b8ee95498990950edffb9d2b8672d414356301506b641121b84292778a79b28cea6383e7647799a9bc9ce23981bcc1314ebe0bd9b1a8a01131b4ad8;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hdb472c8439712dc380b9dd7fb6b3b5a7dcb717c2ee342a5e8d255ad89a9708faeed1caac45c669c816b9cc3b57b60e46f01d12252a4384096f88666f08219547efe860bc81e57951de96c70a2356747c2b5f396c85a2452b3dd4f7ae030f1363230013d0f8d9ad74bb;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h16e92ac3c779809c178135c9cee8895b439b4490975bf3b0a800320b40d9d7fc4a55ccc71130dc97e9bcf18ac6ac95f7717ae00d78ac1828b69587e950f4f774ecc2eec57c833c5c841d91c0b386cfb526fe4b0ecb2c91deec384a271c024debf090eca6994d638cd2c;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h53bc6c5c369718a22099ab23668e5e883467be26d1a9223837de2152f908380a6d7fe5df569912a393e85f9f0f7065683c90cdbe67fd0c3bea365dc62c2821de49593820560cfc78e32929f20fe06621b8d67991fe60a86a8acfb18da0e538b2db4d2aea68da4008cf;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h8264f273f325737aefa4ff80b3cbfbbc912f38d0ba6d4b9e9a126269041c64737a40f712b070cdfea76f87bc2b3fecb4b093d41c0d47fea8d3a7386ae65f6c9fc10b5883cb9be15a2c2cb8ba2efa30e0fff980af10cdeeb363535baf2cc9d766e6fefbc092ce6bb03c;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10fcddd047611c6a13993de2606f56bf9516e26dd5bb075a53393424f7c1a337d523d06b145c624739af5e20bcdec7032634a6cbaeb597af265c7d570cb3c95677b41f9773427a935419e630d8482dcc83a3310b7d75801622a98855a8ef9ab962807cab2b36b5cf078;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1483dced4fca8009a435e575d304250a59af529fdeedd0e31e50bbe1970cbff39348a938441cf529f5ef147eab8dca84067e0838eed9cbc589bb702b43b10de3efd0fc0e66aaa8916d9f9c3ca73ab7395adb1f7bb0de702a3901c53024e65729512c7d8f74ecabb2bff;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1295c05e4c0d45a73a76c96d0ffeeb47b541333353a41ad92294bcdfaf0341e0144cc59597b5e65d1e7ba0eb219ab8c52d59afe2bbe73c9a772c8813654377d55c702e9fca8f016a60adfafb2e3944cbd56bd9638d028e402650503c2f25bea3a16a5159036b76d9361;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h162440a06fbb3f8fea507bf3b95569efa1515d92ba5d7b1f4ecbea6bcdb35d1595591ea294fb83aa39ab0cd10d3b0c2cc4707477d95a8c04468ed45a4707b9163c2ff9ca3f70ec14ea20ab4373b50ea79ffb112c0ef83e41c130e5a58c5f4f0a09d8be2fa9e361564e3;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h18f3aa3552c78458dd5b6258e7ee781acdc535b868580687de3756848c57e6425f653856b8418f0ce46b83034aa2604434131ea676d9e2f604c7faa700ff07e64205c68153ea2f6a540d014cc16df1091532a91ec3cc32141c03d89ef91596bdfbc281285d782681f11;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1614e2507853b4b4292cb4ae1e71a43a6f88aac70b62c21f3e2a9668cca3068be7cf32d07f4399011e2583f2aff9209b6b8c4d3f65d25550b5b687484dbcad60cf8ae5a4dd0452f6c6fd286929f8b1c81baa10033421a29f48d10ecd325ff8bf4b24b38385793948dd;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc1c484aa155d07c61378b88acb48020e5d865bfab014fde1adb633ba3d0e060c882e6714c0f2e6b3f21ff4f02902c3ce1d47c9ee95bd5237d897ae1826cc19f7a005ed030429a47bf06ba6bb545f0dc1f3a368cc1d2e1880cb8330165ae35b9c8bca5a73f186f68bf;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha63f1128fac98af1fa623dfe6cd9be1c528b3aa4ace44ffc7eb354c692bc8f92c38d3dddb8174c72ac4f190047486443161611a60f16fa57a5be57222a62fe85d72e67aa373efb6d12dff4e728ed71a8ac8c6c222c6fca735c4b2d50f4202320a8c3c5b203819efed;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h131e437c768118fcc86780a838194e7530d2ec048f576dccacab77e09d2b785e8913573ae5638869af0b436ddd0c498da06e490ecc12365ffee4d5e955bf2a8320dc554f41b49c1c7b2d84aaa68c0fca4ac330c8b3c27621fbe59cb5dfb8ffbfc4f6d9d40d6687c0e78;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h155effcd7355afd2acdea679099f7c1fdd882bfa62c675198b19bfefef10ce77ea45195c5125a7ce73d4d9865ff06564b8c6d8878b276a8121d2d042d35fac438de74db35c4934df8ac4049f8900dfc346e95fc9d4325e42f81a939f77cba4c624c4cca46647254fdb;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he71fe6145db22081b675d8cf7ad5d4b9c4661c06f3fdce6cd4d870f5a2b666c8814141d2641607f96c84dea4ab6f6cccfbed35bac78699384767a0ea83520851aa2e499ce009401df4aa4bed2d70309da817178f13eb15b32baf8b69c59a238a9046252d35c5a0c509;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h182e66eb895a66a469334615357717716ecf3aba5e3e81e8bac5bc1d7b85a150dd34bdbb2b6db6435d73d706fadde2106b960c8b892e08cb31b8694cb09642dbdcd59762ff612607c5f3c777d38e06d491f16c804a2aec6078f312d5411cb6611da8cb9b03f0922386c;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h14d129a5a6671472aa0ecf2e8ea98203b85cce8f56bb1a0ecd227be36bedd9a19f26ad1f5b952aab5d571608c709d1f325af2417a77f94bc3841c46f25a39629a3bae86a35684120d164f4da32746e6d2347469e56c599d200e9bc9f02f83b7f5a712e8c9c40c956739;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f6e576ddd67e054bd8c005b30fa6f0dcb8c83b375a5b52bab352bbdacd9cfee7c466db36b461cee1f551586e66441b29dc2605ac75f194e0c0d4a769f7dcbba109b11fa62e37695397ebb61541678458eaf60cc5a493b608da1ec1cd096a142022001f04ac10a6d0ff;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h19caac74daa30755e6614340fd3f554c9e505feb59e11aa309a940836329c4cc3d40997b225ac24b996acc7b8553925b7e32f0a6f88aafaa59968d6d309cc1a5c00abd201775967d1b3ef2cf3d68f059b7e752f7322c49321f630f396c12e6450281a939948edbc7569;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d8ab3c6e33b501fb2371e1b2b0c8d1cdc49261e950a49261ce6321fe95e0e95d4d101fd09d4640f14eae76d69f363de4e10d9ec435131f3ec51c089e878c3eeeb1d623ca74de8315677dc7e75f1fc71ff5541447e3b356d72db1ef6a7c71669e76ccb246e9827c788c;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h231a653656f94f708d5e76e99b2939db4d9d6806854ab2324b7ff502e849ef2a0f50ccd03df3ea12c4463c9a6eca91faf4e05435889c069a16213a8a7887d42be36c695d2cab7e72ddb6c903b9f63b5930d3e7dcb985f5c52c07e32fdee5d3b2773e4431868d564033;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h6134c8cf3ed4728fd7c64dc2d4a725543c8ed7d297b08325471790d3cd358f03d5232f1c56d16f81af472a52c3907ef59abba7a8daff0b879e3b45b50332e621400534b55579a78e7656152b334731ae2103b3df3992b18fa305f746e20cb7dcf92a839c4a1576fddb;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hab4efbd8a0036ca49064281dee9fb1bd3a111f232ff91dbad13602b9e5135e01c33f0a466f5632f74f1ee7578f8a5b51dfbd06060948d82c0d800e2b66dfd81b462dccea18b473f949db78b1fbcb1025811e8a9c04764d7c7de9f739edc75befd9b7a24e057e16343a;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c68a8fecd2c5468f099145a3916d272355a716bf31569c65568617fc19a5a1664d388666050f5fc9e0e9568d75a3bd0485bd32519b646ddc3cb6b9ba3bf62deb16613f3c93ece47cff08ebbae5b076e5575e5ba35b2e615ff0d13eb458f7343f45692c7478b736cd98;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hcd9ed048dd80a073f66b3ca3b2d307aa9ff3807f58baa963091acb5a9831907841e35c4a349ab0681c07bff6fd2d6a89465fd49ee647a5d2576025a6472345ca0cb8e52d28ba6ea586d791d220fd6e1b55d09026ea5a54ad16cc97bfc44c58e413446cb7ef3edb7aa0;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h123d13c5885154bc979da9d09088cc42db9af930a424a2c455627ada0a7a61a254fe1c3a053a9aa03662ee4d5ba070e47a5749816ce3697f1dbc4a98bdc4cb3b75095667482c2602aa2c95d308b959d5b01de792a3660a62297a51bfd0122735ec207410e776e284839;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h6720b730ca411bb01611bf96900ac919c2a1976138d616d98c39a9cf567c140d6e3b0be0f62111b2734a310b324408ce47cf12b19d287a5f59bb4f51790608f88523725a82f7c2abf0c7b2536aa9814c0a33809026e8e0421e89678cf1860aee6fbeb154357b2dcbed;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h8b323a249901669ad743a570570dc503a792967d956071aa15d32db563a1adb24316b992a5eab6de21e2b108d5d7e093643673850979d156951be8544ac43f60003531581c9af88a12dea7b237725ababdb0fc23dd10fe67df4de2fedcf8814917af01822269732cd1;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1cba5b70001491ba5f1097227ec1ff0646f1f2dac27421935a19843fcddfcc3ae6d9571174df396dc6f0dafe09a8ecda8acfdd50f978a731a7441389defc2e1e4c7a8340106ac3b60992a066cfa396640788b789f4de9bff0bb251cefe4f9f6c656907f3cb2cd83226c;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b33084473c5f0e9c0848051b74e564d96b2eabd4a72dc7f41b27788a8dc2898166ec0e3ff87dfb38f06ffffeac774910bc573ca85b2b09c754c299ce25df2b99c983ffc41daa8b75c8abeca02751f382e17ba25df6226e0b68ad8e10b232a2b431f1b5808f3db00bf6;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ef6b17aaf4762dc229c800b213fc8e9d987b67cf23ead4f6df4a3a8217e3f49ad640af0a24046a6baa616794f3374dc9fa4dc83cbca5b484c63345fb3937328433eee56dc7eb30fb6b76f188eb4393983926694526ead047d38a2c0f280c85c833b366da82a43cd97f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb0e45eddb388eaac1c3421ccd559a098a5641a079ade5d3e52dd24e6735ebb62e675aea907a2f5677317b4d0601189154fd809aef21829fe519f745e0fc70174b5444fc7c6ff17cebc379c822cf03b4d75e1bcb12de17e2211764b9a9e49165b3d4c1b8e87fb94ba62;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h108a113d62bb3b8f556c55234461b9ed3443b79ddc0e899c56fbd934865a0b2d77e319441038ef0100161023b23cb4462433b5cea64078bb85c0c0d0ddec127a472e0724401142bccfc0107313010d25b0a3b3cdeccafc9e5a8fbd6da97c5e5142eaed1695028ac5956;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h149af05de5d23b66507df359f43b680a9b2f793d7189c448d2038bbf3774d3c6fab5ce591e18b91ba16bebaa6f487e8fc12ef8e8f53c5da295003756a0377846af2899b68fd8b01f2d86ee49f278c13e5ba8eace40859f5d47ceecf55997a4039c28e32ae7537843579;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e60770f5cfa3e1905d5c2941a1cf01b1e8375db965e4bbc4515427ac21cab7d2336ac2a6c01c8e14b7e5611525395655faa9ebfa5e7f0ca8154655288b954975331ebe3ac4d1b3fcdc089119c92c58191c32c22093801520ec0cf0da7ad20be99c7995d6fe425aacf2;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d61bb70a119bba9eb2c6b305ea612b71bd77ab316c510b3c9af1bce06596f9f265c258fdb207a50be21c1083d1d0b596b56834f03eabf8f4e93b207438163f5233d7d4baf93364248697f2472f6d1c04ce01ca94b62830e6561a09118f5b8b6ab46c389dce76be3ec5;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h111813bdf588a8e42b8742e2ee40c38485e6226ebc7c2f274aabebe66095855f87fc2023129c11170e2e0e0b39b34e66ca165822cead6564705cd12bfb6a95c0497f29aa645432b60c3749eb967f7c9563ea8201e3a3305db25b652d5bbdf87189c9e03fedd27a0d617;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h13ec014b363b2cfc966cd8375e2bd916eccdd88c64b698a53756f2dc76c9f8c4e68953f85cfbc452a924f330a96e70177dbd26d53239d1080e31dd0c1d6bde5d527db5508493710020f8265cb635f79453b60f7fab16ce37ce61b6f303dee36b733791bc68c1abb4705;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he2e5230bd2722159b75c1487f8e1a9e8b82009981cb6c1171b2986e3cd5e15f1dc2fc0c50d7e64c961c16d282fe755aacc9b65ff6c1bc01f067317d36086f16b2bb72c95593db0c4ca35220a930e875a89475833faf7707ee2517706440191b2a6221f3a829458b5a0;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10364f4ac1ad9e8d248b9128d3a3bbbd45802bd83f17e5761cafb8e61b9ab697e41a4a6a3bab3070611e1af4faa4ea6b0e5835d0db6a064ec07415b264fde4268d624ad80ebc16282d0b72b9adab9f4117522f33d43b3d43bafa5fb4b1235349cf38f14d9b34eaca539;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd817670a8365a8e0e095c78b1b67578c4b9f1cdd193c31cb5c98e3175ee5cf5ccb29296a88c044b7000a4669de12c5d3eca9062056d83afc8185516604e61d3b5b90bdd2a722f5206907d6285d16427b23597ca1466541be1ab81123dae39446aa31af65ebd1d33b51;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1597fe2e06332e6369c9e67144367c8a1e5cb7c848d70df5b7e5694b6a9a5610eb3d2875dd87b79360692e3f0480c60fea2c39c3fad24da1d8a5903341d98718cedf08b2b6e31880651dc78da0896e8c27d7b1dfb0f8f76e9756ad1a8b5ddc52100f752ccd96d97b6ee;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1435258322111215e92fb7a0d66321216839e17490f2de1594e85c6a9e123ac0c1ee3444a7f52120237c26a83dc0b05d83540d23fd6030d3875937d9f0af80a62445a07578b8581d5816da09c8290e579366b9bbc000e00e762823da7e1730736c95597a5b03ced2ba9;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd40e33ba16d7a55067ab0d3eab45fdfd3f72746f9de01fb6393683cb64a51c2a2a55526a8b693fc0033fd42f0620a3b52c4e3cbea0bc422ef2b40835273f551831fa47c55c08dc35a8e8094222aa862bcafa9cb527fa7c91a9ac9820dca5ab489b468e8466d7682b7d;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d47248fd33d7c5cac156a1081ca690a3113278b5bf658f0138273cb234971676c269c0757be8f8f8419769b8066b9e0b54259736abf22133f7dbb5b66e47109e283d8d4c039804765062e8a97ba0603fbdd059573938b617c27fcbddefc1fcb54e144a0a11d73d253f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h14b332b8f28c21f7ed76eaabc6d9b50ab33283d27b29bfc7d0994cdc985b78645da009bcc9a97a758fbb7a0209e9503158a53c2d36fecd14db81b2dad0fab7462f3b85c98998a686f1660abfd3807e799dc79f867fe24fc1b021c36a01e250bc3f1895317dc5dd63f2;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h19547fb8b3dc14fbb50c0e720a80e464a8647be00fab15782ea932098bd75dec607c3df60e9cf4cc1f9bda66487f0baa608085852e77d945d99a4f58d5790e5f73f0605bc3ac5be1ae50033254f29d4f5d9a6211f443a83a317e53a03aca671e901bcb7925aa7bde2db;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h238858286a41164aaea505e7509d18977459e25fb7a6a9243023fb3aedc7b271efde80b54a8fc3d7cebea8278d7763d7bad69d9664aa1ea0c207792f78e39c93c1439f3509c320f2ca9962c76ffb3bff647db30c57f69bb0ac786455a1438db3b60846a64257e76c08;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1351cb0cf01a43636d9fa479b8bb3bcb47ebf131cd1142c575821ccc13022393c75dbffbef3434fd6dfdba1acf22721e93ea429ec23827a03f074e4633eaf70ee2a7fdb1e508a0ef72479a4b6fcc57d466a6a02946066931dbd484cb21d74ed1b972bf60c2a1c2dc64d;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h182c8c7b88b420a44520eb43e1bcc8c8884158085c7ff5ea5e3e368b537dcb3b1e8034056148616ba9b677736ed5ed5d8145f551f7e9de9b9893acc86b8a9cb4338b75a7771482fc58331ca87c7865d65300a1bb63a9e0d2e9d625f68195a54bc84e3e900ebc4720b44;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h14b52129f857b3b3b20e9c132a2d9c1bc5dc90c9373aade7441770b5b8c5c66d559ee6e1485ac586d8aaba64f87feb1b2f026f86ee20bffd93e508c256e9c779eb5bdd1e77e033bb1501e1861bc5821ecb938cd721b4b73b4bc690b3c6c77dd8761a71651367e423d92;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h13b1dd62ba61e86c1007a4c13fbff2a6f105f9b28f5668259c7d8276fda48f92a50c7a30524026f485c931105d7e19e73e2abd23830003e832eec443ab8ed984b0ba58fea9cc6ef3acdbc88b18bae5f779d73f459f0ca04431f7097460e1c45bc6b85e5f32edb118c7b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h5da4fb276ea0a76dfc01c1eac275bf90837e942a6e8542dee23776dae62656c04f12d209d410989c80a62167cdbe4206a192b7fad98b528ef23b01f8ff9c44edd9d599fc409758aad53dbbe1408b3d7a146860580561d6fc4fbdf54879217fa7169d71618ad315830f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h165e47cf8c4cb76dde55e65423548ce762387f5a6fe15347946edebea77ed2671effc2e58db95e12d3c9afd9b809a00e392cb044db7a64d4aa6863ed8a39fd493034e4ac4af5993719231d8553985bd43479144c48516020b6bb594316ebc69c3348b0dd0f5e3f75bbf;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha40b28ced8756d05eb1bf5ce8ce726535a0d217f04a46e07eb14d9e7593d2eab8d418936811e20dae4e5d0c1dcf9b741db295d45e3ab88a0c93318e26f90250c44610d7d7eae9d1447724a2bfa261e1c122473321b244017ab48459975cb6c4652aa3c3f1d6b77674c;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a488d472e7b60786632a4439ed2a902e0b2f0c55f48b2c081ac669cbf49bfc64d06df265ce4bb20b0f77c0c830823b4bfe9aed869942c73f3b1a2a82a7bcc3b0a676acabac7eb9232d5b57039cfb8b557d62189712726a5d6d826d4387fca4625d44e66820952d22d5;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h427c9c39bc55b25d829a1a5498d3d6ff7d5004fa3758c84c93ec8ae23db72a2b7fa8f1178a4155f966a0de09b25761d567a3a5355ad55f807ddbac9059a8aba0425307f56aee045be6ecc45a31065dfbc1ad2f28f4d2b951477643cccaa70e10d3c84a69e1e5aa6c74;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h308249cca0b37d8900cfb5e59d662c1b94d4bb876e5152dbbb1f91ba08f335451fad81c500f35c0b993fc270169f71b345b308c1c31e2f17293878953e7737bd03e9d58604aae5f664660599b6d0edf8cfeef1830f49b572039f383f592f16bf54344332f76b336fb3;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h3db66e5f89a52d6292156822c2b4c16700b185c5eddd01205f0ab7dec3306d5bdb59a20d8f0993197dc4e5ca62e82631659dfb7763c6f6f2fede5c12c111052b141d7a0a6d4e0ee0f3d28f516cbfad827ac1916596c509f4debe24f68e80cdced0444fdcc26c303fb3;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h80429fb89fdc05c3ba52cd4e1e79087822b3ea0ea5bf2a4c4574368d32e9d40deae18c7e2f525366b1ae64eb4f1dd1100accf405d3a7d499b67a8427019ceb607f2b74db94d3a771457867e67c801e19d8feaadf735e0a48d14306944720634c66e6d616b730170cc8;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1396a319977d6eab54898d4ba9c746973082cb8406e577772cb5058b177754d4b1c5174f2cf006d1b16cb1a08b23c20432c2da8f9f067bf5d677abea2e24ffe2c419496f1b4fdbc425780d76c3960d24f9e2fd4d10cf163bcdf26e030342a93f9a8538af305919925bb;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h14539635f59e3c06782ebff53c9faa968a9e4de13a424a595a82bda56beabaf322b9082d5676decf03eff2e9b96a6b96eb5a992d12d3a581e7744abea6bae9f982107f62ffc3d7a396a7c1d4f0e0300df0ef9c24981514beaf2b8f79a2301950ffc62655b52dd26932c;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hdfe6f2468caebc95eac1e0842d29970ef03cf0ab5ed8b86b76f0af3b9ad824ae17a89d19bff152550fe95995b42995934b0932d02db663fa1bac9499b84108bf8ef0cf7180d911f8741c9b0fde69d7aead63ea54cae5cc7ff89ec1672dd8c7dce4c53328d6db3283e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h113c99e280abb7c27de98cfd42bf0d28112a905bb0141142ac98ad21623f6f43a4a96440d2d1e113e224c183da9482fb0fcdc896cf34e8b3c997dfbafddc90a77a51b2634cc172881322b5efc526be7cfd87197d28045479dca18bf131fd22a3a77ee9a11f8a1d5fc26;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd8292764859db74e6fcd5cec8c6d4bf9b6755980a4446eb84104fea040d18e57e2d8aff08dee71288989ff540487414577b6057fcd1979aa1236a2cd924cd8202c9611f62b6aec9b3518c166542fa2178e29ff22a89274d6f0f07b74022a4bb78877a431b7eab5f0cc;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h44ea020ecf76c5258dcc7568c25f81551eb34610cc4a76a5f8924a4fb74c31614635df0863459dc8fd1c96474a1f240641ddfc51fd8935f774a556e3c722e02d6040fac643ccde456ae36a09008d836c18f0965e968295c4fc9e788e99d9201a97c760270801283e93;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10f780c0c93e34603efa3ac972a6da16b9f71840ebf22a9598c33430fc71b13ff6b3d9179ce833f4bfd6a33a26939d0cb6184064fd008d031eca9839782f99ed360704626740ef05982cb362ba6cef8ddd85a6bb110826ec229ffa1733c608c2a6ab9975a91f13cbfd3;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10301884be96ede5f08377a571ac35b0d8753c0a02b918ccf46cb915a60e70a0c18c9137be861e2c218fc38e6dda2b5c3203def03748bd2e112b806f23ec8339b6b1680ad85e29dd5b12fe1931ff2e1f97ea1c444fa8eed3600008d33a9d0081c61170b0ada0c681abe;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h56a3587ebaf8e61472c8b949dc3b95f1488da8c6a39db848720e5fa32d0f6c0f8dd0eaffa9c9baec4ffa3ad9fe31bde12c1ed3c37dd06fa330b07d32575a3d50839db06bd08bf3dbabe6a4997b01115da71d5be8135762777f77ef3f42a044d0d20f4af7e9261771e8;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a3dbaf3679538d0b051f606660cf2e19ab19499d3b0151e559ad94404d17d6ca59539e34069f67792fcbaa35fcab6a2d40e0b7abf3d39a5ea4a90e87fa529131fd6c6a5b9ce8d615102f7de9b94b7a58b669f5a98e351bd046ac8efa1ad61041a75809432f85b6bf8e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h149a698f491af5bc068f21996c5df941132dfa82c6b7d7bbce62828cd985c3481a67fffda7cc15c5408cbe5f53d29b851941c2a145486036d6b327d4b7c1f2e9cfbb07303c2049bca325804680c54c7f7784dca2a7aeba8510d2427301bbd13dabcbdd64aada09f280b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h5544fbc0fa14f0eadc33d80f0c1ba1b84e0be1ec02db21732577bf32b3a9cec3342aa1b5cfefc8255ed6a706c827b287ad4d3526d1eb849a3c547a63a06d6430b8e660251a97713bf85de0dc02df83582a2320536d10500e35b3d38619aa7c689c8eed818eeaa7d1b3;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h93e9d345104ad0f8f46135407881e553633bbe6cf4a1e0d0131abaa035f9374143b52872728276843fe46ea0d7bdc07a9a5163366c8386b9d07da400fe86dd9b026d06b498c3deadc157af5f28aa43c27d709241d5c8741867a08996ec8e5832d37e364c5188beade0;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h21eb5cfff0bc968493bdc337d36436f9c74cd0a46a75682753c5053e9ac97a34457675f6c814433a0a901f89bf085b969da8b3b3c279f8b02733dd3c097cae0d9926dd5a3e40b11f68046453fd3b0bd3960e0a9325cda73c76ea94a1b5e3c6760fbfc5dce90d1b99b7;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1caecff53f551c6a621e8826bdfeb9a05a984678003349f4317e9520e42966ed3cce27e175958b2152db930e71741706f026500b04017121bf181d130bba05920c62d28202c4b876a7ccfe859983eb1c6d87b1612b621cd033c8d076b8f339f1c90843fff98389e6dba;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h72b981669ce83af6266fda04018da5bda9fc64aee295ec18ff503bec8672510fd7ecf8b5394e075306b295b7d8c8d6f4e63c20b20dc9c673c1e6d58d45d65abf2b1695cd9193391172322ac98ee61cac9409ed7a0b165ea0c8a9e7eae42b8caf83851e04a70f4b56c7;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'heb46622c7d30baaa8e4c9c5a0df223cf713bf5cd20259fdbfe5560f7ac980d76c4f4654ad28328938c02f2a8ef1b654e60c1186a67c1d4ed1cdec0ccf28403a949af9ef263d5d363381516eab0668ca4db777c3876e16650565ff9d949ad0a1ce57da5995003b2e2ea;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h34ede367b5d2ccf571846ff649f4e600e72bdfe6eff7ebaaf437be4e5309ba0521a7213c65b84dc572d9824e8a0bd894386a82805c1388282342f006b198ed810a6fb49778424fdde24c15a6ba809376054d6340b9bb124a73f72880c01b4b721228f0491d78f8c02b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc843a30cfd5923e41777e91439b8f159d088af5adedd9ff01be156c5278fe97172853d796384c51d26d19c38811f3e70b3c1ebac33f2225cc81ad23c3061882d39eb5eb2ca39f72a372f59d4c7173fee4d61d2dbedc83c54d43b033fcf5d5096a88eeaca02e62b7da8;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h19821bb0a2e25935f3a3d0894f0470d72236ab948fb5b5ae1d929a5876b4f617e0696362e1495b1f27149ffd57ce39206382b890ed588386ead057840ffea5a2cd25f7e55bf04d8f1221a752c7e8f590a20343cbfec44843becef3642631fadce86d9c1d0b79edc8bbb;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd0151c942756dd8e80ffd4e3235693bc9f8e49c938bdf4d54ea72a94550397e439fbbb10ec8315ce50e8e79dc413135dbbdb1f8a26ad92a3340f718e4883952f352807bd318e19e4fcec446a06a6e46891bc57c06d5f17777cda90bf8290790a15a4e82ae16126e42;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha5dbe9a65d34b55a1094a42bfaefef606099bd356fcc41cc6c404c6d87b1f4d2aae31fd16d3c73e4ce77a795fa1e5c8fb1fdfafc4cc74795a995bbd87fe06a978f00ec04e3bf914e21c6a8c95b17860e01e49736ceb3e1ffa00d2b1de46c3f2f8cbb5ce094cbe1dafd;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf03fc08355f987423256f5d385e6bce18d8b807a98c67d1064fc44826ab272d322b0df7e41c37dd2f7d5fd15892eeb187d7899ff418346ec4c72850e7ac9607ffdea6bfd0fbb5194dd15e603002e22a66cf55d43a8709e3742a0774934632f7c14ee12586e4ae87767;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h13b2db1d66eee0ece3727b84c8e95ee697e635f1725f959b04f71aa4efc150ccc103e54918f84de1adfc31e6b0453d8ec153d04e9c9bc299527cf2da4f836089e4bf59af3a066781920de7a6729bb1ca338210505466a17e00929281008085215e2770910555d4b9f09;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c145e8ec63a8ec876e810fc57f23fd8bbfb29949f10836483e52c2c65fb4f66145757006d1a4704cd852d4062401353cb959216e2558d9bd5482a151d781f287094425d0b74d5b61c679337c1f8efbd5837767214b00d37fbd15a2c40c141b93c47b96b8599e8475db;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h64f37f9c860d36368d592e178fabd48406891dd5845c1a1699cba02ebefb498276f29b44a61e1e5c6e9740de6aaadb8f1971ca2054a89c6b936e0b977f6df32cdb1f3e42f755f94e3c63854cfa1e9ea5952dca8a4c568d03f6ee29ea3320ebd4c885b3fa9c6771a3a2;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h2f34e14cc4e05126132da70680aad792e529f79b9c6d1b25b220c901b1f71c9a3d1c571a0f7475c10205b515ca353820bf1759877143b83b1aeb02634eb0b5383eb382ba89ab5de1ba2558ad3506d00520610a467e20779f3bed5a1325826036af3af62dd46bf45531;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h460592103a4fbbcb16a6af61c4f5698e55e41aed63cccb45e472e3dfd84b95ba2d3e501851601d96b6709b844e12e11605bb996b420ee480788e5bb6c4c2f91630b79a40de770006cae612a8fbf5df3dc56d9c6c36bd734d1f7f009074031ef112f2d0915d139a7fb0;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h17e0b2472adb436c1f9a5cce810e214ebbefb65cedbf3e6877054cd1eaf9203bd9d042f5552e72bd626eec47f00aed91e2268671f72c06ff35fc41ab07ccf26bfcc070cd2acde6a668c897279e95319016c9efcac57154a199c2ab1a910df8b7c0905036dd6e9e7c1d1;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h427a4d6f1d189bf8f616e3307ffa790cdd7fae0a75c9eafe063aeb25a7872f1b522e2b964b16c8e232d05d096f83a8d17318ae33d2ecb45bf979f6100482db6728cbfd91678db11b78f8ed2bc2879f850aba5667cc8b8b552fd1a62b13573bf3277085c51b0832d8ee;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1cb89f5f82a3d1ec720359a5f475217b21a129fd8510995106ac487dc7579edc065d458317d7bff97c8af71f3d46e887f9a2db58d76bbd7a8a273f21849954fe5e3a5eff24ec02ef4de037d06b46c4fca665c590adacf50b9b8be86278d63883fbd537b59ca05484c93;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h45e78ca6ebd63190f7bc4fb8d3cdb4f2f00ca60bbaabf84e0408b883138247b0a0df5a85d2f9b5a45eb0319559e908a81365ae4aa76ab6c7f09a938ff55be793e82e1f2ccfc72531a53fdc9f0a241a1e0f8d0adedf3a0ac3390ec94c1a69bb034d6f83209393a259fc;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h11a5716d3a334d1b12ccb45030f6a4c230be6904d5f82a38b1b8d2d2d306a1e6a3126ce42488ea6996e1439ca0f0fbb5364c4dd39ad8604aa54f0195f6e381d69a44fd751b4f0c8ece4288018a768f0c385bb868d04c0855382c0b5c22bb20125ae288a68555d24d26e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1933c593d0ab3896d10e832308418f912ea000e83b474e00aa6570263d4118ddf43fc94b9dc449329f58d16c92ec4fb0eea4d5901f0f6afbad3d146aedb68c40cd6121adae7a0c1ba3dba92c67d583649e1caeaa0f3da6d8b2fb779aedc1e24771a76bd735b5535e7b3;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e08472d268286ee67dadb121a8c00d13c72fb0096a0fa9ba2ec627fccada1239116a3cefec81b9e61573d4f86b2329b003aef8fa9d9cb9593261a5d5ade6634ba9334e23e5d6105cc2b108a17e802ebe59ce09d3b79a558e676a136a9854a88c7f948b7809471fe27d;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h50c2ccd852134d85144b78e1b3889ebd73db486a415cff201e896969bb6096386597f89a9f37b494c152175f33dee68c4791c64f428d8701b662ac335c068143888caa09af21400e414143a532ac9751fcb5d6396be3495ca6b0f3d72a3129f7f0e4f69270fe2cf59a;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha880b7e058eb8af5254d23cdcf4d7a3b8ac7968b0e2e07ec974bda0ee30450c91ea9f158c9cf4130315c80b9cf2a545749106b996060ce8e4195c384f6c482d94e23aef75409172cdac8655ba9b1b9ad5d519921abc5ac159597f14aca904223201fcd12d6a680c8db;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h14cc67eb866381b629024bcd96f53764444097b3ca603cb5b35567f3e2dceea265e84ee8692283bffece73bf7ae3cd2661251329f6d1fa109b8906eccc9ce95c1151a69245e70abaa23bfe1a70bf5d80c205f38576bb005c1a58f0a46e62673b98bc8e8685afcc342bb;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h133ee3fb9d92234fe40313b1dadb1d7dfeeded57fe967741684cbed667c4e9cca0502944a6555f4f180f5025ab95ef74e3210c8e32a9c434474cb02a76a3fa2a5ef1b63ae286cc5aace3226de1bdac17e57fdb09976f88580552f705767bfc5e0db3558b9c5f3fc3501;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf970369d5f0b4152a7be3eb7c99be70d2818819ddb650f90050c3f4d081d1c34d065b3e2d8ba73124008506b3a6bcace4dcda4215c297c121198383f5c30c0170fe8adf5247eb4de29f0aefd4a0974f4ecced8a90c01d488ca80049d8ec3a0aca9b06e6754fb796298;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f6035471826cc3400513f42765c61fc4d1ff5bf8e1f3dfb7fdd6afc887acf72d386919d041a66196f7beee386a3e130f4bab9a86ccabc017d27fb3a7591949a6d3b7b18d034be1ea2355d0234e71bbde141144d72d97afea81c6bcbe7137b6857a71f063c01573fa5e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h12ef0a437eb0d5d10e1f55567e418f5383b2576ff4679ee8c38e5e65c02770aa8e7ac2a35668ece9ce45f1a91bff7adb853b766480232b1441c1757598c3caa8fe371fd44a266c319582a1052aa476a73d77ad162e088aa5bed8726eef22bfaa4de5c730f2706770e7f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a8f5f089d1c23aa90f12fecc17497c0708c6b0074c578822ceb700022374ff21b1d21ca1326a45d08022bbc7952860ea816b6f05ae0c4de9f7321ba99f0b8dbbbd02db901de4f5097535a308f884b64dab75bb1c54f8d8e14cde35b33a74654e8ab1b82ae542b528ae;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1831e91f01bd1cd6e57b945fb6bfcd94d4d0092437c21a02950daa49f10e1ef22e4c6c735feef9603be3cf7d2bb4dca94bc70fb2cbdf301c346294c2c10f2bd302ffac56ee8545b2dbe6a99a0a8c4e56bcd7f3ef6d6375230dee1238bbb2dd475bd19811958e82bd18b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ff2d5c76fb3d64b1180b9cd9d415534720d1a4eb3694ebe622c4b4c33eef20948daafd3caae14ad9e912d2d83306c57f4ccf8789aeaf5535d8435b8e848d2a2ff85e724b26243f66dc81eca00c55d3510114f04b2c093c015118b192f89c32d361fafab234c37218fe;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e35c4354b65721941e898e02c1bde45454efbefd0ff5ac9a2c4bcbfa74a2646abd14dde8eff6a1ff4f54d61d4f955955078aaa5e549e040a8ace9b1be2983b309cc53ccbee829ef77bd1db291a83ffa30e203fb2acd96b7fed813287f24ed0c008320a3b32e3c973e4;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h67fa8f31833c1ac5fd3b63364254c1366b06584fd19cba60eb1e99cffa0ab1b4b6b4e14a037a70ac3c6842820f4b0f90df2d3abccf55ad674bc50cd74e01649d76bca3ce419b1d011576e50a586831d0dc8614fad56114ea133d4b82db9f3a81404320a851951bea43;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h15ee85243e182da675e3c3bb75dc73ea8a82a74654552177163b8108a41ca775dd735f30ac177030c7406f283e29111255cdcb5ee6cee8c96f01832140821a4849d5714e55927864b6f5221e9215b2c190a87d8c9cea821ffd8ecc2d878a914f2adeb366ae3bddd66a4;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h18eb350d97b17632104596a245d80b991b7bf35874e834e19ac465059fbea8aefe4f5a6141bf7bcb4c1c3749154fae73c20f312ba9d41cf1b1845bfc2c6c4b845bf10c3a72ee64526e9f7f3ce858ed9b22e46ba19e552b9d8fad7786b5e27e6aa660e8a5b0847f579c1;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h642faefdfca4d252d323c45288e5a8e7521dfe8d0eab912a557d61e05166f5e7edbfa0168ace5fcf51566ce796d144bd2241f76970aa5a130ac04f9e763a004722d24214ef0f7dd96076f0fc8c3df419913eacd3a41c304a80d6893501a8d5354c41e152023d4fb575;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h9000a663306ece571f84a30a70205522503911d46e558527c3efde4af1bfc3db3e0100062492d08ed00966e36b3cac30889cec3266e87a9c3434959421ce62818518029669c484792c3b47256b6e828670cf22b5c973b7d6ecc4a9a79a0436ea4c5bf334e832b5f93f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ba1a58d8d00bb3103f89160722d1cf43ca767f7337a8057ef7a93efd05fbe0de7afcd648fcd90814b745c506303abbc97774cfbef45f26ba50641a63b694673094777fabd9fb73f4d7c7b7441d64484574b788320099ff45c2e1ac6ea204763c26ecdeda015a97e96e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hfdf5212378cde12030180ea85d35a254969683f53fc472fc5197382558513236ebc6a8aaa3072477f8ad45936e6ab6b2e0b59f3a0ffd696947ca99f144e9e3dd58bcf4c4367f85890eb8219ad6e3bdf025e7cd6f07a4119a5e069bf352fad639c9ec923df4549c59a2;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h17758b77a63eb3bba79b15466ef94a12039f7150de5f93ac522cc8e2bcbada602f4088494539725aa3fbefb0627f9ccd171f58d16646491e6a646e48bb51c5fe96a2b8b393723576ff8a93d570fb63310dcbdeb732ec7abaf3ee5a1ebb0c4068722540e7d5439b52e28;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c82ca7871c2ea795da3f38ddb0bcfd99ec28dc10d9a3dffbe47e8ce9f217e82c90ace2d654770cffa57043d55c151f4f9a423e578b2d765b40065d44373c6e59d23844ba35326216b111c273f82ff43e9f968170959aebb1426994bb10e266ecc69dad0fa6c1fb972b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h655a8a9c687ebf0ca33c1d83333704e12a728b5055e77f606cf7d8a3b1d7af2f89c1a46191526338e8bc53052275685056af30ceef13aec2205b78bd99dff83270635e5f5668815926ae767af35ec05acad990babec90ff5eb544dcac6c06d131db9ccafe25dd729c3;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h40bd8db3358aa58c539b44acff3b38c85e769c3e0f589bad7c1cedd3f1df286267a0144f5f30df62048da1f0743362404343f8853c3f62c1cfccd38f1d6175a6c472990b58cf2365b31e3fb91dd0c933c954d64093fb2d29ab8761379b34224f66d2346735a90d3e0b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1fed92f9590adf4fce51838ee2fa5661fc77f868e0176cc253c2281355c4c4e29a42484004c80323dc1cbf8546f57d8d1f4eb3515dc581d3b84436d1af60d4377250b64c9074f7d1e64f961bd880a7a2092cd7112fb359dcac0509ed13cb6da319436334d7b37303425;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h9e0bf73abfe9d11d03cc34542130b31a7f9cfe03aaeefb97db0019863642487d5714646b046d4e6be3adb75a957b2cf965c2518ffccce3127c6b3416d0e85b7053134f778fadd8042ebbd7027e1f0b63c34e687c3ccac9435ba6f55137bcf480d7732aab2a480171b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h14c16c8a526e25e5c2b57665d2bbc40737d9b4923d6cbea8820697e0efc9f7f8e02a96d7f9cd13034fe88b5e67a761db417da3c45e25dbaec7f8bccbc1ce36ab492bac97531fe4be9104f7ac178a7bf76276f07ea39b3b2fb2161aa4caa075bc8b7d52e4b2fa01e48fe;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h859e75723e40dfada7f8de0e2b6533a9a769102116908860e0ae9c793c22d70885778b21320eda12b75f3235ad80157b44e0130ee57819c46b7a0d57109b0e5536f24fb0a001a1c20c3dbe6fbad6f3b5fc4eacd9d84daced56b4d93e342e8197001accb96a4eabf789;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1749760374f23e2efd1efb4d53e0d961f8fc71c3bb2a5116b26bd7ded2b39cae54ae9e06c1b8f79cb5a9a048e6d9313ed745d77015a297c7fd56a55e96b1afc38656906ab5f9b5ef3730dc27fe7aaf11ec44c4285453307036195bf11065eb4daa08a11180a2caaa807;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h7573c902bd4450a8b7e21096a1475fed0e2080f60942700081bed0003962ce48d1c2efe6bddea550633d43a0c1bb6af9d575cc70b68958d9791c7414d92d4451e8f4f47737ff3fda21d60d92658f55528dc4aa285b232716f3f1b26964080aec2692cea161de5ccc04;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1532c5db662a49a2b60abd7e13806e9fbcdc7c311f2b6e1bddcb0cae08255318bd8b46f9b8335a47ec9c3d998d5b2e0f6a401a591c32faa09c0db30f308b11d5a642a7d6d0f7442098f6575e5263e7affbbf510d11c58568133f9e2cb58eeadee77fedd49a1b4795197;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h90f01d7f9b6fead9e38f1a5e1dcd8b8c5b6d0ba36579ebc55d7d406249b7d43f2872169c027840b2b8de932f16b77a9ee1768b861e432d5fb85cc6aaeaa694fecae09d7e353da88549d8607175adeeb24791f6240b13fae7280999b8af52d16ee86481823688b2bcc5;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f5a06c764d6d495c2aa7e0b1fd5e5826c7fb8af0ba5f76be501838fe6eefcb85749dbb3780bcaadc190748ddc6a80e9024292f8b7e2ac75ee6e52d5a6a773b0edbcf5e4857c55adcd4ff350b281f88d7e82789745be8f2d9c5de509dd5b7dd9fc66c3f6274d4c09589;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h177d1f9dc9b1c8c74b4e2a4f16f1500e685312df9a5be8ea08f7c7b4991c65cfe7f043f7d4359e7dbc376a6750419cca1edd0a10a08d0f7ca00f3441af0c9eb8074d6395509e91f248160903e1ec13725be8f91e318cf8bc2c68d8e547e36e2eec2e2f7bd6ead1da4e2;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h2ccdfd4addb41e19545dc857d654bcdfe827095495831749c48c9c7b720952cf0241bfb001259150ef0a10249ceba30eda44e215805423d48d1758453828ca227de13913f8d0cb0d73168da0c115f1e85c6550f35c5c23732b2f3a59f37f2d19774878e4fbe9322863;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h78fa82fafe9b8a36898ed44d5004c571d5966f5d8b8a0afd1f7d38cb1c939118bd3a778de969c67f280544cb094521e711864022ead58f621b2a7e86e4978dba9508b268f2213fdab5d54f6d4fe6222b47f595f1af06dcc15d3e5e0437295f9d4a67356894183b5133;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc8f36ba8924020fe4f8ed50c5f333c45a1abce0db22f9f20fe377e8fe99bd1b8505e8df6ddc7c3f7923a38637dcc0cad6ea27df0e8abaf11da6f347bc3980f3e97c9d4685ed0debbb6c5b42253fefa63755a170d75b5bdfe567a81d838c3fc26c5d7765c7037b53b19;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd20335ac9220da1018f5b49738ccc87eec99720deb2f34481683dfb336d83013c7304615c498a29491e40591e541e2feb790f0d5f05b85b8c89d322aa09685d7809d8d9f4600fd197205a9e4dbf8aed8b3365520536ee8b7a2edc7a43e40f57508149f37e03f11c8ae;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d3dd8840fd28e69b59bb95ba1161fbf4cb929552aac0f5e65eda67c290106162c0fe3485d406a90f7afa516a515b3ca24565bc3077cc78960f835a1ed1df1a5d72a524c6585b30b3a5441c486840cf88189e9d7c0d3a901bd7ddbeffad3e7aeac911d04a62a14c4680;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hfc469079f738a53f852b0bd525fc95054e0f3485e2d124eb5c7aa1b08bc64eda47b636318d3d184b5c03760a3258748a39582f6115b81ef08e45b7596b318acde4fd04b5708eeb80df1b88ffee4c1799e4404f473ef662fe97c49c91866dda848ff052b44876890202;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h47b503c2b8b58886aebde7c724dbdbade771d030fdfadb8c89b24b24246104841c9cf7224b6a1417d385fa6ab53d9659e52d8c8ca675e3568cad686efed3cc0bb6e78d071e499ea62d599c60e06641539ffe7d593ace4633c06711c8300c85bed0035ad56fdfe2a675;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd1417c20cb81684b7d8c669340b82052b653c28de4eb2da2b26f4f00ae7a3b6dd02e146dc7d773c2f8d3594aa7345f9cb9ff49bb05ce896f28ba9c43b57599243928328ef853ce2df9e7f85282a98b471021d53301dfd0ecb3b4fd7866b5c5b8adc1582f9295cde92e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1bf6c0b3fd45dabe9c7780d2f6fadeb1507859b7fcca535fd128cda04966c6ecb846b67eee77a4b656cd9c696b93eedf8c5e3ebe5a5a96f4db4254f8d90971b9cac7333e861b25ad5737ef0ac9d1a8112e0d210f2a2062722b25dbe231b899acdeb8521605a641d0650;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h83608f5bc0c71596a2f1a321a2691b843dc297702e433ee48f248dc706fa36171e6836b85d9ac6765b958b676a3e52d9772e378d2cc4d9e941ba8f0ead97601ebbff9c482967dafe63db59e10665e9928349e11fd05536322c1e89eae11a54b69a9d5ce3c2e2ec0b7e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h958d5d16cf74ae26a86a3df201c7f02f1beb77b4b4467cf20808d0f80517fe9dd32efe84430a74131636531614cb9be3755fc1ae3d7d15dd4c330025b6dde77e5e9ee2ab65c9b7289dcd9c951a13c2ef24a1d5df37bad1e0def8c5c6c5a704dd89eeaa854197f3c598;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e4aa87de7712e210ac2e0191386b31a62492910d5ba2224d03bacc348fa08b11bfa11ffe118d790b7387057955d7b3ba96bd284a133a75b4efd7aef51eb8f05e23bcb96a44991941f8b198f499142b2e3d7f0165f25d3c8a80c6e7afe2de2b6e70ac8828f0b3794ef7;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h63d2634737b34c5151894d0b746725076b9fcf0b0231a227adb57ee15395af636f2124f486c427abafa7b83e9779107bfbb50e626d572f282c4ee22d34a2001c095fc10b0d30c34ee44e1f813ee65003f4aef70964f1ef52f50b92e26183fdc92dde4c7bd6bca6b738;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h12d9adb572e55c226dfa7ed0218aa7ae0cd8245688a66747e0e79e256de2bcd1e281a5749d00d0bff929c285b26f253d1a2a5608b58fd2ec8a5a0d0e752bf47c02be3bf9578ce8b395590a17487a416ec83a2f99d8ee098d95f8c7870849bc21c022e95051ed23c94e7;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1deb555f3ea2df0fc9a0740248b7c41819dbf8ed3731128949414e631618a9c43ffff0eeeeb3b9be565f4130fca6f7a08aa9e538f44c94c10c8fcc09a043affb66028bb96b7550a1121ac90b44babec11ebb031816d77643c1017f9ef25b7abbc167c8d12fbc2d04c34;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h8f6008535c3e96e3a12d42e42ff9465aef8dc10b0cfb6412a90121009f30e9a03402608fcdb15a15e308bcca97d0b89426311a6bbf9470e9de4da4a143740a6f903dc2fdfa275b0db0ce7c19fcca4ade71a5319efa2b780c95a6503c0e7ac176dc3b585e41b5a77692;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h13e4a8b208026a803f4942901985fdc95cf9bb18e9f7ab80a30d06a59f69fc5740fb0286e59d7d9e944ba95180592f4a770eed7bf67ac8080bcfbd67c81b50aafa544bfdb80113be242eee06e33b9601bbe92b7788523c6054666eac3e01c122fa4ac078fa490bc21ce;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h11a5a55e71be9d9c69869fa57ad44754f6dc96deb63de97a02b69abfb59c705feaed6ec0e85c924b2b8be53afe9e75b9148d66f256cc6bb6965d2b14f178e685bd27c53735b54695a25502d26ddfa2f014eb21ad8799cc941ea34c1aa421f1534325f808124f7f55d82;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1fbc6913bef3063e6402d9a90bce583aaf9b6005c2e0b81b577baf9c06f0f02b329dccfeba10de30ba8839807fa9ab8a76f9962ba8c73231a2fe50f2f29589cf2e3dde172aac3cdfaf0670bdbb054f36accff84c51141d0177364b2e7f0c580cebde4f888689f0d3b28;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e7a82f7ce4ad3fb44687125f1476bcd2d6c3af5a06b1b2567418293bddc9ecd0cdc8a59918d3485eceac86802a534ab8d9f66539afae60607d3d8468edb4d4378f49d1003ac1ccd98af72753a6b437d0eb694ebd8536f33f8381b173634e57336466ff47c6e6e8ca6b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hfafc4f99fd3a0b476f2cf8d7f2ecfb4d8d0ba124eff0189c70f46824a52c157cb2462af4c2db5db08fd757242489eeef7f246a30fc00d27f588f3cd8d55b97956f1a82f5e3648742c5ee83439193dc76b1639cfe615d9a10ef1ab1f2aae1c52ef9c9ba9acbefd4f70b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha7bb6df3902e22b7df5316fb1eca0d12ad7b393e9d8008eaa6ed61bc7eb3e1a2860efd37912c22f41a6824c6fa8212c6632a0c151aaa41c38accb8e5a38fbfe1fa8814db3cfbd37fcd8b1ca1310a5ca9f17ef4aa6e5e3ac4decd879b35947d5f60fe494430cb7f8f3b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd3c03a4b76f38abdc2937059fbf0f42696960b263fee1a7dacc578f9e36087931d7ae7ab99d7a1d0ab5e94a28f6f9f3d31f41d6f6b40534319d14fbf06f73aec082a5ad30708cd71a69b43f7a390048aa6731530a836fe97e011f8f755631d4a65d845bdd7bc358ee0;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h7a15ac6e3dd37779434fb56853e724b6b6355e82988e47d7ef1d960489d31346c4dbbcaa584ca1b1ebf2be97d86792db4cb5d194f7215ee397771e42993054b08d3ad295417aa74c8032c9310e553359346f143e18615d0536e43a06d6e1990ef955b367396fee47f8;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc948f68c7384e2abfcba2e68afca381af374388ae3b1b3c4a20e5ad086d0247ca474365e831fa677d82b49f312e4d51b983155153528f78c45a9e43d93539562a75f2ee052ac5c6fac65b2f01fb22705bb95a1c2f54a7f9d12bdd5956ca374663a24ba3cc532fc2ae8;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f769c9c5dc39da0e1ba3c99c6c1b4d11b233f9bde62771a91f9a9d6a0fc770d74d9f7775a932adf45fe579f8feb4d745288a4c83f6eb68bde21175473ad9bac0edbed78e021f87255de744905a2be40833a5465ad206277f9b2014cffe71be2324af504b955062981e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf01f634763c83eae65d1123d01f8111df753521e77df088aff05f2527d57cba4c9036bd3d342b2bd32c4de9e49c7ad0204dbcfae8202fd42d60479bfb6611c78bcb95dfdd742c3bc65cab578483c989763f755d4c1f4c943e61789f5258270079d68c5bd07a85086ae;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf1fea05332840f2c825b291ca74cb9c9cd8c7b62e8c95fc25063f5aa04c721ef3feff42b5ecc952b901be7454e62b2a7258a4855c3e4bf25af2d3a63678522896f8dc9a0b2077dee4e052a1f7fba1007caa05f45e79561ce44703e2c706f3db48713a091dcda5c314b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1af809adc3b7f698e2646b2978b68d6dd6dc2a3a35f8f16f2b1b13c6ef18055aeae6132ed673512251cb08974cac73e8a0e552bd975162e0cbe411a882d4645f9fe315b6899713734e9d9fcd69bef7ce8aaf2d83f5c7fd0b2b5aafd97f24f8685d10fbb389bc78cdcc1;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h163caa6736f73eb37b3037de22ae774f87b15b22c8725bc449850f2e8f6f3232a15ba0c4bb8f6b8f03ca8841407c2b1a987fbc13da5afeba0e8e825c41d8f2fdd372c35ad01caf1293aff19ece7c00da00e2362e3b01b9e621fd5d3d6f7b8c7455f07735c394b865f7f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hce92045c37c2277825b92c5952f1e687cd9e3b669fcf1213a0ea389ccf6a5340d747315ff68414be02f1cc0f55410f2f89d1ba543eb957a4c4045649a7fc9d6b4b4da145b2f231dbd32c3cdb9b338ce1ce1d22056055c9a982b18cad5d00b13e2447f4964d817cf973;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d2a3dd77e147b9ea4038ed4f899494c0b6b3f1542d93a676a74a4d4e92c5c398208e7bb0cbd601ac199da559f9446aa8fb74b003f0b93387bd55047c585ef009bdfd67d073772391110b8aeedb75f166345e5a49b4897f7380c1d00ac65ed203ae6a32a4edc9bb5546;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h19f9d1b8f64aec4aad41455cfcb8131afc102935007a4d0e15f5bd4d87efedd9df3b38b08a282a57f6c58f90a7da1d183ef4ed481312cf1c59f5b8ba99295e21eb08f5fda126b4f765aa01a666314006e704effd150dfaadd568c9ca3355f15d278feb421f3de13029;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h12498907baf2b97580f842a637584c9b462793a549581fb882125476c4c2f4213829b5bee91ff6488a7569751a47c49abaf83373717d6633484477f7bdb12a7a6b0b17e298cb3b5f8c02a2d0fa677a5ea62ca7f3037cc208c51ac899ef86455b3efeefbd48d0aa47b1;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h21805ad961dbecb8bf3548532cb902485cb4b80c8083e9e80ea95123eca530ae65f32dba7aca3d50ac3cf8ccd13e41d857df1145ab8ec607f1aa2a9793cdf59f52b1967bf147e5025f95c14a46bdcc7c2c080ba71af9513ba51311639d2b80362801c9152a3f84ce41;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he52766fe6f64a5cc2b353b20ae6b47e3c538fe04a41ff4da122511b6d936bcedad4e3e543d68b4ef8e6712e798c4d0e307f68d6c890804fa3af36017fecb8e68f7691443e5a5ee4d3642b5c470e14782a8445d991fedc9ea67c1375e57f55e747098afcc534a1c9511;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h122bec590d58bf024e455f8592b28e8f8044dad5f53e5479058a953c58c3095efd37cf13b031116502e9872d5c0393cd2c7964c6246c60584aac8b6db8396de21ab95a95fef2980d3a262ce0403cff752e04c189a694a6383dc1dbfa160202bcf97bf14595f9772ff84;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h19f98f312ed5c73b884a6fa9194fc49ec08954eaae4ca73195c38dda46964321c3b311cdf4bc125108a80b0fc06b748db55283a045464318341e5693c2f2473948d442edefb507758f19151118c0856c5444afb591b9a2a711413f794ef4ace1bcf1c9c0a25c9a1191e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b96b86d4dd1b5f505b45104359c4856aa1165078f2042f0280553fd5b908cb766d1357867f4c2cebbbbca0606fefc27ec83d3495701f0234bb9a669b8f293c1be34dfdbef1f00c7b1f6f891fc18fdb0c3aa1439e2eceafec2e1f06738a945c9cb6ea90ec61c514257c;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h46e980c9c80d6c23f7498c58bfdc48e0e5367b452822e4509b4e07d0d9d115b4f511ed714479f037146badeab186d42a94e2d24fa396d561b317e0a027a1f90b219d6e29a18065446fc8412fc2603fabc42d4a05e95d89e545e6dfc5218ce4d16e4ae2923c1917fab5;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h119378cc44f0bf993b93f25ae0165e91b685586c52b9139c2c990e21b77a60cb71fea02ad622e5c63e16cccf438e599befba93304bb319e1a69177c018181cedb345455b63a3a05e78c063801da5abb348f54587bc5604429c91f134feb3490ae6979227e92a1511fba;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ef8f1191ea34780e856da3ec3e4ec9a4947b6f2c3818a285468d029493c21dc9aec29d28110f972bffb31311da5ed23a6956088844dcfdc759bde5c65be77fc69086a15eb76696dace5ebefcda2b6912b7961b89ca438e5c62b47425f9d8d6058dbd8153c6767d4648;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'heb21315e413eb7adeb4303b46a69b6faf11b65b4ec55d52758e0d99f2046bf235cb6cfc9f4596d7051b22299e4839247e3087118119f4be27e8259b06ae6ff495a0dad4c868923fc56876ee06299ce4bc839f535d864a59cd8e843e13c77a37003bc78f2b4ee586d49;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ba42c75f3c448f0c6c6c12e2da0f2d45862079eb7b1257e5370811f5eabbdf5bc3b4501287973b6d8267bcbdeab497b58c14d90f35f4968546207a6dfbb3e4f2ad6de05538640f9aff81668a423aaace0679a16491fdd875771261e45665a9fd37fc28694b167b402e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10614d7d2a8e6ffc5112c9ec4d4ce42a0276ad16739b569fe7c3c7fff0a5ac5583ae060f1835df2ccf5a43b770176f121910e18b53d4cfa188dc7e97702f137fb4dcf5061f938b022e881b8a862aa58a1a9512c8705dbabe0479598a81c527804ac102e466de60136d4;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ab29968b8cea5771c0b28da84c18a626397447d99f07b85c4ba337f73df58a068b76b426ce1941a4844aff3ccffa7abc09a7ef492c343cda015c401c91fed0a22cef808b43f3a2e09b19163b9f9fe4ec7ea1a3adc9f2ac45132d6fc0c0951ba3702aad816448668e67;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h8305c3209a053e365ff6bbef70fb5c53aa659d68c3a0b7d90b5cc532082b16a237af23be448407ecc8cf141b042edcb53a48a699dbc4b51e43b866b6551c1bd0607cf29c7ca033aa5280550223e452e2e1531b0804f0dd9cedfa1898ee4c8511e3b2e603cb2d7e1a5;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h118518a9b79dce9a856c387e541cc016b97433cbd2d0439ec4f51f929b2ee350577c3fab8fd55239ade91ff323e7b4cb7a2e27398dc69b683df3db523a8c8b5468966e6844930d757ac88b6b3f0cb4c273af473f90ee29161e0d19131495514943461179770d5bcacec;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h683f6e6763eddff588e492388c39f5782c383e09a0e303d0ffd00f3041b04224bdc4ed09d82c4637957def0f3269bb6b721ed9e87e6391d00aae983f0acd0def7f0b5244e1abc5f41a58ffca61ca87232a0aae7fcbabc504fad37071ca9672f82eaeb4ecb27cdb4839;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1827707f361da6225c9d1452fbda175376be784af8a812603b0c56f26a704b2635260bea521f39427a08f8a5ff5376c111c713ee82e970d4814cf301c6d4da1f8d499d48e707d3ed04e514dc8567319f4ba4d05b160d14df3e5872eabfc00ccbdaddd5c28daafb0ab04;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hdbb019b26d0d7934d6b302d64d75c7d9153f41bdee37f77e77d69d626ebeadf2a16371091faaa20199d4b264b8a22e6320dcb5fa46166e67c46f7c056a4d6e2ea654e478a6030af40656cb6bbe60461c4e8f3f75af9740acdeff6ec77311f4420b1674f297328d6da9;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h357cfd88857327c1ef1fb43bbbd104b4114cc655b52c20f39db96c69a0cd4e232c5aa9bba296e3cc0bca8c8dbfd4dec308148ea140cecd1318e3f49a93f11fb896887aa5ff6dd1e42774b6dae291e38fa66daa5eb382e6b824465abb89ab74ec0cad6b9223468c025e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a5f50bdabfbb1e55c903d9af2b37f41686aae8eee0cf509b7843bbf8c8de8869e8287e38ccc80ee293537d06ef1a97bf58479810816ea832ae8ec011890bf4c322faddb10ecc5b86d88a79d7d056f1732d74251926c7d10d483d815cdea11752aeb90f5d7e1dd2967c;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h4275f2ded41c3d5dd7c5c37c8573ad07e73790fb8e0c3d902326eeb459c63d327a7358820ec1ea34b8ced21382484b2cc1741927e409ae3414a614edb8c7736811bae86f6c58fc829306f6645d4ecab65fa079e2b8b42de590f863a38f05c132388a592d01f51e9d0d;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d050fc16b8aaaf4de59f383400cef2d4c7ed6979ec898213e5e4bc414d38624fd7e9b3835bfcdec8a2d73e290f7e30222bdf1b399b1719724d84df42e94adb2cd1051b641e5ffbbd0cfe73d809ac045a90bfefa0490206e5ff596744ee74c2e96216ef90154b0f6f6d;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1203729c8186aef5fda8980c47df96ffaf85a6ffca234e4d2e0f072b6314229c05a8148633b407efcc58085d6b310c37a1b51efaba96fdb6dd7e5c4dbd765b887ccd74a3248eb8e9f5ca96836d4831aa63a5888dd32119aff3702568a9adc6eb765e0ddb1db5002ec71;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1738e45f3320b6ae96a82f5e944e446887696e9a13d82f0c6ef1a9ab207da9d7ec3881c092dfd8597d8aa65b59f79f8caf03d19a372c77a9dc993bf84f324271581c96345ea26d28fac872696335db0ee01f0d5371bc8b74b515275c408bc1076add210b8dffae7ae05;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h190cbd1f1248c850103cc08fadee84042589ffad39dfd496d0cce7fb170b9a917b286d257866d164c2c89bc9ae672ea98aacc41796cd27cc162be8a42884c9de1f9c862e1232ec8dd9ce5ec00c6d72490a1c9125bde4cbaaf3722dddcb8805899bd8af46335c5834e65;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hde1bc1b708a5e010eb8b53be74bd94b8eeb3be02f9344c637418648f1f5fe19cabf84ec7405c388ad8eeaf41a52a33a35f83556999e0cf95fd34c438449ef925080d6004a231f4ae92cc65e8201dd314f62224120d3465dffa0f61d1d5d19748c9c470df82ee75fdc1;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10d469e78b4a0ef0b672f84ede13ed1767707e08fd1d3e94e5e42ce121aa12175b9bfdf6efebf95d9450f4e280229f6071fc2fa9f085f36adc1fbcba014449d25aa90a11a557d4c9237c0d265d00f48a5fd2b1d52bc32840468afd272df9d853df66a61a46b9ff36802;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf4d25606793463d5820101d4b001c30c308ba19abf7d16a2cb5baa96e78fb34b12e3c5cdaf8fc46828670bf850cb3c42d307327c0e2e123208569ba65ef81a07533356100e052184ba2b3866c55edefbda7a76fd358d95ffda0203bb614db4b24434a66c2187631b2c;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h12a2a6642676b42db51a98fd870b0597ee9ab843aaf8995a437af1f36721ad51bdca5d6584d655f1e0a59b6f27ff72e98b6bf880639058a4c6aeb2b5b96bbdd4b5d3c21e87b962e141b6445227d8c5ade1b6464c4b4597ee01f04ceb48d5f5f4cab0b4f9cdb95c5273;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h164a188a3530275c6911702355f341c23b05bca633a886bc54b324d9907f1d1ed6bc355b188859551f3c30fdcd4cda4bede3cba96e76d1ce115118478ef72c022b780f5d919ebf42add0df85afb7e30a5e83016c1daed0c52a834ebaf9d9703c0f9cc15cc1bfefa9cae;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1cf0ddb35040c0c3f5c1a27e962077eebf05ab8c14edc1472029b3147daff79cee900fa358da64c75b0c96adcd7f79aed3f4566888cc3bb23daab0e44560ea5fa78f2dffadb9582d18f14ef286a7b431179034675235fe4539d2045b726f851ac1c7a7e29bd62c8cdcb;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h12125ce280768006d1f4994250cbdb0f098984ebd168bfe831f34f8fcdfa21c22cd7eab119c2195295b5e8e0a13f0653ff812f4e775aeead72d9f141157ae6970151f510bacf86539c362f48dc890417de06c55e9d6052294f6912ab5651ef3639b9a33835aab1bcfc5;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h16608dbd3f79a1350ac9d4e25be177973b288f730a37918e60f4c85e1b27cbb05948bc79ca5e2f33b64c236a195abfae492816bad630ce9f51302b8f92fdef8277ebca4c6724e1cf98a3df3a27715afe6128c773fae0858e86d526f9715e99f8e3d56f791bb536d9ea4;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h14d4b189a541f3d78115cff4b32517b85c8e03c8b020d89b45ca405da029e88215ff12138843f5fe27140779d838fae3b126f4174512a8e3819b7dc2eece3e728a8008f94b0795e96b8d71e1614abbbb335ef80591404c4cd87fc617132a9fadc10fd8edb9af38269d;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e27fc131a62df5715083b70d27f36ccaa528a9cfc0181817bb865db4d1d5b9a9881bed4dc3481dd0b08fbf4f27f7b52ee31b24ff5c940bd2c9e81a53cccf0d9e8f623c2db3c4d7a31d282da28bb630212dacc3b7b40dfc0bdded1f1a396338f3483c857b47e51112ef;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h17a222c17c6d8294bb7a6e6dee3ede9dea18642df9815bc86c9293da08f07e75f989d6c0b20169fea04ee57d6b80f2dbfe016d5744ce274cca898b389b3a65165cd075b38b553e7a62115bf0ea529a5f7027701507a45a99e415aa7b22dbf9707cd8d2544e8dee7e650;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h19db57c7d2453e5a9550dfe571bcd402994370b35d46cb82751b9bfa7cdfac2f6744010b81cc3e42c4307c317f3393e62ec09653121f7dddf155d2856f96877b2949e4552708419bf584ab509860445fa1d98d775762e9e3d11f6104be3a184014c564af71e88d48508;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h37ff844002413c951ad06d4763120be02d37fab9b26d8bea09e823d0157e6d5706b81b6c0723650884ccad6d11b0db2063bf91175a80b0d0819ee27ea5b88f72b081fc3e537af0b5b8f6c943049922e6879d3657008a1fa42eb4ea7cf23a0c7a39375609549e352b64;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h148f4c58a3db78cf691a7b9a9c6af2ca15472469215406e98570e5ab921340e05cd2be34ffdb7ed63ad0fd676787ede2132ff97dea3a04ab4d5590795e21af53a9529f203f40c7ae49ca555c7db16ebd6b74c5ebde6a3c946c98ffef9bb3d7e240d70a84687b2b99a72;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b30858612040fb35732df2e5a8102ff6b3de6483d74b721f682c85351f2bdb5f6d15485572d8f128d50f5238d3a411b15651aceba6f1b1cb6068231d8159ef8aabd6f7f9dad119c1456db2aaf05c4e24ff9042ba9467292a143e8fa56ed4c353e277f13ce85d1eb275;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h293bae7180312d28f09bd0666ed1d4dba72766d55967955fa6dd1316ecdd18f25f827b9a49cd871676b04502dee36c52ac9fa119a862625140c225edbe585670f9be481944fcf26853098bfdbfaf55901d983dff5b22450f7995473dda2ceb8292478332662689d105;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h3abe0a7f1149579806a63988f180be9471517d9aa1d3d80fc07626684d239b87c311d482847069fdab49554e27ad82bfceb8fab70902bbecbdf03d370ed00f8c64c5c7c27c0a4a6130f0be877ffa5622c3f94daed18d8b964f9f1060c8dc6a33ff4c2bc5c7554b0133;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1887c6a4f1e48b86bbaf1b0ab85b97446cb765aff8c7acef2fcb2b540de4dee3f0b4e5f5089675b36cef07dab6e20797a7e8e9266d334bde3264ebbff7b7a3cd02e2264080a0fb35bf89251b7ae66662ba9860c03e121b658d8c2fd0be54ca0d7ce3d107fb5cbdb605b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he597b2054fd4bf8d1b1b590951a419596309ae96d4a4820220a487dfe68b991d4f5eed21e8965eb93f88f49cfcb9f8855065052522e0382d0e36d5ac1f91705f0e0bd1c9749db5db7cc764eb12ea83691dfb534eb660321abd328e651940774826892eaef3c3e7fd5d;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h12ba06bc7ce78e68c33180a6846eb1d5ed2d4cdeb5478411f5522b737372da0a0592192f6038043e18d06d9dad35f012e71a8962116d86f4972c6b81f74cf145a2111e4693d2b116851eb81e2cf1410bd8b5dcf36565e58e78b69cd773a9d6acd7541dcb0c4148ed10c;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h173463bf3951b9014964aadcf452ae1cc60def480c5f4e32d6531bfb61b5daf16ca86104b14584a9dbefa8490732ac75dde51242b3e2559d59deef1e59d42e431aa89d02c5081b783e0e1a0e2b78c25fd7ff4ef3562d67d17d96040f3efd0830239de19c13702b66452;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h117606738e32e829de510e0a5b5b3ffdadb80c19bff6a1bbdccd655aebdbe0cee26ef9580bb74a767848ff185dc8688b6de31db740a57943dea27652d6b260ef773e9ef63187bba16a1a94b6ee26a640aa71504627609987cdc4c1917d99d18a9d24c4a2e245283482a;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h3039d1b88444bd8b6279d636055ae41b817fe1a1c992d8ef166280b63022cbd0320e9ddce825b5b0dadfa2beb4e8fd205aa4414bf0fd218a8441e3f57c5ee426e2a6194662895a15dd1828642002a7252d6d498205baca017c95262ed774357e1940c7c433be5bbbbf;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h35a753c9b92e7535b5159cf5e215b81cbff784479973381d10be3b98bb53d6a5078b60de248f624d93d367a3d44d454b12e7b8159e42d1510312a69323b75944376f31371e0ecb50cb879ff2ce3eca3feda64d08f7121f39ad6d9610d9866f1fafa4ad273f1d8b8bf6;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e511e4e395614ff25a44c9ef5a2f84e2f5ae23f8ea4c7c1f2d44c5c22fc4bac8607eef115e1227cd9340c11a959d8c28cd7e094d5585b7825cdf3104c89f730877482c6d420acbe41e39c1594d80aa5044787c718d214cac543acf91356b11f6489ad3509b6c54974f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hdf7bd9eca6298376b34c3707f6f0b253a4c7cd89d03eaee2001a108ae33f3b3564003643a40f71b99222508668df853cdc77df2d69ec387fbc379eb3502a9288e450dd76a6d74212b063d1ab020fe2dc3593f8958ae5eb93e622783d5c69e68641bb7b7b96e765f916;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h134f0349c1ad45ac6ab8d91a36ba7ad453d58bcb18453abf66464fd59622fbcc0e5297d67c7134a789bf248f1b302611ebbcf4a7b1ac59cd4a5c0ca21f8fa3332f434d91e2fa7b61bd9ba2690204bc149c7c9f0ccd39d5fc409810b492980f3f20c2ead094ed611548e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h19b15ca6611efd1fa37ef184344379a50a30fb43e2a5ef69a0ab45195ef1b69776f05627f1ece232178d43f035631822b2b6907f618bdd0143aebec6d690abf8c3c9992117e41627edf5d0a17fe8c82ec17ab10a0a02bfba82c84298afab3d51fe263aa044d387d7521;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h9c8d315334bb2b785ca52a5f158fbba922061c72b70b5ae8abe4003bb646209b39fada3fd6d22d2346f1e5a6fcbb67ba021ce4181dd429c16046b6faa11a8033bafb3cb52b9207673b893d6ead4e16b03a2faefc12797fb033884c77122525997794e55468f390d759;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h77c986e9b78d65fc94f8df592bf2c829f1f25d43f68291c0ba6d384a52f8a3e50a00b22531f8677b332c23bee2f6782da0452799f0b3c1d96e949695f1048975b23c1c60630d1868f2fc2552231cd26afad6588c5dfdb20f43b9ca4e3138a71e196ec3b88ade19d65d;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h16aad05f849169767da21c8d5e169fa184492dde55117b7b432da74d480e7aef20c6a07d9fd0f52603df97aab606a297968beb933dd758cfecf3949ada2ce6bdf1c86c71c8ee60c022da90c225b39cf9862b86e1a6c4d8c3d02baec520c88c994d441352e87bd350823;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1319b45c7991395bc876dc267a1eeb0ecf7df2d53fb1ce332ff3d48ce3c2f20b8690af282ab0b879492992b22695435f47d06e78afb0a4c771d72003737dbe41bff08d4df8702a6178a0a77f76a471870086a1de5710ec9b4a837fc27fec65ba0076e25da6844c99433;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h351b2c51a851cd0cb4096164963887e84cbdcfbff3b234534332b34c0b2fbfd023c15855a99fe6e6b52c6b9f25a6fe42d641b16a0ac41e9ef331d5575f5f74cd62cb21ef5659d16710bc543c6f095bdd7082637b97d018b47e8318d5684386b5ef63edc69cc908722c;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d9d4f00ce1f9b3ca90623421566bc2304bc48dc87da3d8d92a6ef61d34ba3253844cb01200004107ce33098ee4a54e3eec5aa916ec4d751b05d8cd0837c4c61815ec6a66df4c648b238609d941757517dfb814740deba4d30cded8597749a5972e189e456293baf6;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h56eff60f9ea8668fb951fee95bf9a25cc9718e691b0d493dbe425323e2325e2720286a4b8f9ea4f585e78417a7952674de1709ec974ed7365b3a4874019f90909c340762d204eb6e27c6e3072071712013cee5a3361c3eff7a81800b5664639feae5dfc0ecdb8f69e6;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h9d04cd84bb7691ecb663d4f2fc3174c381f29d2995cb6ea53dc213244d88760c98624ac2cfc5aad8d0f25546de3522de425e10abb6defd09554c7501d423d3da45056a53212ebd2f7a8e1547c8286f8762749909b36ce657d8fe13e76c32a7a4918128ddcc2295c50c;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h4e0f80225a11958eea8306184a931397515224cd7927542ad628cef21b401c7e5c18b4ddc67155a00c1f019193ea5750e0ad7cd1051b653167be6dd020b5873fecd420dd31645b9e28124cd03e465a7cec12b590f2b9d43f93e7d633b65c48834e285ef6cdec8b7e13;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h15233fa269c99c9d36221fbdc3c30bd2688ec81c4b43d890b78f50868ea97ac9af5e7aba8f949959d53d11373845580df7a784a4322105c4c73904b092a46b5e6d1227f97efb116c1e7d22a4cbe8440fbe25d1ec9de859092905ca6e222c7ac234fcfb50bb2ff5005f0;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h85e7b1f0195e018c7b3ea157615dbaadb16882e4796e7c005b215dca3e284711df8f51eeb0fe499d4e767678cacfd6641e5883df4203143faf67d1ea32d71675d151284cc23a3f992463292f4fff7f2643aee2fe41ad5c29794110202a9bf2f456dfe5d6f1ee2d33fd;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h2ba898e63ac7cd7dc41dd91a442c340bfa930dd07151104051e57c1c431984480dfcaf321272446914c927b0604333986eb08bb2d8b40fcaa1a0502c77862c438b846249cad772e0bdbd75cbfb8a98c315c159906c1981231dd81642c6961064435a0fd4d7ade6391b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h103b9b6c594749fc6c0b4177285b53143989e25bf0040c7a761afcd2dbc0ccd2e20e3e040503e7d5a3664eceea273c29af6ecf247bc56384f74bf2587f32b74f8095a1e98b35a30b9513bdb7736d4ee474501712dee9b43c6fc4cd78d1d7745dfc19c171003e8d149e1;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h8db0eac51f7c834cfd61ed3c7d0e7321991fe970c6ad4358076fbb6e4a3fe193f850dca6e2eb748e3adb21bc67068d0457e50b0974eb070b8f039ee941a5d60f3a8f3906af8f8071f1aa9717bc531e4df14b9c57f569139059fe9f235ecd1296869115a575b3634702;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h8866ab81a8b411a1bd479c533ad1f167774b07d79daecec504f6fe620024029e92c11f8f6c4bad3a8ae549ae118ea16c197288e4d1b639d3e9919e8b18be2e4fec305f06f115881dc30c6837b41a8c51a8c801eb11b88b893998dc964bca44f8e7aafe7bc6d4f0bf44;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h177c32a8dab85781c763194317e5191f75173468fa0362afc0b3d71a2e9f90c46077194ee5900f302a4dd42285792d358fae5be6d5ae77bedd387e18e9a4a89fc32bb8376f023b369d2f4b26b15b2224c6bd7fa2a63c2b76d766d0af65a07f81c20661199052d272dfb;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1abb490206ea03f559ae065d598a6825b314a037539fdb850b4e1720abcdb56f0447b27098f40fc8b18f39fb3e0c7dc1708dca6d305e1fe73fbbe08d9ae0a9198082147a2663e92b7ca01c25ba7457ca927254c72522f3a5f551ed08e52c2a36cd1129ad7054f33f397;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb616ea0fff84f6a0f82f70043e5a215c8c1984cdf23a3efabb3a3c6198a0a828630958043a0d333bcb12955022088e5c1aaba88e3866eabb712c399223130d03d17d4056d1fd5f02bf63c459363a92e84778d02673635e10146457d8c6959a071f22bd76af2cd6f631;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h12c443a371ea38102358c587b06ee8658cb02c34e67cb84c3edbac8ed3781bf7b9414e1afcf92af9af0a1a05da8f28bf268a1874f4a040003a66f19cf8f31317fe184e071a62afdbf4468b5689d665dc2a1b1a1d65de2ca540a4b570bd0c16d278144936bf7fa0dcd3e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h827d120beecffce408b94236bccd386b248f671edfbe994051e1c9bd0e69a2b4c840a7f9472cb20cf94bf73ec6d5a5548440002844258d20c145613b3df095f6d032cd5a4c4f4beac0088de06ddea8a54be6d8cc041085161d0793ae774c04d3fd498b9a67cbf8e9e4;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb0fc4d681f58bef12544b534779cd72f973216a1a614c0e25f306a638136e64b29fe1ff73a7d686427e78e563c008a95f1cdba587b2d60b5adc52f54e768c95b0132638748483ee015e1ad9961cdacd6f7d66f128414ca0e607146ed1e35f4635f758b492bb87bf7fa;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h103783be4337be19db596a73ed86ab6fb0bf37497bb17488b6d12f14eeb1da3472b857d832b0994480b21ee74c55ad99e8b554a42674fd90ef5c607bad6ceb26b8f0985af03e2b190754afbe98c24b47ca03d355cd546a01eb11a5965ff5a19714643e6ade0e6d78063;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h19af0d472f278a5bea51c02c3bf257fef65cf90da6d4c7855822fe83326a4ae43c622aa8b301cc8d4027833f564d9cc5dca53e04f4fb97164de7174fa1dafd1b3543b7652b711e0ea080311802c32e0788c6e070466d45ccc7653e364ac2c6f708fa4794a8c152dac74;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha33553a575b104888fa29911fcab9b71c22b48b433c38d65f194dc3c595b86cb8a27cbb1b3a9eb82fb014d7bc2a05471d92a64797845e1117bf9cebd35344fa791659a8929227a4876f7e84f4c5b1504dc93658aa640126b6f03be5cce3be14e920276660032d91029;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h165c1b6549444c1aeb714d3c1ae129e3cccd9b0613109d804c0c624580fe95b0af61eaaffc1f48b169f10c31547bdc06f0db90b3222061a35267a4591c2d2f05d898669859e9824e57c0b38ebb9eabea24e2ab7b71de3fe3669aed878b0c086608aa8dd870e6c91b5e5;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h130d448eda4cd6bcf2252bd03a86854794babf36dfee385a343e92b29075dac7e60d40bc39cae1ae22b1ce869b1f451e60241591675f91107ce7e6705495a62e444b2589fc9ff475c6b9333bfd3929dddb6dc325523deb025d856efd3cf1445579348498d284356fabc;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb13510e832362db6ec3d8f8c1923fd28b6b7cf387c72960d9c314a82e4efa0375be5284a9aa91602b710da51080529182458348344fc96211b49ddc8db3448a7f97c1523c9f0475061a22d0139627441301a568aae182ef497ab06f9762c85cdd0dc2f150b6f01a23;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h3aa0e088b0cf864baac42be6854f431fe8fdb0ce11c0a9d97848cdbf6992b4abb317959bb71615f7770854ff90391055e42e3887f99e7d95b13ba8896b4e7615fb03e33b588c1b4aa25ef6686e010439b1f714fc7ebe7c34889529409394512c33cea04b43e4457796;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1af48ec3f488c40c8e5a50f401607182bed08329c3777a48f83001c77140d75154fb3ac410128eb3f6eea14567fc4a98859c16b569d664b58e7c83ea48969843ec6c4ee31ca582e2114c23d4df75c8816caaf0ac7d1bf8e56743f5fc9188c63777f002580c14e46a50a;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h141dca155df7d92e1eab3a3391725de3243cb19c583925554023247dcf2e8c792e45169d3fd0b33cf04acbb2390f015c7766429a4f9f56bd9332cf2d7ecd6543f04ad254270f3a7fa7e9fd9a96809080b563098ef5441c6aaba08a4bef840a0fe28955320dd3892f49;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h191923350dff2b3e989592c954573fde937dc783c341e23598cd35940f6eaf47fba64623a98b24eaff24fd45d9a26a79c5c2fb67139d89c47a482d2e7cf8b90ce487c1e84f1769d2765f7bf8c7d20b5310d09942cf3eed0161dad2766db29d08e234a3b080fd67b8fa5;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h114e6896fff4d8ee08b412434daed52cf48f32ba3987212ddff163bcb6683ce87b5c4527c8a12658ab55b8edb70b22ee2d55b32c6d7ff60788ec9dd07a10099c85ddd0038e7eada1a1b5688765a036988cfd6327a0df176aa1f88513eebcafda740ca2f21c478ab2c5f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb6b819749a33e10fd919cf45ab681b0505385699ee80f60c8d75c5f9007055f5d030e03adde3aca3c4401adc772ba125dcf0583119ad0b572867d3b476850af9d56109f8dbd8dfee6707dc06221e1fc4aad41ffcf14e6305a751e5c5c387a71a6971b2ed7b38641dc0;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h618f17ba5f104cfe542cafaf3c1fc62c4bedae38cfc205715a4d3d5371cdd1062a2c3f1cf819888e7c1b4e2db5f1351dbaf4a31d579b75fadc5bb169e691244e025252a9e23c0c2671f2eda3a1f0b3472e167092c0a70c843899c61e4fd45463bcfa53ec0efd05fd89;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h13f42ccfd84e8e60e3ee9b595dbe9dadce0344a36d5caaec99e6a56643fb3c6782312294285ca07775e9dfd049f61f8d76bfabad9448fa8c3fa87105c7e65631fd08076b1620f452d9f8516f7777a17a5038dd7ba599da729f93dae059941ac30b008593f173e2c07f8;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h63ec60f7c447371f7adbb98bf223c6817ee50a6aaffb6b8b28bdceeb01d9b5bb3cc9f3dca939d7d5a07889bcd061033a09503d2050656287c4e38c1fba263115abb0e7600ab8a0a5c87a8c75d6579a8660d14144a97f5475f73f629d5b2548e187121db54e9f71650;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h16ba07568b6528c3378dc4eaab450cabffe6e563f2588723bfa42c138e4931bd3c26a2ba15a87c7919b54ec631fe2a8b99884baacc759d7d67ba80d0f6f54ff4769df42eb75c5562e3abf016ad4cd911246b8d4027b7037cf03457962cc58fa9878cd00a3a986673320;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h515c7630e79b963a621841ec9b635823b23293fc5e6066a9364569ac1cfd01f9579d808b40100b2029072fb767e022144fa7710954c13d572c01907f9025018047db8878a560e8631e3f9d7389fcd86540af0bba69e8c97b7e94dc2201ab5e489d1223d380c7bd9c63;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h159ec90dc1efe3e3b0534375aab5d2046999a5d199fec4f363565b374eb089090e9c607bff8819daa454e94fd27feece09c6d972bec44bb4f279a8fe220c580775b18df5600967023deb0f6009341054e375178c7440b165df1a4d609c13714347e6965b79f5c6d3ba7;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1faf9e46dfeea1c276f5b28d676ac5f4fad63349fb95474498e5244d7482ebaac5264e70ad6a12b8c2d38662c6a12a53b23cb3d5708dbaa713cc2edf22ef0405ebb8f719da1a6bee4bbafa45d25e758c779ef606c537f1ccd64790a73a21f9da9a4be28f30ace6372fa;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha635c7228abec8e5751535d0d22a189fbc0c90e5040cecbed12b3da25235cf67de704955fbfa3aa0ab1db03ae600f89cd3c181554d000ce95712f54750acb9ac77931d136aa5d63748f77262d849f8d202f099c2b2dc92f733bdc316aa7b7d6a7f21426674666f39e6;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hbe70e5e8f3f4694f0423d7e57e79dc44fad22d9de22b6c2daffa8881b8280d9a1d322c0ef2c1b76e61035b527ed23a85df9f1a420038e7f43d31ffc07982f7cf5ec7ff49c80c00e52f783b777b1cb706e06c628baa72c82affa778452aebec10a6cb2be18a073290ab;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h603cb195c37128eaed5093061454fc049a7d4a38dad035ac688928036e9ae465179c318a8f28f49c0766d6dba7f45a8affabfa0dec9f1cc7755fbd79e6a51257d603ed815a5ef3147d0a058be50b82eceeb3f506565c3892e94cab3595ec0848f10ddf0a5b94c0a7;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h4243c5ac96ecbbec913babb7bb3b492937f25cce19408f36a77859c753f71306d99cf370a2aa15c4683c6ad205aedc150278d1506c26b4b3b6e950cdf4e0f50cbd0b50c672f18f19a8dc11c7aa1f8cc71ae44f88c822c95cc7733238ed9b83f3322fc5ffc24b9f3ed9;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h126509a79045993a7d85fc98c207352dfa600b1e18855f9868dd8cd553be9814a8ceee8c7d6658403b21ecdef8fe3d02b67e1ec812081e0f6f720cea930a9fdb2670d23404c43336f08180f56159dd769b7cdab72b7c0a3b664c6ff71b4f104ad95d8e0883585ef9950;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd14a12fcaf4e3e02adac90e19d806feacca0385e5c612c718515a3cc7bd986e4345078a7863587654efbfc56ee6c88050c5097a39bd87127012cb81d79c78718e6cf6b3e499076016c91ddaa120b944909f041f6d461e024f04889263838943a0eb88c3ef85f61a1e8;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e098f54b6cc47454a29e87bc93e1dcfaf848ae3828e5b7c7ebfc147364040e7501fa65b64f063f630574941625240443f02f1181c24ce55990fb590588decbe31a6a29d30efa2875cf7caa28281589d7642e896387cfeec09ebd263e1ea5785aba906c3950a42c4ee;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1940ab8d754ebe4744a0e50de0eb0be83469c4ff6faeddea668c43652d7cebe2442990c8bf8c91f75e6dc3ad1d111a91b4bcacb3f89ca35cd1ffac9d493fd2304f1e425fa5a22ffa812e35e33d9da23b7bf2bfe5da8487b9f6c83b979674940083204de4c253242d84e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1de06ed890bd104561fae903d4bb174400e0948f896993b2f679c12eafad1cebf92498153cd11794c24f13afe1125fad15d418f22329c6c7c195e307f20053a220edffe7ccc771a1002be02e9db844cbf3c48967ce451d176561a239a11b7259c66017d36e9e624bf0a;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h61b94afc3ef488766ea648917876eed766f27a4eacafd82fe07b070b75b1d679fec929343d679bf340a6c4f7e6da4cd1a6b060702b12fbd3a9cce304b5a18c785347824c42f2b039fe026d50a2815724e6c48e6f982252e158be6ba035546ac7a220bc8d1144273501;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b735267af20b2338197335f78cc8e879fb9546719a5770a51fc3f61cd55570b74cc4fa7e5384e72633dc94ac4e225e2b647404cc0a8616e40a4992abb2338977ec75ff7f3e7a201d7f107d724e4d6c68c132652831b95a6ca92d275f899a5295fef7e092b395aa96eb;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h19946281bdeed3fadf00d751de36326383933e54fa0e0c171526ba10a81fdebb075a0a8cd8e226c787c8181d18624bfc125faaee595ae93c430b6eb5b25b63efb685ac6ec639c3e3deb9e85d12570655f023bb739779994c92ee1eeaf12e2fd27dd7a68a0cea94a74c6;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h38f44c0ca959bbd8f4076611d73a02b301c1ba3624664d5746b8f6df2c732db9763fb85c0482d4bf583201c445be232e174fc4302f93da917949ad5a5c981b87ae7fed2ce766587ebf74980826d535059782e33c41a05b379a212753b58f22db659030f56594a84d20;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1299fd76dc3ea7393e107dec7deb7e4cf18a36a7d076293a29a7691eb1e889d5b9babc3598f6e29fe65f1f58222c845015102b102de1de7d4527180a1320137f36ac5204a1cb6b7adf59dc0bdeb2a13b5e69c13d682665e2c587a27f9928b9390f1f99c3c1205368bf0;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h16b20c9998534eb2200e174fa2bcef4e23827ebe7f0924e4f815c3fd32851ae5f77fa8066890e511de4639f6701eda42e4723f7b577327fa5d6f004d56cfee36db54ed0674df6f1220386a2e7ed06662deb08a859ca279d1c333cc14aaf7100216d9274139b15afea54;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h5c775fb1bfd36e8fbe60be422547cd3a5d3d193310944d1b30038f7fac063be35777b88633590215817728a6e4809ed2a3efe46f4afeb2eb6ee5627c3f4b8c3ac798bef2132e30686054065708f377ab7f042a72041ed404f64183daf6025888dc2163febc6ffcc5be;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h71c6eaf33b49022f1fe8e958a1cb75f00414b75d9f1e67c60ed015c0da32ae4f1002a768386edaa8d0930457e5ad38370df7dc7bd6e05d5bf0fb4161c71f07bf5a582e11759f1646786442c92533bc37018130b202e09daf77bb5a1eb73103d14e1815b25fe2220fc3;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1385c79d5e2b87c9664b23d4765e4e0c27a76c654af9cd45078c378790043d2ef226e8d8c749feb88bdf71228802bcaa5590d7763b92d8def8ec90e33eee95894c16158cd64aad6870492e8108566f2d00cb2fe321c1b3f0dbfb7de096ed995e69c32bc1b2f455f3d9d;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h179624827ae40d6afe6673ee6e92fea46b30f83d39cbd74206af30a7d9a4c0a9b95da1113f56ee26260f62ca95f55177ada176d1d8bf9d6e111570a8c0eb54f7b91a2e115d14800feafa947bd335bc53d2b417587df90c5c56176b4bc3f0bd8da0ae3cf39439bb82f66;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1cf285f44c6b30c88db7cf2e45732970ca5f2bb94c3134f59cc29185466110edb9db8107ca7caba927e72dd7ce298a60171a4ce4adbee73383ba9af3623e2f4f97f289721c3d5a4c02d4092b00a7167d413c01b2a38e70568ec5d6c6c9cf8f032a39dd9462a1a0c386f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b27a8ae6837d22f2e100f938650558d9477a1218b86530758c8e667f9a854a310e4bb1ab4d29d2c03c14e3243b085a0458daa91ab7615cc31b4a26b170d41caf234e3315a0a1ea5285cca647c5172958e5bb381a4094f39552440f5b3ba54d0a35acf9143ca6e975ae;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d4dce9796071dc75fda551765255a9e92fa2b0a74158c30023f061fce0df171499cb4e8ddd013564b625cc0c993f2f938113a4b8d64ca8de8bc127b865f4ce4944a97cd665809a3e70460a26d67142094fc2db5fde1544e83bb06141ff35e3c314ef9dd80e8c1b5634;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ac68c434d4ddc3ce2d060615ec2a4142a8e2bd82ca026c5383ec5807c12f482c22b162d86581740b0164cd900c44735c7e7d39357263709ca54726ec5b5c49a81efc987f03a6c8a77376878d53575abbd737b74a1a79bc4eef9dd6657110fc040528f23d91fc5d4f45;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h6298afcc544c237ef85712254c406d143f0f364b1b6ce2a6103869690a2563887658fd089089212dba223834d2156e87ce1ac6f7267cc737cf62cf905b4f564992974b68461f3b33b1a537f8f3592f04ff9562236f1a82a591326db769f18fda35f8017e70326806a2;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h11d855b8b3e767ba70934a405c607e9c7a2d45ec104d2c94dab46a70c28340664d11ff626a93bc28bd022bdb29071e2d6d062093cca688cb1c64b833e304ed2959a589426121aa07c363886db0396426fbc45ccf2fbf640e59619190d34759f4af35a48fe8e5e851964;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h16bb743d646f8da96178166305b46b6bfcf132bd9c0eb048eb9df874699e8f38ca4dfe3dfd968e7c508e6920ce6c7d7847c4a6197dc96d32975e5680e718d0e2c3ceb762a5fe7a825242eadb7799354094899be6c3beb78f081269ffcf62eec7f9019a958bd453230bf;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1636957d9909695c33e68a4548d1e5de9651c86fc17e1fa97b6ad44d3a0cd35dc6c34aaf33012850957d26114d8ef707eef962bd6f0b7af9d443d73c8003a46531f45a9e85f13538388673167eaaf7c469cca6742d7b3bbd12658572975463e8a186c8c5c3d8e8e2b7;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h17bf860e90665d11932983f4149c016bdff3a55787644153ce172b6c684d04fa870a650032d6f6e685ad85846c51e7aeb2c12da15ba6870bcefa50be1937d420ede342cbca7775ea2069aae52faac016d7f477255e456d35077c32a85fa28c98739b6b6a3bedca7d10b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h13549df7469b81d6abaff8ed9849807f9f158bef2143cda210c448c7ad0523f37a245c141933b299b6ca6f6ddc827256b08157905f07c5c6cdd92769c7ab9014586b25caa8a4e843902db87b8b424ef07840ff222e07f90c0e04187686c05511c0dc3dea8038c32c0f2;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h11c2ef839da960b28d48bd8d7f1216846127ede57fe5a15c39ea5ec9e02eca7bfab7922953ab29d4224285121c25217905fe9ef369cc91a1201c2675942d62a608098b3185ed048fab32cde43b8b65758d068389213b3a4c564f8599b74a020230febbebf5d5efd582a;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h7089edae0d13e33591e0c51e1be77a814d111dfa660b8fde52862cfb1be1b59946989a10cb9cb45df46c35559ebce2a7724ab980a75e6c944c5a7dae82a6a84b80461924e023c432ef297b2e134a8f67e45ef54c7e2ef2c70ee6b2a08e208de8fd8af0c59975b11f8a;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1faefc8afcad974f542c34dd2c56ac0a4ca95863b73ad750578b681aaa98726260b0eac3a31520e23819a34983fde6aba422f95d990a1638a4da923697ccfb20518020ee97b78efe07013cdda9e01e3308d96152ede29d064a597839c2c7cf00657493f3048e01cffcf;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h197aaebd1ef16b85850d3c0c557b1e487e72420b4b76471d66f403a54c79d399c59effc73f126b52ce7d9c140294d6b12da6032ba4cba04227a7aa6c12859871da079163318c45c925593f39ed572f7d03bf1b31bab41e2647f0b36689ec724ebb00bb5149be92fff83;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a349fc8b00520c4eed19cf106c351a00a18437bef461b0d80b41c8b9b7664714c5ca9b8312b8bd9c4c7f1408927f5fbcd241317d28cdbb2a8d93de328b34a60dd422b7b12880cc4adf3838ecb4a939e90d828d4e7d401a891b5f6fe3a58b645cdb71903a3c88ce7917;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he736135962b124a0ae34fcc00e56906279ab238d9b3bf32ae1c830dd3ce788c04c8a3cd2a006e7ce08556bb523d31e8cff47ea5190678c8c307845bdf750b06ec222773714095cb24f61dbabc7651bd229c27bb88602c52d0455ea4e6e8c0a26598ba0509e48fd7f51;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h172f789e91100caf195063530603fa2e9185ac5ac870d2a9e1fa832d501d0c86bdfd1d446db75bc19e293bf765a0056573f13fa53ed978f75a60c7239f1b676e2de1375d0f44f933289c6e1f3f8d07b6ffab0e38e7bcf135e74edc81d5a64bb4cd1140a204094a9227b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hbb6b67713efaab44c3920e62e4f09ec7d6faf103e333968ae5eff392e9a078b6dd3a65427adbfec39563dc3b71bf07e871b3a52fcb1b38ba4fb4c636e204604d8457e5b83f1d639438d6ebedab64137c9ee4f83254af2a2eafc5636c176250c05f3d76cde726b1e316;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h2fb73a9ca4b59fd5b394f9013bf5b2c34f8150df1dd81c9b3db4352b804441edf7b0c2a59ad441022a630d22d7ceb1c00c3e84149ffdf1a17c23839b572395afab661bda93f46ec120810b044cea8ecde5d3f65c58a86e2b68505b5933d1d91101c8d8aa0e244f3023;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h138baf24b4c58c4cca36474f7824bebf72009ef9c295f92d721d3988de7c991d744f49abc68f58ffab6654b720cd721f8fc41e6667762f010b53eb64a02837ad4304cf460abb08925c2f718cebaf656b5d49a43e2c8788ecc91f8fcf818b43a6c63be8892db6ab265fb;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h3b03a8234a3d713746f4a1a489ff08634ec1ded281632e62223a466db4c42ce1abcf9cc074e1e0ed7f46b023de1e8ea35964b7c12e98412b876460c24c0d4f0cdc08656e11fc6d1c4f98f9d48f35245f5284e9505534cb2c260397af495669610e252e6742d66eca50;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'heafc072805e2c91ce31070ca3efe3d504454054f51e307c719bb42bcddcc178a4fa728823934092d417f5197eb15f86746d707639eade5cd75fea7d13ccd87d28f57a00b34ee19b000c189aeb70a6d570a227c1f801cab94a9908ffd1b11f81c9a4e79ee176690bf57;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1123e024dc650b24c89ef73abcfad8e83f93ae63a1d526c535a06574ff15c100e1e44bf97617f295aa8b33ba31d07a54ac0ed34e035e9a22219ee74b67cbfb4fb0d9527f1774f3231f370b78f05ab13cf049eaccdedda5f96c41c25f4583e6e6a466135e1e1d98b4a93;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1575a849ffe63cb784ed46e61532d19c390f2f7518fcf5d1feb3eea1556ccb5e41ee43451281351ae8e1b5f56452512cf0ec75ad476814da14155feb547486f5bded04e771324077b4a961a814483d6251dfa185c89dc35b592e7da9b48dd0a1293aa43132673481020;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d82a5d02f2e642014c197bd8de426c5cfd059c4f2bdbd5335ea203990c8636c3374300d133a396b3fc5e7ada7449f24abd307383216ff0a8f3cde514be447ffd332755408d018bca5d8cd26712a2a28547b979affcd5a7030a1f7cadc8a44121414f1ccfd01cb30d78;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h150e8839553e406077f3f62d1ff8bb5e13cd419d3c230c460443b9f095f07ad50e602f76a115ea11d2e2ee6eacae6de05125f3888da0fcbfab742970fba915894c217d332ed71ee2aa09c482b131405710903505b6d5bbbb84a71dd18c1289ff4c0146dd75b0876c7c4;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hffb2520354c7765e24c0dff7b8a612e9304f13c5c9fd6fba832d8bfd134b6daeb032ac56cff5dccfac320c874df57f7392a2f012204e73bc0ec2231ceb1e596673c7ac6906da5e7a2a1fdbc3bc0542359fb953b5d1e1b889e2d67350e8d901b604def2bd3744f537f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc3b6a1f3b676f43860e2e667fc78a9346f863d0215ade5b978289728a050cdc1e33f84a690d79afb9416e02e83e171cae465eb936ccf81d3ddc3207108718ac94fedc91bc6dfea5a38a83904c45b4f8e681e5d6ce338340a1d994a086824e516410f3e8275942c281;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h16b23a9eedfa1eb3431efee6ef4f726838751b9b98a68a5abc7801f3ec36a72f479626d6eadba54d824aa6727f729ad3fcb43a7e1d5b9b6db9eb5828f1f2e37124b591615f03adce183e4deb1106ccbda1f6973b1104e91d2f3c323f28373dd7de4d717a312a0c3173;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h181619583bca77154c1bbfea4f53e7c0af76129d3708c950c0fc04b83150869c73a405ada1b0aa973e14e240251129bd690d2a9b325be6b6e61192eddefebf502aed0368d2ba5f0e4f4f9c09c93b8b032c2d49d791b801b80a2fc15f2a97ec077b57ec27de38976fa2e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h39e1d41c09c2f2d39c5307d1f05106d7de70097c0276092e074935294800df44c7d9a92fa3e7492cccb704bd0a8e911ac52a6458bcb41cd2e2614bb9abf66008e17fded666268d2765567b13940a12546e2ad31d1cda1910b0853b109ace4737d0c557efde9a283b39;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h755d0f57dd6e0b8a88991652291f41b19c0ec6a525a16dd305e23d81a9b1f38a89bb623b5981bc147e558fa040c46977a969968959d865fa74670640449d71db5eeb1ae744545d3eedde383d777ef682434fb74fb8a733cf10a34144f52eec1290cb680194d956ceb1;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10f0568f310caf02acdf9f737f4b2e82c75c3faf4637faf47d3fb68eba1c1ba5f070b3c5bb150bdc08219dd0b4478fdfa67d771b8e95ea224e1ae3466f413b9a80d8c156fbc63134f7e261240859eee2ae79845054d112b1275cde8955dc9e655f4d61b600bf563719d;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h66281b445b4d73fd347d76f7ee96c3c64d104e20c564bb98d016b8a8470f7e5ad9cdaf431f9bbbbea1ea4a57b1d81579b48d56dd0bb9fa03dd4ee14819ca33df5fe5aedea1052381f225b7ed68e15e6dc90fad29de84974994f6a6741271a12e25175dff99bdeca568;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h19a6720fc4b9138b51231262e8acba6242a48f3a5ed67497afb6b413d97172593816f1a0c47ffa945d632978dd4df3d4a5fbd01f14bc9c71e5b7c0cb573eda7df18ea761cd6dd099773fec49476ce4f8e0ac7e2b28edea57af2de678a12096e70d29cfc5b6ce5fb93e0;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h16a4afc44a41f61b6756e9bfbb0ee62fab41af80eab0fe71ed5e4907007a1ed56570f32455d0a3735469eafdb4e95ca73abf5536200ae9543bbd3172dd6acc8a2499c1de828dad581b9ec3c88cb2e5243c554553b632d940b13b13bb3f449c71a25097acf5e5ffe12cb;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h7fcfce4a35866bc12a2b1f001a9fddf055f66ce1eae4172badcf9ec607cfbfa9c01169c8fafe9dba847911e0456294f5bc45063c890efde87e0b3f2a250569f4a712942eb2e64e575ca46ed7bf003a955408f21d9e455dea995ae74ca1f76bc71cf242a4ef097df70a;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc8efae0b798c12dc2e9980d4dc46423a9e473fe8582b13aded7f5811d67b7e64e844e4bd397faec2a9c70e4d46208d59924cd745f1a6ae4957e7d6e8ea2d4aa79932c66b5bbca3a557631e64bfa776f8ecc78df52feac53ad3a97dc4ca36935844ab1c444bab3de4f6;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h19f0e315f212727122fed51c56a21fbd6b31b02e54f5ef5f63a25349c8c6c0d273a9de6971ae843bee2b08ad599b847ff1449e462a2d70f1a54a6ebc45857e687059be15e0a944fe2f1fce11b47f684b7a24905b30291cf4a9972f5a271c51700fc17bd7100aa319a13;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e06b319c1284da2a8b9d9bea94f8d90ec927b2fb0d7ef311da2631a271a7fa94dba322541aaa4b6cfc0d530f626ca242fffbc91796284f442d0691739789e1a5fb39068965faf67028aa4237cef9c8c97cf88840eaf6bcba7771560ff1b703a85951a0b70a0eed6adb;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a6fbae8bf200f2ae4fe4301824d9db3e59c144f6666dd192184290a2a5df27d748f450e0d22b652b233d41e7ebb8062ba297e8c7dfdca9bae2b3b0753454343ce07227004347b1dbac39f724d440fd650ffd1397525351f7fc4f738782604365ac82e21909350038d5;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hfab6c8314a6d8ba711173acda9a3a77c0c5f626dd365a14ec1222ab27d7cf624ec581353fc33d6f5335313770a81edb20cd496ef30030b8e3a87f35e74aba857bc0a9a867c4261fbbcfafaa5bb4196af4a4c600a1f865ff5f39ab4773104dd1ee3ebc3251e8e81fe26;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h26dcb581d1890ada109ae41c599b61dbcf460b0f4659127feaad6cc05fed4496efca595394f3d55878330d71c775286f1b58c9d0afe31e041a96e7628068612da5ba07281cd4ba5976c1774f86e712fe3451a2569f52c12bbe08e6a4368d6f6797883151b25fef2660;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ae20142e90f1fec1359057df970079f1e9f1de55c014cc028a023f550608aac382bb553cfdf3ccee350537e6fb92f5badc4fe4d68e0720c6f8a5471285cbdf7f32249c438c6ae1f733e2c76e29565a364e078eb9192040b76acc5b0585614d354d9c20cddb303b9017;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1cfa8719cc9b44b2f6169e994e0063933e278b13fecae5062fd12e4cc97af38b703a735d12d577f644d72d95d2bbeb0350ea37b36ee2a3062ca6244565f527fcf68d4436d285f73f801538acd629478026d21e708a10374f0bb2c9e5a569bfcaa0c62e3abcb9ba58951;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1bf0ec6ec90af686746815c0ef3e3492021aface52ec8f5f354fb7b5339df6046d48239ac83289d42b720b305a133e259009df63d6a3052f6975ee172a3fdf7f3f8ee8ffb2a033397ca974951705a232d9eee7e7e06f502a630c6e52bcd3cf34fc5708f9fd36eb86173;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h312b47ac9b3bd95706c342407bad3d5be2df4cb7bacd68653b1e93b8e00f97c208b422bcb0bc0bcbe7eb744e367cc42868ad5677873b869c50bef3c44e6b85c4cce973aaff5cec72914af1880de1600d8bcbc3864ae7ead29c7ef996f376d70160e329826f5837c1bb;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h9c2db25f142391b307a8b864394fa70e46114c03807dc0d3a7fc23d9b8f070a3c73ca85aa1a0799cc7ece6740b229aed4a02a159b2158426531924a728e1bd405327badffcdb8c3da601d25a67c35b497a4d20ccab60e4967fd30fb10d80917299ac754053b8addbed;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1fa5c6402cdf0aa1c99bf701e4173e492872f0093d35974de9c4a41dd5dfacc275a3bf8c8e8469a5c723bfb9c8e78cbbe0dc68ab7f4f318a086fc37d408f5c896c0c7c5e9b14e1a6f1af7bc4dd77f3b3749426662d0632843acf69d1b360463b5db7b74d87f5ae873e3;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h62a442f21673425af6caaf72aaf9637191b107b63dc4b09f5049c0e4e202662919b5f0d1e40deaa94c3379d5407d378c7e71289da111169c61332ea0199cd9e17e7c399e539a6635dfd54f797528cef9ac2f8dd9ae72241c7f4ddef0b9f7afb519082bb8bb7de08a8d;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h18338ab7dfc069a58730557de780a2e2b7aa978cf7a4a8b0ca2d414c71e2604e2ee24847e4ff30ffef967c30ad23b09d23a9568e0d433c3b22c209fde8217734cc14279a51d35fee92304d0e964fd697772c492af4230cc3d09f554debf0ac4eca751bca524de5f7d7b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ab49e4126d4a298b8afa7216a4ce6675e29c6b1de2ecf04e615400a6c0f8a4325e39f13ff6061b3748c85a8ed6c52d03b06bae65103700de5fee21aa34aa72ed2e3de7d039921880d08cbdb4c1ed987eb8e02eaccbb2d58ea9ccc6801ac7901b1fbc49362b6eac8a;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h284cd63ff48f20a8440d7d03e126f5824feff64662a31b7353041dc0135f9c99f8e66b5b79569553e2b7222fb529e337f5a13b0984b4369f9195f1e99e98d2eabff10f0c6812d88821aa83561a6a488b5c6d8df3d81cae3a31182af18ef9ea1ebef873abfca42f6408;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h13200b9d314b79736ba20b190dc4c6db1390b051b8f1eed83c673b61fac247f2e8e093bfe91c82718da4f21b2d5537e8f9b6a52e35cf2f3ad7d1589869ff230d02c958bc161861491f06021d16f4061f542b2e9843aa9c24d6e0755c27cfa5b34c9039f5c1d31d7fd78;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1cd9bfb8bc507e20bfc00624e4f3be6e87d2216ecbe7524b94381076ae9ce69cb8df0d93bd0c71959bc3ab5a46492d73a4b666ca4b2e781bccf2cfa88d0e22dbf2d030bc5c25ca8bbd71bebdcd740561e1ed485346288b654cd24737bb9ee75bd2e28768ca4abe08d79;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1744b29cf046141862cc87f97b02fe22d0237742d7eaab790442e8b774066e7276a0bece6ffb9d18b202f9ff975e03b5c7de317496c25fc5376e69bc725e2c20205b4a19e9bb8bcb970baa8fdc3e50213824c2a7ba52db2d12e401a78bedf7791985cec0a416d6bf292;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e72eadd3d6fb63a2855ec230f6aadc6bde82d078aee1a12c996759d5b907e613cf226932fa7a58319ac346e5eae558a0e61a5efb653bc4c860198869c1810e91eae65ec94e4fa67fe954dc37c89fd01b1baa6b4591fc82d8a6f82a8b46bd1af0e7886e399b07d562d7;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hdf63d613fca52e88b746c19685924c61ccd6d394a8c0078a45854869b5fed89f45dc869628a3afe58198959827e6f63ed3af3cc8a569933fbf0898ef39596c8f92a30eeac3952278e854b5f1e91a92fd18b3c8fef9a55cbb1b22d1b53ef43c12dfd36e1166861bc08a;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc39d4d2d4af3a8a041757955e0d655dcb2d78ca0c067b6aacb4cc14134ca05c1d2d1e306256140a3267911f195bd7a569a3e7ca6aec8f924aa9a50ae885306396f7add6d7aa30b5259277ce47305a5db61298550b656c9915658aba4486275c2f23535dbbdfc376229;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h11e24ddfcd29ea60a3984d3077022a813b0ea6b520fb9354782df877c5a0f8359855a330a4836d85a096c059063e38837c6ea496a6c861e403c9e3760086fc7f2db517d55b48dde356a59ad3d5e27dd6f24767094e867bff4e74efa784eef8be114c4cd9beccffbe7f3;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e8834d89ce2cb1d41ca879b72676d6b9cb5aa8698500d7033edf59eb77ab92b9cf5dc80a5528a79284b05b0f100b6db8634b3447568b8f25c3fc0b626fe15717917985724269a98b0eae57931fa9e0e0cfddc6b3e546e82e9a15074eb2bf2884cfd68a32a1d44f97f0;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h2bfbdbd82fbde447f482b2adb980ad5dad6f110b6fb268e3f69e4b0cf16aca2883bb5979aeb0b293c29568a026a4ac60ecff3658bebe5d1aca642f2e34edddc347b8c3aa247ba5a8d19f8cfb9318ccc812d700e36e3e48244357626652a4f6547624a13a98caaba9e0;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h11a2d18c7ff5a551cc3d67ff679c560c18c79aaf00a35485c0233c7eff409ce78170eb46344c99b2d7db956d1e60e9d26b0705ba15eb7ad10062e6b081f517f24b4e55d4b0ab5645a633d07a7c1f11af20e235228108bbe60ff0d8f7bd0cc8dcf03f20a9925badef409;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h156831b71e38a99e52589acf40b7410d64ea7e1ecd69fbd11d2b179db62abcb2c1661c5028669d65d5dc0b88fbc404577b908be4ed94a2e40cc3673f899b0e807a30a3c30ea731b44452913f712876a8d5ef0b9d94aadcd22cb4c983f530ea917024a42cc6521b2c8e3;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hcc928c8205a553e6fa0e051922f76b6fe611e1abde3bef7121f13abe26f622f0724f6073d1c5a7ce16182f7200ae83158532789477dbd193d6adf0386ce8a537fc4de2b6754513480710d0fc1a5f4ff98e3cc6863a472b6305d97fd3649d77a0f74d43d9c47d9dc06;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h182290bd157845af141d53e0b3842de017f5e762b6946759cc5eca72a6583acd58123c82f5d294f5e24b709a7c26cdb78d394630bdc2c216ec4cf93e78a34962ebdd7406323706c10af0ee26577e97fb2f9a6d0bf4252220f8c1ac48cc223b959e951e1fc9fa6d6b998;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1eccd68f01feca486ba7485ed6dde46ba0ae161179c142eaca589f5a964363f3ce58f23f36746093f137465e876971821864d84987016638cb074a67418e824acab6b773c9422823bb1578eb6c5e6e680b27a928014f0c63f1236e592e291bb663c1d1e1a73da2125a;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1da0b039510c97f7271de706db5a33822b51e3488bd8b3012684bce74966571b0ea3158c05525adf0ad14f9d52be5fe58e3bf60a7ce78589eb38f08e4c54a3dab2503cb44893e5297f0f2055daee72260c870f29115b96796d32fe1cc88a4ab77d8549783345a8b0143;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b2dbedbb562e9dfe030424e0067b9be3153c0b4b7c3eb8bbcb6e68a6dbacd0de1905f0efa6bca36b7db34723c029c741f7986af99576ea1d7b1b9e82f6faa0f4bf2e29e9ac04d61d2bf7accfa124756bed4a0d07a9c1c966d33bc64aa5062f9c4e99f903bf11ce1090;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e945e973adbb1403900cd07713c69a3d634913c0d154a28cf29d26c27fbf4349dfa672a11dd4dd229b4591d45cf19155d5a4a2fd72ce4ed4a515b67297123d8156dd72a9850ecd40b3ac41c4ca4e2a59ed4a78a3075c4dafc91d86f6de22be629b5ebd2ab3261266d9;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b2cde4c7f66d0d6d73ed1f760661675a0f31c62557bde1a859b652a410cdcd033a6a3094770bf5619a115cc863eaa5029b3898f579ebe6c28a79f23734899eb9a4c899d6df1e880c0f754fe827e5b6861596213fc899be931408570d36f19935ce776f1180d0a94b42;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h4c263b9c1604eecdb9185fd6a1cba5d75024459bc6ff0c34d289c978eb5130ed2e293ecb550ff117cd81d8d5667d899ba1a5c864fb00c1e4b2c472313856cdd098f9d1e34cd13bfbaf81245b053f678171fbff27c15f6bb61ee621ca14e49947c7d68f4b0d3e2f1a66;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h987c5bbf57ca2584bc7c1e5d0df7d5bd5c7ddc1476cae5f272dbe21561375c13eec7c3bd9186a519ebd1390f911a3d1b53be9233c727af504c600aeb047031b2a887f8b76923b487d599c8733796d90c7b79b5a9281641bf139ce2d91dc97cc1c69b0ff987afcee705;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hbf5c9d633b4df03cbaf66c540a14790a4973d616ea20216093940deb78c24e7adac37dd17448420dfedef91a2657168f0a10cf06fdc0d7f76979efa7513a6e02d884862af0f414866be954f32a646974f16d225a0f8382bf4c046cd71db54ea81426d1df3625f8d54c;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h4fb7ae96e8642f358dc63b35ec7f09d22eb3bf46f7f7321de1604daebb27467a964ba5d99f87029adfa88dcc4c2b7ea76e39dfaf304357c23f3b3d4d1553d415b4b485606d2caae31c3439d35d884c320081dc391ba83c3f0a3f22d773ada22dd37b73acfb7396e6ce;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hbf3363c63228c4c5bf46c10f1dc33775f612248f652c178f825d56b036668527e8b548ae62e0db8b2956e0bfc4ddea5f0803bc16905c3831a2626f457667973ac5308b8da1ed6c4ac7554dd6b401d7b3d5f4762f04d13cd2e9070f5ebe4320aded7dfb6f1dcc574309;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h33ac998b68d9e4cfbcb5b71fe63a7fb77ff15ec240c7e8b06c000043b74a42888036bfce25786351fbfdc73cdbfefae534ff87502b5831c9ba1aa3601a8f8e0f2d501a5f06948fbfcb3ab7ad4821d9608d72ca750a6205f6ef3d76c9eedb67fb8b868e30d510681919;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h126491f31a9532893d3d7e2e9ceeae1fc5167b335b8aff04682e8899353f4c417e64aefbdd706ecbbf34bd5b0c7a082740177fec6a2d502affdd031a41a81ca1841b2e181502bb8e493d903c2959664420763fc155ade446c907f1296ec51f20f469df417068188aa69;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'heb5527a7a5708b6d10a3dc2c6c38b162e69e899df25f0e0a754fc810a370741161842e0d3156f801a061b2f589cd0f37886fdbf54fa065e6593c1b1491682f1c3b04d7bc02c8e9112e26fd71d778ad71906e2fb0cdde684d078a7d46479853e8374e224ecafd5da17f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1779a79c027a13bd99b53e0059750e0ce486acb6f90385b5bdf071cfa4f9a1e45761a77006b60a1bcd3212667367ce786b80a69f6266f53eacfe1bc02dc287e1bb86cfc747ab18587f56f1c7650e3536030dde332575754f876c144db8e29ec8c92533de4c5f3837aa5;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h9dbd937bc0c375ec4c790aae80837ef7f4081dcd9c01ac59cc93bc02d0f5865dacf8628f7633bfa54819e1d3f1ede943d99254a088dfbe647efb960388b84348159b7d0674aa720fff9ca58e909c6a05c515fb347aca4e4dbd546a4f5350305be547b5de3de5432a42;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1626d24a9520b80a5ecbb40a9d2a6d14314d977b8045c147d1fea0e38c9c7d7cda0caf03afe4d8f6a250758db081c8ae6cc6d30b2842832932413709b8ab34116b1e18721c0bb5aed0e7987edf5f75325d611dcb3e78c09d0ed24acdc4b2ffc4259ff5060d3c40e6cc1;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb5d83978225a7228fc02bd9b6cb7dbb7b0e9f2b59bbbdf7580a6fad6de177d5cc53e0826564478e66014964e6d55beaa657c0d32ab4324b65fa21f1cd11b4be8b968c19ba7b309615b571706118c9086aa7eaf869507aec4cc23a4023b525c5822e57668b714814aad;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h44f38689fe6133c56ef8acb00a02191b1c2f39bcb04bd19af30768958bd234f16936815d12c594884c8d9e38d14e0ee9922891b6967eece96c70557f6c70aa6ec8f3b8e5b412b1d457b786f300669aaa65fbebfe9a969d2a79bce10c512adaac73f963986536b708eb;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h95698b620b93171707c18ce75e31bb4120055080e06611305dd47ab981187a788d75d7cbf1224978149fddc6a550057534331c5e18345996b3870f23a2d18775e1bf5d027529a79e6cddd3e03e8ba991f4217cb2f6ba9d1ee7af93ddc6ad8b2fd04b2e427293b12fcf;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h6dc511dc75c7b6c50943263d1f05f976f58d77275f353ec1b397c138e2dd08cd431fdc9cb3182f74d72418a2b0d2126bed1ccc030bec4520cb7c8ba867b6cfb213f5444c0042352c0e1a5b86d3067d049e072fbf12bef02d0b2f1dd88b8119573493d604bdfbeadb9a;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1036d226e64d139536894cf27544fd8e181c8ed9021743a41fc274db126f153d82f309109e06b1f0cd63a7ee83aa04c93d70a50d292fe4cba5a1d68e4614fd0c53fc41c73092eea4c5d51cbf2bf8db263d8e0243e8d3e4095bf296e4dc7d45248f72cd0bff7a0ff45ea;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h78f128e464e67dbfc1c2860d3d47569d4eb42a573cb1204ac828aa29f3f25eb2dcd629ebff50baa87940510a59a2e08f8b4ccd312251ba84a1ba9a5e2f9404fa14d983d4f19651302dccb17aef79816b609e50b87fea2896d822d13b53e6abb630f4e85702d78d7372;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h2dab5c1b68a393e868c209f3e5877ff506ffa0a81615736766bf7bbb36ad7cdbe9e02a85f64764ed5992a59124b9aae9965b6f41b36e1a83c5343215d16adb74985010693320502eb2d26e11754f7baea0811263da69b5e10f9d7ded38c36bc815259c3b7e309f0e08;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ecb38169a4c6439292e93d4083337a3e23b843cc501bb1d128045872fb75e0dcc83dcb184b2075ce4f436a2c05d365c0e51b73c8e603caa3ef3f886a4186f3f72b4e295ce0955c6aba81fe9d21e52b901c5afb248d204bde601e95f0219d7809b604a1949ee5d04a67;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h4475a957d3cbbf7f48a4df6dcc06bbad0f3e2de59f1c279a969d761661c92eb51a86e5d21c8e1c753ef322affa7496db3ef34011709b72efa96b45a31659026d9f63b77c42d6294e5806193203e4603cb248fbc2046c13333474cc039e7faa537b69cc39df893cfd86;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hdcffd8c472a09be50f8e87dc41cd98dd182fb9b93a0f37660cca9dcbd072a5f3ac3511a1e49a4d86a2d58ba44196f0026be6e63d2f9bd406ac0a7f2b53e63a9eba76f4734b3641fc7b4349cb45c9819771c8e930900cec84a1a6284d08b615bdb41b2d37d64c47a050;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h2389f1679ceccda41b4b670638a190d08614f705ed9b1934994170822172db9b2296b18ad197e06e33261d1a56935933c40d632dcabc6b347153cff4f6a7406fb2b4d5c7b7bafbc94f1e48da056a6cc919f20178e84198eba4553057847eab0127dd807ffe3ae838;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h729f4a33879146e79c8625a60606823f6dbfa3c58c34a67064e61f1e2b0e723ea921d8620eb543892ec9637b8e5e636a5d64b30dec3c7248e1579618941ddefc6663edf98bebfcb7a9865e0a3102790a6ded515f78eae5f7e56204c004d86430bdcfb424758a9cd9cb;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb65357d3ff8a1fe4f7adef9d096db212401cd9567ce1493488cc00e26d9fd99e1ddebf3c0cd433c397739393ec704e012ab51b9e6c8c87077ee03d8460c73fa0d10b28d2ec19620ac97f6c2a59f4087de049b8f50712820de8571a1361f596dd6da79fa06a55e669f6;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h95429aa928d925db43f40e980b46fffeb398fe29f052806c4968c7dd76f22a97d357f18096cb62985c6d57436c5c4a9a2e9e52585b60b345a6573682d625b233f20db6db4d8737504e0837606291415dfcbfcea13416654da2dd58ca5af714f01b97e43887664f5ec6;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1dae6072b1497c9d87f8a8be3609d9a1a9d0056856c5f693811cc47efd7cda62c1b344967ba94f0185825fb36fb30b86f498442ea488f9ee0c7b3a93ae277592731d2ad01758809cb6446d1c9b33e16f376b8e9b9a11f57df7f248c362625302a15d1c18c3348c8ed0c;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h69a40ec8b0280d6ca1d73689e9923a297d771d9d64f7a74615707fa016f4ee71c242add5df44f63da7a1647e6e2281f122d2ae9e8a0018b7873fa18f5671432ef964c46308fbf7613f9991f4ff9ecc915e709a05d38a00245dc73c327fa4f0f95853a082e31ee249c0;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h6d0ac26dc6422cf4a894a42fe03cb930106d05dd3eccf69f0171785d9df5033a02811afb3cece7bb692df930c54ecbf112639778407dc97a6210e3cc9b011e73947249702c1672c5af31e338228c19ea7aeed3567ff7cfe64aafeb148e0ec9c5933295399b54c89d90;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h9921b420bd3df5998252573c698c7def8a824507f0a7f3bac76ce8b0835b23787e625167a0b2ee47ebd0986350d4c2f32f88a2975bed5e0e73fe2e12863fbecbbf241dee7459c7fec20646df7c9bf58f4760c4ced6c51338c8f3a7888305e62aafd09427aecaa363f8;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f22dd4551a22c46cc3e4245f50f0a5cd9cf9b66908e4d00f32307810aefd057f4df11957b89eb06409c2dbf136ecea15273dc4133fb5c3f0c5e0e671042d77542347b37da02e0300fc8dddeac24480cc4cccdf7de0add3f0920ac00745e4cdaaf7b77576ed68a1b674;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb7077b6ca18c5ec851790f357b264e836a7ffb0a844262e2a39a28ade60bc1659ac5cbe8ce3956c977318bf3f0292fbdd347fa1d2fe8739456426176736c9f44c0823d0044e1f98ab6fb552e9d47b133dafcfd202b793fdbd9e1c39781a02313d21d096d3ef88edb32;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h14711e2ef8fff82d0d20f56406912efc82ff9b3fefb934ca5f592b31a870961d46120ff897a5efe2faa1d8c7c127677a52c28e4182daac5bee27a1643a5d1e590a5b5bc4d7106bee55954b0aa1b078ed582ea2dc1cbb42bfebe6283c294fa64833d60f9e3495545df61;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1cf38369b5b118e3c34562f21331d84f37b2f65b71e0cf1f6716aeab0e5e1dc05a8d920ae3f9ac220f1cc03724ca9c12b777a508d7d0b305a46dd0206267ea90352ea6ee404e467b061d7a220bec5c5e7993c4cdec68f4c2bb3597eaf91f0f1c76b9ef02232815c911d;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b6e953a5b23467bd89bcc3c7f5da37ddd9538a2e51214f1eba88adc426800bcdd1535ddb120ef5620287b0e3c1346e62d3b8fd3a8d0f8f52e8d08385e68114f36a3aa8104bfe0a6653799bfad749bec69f4973ee2ef1a4a511c20877bb3a390370a7d6bd9b8fb34854;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c1dcf24fe4cd786e80bde065a4ad3b79301fff8b656f0445254b73b9c8c6cbbe9fe5578a891993ace8aba352353328bb273ec49714f7971074fb3e84bda4f1269f9d7edeb6bfdb6bd611b70a3b2a39a50717234a63edeb8a165d5cde689256395abefdc4168dcd11a3;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ac014ecb52e8135d7f42591356f1cce179d2b6ba95e342324295202fcdbbeb7a3b43efcde2ef0dfe31d4b7d76a374415b3ea1f3b62ef7bbc9553b567172a9fa06f04507511a9ac5405a5fe0139212ddd9f6fe859ddf3be4c71d33ea9dc412f847b8b47d5f8cc5d4eee;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd5ce2d5b880b4b93b422ca0bc1061bff51923d4892632b7b9a15f9bae16dc3c6c9868b8f253b9157ec648f692e915421d8e834e39384d3240f4f7957f78151000e2a2b57436cc821417886b1ebd72cada1538c74b87ea6412ebefa90ce9c735b14c45aff3475c2ad1;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1159d8188c530711ff8dff76d402b57e00d3d4f79146ce1d6f8f8ee839e2adbef66732c1926369628870fd6239fea675e61a192c90b00adf96cd26711b7f65eda8d47ddd433ebde8ce4ca2cc27d80aa7b5f52cf9606fac07c00f30bbd541f0d996c9c93936d1f43f74b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h106612bd39028ed7194c1adf60adf3328e3fc8b291dbd004c7221ecbec1685e75e93a28d738bea726cd31d14e286ee5545d82d24abd389693a4d2305c6cdd8e0bf5b7e3c4282e5cd6132b6f45e48c052d93aeb1d3aaffd49c3ed68f9aabd9c6270aa5a2d4032a430114;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf82dc5c1367d50ab2bd0b634dd810b9c7249024f99aecbfeb1374fbbc2cc9773f176c848a63f95aac5b21743bc7e48211bea4c32347623189e41881ff4757a6ac56803cb426d9ca4464770e9ab7c8e0c674c251560b473cb1ab6df673b0a2b9bc0fb2a107c1f7f8d3b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h125ab0ebf473db1430c49cd09eed3320c410f15afad41873131992dd074ae19653ded15ff6a31d5c06ccd2f3915370101c047c9b18207c182a523f54bab8cabd518d1ea6731ac1792c8bec222bf3c6c5a52572e0d6a2fe79f4c8de5167532052ccba4b235a23a1edad7;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hacc7f959d3f93b861d380bf431b8b25edf69fe349a9bf2dd44032be24e0be80c54f3a1fcd4c253d8a4509b44be97d863c597d2c5a7bab8b99dcc354333ac9dc55cab013a510d5d0dca1f862f04232bea4333d74344fae3706c312bc9333090a7113c47ec65459ddf8b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1742e8cee28b89cebcda5979df25a22346ed12300fb0471629c7a682d11de1b6e123ac5aa191aa5d77e9129d3ad88cb05cbae4885e53d0101fa30b810e8cd43350938ad191e08cb9e5ca9dc32b289b2c2c8511218dd302c593b37ae1c5d6577073e3170c483ad731048;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ea78e4ae661d3027c626afd5962470d6b805a8a84588225f3abf9c61706724d9ff81a55cb148c56a27e95fc0501c560efabca851cc675ed40d7deae4a8087325e6a263919cb54797a2e27acf30a873d778fcabe112e4f0b220db89b3add4f39c071880ccc166af76b3;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h128a208f9fe38c7b902834bf532137b34460e6b40ded7e413b09bd822b0bd69020d1d93b76b171f5ff4c44eca3b638486ec5cc530bfec3bb4cd2389fecb68d823b9a564c21134fbc5c4e093f59d87cd3fee87524ed1ac1b4ac69f13e091d18b8307b060d6fd3514f91e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h65ddc685b4c8e22791b9a42b2d23cafe823d01b02bf9f42ccb79e44958ea4e771afcf4b5f1563b268ef8615f8ae77f1cf41fdfb4de70e3ccda15f0fc30c276b9df09d1fdddd8cb7b8e17bf3f0e41e0e2ed31aa0daf44113bf6046ee86783875d5896f13b39103c3ff1;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h7a3cf3e61e26fadc2dc97575d8836525f2684beb2f4aae36807faa10853b522b8dd602fdd68024aa05b2e51ed5007d281f960a79e2aac6e321c2f72694705ee3ff0ca31bd0cee5e8b65ad899448eea0d3bd1ff6bf1f34d04749dbd7f0af8c26e5ff98fded4957d6158;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb943d7c6ec73d49c876b638a37fc78d758a867fd0b47776981740ddee84f8940174c97e62bd2fa2c96bc8aa3a0bbe38c2b14560b4237a52052a15a0800d618c23183c54d7f3c3ffdff0fb6f10db11f9432a2972c09bec11210ee284adad8f8da2c8d0f4749c61b0493;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h18f4a69ff464fff2d1aea047d6e22f2ee6cb891afa88c9f109d3aa783537fb873ac97bccdb81bdd55bce8af6027a4583359881c750b024d6f0f269832cde40d27ddaa9bbf6fd2a9020bc09ff835930be7033d9970c2c44dfe10ec4f40a7c7510aa2c1241ef1a9ee3108;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10bf831b6126ab052e935a84e19b3127944e6aad1d0e942a4400f5a836fea53ef772556fa283468dce82afaee276d80ce6615a75b58d4cb37c1499ac583b75a5d71030a22b5f530781fa9d13663ce86c8890ececcda9bae27838a824aac02a464e487114d47e206587f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h2a0db8cfefbc3cf69dcc5a6ce5de64a0d8f00a9ca8ead277e414620bec11762d6701930d714b856924943b9b74ef1faba541f9ffdd4082f94ac4d8cbb4073a2d53f014ca31b28e5af93bc161bfe658e8d11239b77e989976705d991e7c755f0985c399132a4f78d209;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb5aa828e824c90038087b92935435a7dc0e5fede3bd43d42510a1b7f7d100457725dd31bc16bc08d42329392127dce4211f3d562a7669193ea74235e6bdce051d9929261c627ab9894a940bce2ed428d7a85dd9759a09007df5cbcdbb70315c11619e86726f2ec2539;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha16ba0a59f4f398283b65e8962d263f1f8165368182ebb9a5d531e1829069ef149a5f4e8a50577e4f42669300f49be15338f881aedb4fa6fd8edbc723014c07821b9c680f0f269719717b3b36eb220a976f44b6ab96db443d9c2fa8618a2b8fef87fb32245c66a478e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h16a9f7e648af5aaabd57f47f5717de41cc2e0ecc6f4fa56be093ad206a4e4e075835b99b9828b81ee6c0b4f6471947ef81235700af8a78e56d4a59a1cc581c2046acb29810f128dd76f3531cf40a7b7b6382e36bae3e16a0ff911ff785320713623d7b1ab1732934564;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1da8b0f53f5aa21e5f7f69a958e05403d3c2b99275c94459df4e89b04cbf91ea69f7b1bfbe3837dfc5db794e86cc319651e6a234de3969c1618248af500e00620fe017e337f431c3beae6b20c155ed11fb7f5baef87b1df89296e2ba2bdaf7fc80e4ea372ed6fb22fd;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ac0cc751f4ca2ad3191d47b90f2ed9dd6711235ee387932b04baba1e45334f8841f666dd1386bdad6fa7664edd727194e3095594fd8341e2687a0c73a5f534da7ea4769f68bd12985257c52b7fc70d5c5b99d4a71fbc2d3541b7def87520527da2fad7e4df98f0b5da;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h107f293a908c981b723e3c15ffd96564fae79f2a58728ba928d49ce73f00cf234677fbdaf8506ba38432fa7a11a35baf9a052c3c4fba3b44843f1ea6fcac5bd0e04ceb944d22219c0f0b3e66d9b13b14ccfaa916179fc68c8b97262067f3a49b8110b4af8731e719d6a;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1082cb8313f4045605e087017b73bc3cf1776a1af3670ff8537907eccf788c2810d6d8c7edcdccbb34680b5df85457927d2253059e4a4dbbb0fa61fa690c1bc0eb8c4acc1c49432a5e9022d15fa51545dc33db48c43e51b9b29b45a43dbbffbe6e1cf2faf86d4ecb44;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha617c8dca2969540db76b002a3d504600ce53f51d143f5dbefa5a7479f7c922198163a293b71af6b83340dbb43bcaf078262fb79e13f12cb1f099d6059b2a6706c03beaf55fa01e3959b65a5980919e321b1df0f1ae8411733b77bab70d61c32cc6a7ecbc26e287dc3;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1cfc253e7eb583fedf471d014e700617b5af66b2652e0713d7cd022685d3f590acd2881c0419d682dbddbd35cfc632da5bfaf26669930c14cdaaa4845340f1f2e6d06456f06e8104d3f3dea704a6adda76bb6ce7506305330e7b2ef911184b44210c58f5fb52ff4172c;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h125cb2ccf94e5ae73095d8bcacefe45db74a89653b51e5b1b7012f27d59358c21517e460a470733ac504a4ece33dddbb21d0ae1f75c318b4b49c1837ad37682007cbcbd8f43ae9c1f44d62e8454e88502128ded9d133c5d578ff06a66c55a4485fa9a14089370613f7a;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e20e5ffe9c908e1992621ec3e90d1c2c9c1447000869dc500b97c1f3c0a6771461fe4c8116bfd40f1965723d30dc3c875c4613794a305432fe4b30f42a5fbf15707dbaf4d56fc6f2d3c59a0d28a9da3a57e6e02d0eff336b58a4cb41a33740db47511593d5bed4c8c6;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he3d9825b2d2a8918f654cb260251de9866e9ca51c3ce671c13114f525c88d1862c4787125da1ea7d26ddf5a1f772c79bf1e85231672ca1240cd9b12a14427ce3b44774d03d18e1ce76d3e4ddc73039c910216ce60b85d3f4db51bbdbd0ad7402778010286a8612b47d;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h17437b55e87ca391f61fe3b10048094a4bc7a2a5b92017b4e9ed89d3bbfe00964c7b26c6701b4012c5c6682e1a5321ad30ea627973c0cbce66b42142521292cfd76b1707376730aff83c4f7de99fb90cad446b45e2e4809ce67bcd4f99d62428df21c3079bb185bfbd3;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1dba7f1e2ec4b36751d3e644bb3ea79fa1a945479b9e203a89c0d9157169d80ae7dc273fa68e462ae5db68e55e80ef932ffd80926ffb08b79426f8050e38a8f7ef3838426226429d992dcdec97bb81deafa47ed700b60a360f925deaacd2cf09f571d30dd0704d45f20;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h150cb9db95309c7800231992eba4fe7f56aa87f6bce65d255f9684d83401d58e56e9d9d9f2ff8a80e194736aa452a5a9a5371ba50060027842b39db07746f0ff61f5b3833196824992de4436f43058b5ffe58f69da0864b419a2b0c41da6d10ee29cbfb0f87335c4ddd;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd0b92bbd1a499ff7f773d227ca7f0c4419880f8985449ee8de50e4a3cdc152b333aea1c2353a69f05acb91d18af7b3d9049b4943ac1b2dec8ff532dbe0cb3b7931abe5fe92408a95ad17d249b0a04517913c4c2c01cd60ccceb200bb7980b4a52e7ea9a7e368e3b2a5;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h16a7d64afa0ddcbb6d785580dbb3bc972af72879476e9e20129c9809ee41be6446a3edaac4112dde0b610b650aeeb260282ff182aaa1882740fa79f0d5116a771686ab4be97091314543b580d4c2cfd31a262dfda5937ed27048c1f43aed5f52971a7605fe33ccf96d7;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h259d54b16bae835ee6da2f84404680f848a287807ffb2fdf580a6e9f417d8cf16120a1e31ce149501f221af71228595eea3503d5eb5e7f1a26603c288a75cc4d867a831e30cef20101245288bc6fc67172df6f0bc6e18326ad12ef5a94c35d7b406937da978c03d64d;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h9326714c2dd7ae2b223a166d86e46408b7d3dbdd6e7f70552e967538702e0b6062c7b508d8a61edcec4d89344b2757abd19198717ca860eacfb546f42ea49970c59fe223738c7cffd6ed793d94317f7669a74d92f0a011b5ef0513b19fdcd566174fb9a59b5bb69b86;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1688dce9a2df0fcfd003009f578581f8b807140968f61083711ef6087d97104d0a572f07e1fea41c1c2099ceae28895844c0c0f5680e8bb07e3617c2913951172e7873fc345c04341c5924de3efb57982df2446a6defeb2d740030f10b57a8294483bc4a628ad6e8012;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h33cc28d1643134ed3e704a4f95d1c0aaba5819d59512acb2925a50472153e367cf6e991f5292c9ddca698fe63bc5ecde366bcbf8fdde129b4650e52f7a502ec299726faeedb83da9d2b840110da501f96aa3b21000fa4977dc0c67f29d19d56347426f6b8ee270ad40;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc115dc953b12d0a5fdad3787c24d7c15a4da91c01235c0ceea23465685239c420720f8e3a633d8d19895d9e29f2c0cd8ef7bc86085718edf4fee09c8034728725b90929cac27d81081b5bc485ff1b67e50dc6e08aba6cb3039abb1fc75c25ca3a2c07727c14c4fd28a;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h180bc5cc470f688b5b551106a66be1bd195894d5d7f59b708907ed2e0c788ae16e0e068cde86a9a9c8e841f31b7d69c2988db9792b930e5ec7f9f47ed2d94b76d0a888bc408e0979c29ae38ba834a174a094ac8755ea57f26a40ffa05f175fb1c20308e755aa898df89;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h5ba4e38f80cac1d03263e05cad152a160a597fcb3be2e4d976edaa7328d7ba58751ddb43325a12ffa2c9da76aac4c32a9d26cbc42ff49284a835dcbecea4fca75426f47513bec79677ee963b8eadcb6c8219c965b556800347e6a9ecb9928659fd04d8620e0d8f7a3e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc9cc16e2ae8aa604a9b79786679787773406640b748e5c2d9573debc5166ba9141e8cfcd6cda95011ccbb6634810b117f7437693e14d32cc97370518b1dae6f25d9b222dc02d2e15377147c69edd98d34d596c01e33795a692cf103e7429370e1710a514b509269e6e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a64e40bd4f0c5591345e84357843174bf5dafd25d9e65539e9497127ad8158fece52886fbe04db362d2f8b8c229de6dade0344eba043031bc4a348fe97d59d2e229a3386709174da52a8a7e643c53c182e472f2db32ee9d23fc52a29eb7110872d79742e2b24669203;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h144581a2de6675f47716bc5147ef85b251cfe3166d4dddfc819f44bab84cb36615d87951ebbd1ea77e8c0a35687ad0cefedea39aa0fff11ee144b3229fc525da7d7cd7cf3bde749d8d0b8a10b3b372feab65a379ba20416807e9b758548af13eab2e18e64dae904a12e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h26213cf4a54242f71a3214fa8a6142bbe16ddc3f0bbccb201560ee5a2168010de848fbab13fabe52972e03657e94ea7833471ff29ec00ba82d6aa1b5bd9f52427e4f3fdb519cd23a88b73aa5635e5a79b7e144d86869ec8941f9502bf36f48a94afb234bb0cba2b087;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b7aa843cd29322d77d39fd2bad581ed79f6cca0e079ff0650322a45afc2e0d08e81e36623fe0f11bbcaf3c042e62ee5d1646451876c39933b3851b63ba108dc100b543394fc614bc72ba983696f5fe9efe4b126c7602683cf4a735fbb5578f2cb36b695689fc94dc1a;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hfd56360960220ad5995429ce3308f5abeca73d9a693bb2f5242a19cd887301144f9633eb262f253094e718c107600fd02d9f9a492ed84e8caf3010cebedaec55d2b9dd4dda5f904ed6db86235b20aa99e0fe8d39c708c694199418f02344b346301d3945561efbbaf5;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h18d47b268439d0fbd65ecf775bcbb0934377384d012ec945629dcb138f9b7df36a1b0772be177b224df957192d4b5d89535bac371efbed53ebb14e049ee2650017787b66ecad482b4092c5b2ce2385b79e42a7236119398e58bfd1d38a4a5b95346d8ce4aa6568d1265;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h14f1b4f7f37b21416a8f7414909f0cfa516f7d73e660e48172bf0a7b71811f381d3aac9f2aae17566ddfe126e3825a6cc1d0bacfbb534cacb0bfb49b44fa1be2f491dc173f6922bf61a05b3c7227ef6a2b6d188a6f8b6f2f7b83901ef2db6c3995bc266d953c5d85823;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h4f86e7a971b5cb4a6e7390e432c08213e07cef5e2886024dc79d7c33b0cf9b7bc35c5a2085c03dddaa415f0bca8b0dfb1def23a669d1512bb24f983bd9d99fa322c0f6b24fd08b0abf8e0a731c16cd6a077d18d436e8d011c9ac6897ee042d6726f2877fa055837629;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1fff811e2d900bde9646e1dae9f0498661aa711134ad1382cde9892d2dba8e8e02156208927b67ebca15db6ef7b3b8aedc3395430d96b5557c21c92e46ae51739819c53f3e2b6692367abe8f86c30f9e16684565cf16fbf6b1b3ecffd7d7c7c1b380dab53366ffff998;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1617eea5549f5ff72f021bf0f3db8c6d8ad3b6cf7c33fd74a854bdc1b3c9021447fce39ffa75a3a9d46a2f951ded848c17727c78785c85c56b6c67b82b6d0cf9a6378d5307ca2ec5ac604a0a3c8672dee8cbb1acbbf3f1abe1f3182c518ccfbafb61de7a72277eae75d;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a27da87c14997d2f522b732ef0c4ea9a8305cafb523e53d9106002158680373ade4fa6419ed63b7147d8ad55b76026ee7dedf1e014e01d8bc46e1e8484a3be3e8a4d8af0e6713e4fd1dc743d5630f66d8507d472a4d2b519e922489776507948e2945a595215379922;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h12a82ecc6b690de2e6a83f56890892289719d1c3472f46677ea1fada4d1d651184f233b833f367e476870acb06e0452e211a1f17639cb7e9e6149ecc82b64650b9d9a7427975dfdce8eef7520821b9c2ea8f35458d5fdd063888a80ad198cb6748ebad2318560f4a226;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c12928aa8ddbe6900ffc294d8531fcb78f702562234e4e83ee10397b571680c8ecd31686d5e52f92194e63ea35c70bf4135d7d823ce9b8361102a69e0aaf3300e658d835567d55a1b09d082b70862117c45b95f7548a2794ff803085b72cd70e238ec92ab71311d755;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf623cec66fde58147385cdc49960da70559cbefc6372160037e95c60ef30e4329ba3809a3160731171cbcb29196245f63076174bec58ab1c80007bfc18fb050aeea9a2039d62c1f5594ddebb620670c239eb63f50f77198f0837822876e73c25265c28b8053ddc9b22;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he8e1b44086417556f85220aa5ed752bde69efb792a0b7a0a2a02b5124f58f65b8834c370886f7a652a92aec5d7137c287052943ae7a9aed065d5ba0e06f0e4638e9c65dc2fd8b3e5a55526ff3e596142663644c39492c03b900d058637d5be547593151298cfc2144b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h3b0ce0648bd52a416509024d2eaf4fbac9940a004372e3381935232a1d8d9f5483b73e1f1db5323e595132e9c264a3d0d7ac209c6a63e97da4dd5c9914bd90f97e4f9a6ecac9bbb319c23623282003a63c675b077424a8e28ca4de9a0ca508df08448cca5e10d917c0;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h578e7218020289ca9a26c4b2dae9d3048fc9d0663713d1ed81ca39144ed900d005b557435a537880882f3acc9596e336bae8e51af3e3be7c7e5520026b1e8b1c2c6d4822b3db137ebf8f3f65c4ea641ba730e84f9c4910002e54763f6632161c1428147ee17c723069;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h6464ea36de922dded86b1da65fc3cbfe255888d5c7b267457867f5fc4cc7a619a44407358de93b27d4a84753a199b7a02b9edbe8e36d4b89e2caee7776766d38f9dbc3969d4ea35a9ee9056866431dd04b374fe574affa6c15b4e12b537d284652be529a294cf454a7;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h929b884188e3c7c97c8fab68580373da1b06b55d9bf65713274fa0f63277165279658ede5c1ec0383544eaff4996c3f4e7d846d6b480e9ce4bc64d6a1b559048d6572e68052784192d4c4f9896ce6ed527c207e02f6456c2316324e646a7184b5aa1b89670db1fa7df;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h70cfc9be7c91bc7a3bae45d3c72a8235cb91175874c3c59d94dad7ec109e72b1c162d79549af12a4fbe016c1603d0c333a4da623dfb9b13ea3ac9ed3a9dbc9a7a74f5938ae6d68cdd9451dcc92a3aae9c31facea4d5d8418132c6b91617b81a1f787de4a69d9ffd8d8;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1fc26f54e16e5745ffc9e9ef31f4ce6c20ad219a635f3a83a4a6fa896c992512b323102973e8415881ab5de47e719fb5d1a5244a8ccc3e1dad59efb76870011eaf42797a8d5280dd1df38ac9a5c4d020fa38b15f16b8608e8b6b039c5a953f9b043bbdeec0f577d8504;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d81750b8371a7984375fbeca7f21b52c0a4fe061f594c22fe292cea71d2aa9f5455f5024966f163ba2653c44f4f9d67f5989f63f4f878c9bfdb86c55ef890f779ce93988e072ca77218491ca381eff66d32a44478c0d670d141167691a71c5baed90a12ac4e4bcdee2;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc519b71a998f8a66ee52132b4ae93022dabaad1e44a518e6d6ea557eaeb421f2e77fbfb9c29024d51b6d47b121fb809a1639eddd7114ae0a8b4f5386dcc4ea9044411ee5ef02efa6bcd8534fa94234cee62468c48b4cf645eea948713608aadbe0ba93eb0db4078ece;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10909f94d4de4973fef8379e1defe1764a017870b65ba1fd03b5d2c4d327b201721e3307d852ae0e66cbb00bb63ad9f8b181e286e3a561e00feb2b73cd23490a82965c64a484eb28576f38291de96116cebaeee6ab01cad02e057e612c838e08c877fe7af3e214f78e6;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h3d8d62571ee5893008a8b58b714a5bd3a13e7b03d6061fe8d2b9ecb40980d5c55bd9c7903a752ce02ffce07b61f89c0aca1149c26d36ddce6b9e1a5c6d3252fb622ffa41b2ed52ef3e0586ad9ad9232ab88d6ca1b895fc68dc5bc845b9a48dca1bfed0caadc910f3b0;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1af55fac41d7c62ba4e92106671066fa19f0e19260d0840eae9c1ac84c8918eec020dc955a02504b7df14b8cc089e46559e377cb3b4928942cc9c3f0f81df46ff57a8713f8035889662f86b1fc3bb23b2fa1de8af73833b9168f796674db14afc31c2c8a38b36f734;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h9abf452059a239a2c0c2a488a00215dad4c679a3435eeff5a8b01372a35cc8d70c8066e135807181fbba867b43c77658df0ae969d8752fb76f13c605e147ee8294b27a6b4171c4ad4acbcacfcfa6d0eff7b68c1b47bdcb2ec0316530cc4dd24942b474061584bd57b5;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h19c485424c99fa43da9460dbeca0deccf008250755d4e400b2451b96dff13e3a9d85385bf43912642abb2f87bb5fdcb24f76634c0257333b388c4c82e3860e68cdfe9310e26929b6eb3d63e3cd9a6b991f4571b6d58f5a203f86d41ec4bcb892208634f8b9bb69f3afb;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd612c7295ba9a3a1fbb15b32cca543f2ad33a6d166d6787c9939bac900ae32962277c7443a1691fffd6a7f0c2bb34010ebf43bba99adba1b061e793f7380313ebe5ac568ec6ea95a0ea2bd3021d86b0fa12e928136c3e0540966a1b7798c0a5860e6b9246704da6e8c;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1988b0327adfadc5b0beff0ee7549678d988fad311e2164af839a644a4fd5cc10f4e49872a5b331fc8434dcd076239c0f3512ed75a2bfa4df4dfefaaf136f235fca0459dd6291d3f8121279388c645b280bcc199a3b3aef5bd983634d2284f81cb7d4db315abce0a787;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1bc792f3ea6b94cc0fcee12c9a73181f04c2ff799c67668aaa081bc20603ab9272bfdb816daea1afcd4147c69281ba0c2920337f52defdb5f2490fb37dc3757b12114e38b04218b8611517bb7d9911589e15094dce4ddab4bd615dc41d188e3384fdaa6a4d95ab80663;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1afb506c4beb2e364a737922aa36b27b1a320b1e2faa19e553251896c08d2ec3f9c1f1976a38b75718fe5a53827fbcff553ef8b163dc9825cee21206c5141d25f3a1be490ee8c9dd56c44933c14aeed16744e44c8fd006dad33200c023e17aa0252551e3555a54bf466;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b8685f9758a883cf0205e45693af2c1782a18fec17df9f866345d544c6a79aa8c18dd8cb2395d1fd017b7e0431bd5ee57b79c90864430ddd2f1205434b8a9d1085b94ffe531a5a7dadf18e9c27cd83386f20ebfa7904f60ff9ad5170aef490ccb6a2c7514bd8cfdf74;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h5a86c4e58d2cf3991dfe31c464f810ee1761cc91d594a169fd78a69e1e47806bcb5e5993dbd0057b076fd4654b9ee9f40a65f9810773c20ebda41c499f89eb356b1a92f4b9142f00d8bc10ed8c5e3cfb8114f891cced5182ac531d2a34d259dbaefef9b98bd5cb300f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'had8169ddff50985abb4d648d82f1a2b3cf6e844a01a163928091d5d03c378bb95738592c9627e2563f5728ebcff86605977b396639f690f8dc91216ddfcdeed24c0c0121e812339fc2b448785a08d2217784f9b0c51d49ddb3704bb2cf3b5a2249de23722d56852db6;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10b96a43924ece8a11c78253e1c88d81fa73e0031b0f144d55c9caf41800627ee4f5bf7d257fad212ad6e63fa90ffc0bee66b6a73a5b6d1cd2691f71b5f32c0ff3cc415e8d9d4672aad6f08b340c409332bf7d5a44a1b53084a2111c03e326ed40f62620943e0b309a;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hea28c36976f879ab8bcbcce2bb5c9255570cf863dcddf4c7b69a6fe8178139f9f9586c885a05a143c77a4613210b451d3b9d960b3c14a87484b25b06262d36fd821c0cfbb8ffd1409cacbfe4d17153611ca885ed206a86681544c908ced43051c409de94cd26a63078;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hbaa39fc00c8faf65ad4c04d5ecdfea48db08a0c1deafcd006c1b196870f3f22d56087a67e30df015a20032614ccc3e3e1958093a51bef9d96c187f8cb13ba53308a8a9f4fd29f17c59beba47219a4741b0a8d02f429814ea1dcb37a849e01d25574c7e7b501c3da831;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h12500f3b75fb36b38a81567b441299043a45c815724f2e81bd40293f224a4825a26fa035b47190931db7db2d7174566489af739576a8ca99490c8572fdabb6ba5a1c08fc52ac41b0037a7b4bc30cdf4282b2787648ef3c92be6bc9df43ce4a08e5a083f03878d7c11f7;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h11d1213aab0cb639e9fbbe51a447c4bc1e88812f5626ad8dcc44870bc33170b85f410f34cde233db1c0d863aa33ee203825af897c9fd865575a19320f737508452b9442a56a1a133ed86a9b245d6a153ec6af7fae4c5ef8f1dc96d5bf58837a22b6fb27b86898419d51;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c7a0c725bde5cdd9a035c92d9af2b4299ecba446f495313b6733e963f47363fc4905d2b6bf1622c1a7f5ddc9a202641fdd0572a7eeaa19b25d4e22fc4e85fa5c1103fd4b6b4740aed0d788540b6482dc7ec8ba3ddeab48b675ca575a7777fa4970bb14a5a5abcd6b1a;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h11759489fdce66d3797bbfe3df0a0b060d643b5d9827441c30ce81235fb53430bf620a1a19bf87445d68698ba072c3617600690ed85efdd658bc2eb559a218f4cd5902802068ee809fd510b6563bae0ff95577f7eee38c59b48f898a592f544fdc0053fc2fc3c00aaeb;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h16280e1ced11fdf352f5bb661bc6a174ca07f6ae55d633d54dc4701344ab5cd90ce536fdeaad07501eb0a7403ef50b7d9f195a3511fc40d46ac51fb481d0228ecaa56c7f28b7dba960f021df2dc26fee80adbb9dd46e933ab46fc52452b00e8b20a709cced665ce869b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h100bf6b4c870a65d1bb326327b7c014cadc57937b98f45f84118439b92e0cc63d989239c3e486f92f9f7a5ade184f21110b9aa75641a360272326bcd72032a9c2cdf60165f3358eb0240ef110c34f20ce3d0d48eb38be7c1e3fd68ce99f795a7dffefa35d6aa25a5a05;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1dc9976bcedd3810bd2843341cdf5dab4d342cbd54fbc77715cb35d60b135465ff272901e6c37c287d83b15b7572c2f5b8fd34fa1588d7547f5c5b6f98387da199635246b7565743d5eb9d2485b07ef05b954ed049feda7eee97d37cef2c297785eb30a3a170f189640;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h141c7ca7632731d2bbcc720fa2dac537211ef45b503d760c4ced8fcad383d0100420c578c7afa28fcb5feb1de27faec9bb3e034ccde0c25dde193affd3d28992698e96c983a517c95ede06e5987a70ac9c17706abf2847b2cba7a499a0e107e5d45006bae282bea7482;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h60decd2472889655457129b422db2fecc1059d3416579c3491157645cd549137b42032a3efa7af98dacb7853729abab117c6f8dbebd719d5edc4dd0956925b1b1f5f145321b7008ac080e37c2d99783106f40b5c06b03e4a981d854925fed18ccc865f58628a35eeb8;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h34fc1e254ea95e2c92c8d6354a1fdcee46c52b4b796c29780e5a4ed78bdecced853caac0edf3fab23a42b3ff51a5bbb402f94700e3af8772d193a1da843de6659588dab825fff9c1e05a83f8aa1f6d08fc585f864a0f59ce845f42021cd1808f4c9cc539525fa95972;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1058deb6a97b5f30e3ecb38d038ba0fdb536dd8e075edd426fb17b64e60da1c9131fd16e274b1c4e582f55d243a5d3a6d439050223aab3875e46c8a4dfff16ca871da733a73b4bc19875e4733bf15607f70ab946a7514c386bd702bd92af34f2a28d84290ee35d02baa;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h19c043c2bbdada73c7b9fff8a65bf37372c0131a2f72d250d206c6b85eef65f6557f76e59396ca29cce40fd6756340f135575ec6c1e24650c35ae8c91c75cf0b898d052b787e8ce32c1a0d18969a5b764f1a09baa18d0c082d71b524e5a972854352c18c20b48de297c;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h116f3fae9105e84fb402be9d8e2055a93c7568f81b49274ade2da04d839b806cf535f2c330fb43a049ca0604d3814f78b18969fff80a6d14435a76f6c1ad9be0e5ea9efd13ec1c4fb2b35bbb8b4c68a27157d3b0112cc1af6310c345b504e87dbf469cca428ba439a6e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a892fad4e871c7a0d93ca1c90a115f76c56d7e163308151e1afa2cbc812fe6e58d03b0c7c8d7249708bc7084355c9adeaff9c14acc1527de59c6b7d07f59c7aca60317219c784f0a7e90d3bd3a68e8a879a08e8a9887c837bb1a8985d68d5da91c11201e1d99a6ef8b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1dff764af2c497d6c54d1b6f5646763fa45b9aa205d8c324a150eb1a988e86a173d2aa60ecdf35c007ed4009b498877b5924edb72504a570fb93cd8705113c273d1242fc5fa76f7703b4f9f975ccac39aafc0155b2146b513593308f9484574937a496cacd2792d3b6d;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1cbf4bec7dd8421d9f1e393636364d1cde43e0f5e169a90cc4a41cf1fb77210a1eca66a56a0c3f9419b6cc938f47872e74c3e503fa6ec0be3ca0271151aca4ef13676dc4c9951557b36d1bcbda64892b4e553abcb5f890256f3be499457d3309ff683f27230c9a5cdf9;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1019a334f25a2a75187b1489db56c99b0ddc832376832d3d93566a0e9e89998f27cc93438470da7fdd9f4307409c61328a4e44deeaf45470f34df29c03655f16cf63f1e52f6097df3eb512fdc19f79853f525b27eeb3817d5dc4ab07c0647ace3113585efa2c8d08e08;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hbf53bf07a42b674c7486ce948cb699eca956de875a35afb514adabf9da9e34b58090df41ada21812f9cb3ac10711466952850009f6ebc3a5a3f1ceadda25e6070cda609300c63d08af7241782208464a18d547df73ebfc5ecde5f760eeba85e3e98b1bae60a39e3e37;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f0d77169edeb93ff4c65acc04085c1799cf74167be014e8272c1a10674286121aaf30724a34142e4600b2c38604c9e633aa93da8187c494565a40f51a1585cba8fd3566d03ac657c821cc9ca64581f12d6ac93764b00d5553b226d9660de45fccc2ba04d17e65edf3f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h25a4c4ae1ecfa03b4253505dc58e7cc69b794a2c321dcd36c65a449a98194d2cb1b7cbf4c41142991a01c0125365839774f444a554303587fee0a97b3a45beeb7610e70a19d0c09ef21fbc441e087985c629969373bf419793bd605f8e256ea5907302b535ca68287d;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f8c385cfdee93d4ce4145ad2979d46c349489c295a0929fcda53f8cc2123188dfd787d636d3220b5ee1209cb8798d99f26eee9b3488417b2a95bab8735646c36e735f5de8f6d9032f98984cc97d0226f4f40fef16e42d17c47e6649ffa3725f539db23d51a51c7d318;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hfff119efc8d0125e639475ad638e995b2d1e55099973fa55f038395eb765eab3c5863afdb2bcf885c216c08a7749b9ed2e46ac27a9381cee7d567a0711cf47442c3139fd0479f8598ab62775fdb7b87b9bda8292bc9ab4ee5c8d601e10aa3d59a5428498c66c394657;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1265724d59af12957153ac6553ea9c32d5bac3b5f48c98034630abcaf07dca60867791f342929644131aa37a82b49786e4c68d1be4a26868544b61f31ea3786d5ff44ef362e983be53d2f219d84abbea811285c4917f8a26d6398aeae93729dd0eaea2387c9bdf4cb0e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb4e386123f03b9183ae2f49e0f8a3eabaed860b25d4a9949bb1048a523fd67687ff669127175ea86bf4898d2fbf825c001d4631813070627491c0c37fb11fdaa732ba1e5e5bae4c2a5b49c7f6b37dd903f0bceb76f24976e3b8532e0d4db153925c8072dc6d74b4a99;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h111cdd1300fbc8ec18221612f6498552755728cac7a47d3f548fce978cf0cef5e2a18ef7a15455e10b1c3e6890df6bc904477a8627d9b78f98b92291a510620cac5d711c1233b7cfb3516af06afc257f98157a4d825274e439a62ed5d687c331d12c1aac3b7e0d3077f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b06e3a7c9c3bf647d8993aad27bf3795526c389c2f1d70e1885af9f728daffb72fc3a3cb83c1ece9d4a7b064f8d7c6645dee981adfbea2529361f996d50b5cab7bb0f8dbbd265dee20f03ea52193f22768f85fe44849ede61dfd118b2518f962a2a6e7852901ee721f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1166f55311830175bc0a716e364aee569fa39a370ce42484bc2632a440c80a36e48598a277382efdbe9093003ced9c0ccae2985ea71e3e5e34e8a2750a18322add236863c03e834682070d4e26f5dbe9a44c6c7c5c0b8eab879ba4ca94876cf439bbc48e8ad2121a77a;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h11f655b6db2637a6916e6bd88373a32b89090fc2c26253e7167c7ff059600ed87465daf9d68200ce19b32e1959b7c1ff9abf9ad189c21c572640d065989c0773a744660e8c2ea16a7ecba953aeb895909afd4d6db844e1496e29ca9a3332f3223027be5ed0c9d05266;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1223e671ee6ac04515b7f422fb8840cea41fb46bb4a4c246a0f7bfa979afa500cedf70e2da09de5c8deac6749654a2feb3554325402939a274680589e51344cd6b8ba5da0fb6000cd2ac5e9f9ec2de7f77237e69df2702cfef1651646665da7bc8c966b0f208f19c1f5;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d1e47215336577020ac9b875bd1e720b4b35042b7b23a8218830add2a1b757fda0f9f35e3bcdb9d1ee6437221efc08a73ca448884881bb57be570b738f748c7ca76f80b0b9a52b0db36a1a9e188387e6610cbd86d913486a298e3a9d326aabb10a692c5928eae4cd54;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1761918681bf232a4ccb0fff5f27ed46c2a10aba017dfe87370d90f326df1a290e23f2d5a93d2c67f1200946f45f4e8ad06f179c611dce8020982191034ea67ea23c9397a80df7ff8e042a1ffe7c435deaa428098860c086c501ce1033af29d5ee4deae88d8664ea360;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h18c326b5b08fa0c794bccf6357ee756649a4447566d60f27e8a1fd8da6343dc1a20a24f44c1c7c3f1a8db819c0124bad497ea1b1099dde08b54bdd49237e781248db2431ffadaef493bd43bb501f759d67d8302e85c95357f5f51f9617818b14d844c725dcca26697d7;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h14563b03080b5b5b4ec63699549f113a705b4c1acc6b7ba1b8bc551c21f5da405d1fa8aed3a479125f29782bad0bb4e584d0c4731a10ecdfde5a9fa9caf89fad791b8c7eba3d7c5c101520539c6e3f24ce5d563f223df9b00f9ab1fb90daee44204dfb68e4ef5fe982c;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h19f46a482ed2d5e519c01a4e33c4667b2b13ce68401f33a220c7972983fec5a992195ca94ef725d358acf092fd385528ce62a1e48732257a4dcef58585b8d0e3c8ed86876a7df607dc0bbd8dff5667f943bef249961f9d2afe3991da0abe40066689d74dec31ee08be2;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h11967b8c14f1fb584f557cf62083aeab71a50659d60b5fdf7b6310f0c15e1024a6a984c1c0ac0bccd768ea1ae78438a75fe248c56f46f0d9bf838de92b5657f51ff7b195b00c2b6a04988e20b9e83cedd7786503887633af783e0b0f63839b0159c4dbe7d797b399b2;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hebc02ed7ec85e5acf3f1b238de0448af9142944df90e7d9f9cfe7dd4533d6497656edea8195502bafbff34723aef9e63568e0679143af99bdb071f60ec9af6004db8300755646708ee54301aaa28923769a0c47c2f5b9490131b8d84edcba01abdad924220be32c70b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h19014c8cbf5927587cc9ff74f7863c8d78bb584c76d1993a98faf0b76b37584990f2d85ca70975b7f0bd46df60ce8b209fdb367f470c2565e726dd21b3f7d946f498f771fe2b52944d76839da35e7db1f58cbbab7f6dc07f6a3883e04cc00b544aa339b07660c0ab453;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h6d8a5aa50f06614e0c57ecfcffcbfead6423c422c9e05cbde31c5bf6d24271c212f7761312bc30e964963174eaba3fcb9072e2e85f81086b70f8b1f31e334534ac530233899a9b48af305b50a5cc6c89ed929b01dfc575398082282c1128af4c945b24827d3110bc74;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h118fc09cb9e928c8c115ceb90cbac46ca4d5399f8f6eacb9b52794bba9dd5f6936a02b1595d80d2fd63480d1cd5e4cde997dfb2490ce9ed7d2ea12a494f813736d8773971b38eeda718e4cb161822ce187782edf376faafa21e85fd7f809ec2b8ff3e9cc39995d0a0b6;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h574104f67715fad1c300d3dc4ec8e42b4e107e448f4ab9c593ac58df0cda2bb71761580a3be8d8f25d4b6f0426f3a4814dd2ee2610ceb800a75665b350fb736b69de18288076266ec3e15cc822db2fc7dcb60fa4e1029ab79929819ba3d3cc134ffcc0752cee424862;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1daca2489f49e5868ea39599d6dd2e3b10ceeba04ca3ad96e2f86b50253074f0e029bd7648d78610bccfd1b1111ddc994ca68fd7915f38a96f2eadb54327a9969ddacad395797cb80600eb31e831fcc0c61ea432c31ed254f0f39b9157194bdf74d968a28b9b5a66e09;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h95fa5a49423e3371c56df39b2bb884036724c996322f769521d9827b4e4f25da8ea212234a873dcbab80016feb23f26b5973a97ef1e442e06a722033377de1b30c47d742fb04fb209fff5afb329dad7cca897a603bd8ee5316ae6a876c4ff536ed8fb80626e40f0a03;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ee1f81c783fd2988c26962c29e66137115138c1acb5510304908e73664575d1776fea6e644f3595cce4522fd838e282e3cf0046c82e5b8dcfff0cfd167becb12879fdd866826b07efbcf9c4eae1d55ddf4cc7d556abaeb0994c3cec4d388b7facf1e1ab9d1061fd274;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h142e66aa9c38e02ca8487a3a00f424760ce826a7c6bc524339e423a17b598711a565f99040d621ff9f350f7d0b40f6a4fd3383dd24c4959e8bb27d85eeab7f37156bafdc251aff9364e56f3989fe8448ff73f6b76e83e8586bfd389eebcc946270944f4f7fb4f873fa1;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h493708ec6ee092e7df5277709c95fbfdfa3c212a19c5ae9270a4add00f10d75f5a8b55afa5ce306f265171c4296f7b5d83a71396b58603f236cba887a30e62813547754dc3662d48bb7a0412c72c6ca5a9797a4d16549c0c202b33e86a4c4c3aab3ab0a7c497b8ff73;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1fd38b7b0f801811df3874522f465df2505105a5d074f5b857b7b2cf65f19864b95181657ad9c549be4908a47f71db150883c28c78538a24e8ab1c155dc1e1c1688ff20b6caa0bdc6594de85ab1f3135cdedb03a49058eba5830fa11194ba92a0baf6dba300718951df;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h15b93c431f7a22e1924e455bd9bacacee4098528370b9816a831c67d6bbfe2132d16bba092ad9458828221d0265b514c6388127592e5ce29ce71eb73da7ecfadbc161eb3fc99bea63068c267318974407278696dd103b034e7df129c82e48675dcf5452efacf2359ff;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h165c3c4938ca12c974086b6b6c236c2db91566a110435a4ce64ad4e99725706ebdcd57270872c524fb316618134cf9c9f6789f892fe75b04a6a62b98090d85dedd55f354e4f5086bdb288537768001497d4aad99be81e7d6083d0bfbef6f8cd0a773a950995acba36a6;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h4f3cdefae0efba79316e6e3f81189b187d0a33a72d2f5efced45b9bc3bcfc3cf6dd3956d74684ae6f5fc9fab72431faa807162dde098b2f5b3947b6e9e58c19348ebf019482492132e6b7edced64e1f630194d8b5c8301e07f7d3404bc9139ada2cf75477863472c53;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h16fb15a5ba81dfd9943c03faeb2a131cfd302c98941fe6d19179065a67cdfc9fddcdbd1f97311056a59e180ebace41b958d918e418ec35abe4e9b026265859ea139384bedfa46835b2d5b396cdc0ecd1c6a0ad4c8401f4b558d3d4c66467e69eb3fa37e664de430c8c6;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h59728c29106c1e2668e9335f72db4eba46a00349d6c54fe674c02a48ac4ae9ea7c866881069571470fde098e7f6600776fb2aba3294f114768da1831b075599000e0eb1ef9e13cabe95dea853407e4bef6d127bb5fc18042f84f8e548e4864c365fc3f63e17f316f86;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h133d9d1240843d27a8b9b7c77794a584f36a28a5527a6bbbe855ca31a0a4e6e08f90289e203c05616d50ac4ab63b9d00e12bc040399ccff815bbe367447993cd8dade0c54685571281a3b61cc265a7f02db3e59386d4ac3773a542e0c2f85238c08f4b906943e3e7fbc;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d42cff748f54e2ddff0baced235b1116605e5b97a89e85c77d6e3afa2718a347594b4075bce96ccf911b1a02481dd54ebabd36d2ce9d695c258d5b01d6584987c5be5610ce154935e72534eb6cb9085e77b9d8c5c851b3bdb73fb0e69737ee88bbd5f1c993ecbb68a1;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h84aabdd89b0eb0c8e490a44acd1fb6b023872d57b2b849509b22f7cf0c1f79af7fab1d79455ecdc8b9b8310c9df4871c29feb55db547dc0fd7992819efbbec1013f388772eef9883d5291b6180a1a2aeb6ab33e813296427d418a92b190de0d7b1f890577979cfe02d;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ba604be4af6f764633ab7fe372491ed10feda53ccb55051ff59a9c0f95dbacf27887747833f11a3616a4c25247dec4b61af8d7c1ea5f2994b1749ed962bd056049c66dc0ba4ae5170ce61a38f9aec31ab77976880f45506cf98169057e2a84899afbfc0a39439d86c;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h817bbb378fc28705e6f276f65dae2b8eddf1b93267f3964e47294cd470d612ef39775b55ea5679c25f063237f39d7f0e104b98fcad7da278d4d3f91b3bdfb479b8268f79c1ae4d773a5518033e13747bc56216c8d29c64013c4ae052b7c1bddaa1584b045a1dae77f2;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1211de537fbe616e21f68f7f52808873bd61328e6a2781125f408eb2ed34970a839b0d0de30b6719d88c640e9564243ae14d6ab64b965876fbaacb5eb2ee83e1c1c8093f94c51cb14258360b0fdae3f5e53d95b818d2f622494c5aef9b3744c90a8301df8f30571ac7f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d636e34ef59448c4e04fd83bf8e2466293b8db8ab4b7f13a793815d05de762cf8abbb2f453e5cf4fda582b4666c7ba31b9e9986147e19d8684799c6af1e44d73c2e4453ed99970e2e81bd002e15989c6c7e2c6a618adf6bfec1c42f4ec5f4a6dde19b361fa051f73b7;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h15a15a3b2054d5bf032310736064235ddffcda00c610533786c86ea35943f2bd48a07802c3a4bc83559b2bdc44423173a5e411721efdf7489bbbadf567474478105aac896299c003c8970cb3e316c077792bc96c53026d1f5ad3240c7ce5edc45d5073d1b52bf03dea3;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hda626619a73875d9dbec5760128b30305791a982f2cdc098ddeb93274d50d8980b61dbfcbb77b2643a095d397ea248a71d977c088cc2489f7b7821838d2883ccb0506f59056d160f00f79f7c3c6f6d65abedc1b8e50c0c473e326948c540ce282793b056975c216bcd;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h19646820f551be53b28b5d624edda8a0c8a7d3de08a05a030ae599d549e75bdf5810cb706deec62f75e4e9099fee9f6dec634cdfb53146e296155754adb83c0fc1826cc67dc9a5795eda5ea8c9dce6a9c25ba7ddf90547b44fcbb6be8f041eca98a5a9b18f3320d7dfb;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h863600022da92872c08f1b3428b70f6cc206a6b6a86338635e17a54dcaf9825f6152427b1de59ec7383d50dc79e8e184348e5515d6dfbb7c4fbc6c1820d97b0b505bf8b08175020c17b97a3dd1bfebff08c45c59ec69f694690b09caf024181e856cace6822591d6d7;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf30ad01ed7d1fad55ea0d490c4bc17f203d44180026339934ddb2e527fccb20cf867d6d4b73a6f67ce02cbe7efd5ccd9772ce9084e19cebcc4949ee7292025abd03fff5dca640f9d1e302dcc964523c83f704e3212f1427a8dad705cc4115a04b20fcc57b7a7579358;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a518591e4e57d68e034176ba21e15fcc37db44bfff8109f6cc05946e01e9581b44feed8e10b2bded5f839716ecb0e337155ba40fca5164086e4588a6b2d03e5b2f86f10aaf4531da19623b90def4e36e81d133e1365690b7ad18234d6cc380abcd77045a03a07545f1;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hae8caadaa5066623a843173250f75aeb15ddac845154ec027f59c4aa6d00f01bf0791f461f147946eecaf8a5aa793679d2d9bd3464eff824d723f5b6b3f9a91f010d267a79064c40cf477398ee7688c271ce9d84127459d13e1d0cbba8071d620294cbb194315ec9ad;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h57256fa91ecd9c95e8246ca5d9337210a8cbf2b78948b97d952cb722890bb1493e7f2790d8dfb2aab112181a7aaaa53cea7892a5ae091e297b0bed2dcbeccf8de6ecf95cc512af46a263ad626f14d610aee25835744fac7121ad13495218d93d1c39e55c0e41c7f99;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1fb5c6ed3443132f7ec3c6020104fedc4a2e5b4db6b78d96015cbdeff5b81a4619c3391ba27182f12cf9187a71afbe1f9c8ac995755f7d2d057a9b9b209d1e06f3a7b99b2133218a3a3a5f1ec2f86875f7a0c893c9920a6b4d564ceb03df8c1a6755de24ccd9a5da5ea;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h9dbabb83b93b8e8794f599e668ae6d6b5970841edc9d346ee359294f908b9ed88ed55f9d497ed8b0245d8e7c0993eb8cc5a9c0eb8954a7a70363ccfcb2d20041c2948613a6f4fcc1d791c501adee069043d8d2dc4d961d09f527597813648b67a55efbed433f80562c;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f9eff6b3d5dc971133bbd2e877ff62bf7bc8bb496618f9502bdd09cf93ca421971197f99d6cdd93ae59d81088de97344e2de150242ed2416e359293cb575e9f7ccc3ac0ff9fd0345a4b597c00d48b77d0ce6e0b468623ff207193f6a29d0ec45188b184f215a7e85e8;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hde9109b7b0d8bffa375c1b9233a5237ce501489de8937b6226ff53420612e51c7b77cab9906f9a7760eb5cc1c55768511e3ed2959e19bf17b8bc43ec38cff5cdb85ee81ce79d2104273d486d539eb3828d8d9f809e669c59e02e75cf7b810c4a950887e9f41aa34ccf;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he786c8d84d562e48ebf102ce4547ccb656f894fdb0d7874529466f1fcfc720600b268f7c6a741a14c1cce6a2297f7c7daa1c83b58bf1e2b16025855e8e157df4948b2e0b9c49b57cab47da647b28f6c9c056fa421f1e9f7393f38256a14aec6d59c3c9d13649232c41;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h132aa73270b7a98372b24b77861ce6f2af0e1059449aee2fa6afb08d7a9e358b97df325ad9a3d381eea26ddcd39a661a02135e38936445ef236d6e9f5443dd4b9d03ac809b574a0e334ad6b50348154efdd830475164ca790cfac9f4d824cb7ddecff7a7ec0f31f5939;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1dfa2c091ec5766381200d4c1b54af7e2ed6f0de983bad0ad66fe6b6350dd6f9371fe7d0684eb8e4df56f3d590052746c28a5b36c7c79dd19a59efe80eb303f17d2b90c6a7a0f80b0ecf8e23a894258335d1ff94b1011519ed7c8339458a022b78f0d036020dc04496b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb69117f1bce789efa9a0e362a2aa1be054313336b35a304e1696bd21ef27c294ff6309bf4329af49fdbb159ea69b6f97226cfb689e6f02e0ec2ad1509c39516b1f4b5d22a5029a583e56126b4fa571241235c57898063966a7afd536ed12183f186f7d7e720129cdb8;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10c11339cfdda8bbe65a961ca20bbe281130f5cb859a815be30adf7dc380871232e6ce5f085cbef85cab06fcf4a2390867db02930cfb07dc42b3e9616d869d987e81bc8ef31838fadf309d586e62ba8f6ee1794e19bd354881d8651b13103f27dc394401ba27ae9bf3;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h163f76409733e7742c401c9e51fc77f7d84718594dffdf91dda5b1d651704dc674b724343b8ca2ec69c1ca3fd67f7c28c30c9b81c1d776ecbde6e812368449720ba7270f40527eeb10dbc95bc60d3eccef70e91f060aef6c31d8b6825da7f7042712afc573136ff9d8b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h14fad6e90d64925f06f3ca58f826b18f3938bb4f369764fcaf9986a3b36d332ab1cde070df103ba82186f9b9999e31025e2765d3be6fe78c18ac819db0aa2ff1f13a71eb860bc0cb21a9ede44bef95f21a5cd1659714e38ba0f6840fefc0a6896dd8b57d3cdf869b1a1;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1afc61d62c4fd4a850de637429171ae06616d82fe7d1fb3ce62424f3421c9e7bd244b8929fca278ba11f9324e8ad2c46047122f79b902956b928934da3884d64a821a8749dfa0c188907dfd368879e6f42f9aa4353ae5ea7e0e4a98427c77a1efb107682c2773542c18;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h141bd5ce9c5b56c8b0c510d3f9d5e42c88daebde864461eb694c20045045d5367246eb9d7caff43e9b5e10e413627f1256edf7597e8da9e90f0530a9c6d243ea3c7470c6135f73d787fbf955a4d9a7b10b1e7fc372ad458cfc768573f3c09d717e9f45422e67c70eda7;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h83880e93c5af705d33b58f7e0b28688230721c329390441f9389e237d81fc78212556b19adb928e8f6e35a678f11ec1da1b229b9a98c0b3e1fb1a991c46c3dfeca0800409fe724914e81d3aa0ae0648161199dca2dd16839ddbeb6b9f72a06e665e018db54a8b84bc7;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e25f878525f4096cdc2500da0aae618f3de8b26cb87281e5e95774d94cbb14bf783792e1c5cf8dc4ce2c4845e3f0ad375c7627e17c3383e7cb2dbb104bedc1bdc10b9b89663ba55457bd766e95e9116aafd0c719e5e9e1e17f6fc25217376e7ab79841bb5f5205854c;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1630733c4f839078f48d9a993707cbf8be9add08dc9697fb7f5dd441bc1e9affb585b54e33d10ca827be9dfc648a3d8140f3de6c71a1d289fe2d345a429b7056b8bf27b8beaf275544f4ac8168592b3539cf67462928be5c91e66b88d5a28129f6fb5d5f4b9d14b87e2;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1bdf5348bec42d977c9fb033a8df75756b06edd5b5d34aa4f0669ed5ca704a2ed3feed3b7541bea013097a7826e4288f8ae9347e2fc37b5c6a9f8f33f3bbd78b36bd1cb8b0635ee364ff6c1b2a465695299f4a4fa8fe63284e56713d89dd66f6a6b07c77d10cd95260b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h194ad11f1b906d7972b1a6499705683a06808c3943d97fd7a60ca2958686d80cdb1b577cf877bc8485cdbcfcac428bcbb354a4d25b61c08517b658c7be14308ee3cd16cb7fb3b191b810c26335a06dcc419d5562f50437b26f4ea132c54e57e2c8359d95e3cbddc5f55;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf11efed628a2a5d5a7f5f4719a6da355c484ba5492bc738a37e2ee4a866b38d163eb1cead4ff8a3f977cf54af823e428fb882bbd2e141c9ba19ef833779330c514864601e6b182fd17b9d011b4999b1b169f0c36cf1226f981feee6bd0d3a52c9b6d57048d992bf5dd;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h15775f5b8f7b8c5d1d5916ce436651a95173a3e3d07aaa4a0843bb38370d339dabdd50ca278ec74f759c27cf7ddf526b482c0e853ec6adfc3d12bd96da071706807fa235caed0dea9dd3f68120b189698702868030433a9be14146fa6b7d12ff2b887bfa0cc674b5695;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h19064a660a60ae634768444abe30ecc074dfdb686054163a810ac036a3629b1938d4073fc04bb02a69f6b4183821e106b5e85de54642217b2195d9a66573d8fe5fa2623b58a7f722e1cfffdb206c44abebc48b3e51bcd04f756f376ec25ecd1f3f0191c33fa353d1fbe;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1bc53d432bc218337c1ae8a7c662ad4f56410a5fee167396c874944ea97a1ef3bbcc5be0910580d37c8e201fb55680f1e35113d762dfb14518d9c856b72de50e1f9d38be2e8f44972cb4e2d4d46549132a0ce09bcea582d5cee32aa2daef4cb564b0b5e924b9b532a89;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h54f6b4a96cc0c70ac4f4947e4f504d7de587fc2f716e16c22df457faee4c314d45bb501286b709af7eef6fbeb54064eee6f1706f9aea31645a9bf61ab74cc49e0b66b2e6cd534ebad2451e98377df3bf7f9ec339c7fe9222a5b67f8a321b1b005a0f8842481c089963;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h187d11ca733aa7e5b9b6632ccb9fa20a09c975964256dd34f1aec92e45359069675f2250df81a84659c2173e6b11ea7bdb787196401958a71591bed8421be2bab636e532fdd6f3ad65795fff136e00d032a7305baaf5b212c9dafcadd738bba4fb97c750baddc54aef7;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a5ceebab6a96cf6fce413fd66c903a305220171351bb04826b15228070e713c3d14be120f85f23a9f0b190fb332b01cc8613bbe331fe9cc81ec1422c8b4940bda5df9b93252845c09149069a9ff97fe77aa21793e80a3771759a157873af6ceb2bae90d6cf6b29949b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1df11c6c353df06e00c668f162e82063c50d7cc6958a5df828cfeab48ff98cf71125354316857c6344a01a086a85c8493f3eeb6eac3e2a12aaa69fb6407562c0148cb91aa087b68ba09878f11026b522718c735ab239f1f2b6ddabfd4e0cdb4f3c20efc9432b6f62da9;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd1a41326a4d3a8d5c0bfa21c719a7a38ff25abb4edb46e86230775eb03e6045065ea2234f567ee3207866ca232db508b98d0ba082f46b11ad92538ee1ea51adcd78dfe94d9666f303497b247c57861cbc506b3d226e8d26157076f31962402a73778f006944cf78845;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h9b3a9fa30da157123f0652bfe9a364400c5a5d1f8f948f6e42e74d31a77f7ac9407b9a235d093fb82cc11ef8c0c6550521088babfd99be702091f2944ef69a7b99c1de17c04c71797e491087c8b2dbc02220e1b22b2f59bee9f0cc8dde687c8583a8d8388133b5aef3;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha92503745a3846a33505b56c6bf9b46ed491ad446cbcabbb41279b1fb56dd693683994d17033c5a0ed6bedbb23c21342ea76ebcb59aa2cda6f616de08266fa8a88d4f630fd6c39e1ee4f6edaad61867f5909f31a56cad509451f01e0e2838e4748181de15de4d87b60;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h195bd7dfc94961febb2fd232fbbdd8e7c3031f3b090cb2b240b5c9e827c399b209bf1285f6ecbef28dbe02f027057f0e27d4ee9397b122e1f64648946fcde304bda9012462787aba60d8009946e6b36559ced6174fb94f54fde2f5b6e3fbbc9fcd075bc0d814aa99f63;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc267d01c01b7b8fd4b4b927118141825b506418639b6dd1e0fe11282fdf83b6bba029dfe6c4fc333d8b04e47629c42b88015b13c5f279a696ec5332d32788a49fa6c59d81f213f24cd7e5707cf16f98486036ca7e3d7d9e0e98b781f0c66c949a1684bf083f8e94d7f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1525bcff2c9eb817489d989919a335187d2ca5464cab704519e1202df3ba9bb3f65c8b001993b751c3b38cb113ad8fbb3406b2c879e81043604ab370926cacffe3b655484df1bfaab59c6f47f3f30182161f56ad927c69465e7221b02cb7e3e4b847158d17449a18435;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf072be84abc198a646bc58a8a467e165ee944e8e37569373ea26f691d3de66d3fa7e1d6b3a698fa29d0272ebea385847b504aa1f27811616b715d9aca06d53ad42f0e3a924abc930c6df894769110a88a14294f95ea19a837573dea1b7a5b6d5b1e6ce57c3b54cb4ea;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d01736f4b23b2ab1b622303e5b2fcbe11c710b8239a59894951c3a9894988f41f54ce01d6087ef163103aeec40a583c3c9b053730c55381c8f17bd9cc62625c250a36800e1efc46a4ad8290681741faf9fc1a9b2037cfca3821d1d14416edb2a0ceea1006a2197608d;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h11444f3ab7b3b0564552832ac852d573947ebfefa524eeeffba2e63e990d622fd62d530775eacc2dc21f8ec7f2d255b8131da2b5f13307e546d72302afa68f421e223ccc657051f3f8f785dd0e712c19915df0810621a5ece6e701ee7536ba911cbf959bf554cdee3f6;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1fb67d84e1b698c18758e431ca5ae986eb30769df29487ac28e3b6392ce4d24d45cf232ffddcd41daeb6b61bdb9838df93afb9c9f01b7c53ae7ad10177dd4dc8d2b8e08c0ef96f2564e537bb97a999dc21a90fb56b598131ae36bf465c763200335ee660bc6f44d0766;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h16888dc20377aec099e7127bd9a1087fbb672afde4530fd0f56ad5c5b00ceb5b8b0e2dddaa6fa157f961f2e9766d58543bd2f8740c9f63a884f826379345dd1e5c0a622f35e94fc3d69a3fb9eff1998ffbe4325c109dfce658bb3b9b25903227c6df306ab2fdfb9a16e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h184c945eaef42b499501f3262883ac6f2f94cc3bbb6bd9b47c79b203764b03420ecff5dca8cd175e926320c4dc06cf2a7efc4a7d4e9b9ccfdabf732701506aeb2a3383c8225b31c811755c48c074446e6d0ede9a21d9fcd73216c13c66e29aaf051eee52707b0818b05;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b1472ec420b21ba72661ff0a47d3a11b02c6961fdc36e58eef3c990b90128277e70f6842a2448339267f91e95d3a590d388d010fc981489fd9a5f8ebec11c6787eccc09abf97bd27814cf8d6260b78a261214686115bdbc1cc1874843a0e7cf159aa86094bf8f68417;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h199c2379c0fbafaef41f96d9acd1e0c625ca62180138e55ca3f9301651c1608e5d750b962058f9d0758d95101b4789e640e41264f7f5019cb2a16d9c244c69eac5e4bd352c9943349b6a276aae27581353abd3e289cb4991320e794b6878936d6fdcc8fadaa69dc4d99;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a0f3c18985f6fb0a9118d647b04f0a497bfbecabbbec6fc83d6ac8572883253facf4ebe545366c895aa0c66db91025b12b48dbb827511dd546bd7b841764425073347ad70b1db226b77870c02925cc83f33f0c3e024457a4736626814288efebc1e1c137775bf0b3ed;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ae8c870b4b52a6a000df31d62b4a07c478bc82770c08c1d16d7399c9a422b914c8b18f7a5f029e77093f9bde146470450875813d34ea3dd8d3dcdf5c8a613b06588ff1e2caf1f978b3f4ed73f90c8751076a25e79a15fe32ceb36cb8326b7cd22fea43374890878ea3;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f40b301b2072788db9bc57aa51ada7e808842c36c8d96e6ca0ec1ee8941661f3eb0a41874a2b2174856ebc630329d860304cc615ce3e7c29f0eb1b18492f655c0ceba07afb4473c134de3f981ef24f4f94d09e23810cbbe7467293fc006c49df11891a7d7d0d04b256;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h162edbbd84c4575ef08d081dce674a46455b5f53f24f82da366009d6adaa9e87d85e71349f1789bf8f517e025e9f6ab975a41b55fac319a5855e391d99cd90404c8e3a9b1702dfe5e0ec3564ed5216002e1d3d6b5228b5b34443e1b3c27ddfb09c448b3ce3f660a9d6f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h511f167edea1c280fa6c27ba6d2b3dc3b2c086b87a0352965709c05484583b63e5639777de0c49c724c47addcea97847522d0f30b0e2f4085ad79974c0c148ee895c58c1027371f50643d2ce83b4797bbcaf6705614838e6d0a7acef148d274c39b573de444eacea78;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hcff7bf9c956372c542f84348a5fd1d568c8a348511e367cb45fae8ecd0c3cae1d0fbfb9c4a82136193d34839bec955c425be46e6db2a0df2bfad12e21817067bd609af2f72d4ef1dd63c8a7ca973fc907a953e06f9760415b02537ad61e3c58c11c93bf18e052b1711;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha6d00457cd4d1ed172619ab15385985810d96194903528a064041a3e1b5ccd5352630a4ff27483a0a6351fbdcb3d29d120278e27b6d8e381b4188d63f58695b7e007987a8452d2b6138240d04110d917bc2d5ffaa33460435065787bdff134384dcd0e0af24577b6c5;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h101fb3ac73a70451b102a6be2f6f0db5e477d1209808272f5f3553265b4f9935fac42d4aa4e2617a0e870672f4eaefa28a662ae20aa99aeb257197019aa2e3d5b86178f123eda132031117c2f82ff1e849a300be62249a8a541e2c24b621f014cda4464804f6951e719;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc72b59404930d9a546fc16fc5b65281424c9162715f7783849ce5b1aed592c7021b7f1d0aefb207d95fe38376ab794f05815b15840403aba18c21614e96136e9ad570a9c7be101dc22ff93bbee53d13f72eb595b92490d0ad9a37b6fccb9460c9d64450747f78ee29a;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h74060273d9a04d8e1b210cfdc18d7413f586ed524709ca8fa528a5f78c485b709daaeae729054e79c2e8c20adcaea28524e8c09e4f39de19ed9ffd694f46ceff555be45e31dead41a60cafef693fe0151bbd16b022f617cbaec40a74f5128be492104e4fd20f971d28;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h16562568b261abce57f256ca412ef8a371f572e99d1818f697227894668b9d4e601c50cc333d49d65998d4cc786dc75b46542298fa1be0483da58fb70fc1a5853e5633aa88f8c5e00608b5b3459ad97dc477a50da742b5ca896f07298e00f2cbd726bc6865e6bea8fa4;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h73b4167e48790cc9377f7ba09e83f87e6adc9b1dbd12908e53cc248c49c4615a0fcfca7fb3085600622995fe030a2c6e5c5db919bd3dd354aca372c0966a0d9bd5a9dbba7ffd7075bf6d93e571b31627e7422ada916757fc189936a56cbd5c3ea3a9316d989ad13c7c;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h5ca5f79c5d036a9621d3f7e0a44b0b3319e00ece2a58bc688ff7fa0287c350662499d04c6e1776b3dd124d181ed48c914ff46a14efa4e75d9f9a67c80e73066e47a6971fc5b6c0d124db6da2ac8cb065886a29c5a206f0873a030133f613a330f568531665ae05662b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ff6937e5fea92b3c97f53552176e9bbdff737957e30289e2217e65554962476718ddf6dec8e34f4c06b2528af2b53c4aefa9fec0f9467b82500239ddd9468123e7758d1b031e6b2c8c41cf3290d622af44892fe184f89a8e7013b4582b10027e0c5346870a66bfa349;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf2d1bc1e24e9be52780a415e94b1b6d6415be4f9ab43b2e257040484681a6a970b6009ae10097fedb5d799128dd15974841efc41986203dbedf6f0d0b0c47538cc1c8937d3b7d72b6e2c7064d750b8a6572bc4fe701ce507df0dadd96bdccaa078707b49f08e9bfccd;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf37095d3b95a6c8a64dee3f597385c03843099f8b14b89c7fcc2c6b966353418d0a870e64242b86a1931ac674e500e552f3fa3eac3f2b383ddbb563091405d03720f58d6a4ce5a080544450b42f867d8d01e79879f71c397a017c20927e8bc1a5915e4d6c5ab8323a2;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h152c70b247317e0df1bfd4265f076b3c4a53163a103e2c4f521af2f89a679d22d9f8a1a59313d5bc61f4ade2989a02d6197fbdc4b78d6ccbee294df22a8c26fddfae263562637118ef7af2f4584fa4a9f6e0b390ca9325b18203fce08bf54ca2133a55201b3c895ee7d;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h3c1b96e38033089befd26e1fae9e8c512174c08a1ce23e4ab331759de3d355f0123a3a928d7885a3bc7ba9ef5753b24337a6c9d15517cb398b485fb39cb1e982c6c36141c45abaf8a296c9d18ddab588f42a7f7adb6b61c8a0f6af1a93a5ed59650e49ab7540be20db;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he33d11a31de92b4b74ae72c369b0bed48094f243d717cea586e2b4b644333072d1a1e9978c6356d8f3f257593e537b0b3b93b4feb1841cf9238d1b0208c86a09c3396f42cbd4143c6be243f37ab0fe22f85bb4584846315233b92dd4375e4fba351f209c8f99e8f19b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h36e9373ebe4a9dc94d03e370b1cb0773584e1a853d8807d139ed0bec0e089c30c6478dd499942ed4b5ce4bb7e1a51a51d7c2abae41040288100ffe4bd578c4a701124ac8b7fc9feede1c0a7a49f41f3484783433326c4687c1c3784b0e308e3077b006ccfd3fa1d565;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1fb2336b2591d8014c9b7997aaee614e06d9ce9c6e4f6dd690809c8a7a7856d729d87c433e5fe5e4ef700e841e1a294544ceb757becaf70e001c12b111664b707f7fd498208dd421b68637f5f4eb5be8f887ea5bede863e6eeb6dca0bc43b279f0601f9438ffa74c675;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h43574c7627028172395ac474606d11288d1a8595293fa7554024344d286ecb6e2abc92ac0f28358c9eab3dca6861caba8886675ab165cd642de722d4e9b6440d043922d97ca9e4d19054607b53454b60967e9d80bcbedec241c1420896bbbb0ef9fc48a848a549e1e1;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h48f987b1253c808066fb9662fc7562fccc5511ccdb2d94cf05aaf863be33c31bf71c9217a0d624dc0b8550c96531b67e3641ba024020911dac35c648b03c491b0917e45ec425a6619220cb220b0999229ff7b6c42828007f6d9d2bb791b81bd681a0f9371b3c3c2694;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he9b9e95dfe85cf49d1139ce3cd28e5450749920688adc9a3671916a4a26f3e8aca6abd09ad668b6e10ef392c3607fed6e81beedf50b76b8dd5ce1da3482dd824d79587df82ac9a581863ec5cea98987e0b986bc53409d8fc840415fb895018b2ca05bf69c41b39a8d9;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h283da3c09aa5de6547d4ef0415136f8bdf7deb4efeeae4b08994ac5213b83df88208dc0a0b4aea5da605eda6c1bbd663e58c63088fe5e3e1f4b1592b0adbd3f973e4129bb8b371e5ddaee834628a938051b97bbb6c5fa52d11cb616d70bc12e2396cacc821d2b1c486;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc1835d1542eaa5fb3b5e9f172003f6603cf21a3b4b027a69d650421b5ec4fa10f20b4a293977785e1e6243ec202bf4db649e8b9132b2865b5a51c8abd0f5ec299be3a8f6624fef37dcc064b4be284a5ffdc86cae126895e7c2f1c53bc6f611e791f8933d300942115d;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e6526a1394161d50e863b3cfc737e64ab744690384f6195319bef7f9d129740fe14038183c295a28b676d04d082dda155b0405b48b7eb52cbfc870d39de9fa44046b75b4fbd7db965a3a0617392403ff90a0050dc2de99426f4b8fe46894e731190ffdb301d18b6fc1;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h107d2e9d43974daf82914350a5e58d3257621346295ae76afcb2b96ad25513a45519a5a31fd7956f44a5b9ac9adee85133cc86aba6bc0d8cc2b2083d0cdb32645923fe0aba3a9aba9a479ad852a28fe65749c49ec628bf5c22e5b79798aa44b48242843a049b1aa9d40;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h40d3de7dc105a13498010a20da95f0b532a8ceced95d48e2650cbca1e12e3ccbe68b4cac0a3d4a5a7a7786a33a8546cbf02b2bdc8579de0a12e1f7c9453417add6325c1d370920afd81405b5a5c0df385e873a36b6c86770726b4f60d82b79a887dabf39afce1fa220;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he786f632ca531363f273d4a62437c7fea9f8dc434c221086c5335bd666efb89738977c5b89375e9cf66f0686089dbebc207fe76513d7af2c80d29525064ba37e11322971233c31d83d4be1e924059b8db8852413f3ff113c9634a13e05c889f51744b97267d2a39545;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h7cf2ae02c70a04fef4259a1cfae0bb1880f9a46c2037ea50961e3d79636c29dc133997d92612e8a87a4e24c4b0c5c64696d3e3c8219fba6845696c77b9695a9367b74730a77d1fa4b698e9fd11f1857ce25acf8cff194062102bcadd5923421049f5f301005b5b0fb9;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h12120fc75eebac0ea18ecd45fb348f55acd24a44625db59fd003bad6f00781b9b642617377cf35fad76c4039a2cc474b9301cdff4b659b18cb2afc99afcf574a86198c7a8bdc10282e8c5848dd42f88a6fb254510edbd2036ffb1dd59423cc13d38cb1b6d455d69fbed;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb770f88293d91837e90fc2890d13800b9fdfc9c8b276c851d5c0e16505c23c778caa0be527eb29a2aa01b321a465cbb5a90130d93acea548df1712d39a7bcb3add52b30208609db89c06b34b10dddb4a32656374e93ceb738da260d7a29d7061b94644f2e78e5ed7b2;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h3af0a459f0be2dfd3c245cb12ff4f805f6fbbe551b64221ab2f2ed295549e8395ab13bf325028b11c8e63bbc571602317ea1e180a38dfb7a3fc7f8b40d8ba1e54eda0d8d1c6cc70047f48e028f721abab40fea25b696de2a89234cab425c053c1d6426ac01b0f391eb;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h3101f3f949fbd8fef16ef6b869e81d75fa6cd14b0f5b03c5b67802e8819f7147680d417d8cf03545434bc642d03f0a8bf4abcd9d1adb8c75cf0dac30a1f0e8221e65f43eb8fd93a7c0f0de93773f01f176428dbe7d0ddced50afddd46d195f1d4147370e2d61d5be90;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1262839886f5ce3f1732df9ede66633d2b2031af17af7ff59306765577a42d4b8419a9106ac57cdd4ebde342eada83a60b6a50dbca2466be0d48b035be032986390c6ca63cb59e466300645ece63b2db8da2cf585d99cab528c87c56c86b5ce6f2e4f8c5d7634d6eb30;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he34fd31c4a9419241537edfbd2901695dfb993bbd7592a6c0c9a15ed1130e4863a1d0fee26e7f3103dcfa0e5e38de22da717c40b783747de9956cea6e6bc40869ce3a971fed3938eac70a5e41629992c2bcee5d3965ba96c4a0987aaa33ea09652c76d9b1fd9a8e420;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d8c490e88c87f2ec7a91c5142525f30c225604a8c733c812800611baa66c6d89fa07dd65b9fed753aa54b2b203e2a0d359cca66f65f8e524514b48e4c0d862147bf451385e9e378e24c78e076519c9c0ef67d584bffcbe41ea5dad10b90f5804a8b4bce24218496862;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h873fa19a9e7e53ef361955503ff8e20c5a031ef56ef07192ed8c5ba81eac7c1ed28caedc1c4f4ff12301181948cb6142836f9fe674786f396f1013debc919f7874bdc6c77c4e8c0f7bed56e09e9c35895765f63bae1381d2d8a053372c676beedd02e0f584752d46bf;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h381c398622cd1665735aaaca769cd89761eb2d72d5748dea189a9aff8f4484dff210f898af2821da11f587a9256745f839a468791b652c6ee61ad5112fba9464122566663b340b0610d68701a9de626ce610846a17b84e030c99b608064144aa0ae401751224efc068;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha259ed5e8ce30d0c506fa0098f97b1b3ceddb4519df625bccd59a5c9e461c19a0074f0532d58e1d31d1306020b986db998b3fa0c73c6dcacb82574d747160becc51311612d0de4a871492aef24973a6d5f901c63cdc9b67fdbc8308f94b6ac3d0b2e6239c1f3efa74d;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h15cd37e7ac3f446907e6d9c11564dce2391c836f85a363fc47875263e722d0aae76eb3b9c046d5571ce7cad8a1ebf18f50b420399f949b19bee394e3c26b3e4f1354c788a0ec466b920871f71b2eff20a8ec497cedabd9ab08d26523cffe838fd7810c8e5cbe49f3aad;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h96036e73539cb222bb562526c27de369db76e508e3027ffc28ce9b3c83ac56b8cd072c91292df54869ea9869c34bab11af8e962e9b71444b4486799a549e0f434c816671e32d8974c49be61b34167fb608f91bd8f22b511d1922fab1d4d183783cab621ea984a00b21;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b4a3e1c90c5b64962cbe8ddd001ce7e7b8bfda5c1b2dd675dd99b6a563649e44ed840c1bd8c6f067b107c9eeeea30be505f3fa2bc1a92eeb20a9482f957df2781330a51f2ec4193d831f667ce1de70ec6fe3bde20cfd8744280919d52800fa547f59bd38619bec5cc1;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a8f849d15172f8c669c48923fe8e80cb39783ca2f304b9849fcab9e8e2fcc3f81e2ae5701ec1a8bd4d4603e742122129088f06a7472f9c1c5484a21dcae88049b33109d4f85f5f32b31bc4ad8b9cb38dfb3a1327550fcb96f5db3e5a923de1dd1b28d6e4a377b647f4;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h9aadb364fb0319a716504e93645d6b738e5d6e81502e6f32211e646cd735991a56c0634824b50f1b98c091d9457e3e688a5c682badf5c4d7adea38e04ca0b0eeedab7da935efef03141897890bcea918871c183a50bb19952ad264bc74e5d504f3d5669548598751aa;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h6a65c0c9b8140303147e5416cb4e504393109c01d032bb8b1d194d5304abd33ddaa219ff56af1d001dfb4a6fa0f0517a0e0ef82cecf8e0cd3305638c0dc8e8e5ee42d97804b4b1fa4ec024d2c9880ef27ea43dfb0e800290812e4658524180ce16c5a198b10c3611a6;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h154a98c67e28dcfcd8a244a35c08b54a33f6d3685004d0507162753f854015167d82cdad2d0b3dd1463670a2e34093843022f8756574ef9e93223cadae04dbde9afd105032da79fb91fa46b2734a16baca24b05b1c1f7eae5d352745f38c6e98a32275bec217558ee7f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h80dd669c62a1dcebb04231e3735076dae2897dc0b4f825b3e17ea101766f4dad93c42072b5474147deda09228b783cd292ca7da78203b4a42a7233e6b99f098ad5d94f7a057b0b3083b3e0f158ee95fc99a65ed287aa2327c4ef7f8475ed95929d918c74ab8ff5fdbd;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h13f161d7b4a861c2fb8cf9de9e93900e626c52c90d29f5d89e9b9c10a25c62e180caf89e1cc67baf297895f13b1358a038ee711e5b2abc96560dc1e38c72855b5e246226a78da82c66a100f197243805667b4db712ee29dfaab8677d553249011cea015f0e7334dcde5;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b3d33ffcf584b6663a3afdc33dd29999e61dde0f2be35ae81d1cbef44a159d25cfb35760aed26f924b6308498ab7b4bbbeea258367d4305ef91906b6ecefa4289aa1b41bf4142d3d8c22425319b7841682568d977763763164c0e54cc9eca5498a3a4166d1b6d9e50c;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e6f6fa9359d234ca361817b3f6f8ea961ddd570ce96e44c4326f0effa057eca4a73d716c938a9b12bb087fbdda4013069adefd8930b128b2b00ec75d95f8aec0908ab6fbf23caeefce33e897120d72a6fb284740b85c1c18c3db4c56b3ab060b03e082aae883c17728;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h857d2e21aabed6911e6deb5e6823eac3c9fa52b1ede037c95ef534182d546b6d07bd47eb329539e25767d17c3c49cf9a4286a4ee5446d564115bc60ac88801f6bab69de77672a2d9c560d787e706c74a9c7316a66723d90567660baa8ed9d664790b83ff1936f07b79;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h18a4fe1e34912ebf77ffe1590266fd3125a9dd764b027f078461d528cadfc90d3475b4f5454d78deb5836389e94b6d8dcd6f46ceccf987ad5713daa95772ca51d4a87d423d293aa835128dd3df6cf42bdd50aa198d001c47241a076ffe54f13410c41c7328b3f6cea21;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a426eb5d7e422851c1db68c5b8f180ffe6a726936c4f323505683dc7f1df111d1611aba40620d729ab006074f988bd6ec1760675bc637243660c5d128f7c44012f7c95cda6a7759fe714e03716602c1c591058c27a46950c6de1930e2a2c1721d15289266a94816ba3;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h941714058e977cd6f6d49dd79c12eab247294cd797f365d62d66de82013e437e412f96800b94a7dd57b415aaeb9459ad9abcbe2e7d6123918fa3fe4e086a23c4ae8b7ce7e847ddb43cac8f4fdbc7679cb719872743507e6a9192ac197e0afd1357e4898e0d6a1e1edf;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e948bf2d0cb5e11639750055535553a2c9101c6cc712c8e891f048a6aa41191dff7598fd70886e805bc1d1f36b4dfa90499d3132956cebd1d8c62239cbc54ed5616263f296802988d52f2426128b0c6968e3bbe45bbf7bab8493d5048c7893fa56390dc52a8dac0df6;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hbc5081979b12a8e1626906e46b75e741343ca4548470f55182619879337ead94b5112cafbec139a56e9770464f7296f970f33c72f72f1b8adaece73a65488bcd2a800f736adeb195c835de38e31b3bede7c70dc94e1377d59a9f3a1ec76f731ab0881fab36f0c476d2;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h134822c54a021b2cd3a9f742dbb964fe648625e16a46ec42c0d3788533ec63db76c1770781c8b65b419e8b5df7978f0144ac5b6fcee0164cc81eed4476816ebab5d21c71519dc81dbaa9f14094710dc9b0eeb5a20204840094439fac02d390b90b68a7ef64af6dd50e6;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ec0783b71706ae87935b6cf4d927a04a0b0042ba1171bc1ec06d7b0f8be0ecd36ed40d149da18686c8772d70dec5d69987b6a361a17cc1db3fd7f888d39d12c53c33d4036f4d6faec648bc7f2f9e1f40f78117c7d6ad3c278cdd3a9ef89b22ff3f1487d26cce50f3c2;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hed948ffc1ea0d11014a2076aab9ae177746dcaefae0cb6a0c552623f92fb8633d933083f2a16fffa4bdc872a428d6f6a713c914a19d45d38d4a78bde34dd0e41c56ed020e43145aba29e2036226ed2de3b4b41bee2f1c73c7ec9d88b1acf25cdf74383526eeee1694c;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1fb76aec7a4ac6885c378ca9540f46cc8208a0e36a3b924ec2b6e33a83e5efe2505d6e97b628edb7d0a5a48aad0ef9caea07ad0809c902fecca4718cbdc8473bbe09adaca0c3296997a489963bd925e91e576ee17675514519a0e39541b0cd1f1adc9a9be6484053088;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h14cfeb4e3b68650d756718989f2382ed5c8427e68fda764fafa2391935e70ad20437c651543417bd6a5011ff7f241273f403bce787ffe723496f47b36052de77b6ebd40a4080a61caaf0ce5696e8d6f1d79b5c93228a7028981c115fd3d40eafdfc75b87f22da0d025f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a19fc8985b872542309ae7c6f0f4765fe60565991b1b0492509f188e55c2866d8bd053ee5d49f6f876352908761cd1b6bcc6c78588809e0962ba1bc1cb03dd4c44371ae3f9ed30bbf5e1cae77b69f21ead706710854bdfeed9472d21b74d1085ce219244a5b59bc329;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h191c61c1401840703b5f75eaa8a055b489c80e2e79d316cc0df226d1372406adfd663ae4f68ffa655049438c1475b32e1ede2746d08c2a4808d4d3ab2a0c560a20ebf014177a8cb575e16560028400f10607e4b600e5d61c9698542a9ff2ed28f987b4534319f30c7d6;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h4e650187ac47ae868ec726206c98e7ac19ec64cf8a974878b50c8b0a2338bfb6cc6eb06be4286e87612665e3d3c8a64b022ed50fe6e286ea30de736a54e23ad9f937848a58aad18a6235918f0591fa4179970e8831ee5f882e2491ef123b4d0d5e61a9691f02724ade;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h163ba8334965d9197c620d1e088fe478a9ab24d063d8696fc7207b1712da372803fa634e9714632f927085c2e9145adb35a15b685af391fdac80c5209f7873bb6e736adbab6feae1e14835e172cea2ba9cef36e50819c5b79b14ba24e17c858c045cd43dffab7a3145e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h645443ca0f555db3615deafa50ab8ca4a4665c9ad773f8beb5365fed829c96606a6a26a2f63125f36cd4276c3c25ed5e9910b39efbec3cd1b990be1d7566b12e92e9675827fa46a036a02a98fba203aa3082d04bba895c56b2f707f8d9eb9875434c1e1cadca9c4dcd;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h576d825e90e4d95805b111845a0822ee615a84c96dcbec7d2de444709e9f540d934765e2713d529c3fa95bcf26fee59bd12d02710608f74c63c88135eee0687382971a3c033f02efabce0b096d645e3c30b17ede9ae3d04bbd6172ffcb41005ee06038c288671ef65b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1717d86e9907d806c616de1dcd4739243ecc0365be5b6584059c11b9c8c4749c1ceea176d385e32dcd89b39215d206ff47bc420bee5a1ee0241721713e79375686b71b4f8f1937dc81139ec3623bf3d86ba04830781f442597578bad0a37b0555c70021b866062a70e3;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1fe54578d9c74a1e30e0f639f729f86924967f277c2f6f98bddb90a198ba85f2c2dcc7ecdcfafe2ffc1176ebb8ef3671760e6b9f1a7484a047d2bb278fb0436b78a60503ff3ec16388695d4b8778be00b5bc519d933d4cb359ee9236e614c7d808fe20ce4cb5437f74a;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h113f60bc8bc1f54d72da9ca711bddb3e5295cefb0a609c13548fa487dc626963bc4e95818a6dc0e7ba75d4b9de2012f40dd1df1483ee2764dfaca8c4974758fc5c50fd9660a2ca6165fb4dbedc558153a6d9142723af431ec24e100e059c16aa50826967344cd6bda68;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h12300c82175404b4bd1de8cedd162ce1309a019782b72ab25ccfeea637efacc2be80e5e0d69d448b3b7645d544dd927db3fd195a6b8e048303e51862303892bb9305facd01ce1208301016290aea44cc7b11625e97d90ff1d238fa77a06ea7b61b84bb6c1a76c216930;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1def1c831ca066323b5199a4a815d67465318b5d94a944e825fd0f4481c4a1f0a727318b415449ff6c5f4e97d2005960a4e7555c5b6a8e0e960e773ab55a9dae8f3664386816f6f35580eb31648687d32384f521b6aa7d09c89c1e1111a182366a681f45f98662b6d8;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h7b783646a57980e8bc80eaa209daa0315dd5f233a95f7a26e1bb99e22e8c3a910b3ca475961c21bc193b99ecc743b31da6145dac8e9b14f397c221f7e5d8da2da80d51e56d5842989bde4e28847a4931134bc6f466973d8e6bea313cac4c9e99839b43e3c69c9b73d1;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h20fbc0a99b8dff8ee2d9819d4d914f48077b628d78282f039cb5f22f2dab6c33301da043a3be2cfb9a43ff37fa10b5d02a5f1666d3a7b536a073f73ce33cc4eebb14a828bf8c8e2b4b33a54adab7b43982b53546c5b083bd95a3b54aaac10aa2020654f729b4081f1f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h17f603a32c65ec38799b184d13551b59aaf9f7e2e70e74e3c1154605cbb3d8fa16cc1bd1c2802dd1d35bce70ef36e0abbe6d95c4ae8f01fc7ff0bd7f74a9096e9e9ea58bf79113298a8a0fd1be9401df1f8c1be8b87be5a9fbfd448f28128b3d4a03371d14564397665;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1303568364d13aba3c0859370b23c5e7591d2114d7f0a1a340749d29eaf712df64cb10fb6b1d84b97bcb577e633eaf3a7a0f5169c133da0e842ede5c3e760eca53c337f7ae81167a0512e35e3311fe20a21af901fbc76d58201d12cd48a7c0c5bf251cbad032c319889;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10e399a17e004ad3de534dc43cc6bdf1e2d171713abc7f5348704d90fd4b5d08c6027f8de5d91cb4a496ae3d7ae08c9f89e2e5d54a6205483a45a64ada56dd60da8ca91d00f5aeb3a4437c9c1504548d141afebca7d68ecc041cbd5e1109da0e5ecfb1a542884a1c4a7;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1832b14011cf330fc3bfd81da5b6a3db872eb3c9333a77f4f583d09fd7ca32892868d400c76d5314bd44e85ed8f8f3762850839d1fb7aaa5e5b27566be8ec349434a92fe8346ac081d47fff924bc9a9238ed1907f26e52d962bba9e9a5618dec0bf55c15a6f89d8cb8b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hdc69cd333d5ba27af30e9b40610f1dc5c336ec76a54513575d532de4a7731697f47d3be92c1d301db2dbf55541440eb3f437d8170a71e1d9f87290f8968dab7adee41c3c18104b312d21e881fa0891c8e3aadb5fe00e6f47e57706140c4b4afa62a4526da6d0bf1648;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hde6c05857002e10ae4828e1fb2e55bad0c461c0901a2452a50a3ded5ecc44494155881360528206291555ba89d6811854c39bd4d87eb6c315deac02c2da94a2b4b335c5d230912f140671ce0d5a764984a119bade9088a5ff7ac7e26ae95e50442f4f099988ecf01ca;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c4850b19899766b66d9a6f41ae0a45ad54e4299e8943323bdc042c83460f801ffb7f2941e9a8b117f2b9435e0ed2082610091ed1effacda829ba83a022fedd635a3e19656fd855ea6c3222e035aab619cfa6e2b301adb812bff88dfe3b2f25f300b264cd14a98d86d5;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hba2d46859b6dc167236770f82bc3d2364d1d8c273bfb3f6d3a82760141361a3b7a141c59a0eb38071f68aba23535a0bcc1a9ec19048cd3df7c3dee1c4da7919bacdf0c12fdb864edcae8716581b5a05f70852fcc3e86ec645ac7d0926edce6b2feff1f8fbad7a7ea68;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf4edaf431c4c50209850acc89420ae35d5b3d28044c8bea4bedc27eb6465d18a6a05307730fa0e3ed21e1b37eb631b8e60d65cb2ca743a90d95f3d391e1e76c5817c3885d0e43a80270ea65277b9c830d11be94948780ca9489d82f5d14fec0dddd84ad5a7c9499f07;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1037ee560c61477aad0eb94ceba109a7612f711488aefbb141a1130e8c6e64bda7a12649dd44f2fa325200a924683af52cde58d56aaa1a8c08e48808d88c9a714942654a48c89db16831f362294f9a3cfea29b5fba86c4d2ecaf895b587dd502bc6572c95b0b3e9821f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f6d1021a7c54fe6f56707a8ab6998b019360b089a0f910f5aadec42bceda71329ed2a96788fcaa394a667bf30836c83fb9119c283aaa9fca776b042586519af44bb2d52ff05a6b3319c7e968c93e989285548c45d5fab35e421afd75a60fb8258d55ebe0ac06fe05cb;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f7c075fadba4e39caed9b1b2b1d332c79bf60c7e3594460ec78d5a0da975de558f66dd15e6f4196838287b3f3c00f85cd01bde3e7e8b52444ff58e199f82050730873cb26f0a8d5cb128ca6ed819a4db3efaf7366e9ac0c7ef09e2e6f98c1a40ff9f0aaba1ad9237e0;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h15044bb2442c942eef9be36c51b9f2aaed5398991457b7abc63917aa0005faae0688ad8002e88f85e2906de9d1a4327b65d1eb7c171f7bdfa459858735e3cda287a24a2ab474b93a9099dca613f859446691b310e5afa73f743d687e0446b5aa20d012b8aef39f2d4b4;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h7b15c589b4110d9c6b4ffcb60cd4dfd8fe90ed6ed7f7606606af56b8c3c0bd2e7e0320112fde118f73599410232514031b1cf979faf2ecab26911b44ddac30eca11eac93b78a03bc33c7e9c8b1203b45a4d7356b3d1e645f4eb5895b83e78f6588d41ad5764fd5e842;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h3c2c374ded941870d5fd1d6b44e7a3cf6f1b164f66b516f9388a64e406b481314c357dd7f8179cbd3bbcbba77c1be33df8ef7f0471fdbe368d7c1a92e0ea5c03ea24f0af1db120d129b958d42537780879dc9f22491a81176c72fc858442527bfeb61d8fd6ed88aee8;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h135866cea1c06cb4f9707393b2c20a17c9e0c27d3411ebc56b2959e1e5a0a0c1743f0c9e583c056e7ed6c6f68730d7453ccea081ce7ab00e4413b0cd3eeca22e8826c22aa908ea2c598a9809b1047ad5dfcd79e4b3261e19b4cb4d9a3207e023d04af1e0d5f4fc2eecb;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10b8ac55327cf2f46eb81919a3af78e1911ecae3382fb306c1b96cdd71b635804d86e54d81ab38038fd9405716b18d3c1dfed5dbc7b752399f46b5eb49a2e0803a737d4d5d98d2b36a332a7a671ce4f146f4d18c6f909dc5c97a51bd64a4a5948680171e4334b5dabe7;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h195f40695e2f4dac106a1c2e2ddaf2e025c29a4b58ddc0575ae78400afa15ad2bfa7907ab99f44e53528542c61bf4025d32aba7993f3bf6e141ca0190a45e9bdeb5de79a046417dc2eeeb0d520363f3f92f141e370436ede1af3bcbb6d6de64ca6a209d1f9f28ee0120;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hde1d465fa57e8871d0f578ce35ac6e70102033e3d3599b5de57bd30edb3933a8912bd2bd0ec64f2c8fe20855adf200eb0c322f55aaafcb6c01f3bd0dcd095a6271d688f359ee4369c5a0a97f3c131683381d56e875045d1eb33f86b362e3b2ce509ff584ce01f65020;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h117f91adad6a8f3743ae5f54369fc1f27014ae357d8ff12fba5060519933c13f08c05915489523113bd075ad3e89bd3fff2b37a4e11dc95438d81acaf0a21168877340a67bd7eb42e38b5ffbbdd1354bca276773a69c0fcec504919f0597d37ef1596a8a46b25a53eb0;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h141cc5d609c330011c89605cdc0d1d7999eb7e182aac13483418a8ec44256a877fdccc07cb6fb3cfc919bdc57322428bb7da11690f10539fc6fc351243b339640b66e51f37edfa9513564e63efc448d79db8acd4183242e86611af3825d7799dec36921b2824c59400d;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he263635b657f12e01306c0bb7d9e92b458c5ac04693162bbf05790dd9abd57291f2b4f008dbeaa73049dfe6430f3ae458eae2286041fce79e655c41ef25be024bb037b66f48dd985bc98723c3e118032324c3a2171640b9290fb4f5a227fecd8fff0754689cedff510;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h92d35423b2f67f507431d38d975f215cb66ae5e1e8b87f7fad51098cfa4cfaa8b23f30fde963d0fda704fb9416f498ff7f8fdc4b2a9bc1be068f4fee2544cc62c1661c14f1959e522524fa0b9d30632a2e8938fa9d56dad2691bd8cca3606bfe3842a83ef965e22642;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h167f1d032961c87f105bcb72813457ca9fec14df76135e6c7506b98140f53e42edb2881d724f6e4b1ad33e6c93d20bbb7e57b48ecf5ea208656666f5c8febd23c5a64b0a79d166766ae8424a7333917ccf357323acb94be4c081984b3529951000e0b6cbfd66077512d;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h62c1d530d715cc85704937ccac61fe9c7f8d1049dcc95e39993bac3b9febf88af7c37cb07af9d613eb001803a65f444996f55731dea3db545d4fe7b73d3801d445cc8d041fae1fb6f4f35ae363826948ec5eeda26dc81712e22bb8b9273c0d3f2711cca302b67ee2fd;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hcd0e078a4c1c184486a722fb33cd0b35740ad100604988b6d5f2e43860445b493653b0eb8df6e6394e7bb5c1a5ac189705669c461285db37588e9aa9c1587d27069c2a6d9800531ce0af9f79476b80f0c466e141d52af0099290522d6001df2e87f34c2804c0a12c9e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ee3179e1a1d81e7430d0d7704cfde0a9a01a66f90cc28d9a361344869d383f40a469a97772fcb6819dc6f59dc99cd6dfa5f447c147d38f289ec411194f513db8f1e61a60b55bf47aff6e0e68ec1dbaa9f53e6cb44f0c5adc987b54522762446d9cc18999a01654a17d;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hba6f628d58cd63f81ef425367966977104d7dfeb3f55ba8f6893dc7134e71a285dab63cfa586d8b57519fcf518103a84436534f9d044d6efc7205dcfcda75bc94115874264cc834f3cd52f70e5a4d0e31bcaafc5226c4549b2263423f68ec7e2efa1b39f02f34a0b57;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hacdb034a11658774afd9a646adcc2bb5541e4a9e65df361c37d246785e57cb17b06fb28b4a16f688c860bf0f7d0184ed23452d9e21a31796765405fd3026a696b4c1ea6cc5ad2d6c4f4c3dd1ed9d54599c0212444d86b95850900b11dcbfd68f909c97cc9b69e16360;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc5cd4e4c8b30e0216b7682217a5a01c1b5a01520328f4b2bd0513374989d63feaeb3a968ba0c5b99a91caca2ed35a2092a4ca7383e564bac070578718ff125ec5aaccaac46e36d3c488f55bd9175dd0e9d2716facef16a28fce4e157efe68b9cb835d970c305f598ba;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h11ba2cf2609e796ceacf037e9d7e4aad11365c112b96be619568db0b40d1da32062cfa817bdb2b5c108338dbb24bcfa334b27587a35c40960c055bf61ff5dfd194d35861465a2d4403ab23a2a420581b680aa94b1632ac061f1b3d7920453fa2c5e2e1007350f3d45ed;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1718a596fa79da8b24ebecfbb3982283742912e8561edade4974b8d5f51f0efdd73d886f4c456704921a7e139547d56bae6d277d7b49a0f52962bc32a45a9864235f6ddbf07e4ae172f00265b6771c5ed689a19097277d0897adb2baeaa5801bc809e24cbbe75c0be5f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a81240e8cb70d378eb6017c005c82e5d465203c6e279e81f3e3e0b083b171d92408799e8ac6c72d00c76dc3636f8d7dbd9e5ee2037bb1019e3f762b5b105131d8d93ec64e34e4c35a3a312e87ed726c5ff08f850ef4b2e59c5db449850eab6a030cbf8f708d7a15c7a;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h11b5c57515a4c1223f28d678358445ddd0190b24fc9b45385a8c451171569f884a397158cc7cef9e32de5e89b6f7e1aff1a152bac51cec97391d1132b9d79ac4942911b060895d83b456128859720f9e19f6d10c8267353e947818070c7db4fc766e50fe9d486381a;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h11da5c6691f6bb3a8a89707de7df9ec9b378fa759536b40adadcc2a0f7c39f48c156b79cba1c929a2eb63ce75d7d07c4bf4c8243082d3d721a9ac171609fd568f3891e0132744a51c59e3e566ba00daee7ba33b9e188404fda43ec6fdd57d16dccd2386ed749c60296c;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a8700f965ef2044e088d61c95d0787b8f68a8b2f0c854c9850b4161371c518b00d6f1863223286d4088040b04b4c8b4adc8f85ada7177f3767fea384789ff2acbde003d0331588a04d66670d929b633b919d7b20103e315a1535f9894f9c0333bb5292411a7a222236;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h73f9b43c93cd52e93fef613f7cc14b67d1319dc20a9a190ae11750a5a21f71db4e94daae909e54b8d016b4f5809ed1937e9ac2a8ead01fdff205ac715341ed4e2e0bdb63f635bb72e7602aced8b01ed710955bb69da7dd7c747eb4a65378484ebedca3c8318c2ef779;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h83d4b33252b3723dd206a512e4bd0de41620404939999763ffd8f135fd5284414811a2ac1818f20b3333ac3618e60433e9a61d546e2be1208d0f3eebcdc342245ab3c9059a8c3900da726f3ac3d4414dce9992f29634721d0533f236c0a71bd47a88548abf84cad57c;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h46864dd9b7861ef3226db01843d75b1ce30e602174371823363dd9a1d06a266fb683ecc7cf509b70d80e59e0b55a12227ba599ec8215ba63738e172df22e7f6d29a9ff3f7873f154f10b10233f195422710fcb135b06bc0a19bbcbef870cef42f9a421ddd3cad98d1;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b6facf55d8975741a3292f3c3a47b2b500f80729bba910d072e5eb24ab259afe01cf8083a4575d710054fe3fe749ac47bc2a7c788d0299d9af2f0cee4475a747a2e026fa82dab315a8a9b2ffcc434d2134d6cb7ae0177d76f0fec40bde8463dfa0adf92d6c586d658d;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h77325ab4ad5dacf068d8edd7e3d005ddf3cbecc3c64bb23fe105a7f11ed5916c5e1f81fc8468602dfc1f5a275bb486026fd42af2cba944f58a8df3e085970d0321cd707d1107870a2bc65081d3bd531cc842919b9dde7b08109f8c5df4001f8ed79b1ef30c00437551;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h8fdd59965e53525e8b39b7e9adef06ff466ee35b51a801a2ff51494dc647a2b9270b5bb77cda040b0c36b15052abff33fa26527f511b5c0b9a7ab07ea90f6447e6a2a572270739f57e7440a38a2cf18668ad60c95def337bd3d78a0f8e85c0c8dfd720d8d52f7dffda;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h880dbb23ebc3af1e91fbb4bd435b597a5513e940537c287250c9f1a780748dfbe413d18a008b83e4b33cf6ef6fb3588f60090c069e1b3db7e596951a1849265e56e67f83cbd494ada9f38b42d85fb55d799999713f16502c201791849bf350b685e5b79f03749744ab;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h105c24f0e50888e773edc173a732a7cc2e875095afdbd38f38cfa496861ddf65940c153f83a5a636c8e6e4abdf7d38a9730e600e3b1849fff2b33c099c55064d2f6744f999fa2b37a653948981b530fcf56b73217bbbf6b775524582ebfae19e31013639696f36caf71;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf092139b96a8c7f68ee6e6f8a570d56b4c720f8c11c076877bbd69746c10b5f293158c95d23b3b8acc50eefec056d96bdaa3b89e05113af63fa01fb6c903568a57af3b4d3228af67cddce8d5f285ccf427ac462446366b6a35b4a8f41bc33b6fca30646492dd0fc398;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h39a8a83c2d07be80c8d8bd1845b1996b747ba4f79773b7d8a304a66b8f17d7943a281f6c1b887322d3d50f576b94c2f83d9b8b010f39aa90cc333e88cbeb0706f6141df7f867310821cdf8ed6e6b690f78d9a776d3b7534aa53e520d3ee12c1f65a653569c8fe858bc;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1629e340e514dc4e41be87b93cfc2ddcd0ff75d0dfb20c10c98b7603f9c1711db564943167515c07aac892b9c819bd73219bc7528ddd274ac82bd4f36077654645df4cd4ca6421eb1d0ac073590f22c904aa2a7a0155f4e7ccf91469e479e0c14e43cf89c6cd9b1962c;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hbaa0f7f3719a6c51a0ef8220182d7ad8aafb8dc0e07c72b3cf3e453489bfd0bf3cfce47028e85b1af2c7e5016fdf3acccc563a748a904f0004f8653b28f683755fae525a6f5bec9f59faab8bc1e6ef7a10dfb6c32a59abd0b4a42b4bb49a1e5e1286fbe2dfe6cb4d7c;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1fb0c071c634ec5fa827e6217f96b19868cb5aaa8c12914893b491fc615d47ca40e79bb325b02738738b9f686ffae7c2946b7da0103d91ce280ca6afa4d2bc3768f4843a392aa69dffe90bb79ea3570ac69b14351246e5963cf87551e455b67a30af5facc18dcd57bbd;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10e350edea09728aff10df28306c402a2de2042af10f527aa8bd8ebb9fd7663cba68204b43a47eccade1ec0c7944afb5e9d9f95d66e00a1faa48e5c32b37e947a83ba7f8223442fd59226b3f33cd65eda83a953708168302a3c8de6fd942840adc2087d15291923efd;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb1eb32a9889b0773694824f223c38d8a6e067e68349833aa7b856db729116104ffec04bb13c8bc2f252ac8ae1e975b0043a24986c0598f62a33ce05a52155b18db176b2175932eb963bfe845a981eb73f1c644b6bdca24ac88e9abcb6528e53f87cc810fafc7cb153e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h110a78227b291598378f454feb7993c69f31e1b2ca36bc600a00ecc83b28f122e81aab082bb905bfb7d6f20ee9ac1e8380636faee60294a7e9d32b5ff11fbcb82929429cc905e96c1538b7e17d3be32659b3b4ab55b2ad4379efaaf9e58cac01e7369f5be44c1e769e2;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h8663f802927622a77f140f7973cced7db602819a98a35230b4597f913804a0710ffb696f4c683f8fd0951bd667824a1d411e687531ff21aa3cdfdda3f2af366cb4a2ce685dad43838a1989e9d952e3f7661bc2f5d66fe25cdf8d609704dd8aeb7ced84c41d1ffa8bfb;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h5f48b1d2e1b8cde16e3ad70e5c5f0e258eebae08900606bf01e7ef518f02797909c537f190abf101089120002f34a7d212540fc2c642cf786e3732ecbff13d5519abb15156642d0202ca4e4ed6368b6c19f1ddff78f3e978916c319c3e49f1c05d5a99b1235b3256ea;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h17c25c12159be331f4c805a7748f22b22ca4b340dab3fb3de3807a8b81b84e39053dfa2f47a50a7ecfee83f0a336d9e23227d082b212eba0d3377eb396f69989730862f51ef76ca0f48eb7266a1bc6135ddd877bf44bb53bc733a7bc1b2899fe143755dae114be3ab1f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h16828e26402cb06f0e08614623f02187fb922b7ca8c14be217f2a34c16d9d43e10f6fb7838c10837065e76be5051faf79416f98f2308d302990389002b767f288f7182989ec8927dd28a002e0c3cbc7e424ee5139e59aaeff020aad121614c1f90c138bf22a164a9f4;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h8db9bb2860d73c5aa374bb87fee1639505240cd79389ca04ff34c426702b98876199a6060cdcc47c98cafa4ecdd3ccaf4f6515125ce50932853d59b58bf3f8b116b8347a1f20f4c9e1327ab076919c52339497d36e5b7a1423b54648aa0d60cdc7d58807c7eba81ee1;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h17464261d31d25dafe91b17abd8f4184a20f25e907f804532d42dfd349ca2d6d79b10920e121c9c535e2b55ac755a88cf94adba49e17ca8f12f5bba699ce42e736f88be0f46c9a6a7aabeb890634e7630b04d57e077eeb5486f4d07242ff73ccc515aac700b359e5dad;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb10446b0120a040f3ac1ea16f2f45d0190a74b862a90c052e6eeae08b3ecef3bc869dddfa0343b995367983de6889db76dc18135d8229a3ebb924d97edd536c4071a8c5daba56e794f466ccac910be65fc29fb909e0dcb20d95837a5ef68fb84b4eb90defdad12ed27;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h13a36a13197abeebf7a76d44608649c3336e18d553c801990dc997abd21bfbc926b13bc1b79a8bf92411c9b9a12125836d374960b2a8020d2397e4b026d839056019f9d4b78da98d65825115c348e60ffa700614c0d44b7f55f7daaed6de905cab6ef179d4ae7ac5eb0;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'haf8bc62822d188b51367c61349fb66222f4904d9f86c80b3163bd0fa58a9a08c365202c4652f68cb9801e0f2d84575b3f5d9a640016c81c2fa2b95330956a3d867c43fc6c45cbe1a353f64bb3dfd967c009a3f1768095388e0e53b74c5c134d22b5e9772e42f674fa8;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h5d90816701ef83392452cb568fa118bb5891ed24a394a9079f755829d7569e55c35be2bbf4559315cc0b24b7c5bd5139af532526ced79071296dd300e3b0bac243168ced3ce47c90d21948823007b444bc562e34dabe1e68025bc6c7409fe0391a0447299dec2899ee;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a20bc9e846793bf1a42621e9fa35fc29a0c92439559b81aeb6e659073896ed994013485bf34c9919b4c48585abdd8d8e45357124a143f43a426570147edbafbbd7c39f955666aa7efce2ef49fc4cd59694b4d5ca3c19fcf46f1411429519a2856f3fa3333d6bb77236;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1247415d564a9156504ea64fa88f978aba9e56465dc0cb6f383f4b70edc3cb6810d40d7cacbc7d1a9820bdef3c777ab20399e0808fa06159206daa70b4563a7fa4f3fd8cf224546775d6357c68e6b20d77ba663c0496a7d8c0c5c1994624f608e5c0aefce8deaa34798;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'haa71ade2466bd8cd01181870bbcb3fc51830d38ff0eef53c4274362133ebac776e5b8caa9768bb66952a75d55190b8021995d78c39cd065be5d7a08484b10993c571aac34b1e0bd1704271d76012cf4d6dfcd4fef4e1e067c6fbc6369bec5bf61e1c7543aeb8d7cd3b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h225cf920c5c4b84ca3e7ac628c0d74d61d978ce8498bf96f742f36afd8e86a19ff866da19c69e0f404128736bfad46309fc34623f2458f2677343ccf629ef1ddd141ba7409bd4bb92922e8e354630b9391355201c9f1f898a3c378cfa01ab29a17e5c2d1afa3f64148;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc2a0a58ae74eca8a6bf38ecf09a3c9b6f75bcd41e7c17aaa5283bdf2eba2f8873a5848d4a6bf2236ce7d0b296f9753f4843cf5c20cd15736846f7a38ffcd6d9fccb89c6176920b074f1210f2ac90e15c9c1a2e0ab5f34b75fae0a026d2842e4cf2f90ac45d436242e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1883c248db60b4299d39e72f8dd4688420da00694f081d1d1a78d7cb2061243f6c790e522401dd6fe82a72cdfae04f28cdbb617ec2f0b4a8911c17c827732cfba296a0026d0478c3aa74066692cbe8ec1312fc83806aeff9403b95386e13e6abd1dc9ab5c805227aa21;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1231f913cbca93848f1165220de25478e87836c77b1a68e52edc6ed0d7ba59c300aaf58ac0a4ccc98325f4b6a3984b532f19a00d59656b34541ede10688b037f5f743a1997dd4a1eb58413389bd7040e654d8590e3b589416b985325ee26849819280598360d0fc7d10;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h47acbdcfd0815b3ed5b27274bfa9eb63244e0b435cb578d0151f6bb555c968292ac6c9e3036b4a2308192e968c5b7ea60a6a58651b288a26a27ca16b78bc2432090dd61252f3cc6ef00fbbae5a0d148e57a7fcf6cee39e8a39001f4b04ead78387b9199c2666e5e66c;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h6908160f925b2a0f5ca118d04247169079df120e9136adf1a5f42a3e561af8ef9f719c9d62fcbd3f334b5572872a78b5f51da1ebd8e947e3fab8b0576a43ffd525adb3a4c7bcbf2fcf8c98705f28c88e359cb6b0101dee56c0789cbf9a7cce16561d9026bf4ff33030;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e6624556676ab65fb39f6e9fb3f086c7b3285aaaf96f92c7f80f3825cab7784d15f7794103cf5fcc98cb49827c57808a6203a24e93a4ad96b267aca662f2effdb4e0f40d621ddda4867ef5cabe3c4500ab9383a8822d7ce00a9304006d8b262221baf7fd6413bb7d15;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10c47d1ee917e043e712fb1cec655d12c66b3f796990d99484e04904dcd360935ba76cdc87ba26b50ede603f0a2e9a75d58adb3fefd30b6f18c4ab7c51a6588c23ba89261f874bfd9f56838568bbfddd419483a497753661000799dd15d9ef9a00df83838b59909c32c;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h942b682981942d9e347856bba6513c524184ebbbe3d0f3708a63c3e89366a7ce96097d8da924ab1e9a85739ff0c7e0d69d4984d36fb809382723d1b9311c4c446d5d4322ac07699c3572f5995fe9a2a77e4549de8a98b2a7e9c56de60095cc1bcfdd7c751ae8b0bc3e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha7b837de6748278e65ab444659b44a1ca216e6e650d5bcdfa04c396a02e1291fc0de238866235c699c7f7cc352332968824fa53bde1a6c07e6aecf729409be7d4036ef4d726b48e0068c31271329dc5da2b2d9a88f41b8c275c1797a9029b2d38f683d5793dd826cf;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d204ca3699640e802c2d2b7d2b1181444a5703aa815df3de5d546bff5a4616dac52a21f0e3517d9fbf1233a4a838e66fcd92ff0cea98e45c0ee5c4ec3367037c81942bb663153d18ff5cfd0ad2fb1e286dbd330aac2232520691f35cf094f5a952e48bd3dbaab85fee;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h2e8f204d6231ece9333ad0c2f25c301afa0a707113b7bb6a8458eca660a4d65e8392b8eef8d34c1a86f9e98833995b453e56a730d5c2866c9d2b8194d1caf48dd823a8cf2d7141055d028d9ab038d3b416805d1eec82e0fba1a8fc58900d96f6e5fc9df47c39ec837b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h15f028360618f793dc8ca063f9a9545a3cad09eb811cfde8c6e47ce0d842fd5da2660200e3837efd644a9d1a9c6da1291f69c1d8c0999d669de859a39e9c31d2c88cc5360cd1d7841969e1200e06bdeea824cd6a9e2454be2d7996c4318c7fa751a3015aa316f469b28;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h4ba03a1b4cfaa604d15a3ae57a83bee454833159960291d68364f83c275cff31843a5b69f78ff5d1aa031d654fb4df3c87e651331809f415f9938a1f36f19258d731bad4e95d8d6baf978e1942926398cdbb1f752bf9d6acc332e851d7aecc56015a9baee03194b3a2;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1beab01e1ba3280eb5eb8f920e39ed5f1e97ee1fe56685f15de65442b22d42d1d686120986fceee19a965ab2a068f79a89a57cc2b9f0910f66c4d61727001347f841b093896dae4b145c5b08ce75f808f72ae8e09b98f6f0a5c2d505c2d47559cf5b3fd1afa97ec4ff8;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h4ab732bcaffd4a68426e6de0d1c37df8910305df0259fa7e5b0723e3aab4541b9f3c145fd88fff1dc9c11a8a35c7840b135336508ee8da4dd7dbf13b11501c8d2b5d1354f4e09714f5eb425a8b2b701b0f6de5107c1b81181172d3422b777cf0e8d1496c3615ab7eef;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h14807b09a19d3f557e2236d23296517932ff69b73e6f75a8c92aa5bef49f5b0a13adb086ff43b49768dc08d6c5f3d1f6400b9160a42b02061ec1a90a725ba9701ea67989ad101782a896a662067e5937c645b7773c5ebc50b4f430485bb2ac70e8fd799543e43667aca;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f7f43e549d6fed3b88a87b9395bcb46cfe06cc898647673375f1b8e54273b60d054cf516920144d2d4918f7a130513852991f1cf5062376be45ca3b6f5f818081a73f4c3c06e9e02f6075c61110dad236367a3ddb5892a99b22b176b21f3c6e94c2059237853d7696c;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c4c75f9816529251cf7e94d4e8a1aacf3bf67ebe16ae6c20b7e5279f383eb1b48442fb3da769ef3bb341bc966ac69b56288d9752b82b2e3e5db77d7fbe32d4dfc48e7ab20b1a191ad91d893dc6d20cb79035f3fac88d6f4ddbdaf22bee42b34980272b39d46dc402dc;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d8de640787256b143f4caffafcd99197851ace61d575863b4ee7c949d434d1dad9b6893be20c2690793036c3833f84db94a8a3597d87c817bb8306f4fb4074437faaa001f3ceffbad57670b1c55cd8eac7a00a0dda1c1a38e5503afd27d77cda77784503371d13658e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a59910d71d217ffd05ee8a147b56a65a50fe53d8c3382fa546bb0d4a87b6fdeef3ed361cacf86432bcb8eba423de09a3f702c36d03841fceb11f169bfc2a0f52a827399e0459e296bdddbf8a1ca8a688de20477f5c255899b352789dbf7090b660d86cde7322b6cff7;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h83291d509b6beed5b81f6fbb554d28a94e79df6c7042bb7f42d70b826f68741ab20ad6c384fa2384f14670469d62af7992e919194eb17a8192e4d63265ae5d41bb9c70af84e0ddd50fd37511b89e3b5a9331fcb0644d1c55797a54fabcdf92bbf51f7444ab5b67c3a3;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h129045cf68b053fa0daaa2b6a14047c3f8f09004e92459699b92b871e5c1fcf08f65549c3ec6368ec47a0546b2dddce2e4ab289e4678b7ca47a38b363d656e70ceb2ad6417a309d881aee80c6ea9e49409af8aac25ad034937f18e07066526ddc1e5c255d7bdeedf216;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb2570a738a8650b283afdbfaa302d6bdf2636cf7d0020631b8f2893203ceba833147b4fd548f83bdfdaafb233b7096a202ab7146acdb55f7bf597b30fcb8ae84b926f8220f50c9c8a22937e35c7fc6b2f4e8806d2c52034a0272ef0c46da474c68fa7bf42d2c933cc9;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1125f2c69abfb05959d0e90f1df0b47ee367691a5bbc33d5ec1899131ea1815feeea6bcad0613ca2bbb2e5f9afc9e642d6995f26ccf70a718e323fd3adbb92963af4ee74833c0a8247fe60fa332b8220a3c8351dd093dcb5e0e4e5fba7b034410ce5ae076cf2d4a6606;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h6e7179437b3c0440354cec25a1a7823a025b0e8e199c18e3da8994cd9241c19f929813a7eca59e54d8b1eb9d98b2f2d286f9eec8d4868860bcafa20b4cdbcf1ee98c46a97e0ac2c197289aa554e9418a13d21ccc8c8cc8e20a427670d9c6e5a1dd65d186b23472cdd7;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1997b42b3c4d2c730f4958f6379886f3254c8a0f7cc7b48123f7a4c469dc8c72817b0dd0a87d5510224ce93581b5268a9786835511ce562281ea8f65108cc18e2908a74b2ed47167d6188f3204d3c842541385ed55f019d58657c454e30c63faa5fd4b44fc15c8c7eeb;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h957e4d3dbdd8b1a4f22ddbfa7b82d2d157dee5a36398119dd3080d4fb08ee01c86782471012c4abad22f9b4818e10d2ce86cabe81641283dd6c9fd3d07352b86f336dbf8854fafe680df9d4d74a17d8d8a5609faae23a79821af932a9219af64f5719bad603b3344b6;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h16308ff3c5174687d5fce29bd051c49e07b61e86fce94365d40eae8a8b151f8b20a886c8f38c23663d6e995b66639e25c5dacf6fd56dac381f85732c374b4f0bcb94501316a50d7433c3c9d7000538f27b6e5c53dacea0098e265c331b87a8b7b078d8767ea9928c99a;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hcdabb4cbfdcf382e7fab81a1e125332d150549800bec04be56aee47edb91b24cf60fa9d461a1f9bb5ac77c23a14f38de943a286ba0e76190ee17d4c650a8d93d10b7e2def5638d6386616846ad6314d987dd986a698140e2a1593b6d8b895269ed2317342f24309c86;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h13292b8eeffd3463ec72ffbb1fabc8a424b18fb4a18a8118d173e1f80dbf189b326ab36f1bb72d8a195019bbadbdbb726bfc0b9a200e902cfa1fa4ab1c8b93f39513a82225a7612cbe9c97faba1a275f811cc929e4e7952341fa3a6f8520b0a3b2881a5c7d0c679b056;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb5ddef3c472bd59edc89e024aaa8a835b33d128d520afb978621d22dd87c1bbe948fc1d452db9797867f8ffea976c35062f8066f372d64b5c2fcae87016d9309f000c53ad15bf95fe5039cbd6d037ad2c54065ca1cc3eb45b18e0f7410b3b08414818ff637b2ff3d74;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h18fb7c77cae4b0e02c04ca7060cbade5544dca9d0d34c1e45b7990943794c4cf0afcdda9445aa3f59bf27837787a23f47f7948eeb34541637e1047a4303411cdcc21838398338b6fe6c58ca9a9aac42ed856d5d705821df82ed4e8f4d9fc1ad6c934638bc65407e86b7;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc7fcc5cd7d52575f957285f164b52364103e973668efdfbd90cf6cfc814c5ca15405c8753ab5a1f2f5a0617ce41b26fcdfe8dfcc17219079cf4b309e1cf426eeee7a4b4bd0fdd5d2c40ff51e2683b146bcd5feee0fc351855c76bcd54202732d906de25baf3308cfaf;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h15823a86cdada792c003b234453b0c74cf57e1d6c43e36c73de215e451a24c085761fa5d122f6ea12e3a3191b2ef15ac789dc7d686876505e55357fedfaf0375e50731c626627643c6a80a5ffa8380641ee5213ce2f235dbfa0f21c82e61be74c67309edd26ba0fc1d2;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he254e040f3c544e7517719c543f57f4c2776a6987a038d428536ea47242a0f8dd8332b810d179c8db2c7b2d764d54f1437fb7345ce938526d844ddf4cf92798df1d8995e0ed2d8721bdd5147b6deb0debe7a62ab27abed1c83131be7ae5a26aee03e11e224bb305b29;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h56233d301160f22cce49c8af9a0590503ad1f4ee2a71ed75892154c7186ebc1d25e7234bec7e71f9ea8d39125409cf5910efd3523ffcde3a7715aed6067545e2d377c02d416363e43802e1969238980507014b612f7c9c6c31e5754f8a9d48127cbe08a1bbffb9ff4e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1218ac1b7fce918c93e28294d2c1faf93a6afd8f35872e28a0241886c257a202258ddb49b8658376f06b234fe8f027f4c1cb07504496322bf11a6f6377179555265d0480395e85eca45dc568697951e66d0d8bf567992fe5d7ce6720d432d3cc90ef680c197522e98f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1324a8fb1d04ae0278d53e6cf14535844c416e90d90803391a30fb20958920efa3027e6dbda46dc2a7e666b5e44e7b868ec36e2dd2dc9a89cbf8d447d04c9c9ef58d495c83f4133923dbf3e2e0de66f5212c168611ece438fa02def33ae2eb5073489e09934e3b48740;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1535b7fe44d5989225ff455ddfd9572c6d493edb227e4a85b28eced642f1fbc61091e9404b299ed3ba731792cfc77ca2eb2e5e0de5182b1fc8ebc2ce03bafd76cb89a80d87d16c739ad83da9f518842a7826ddaa8e2b2b423599c782ddc7a09ffb5b412995f9ede8c70;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha0b25b20566f42b27564df68b0b57079457070cb51b341c4c997b84ed29f6607b11b5d27c906e70bc709380f2fca27dd8f122c5efc37c0e8249076bc89b6e7935598499420a399ff7bbb51e67c42b4ca67183daf95153c4e8fdf3df67732362467d2470d1f5222449c;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10c9be14d938f059305416faa55712d9f20b919711584db6e6b603a67a9c1455d7d51d9ebec6b882c78985af9786c28c2c7ab872524fba6c5131401f25de51dcd6421dbee6bc6c365aa833266a77ccc769c06bc40ddba208520a651eb35bb66ff3020656d5ab969e2e6;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h15c7d4d01fa2ad5d59fa5d453a1bd43488f08735401a9bc287fdbde1de79cf6f18964955046ade5ed5bf35cad71210a8e252dd95f044a386fa3187fda44f1aaac3faa9490e5fca1cd57cb47248f6b0883d364209ea767a05696c27a16f95db63ec71fb092b175f9c05e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1828f6372d6002197f5f114ccd55db72fe34b727d4fa43bec69651a408eab787d263feefef4ef654f49d2c743b3d6cc5530e92b21d2fdec546dc6ab53343e0f5d99381a5a18abde4ce62060de2ff04440626af81dd2cf481ba671704a12d1645e27f6e8c7cb7c77eae1;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h42c25a3ccfb6aeafc7f23057506a113c063040729c6252650e2bfc70d710932eac0368d58aa8dd6bd8d840fe8c54bb62ceae5eff5945319b792f1679624f71201c274c981b821a25920d6997f0f17bc43da15019957424c53acfcb9fb3cdd112cb5db9263bd1608926;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hfd991eeb1301ce2e0b9cb2359c91763659aaeb1529f043b5a35c3b8a2632289493564bbd07539456c611d29ae1026f15fe2c414973dd511a7a0c7be8e9201d445805d9219a688c88c4bd5a4c897d7eb2e5ec808234247a637244a4c41353fecf27b0953065bd318f2d;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h11a29ee4b00c7cf840488710795b6228d3e4626295dbf67a2cf9a0b1ccf21e2694ab379524eb9462165aa8cb05b4cee4241ca61176981b3a3725fc82143eb3ae15b3e10f655e3c5d0d3a603d081bf72486be18afbdabd2bdb5fae29999f7ad1f40607ca64d5d94df50f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h5302f57159cd7c51a3fdd4ba76fc8ef483af50f2991898c12a2a5f6fddd2d13bb945efb7435d530760a500fbc1b39eb0a7bfd290f1ac075b220e393a96d67e5727acc6fd45e56a1c1e3071567860a1846eb89af8d55be0bce4b96fb491cea9d49d7e4494425ff38b7c;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h9f2ed49c79be3f952accadd90132b7e7cfc95a65eae783f8e71b3800103f1d82f6dbbd11768e98f9c82f310a8979a45a086e21e1d1b3e1ccb5a4835367757400a3a7d40a2783e747a534556a5d3031f67b2d8bcb6632d6f13e0aa92d06eec3bb0ee1716219e4973942;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h9e16c7bce5ef7e548c2ecaf7e0f1634e9acd3a05e5768a07228d75b1ba1d4b9e4570959170a0f553d4674255e7e744508e39d0900aecd2e0df185c345cf096ce903ab9bd5b1252f55752059c902bf0a21d42ed40041d9092c9c2689ca5ba71669ef6047ad677e216d3;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1059cb888a11d1da15f3c7823c192477717e4613832708fdaf6e0b7dd09fde6c4fdc7716e3c7214b341f689b22b1fd47690eabb390988f970a32117b7a6ec5cf81e8e304c837b01838aa5233fd15a3995be9c4fdb0961b5478350d8f6ecd9ab00dabebd22b28b90e4ed;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h808230a6d828b3282705d8e3ba4e292a94475c942712c9644d67f0ae9eef09f2e8ec235d834ef212260e254f5e7c81ef74c6c153425803bc6c856114c769e062c347ee79870d4bd8aeaa8094fb6df1db60babb98174ea0cd5eeae0ab3604665adf2bbafd528f5aef16;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h106da4b55a08a5832c136861fed3cb438ba0d0e5f7d12d5dee9cca421c9ee2d6b9d82e6f34fcf59b20ba7502141f3bf9ac35be94867fafd1a5cece331846816be157aefbee24f3e30f5075edd091ea2e6c9b3884027c66b3503bf5e95a790800d4dafd44666eeee0ba9;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc720cc913d3d583b6346586ce677c41ac1fb530fcb4e3835e5314d55733f55d873afbef48954704a4d24fbe6ff049480e82c661f7a3ca8b8ebea85469aec70f015cded14c9c0cc391f83e5da8599179ce3439d1f6f3d18889a0bd5089db268de3ae000f90b6ecd92b6;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f40297b0af246eb852fb165400272835d75922d9270b6a09d36a163f87aacde868892fc0fd1fedb2424eb1a94b548a8802789245109e3b9f62b12cb01bf451a68e5cd34f522dd7e367f939ab8ad296c1f3312b6d0bb58e8c80a6443bd2dc6e7b23651892898b3df032;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h5d9b1692b92a1ba79e6d664efc098e3520e5f79a40e74fcc7c5a523b263918b88f310785f3200ef7067db7e9305d77ecb4033f47693af3e1c81e1594c7307feb78e92de6612c85994c8df4c34047af55fffcbe426076a2a0fa4342fca9a6db0217597a76499bb5e4bf;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1434ac5ea6bafe30c53b63f911da88094cb1481e4269b91a6a2b98e633b545dc6473482eb9e457318f9e52009f8e296db28a7cff8e0562afcb4206d409825da43f20b0e0f55e6cf1348513668b5e0581fe1fb89a2bf143f895e0ab3899e3552e8adc140e0b943ee41c5;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d2ec80dde2c80e0a164269ff769fbba256b6fabcbaea1c2f9ada29fe5115def5d71a1a73e041ea6a06cd8d6c1d58f144164efa0a402a548ee615580da005b90fde43d47474297339efc9cf4d56625d61504d94a5bc63d3705d15a68aa8f5def76293a14c3de7e72805;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf76010896bfa2b0bb2ae19a87c4b452ed0ae50b8a691004c53ec34cf833cebb315e40331fb7ff77d27619e7a1d659ae790ca00e63ac0e6dd49ea47222f85585844ed916acc5ed737748968b431b201dbd35d988560fa93ae032856a7adf2fbc3bf30b2251e2e51b3c;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hbd2578565c1f2d359f43c1c78d485915d17b53c08debcbfe0ccaea9b9e40299fbb45efb9fe866baeafbed6fcfab2108bb40c095e7588ec4bfb0e9b294203984ca9bfea512cd72d05f37f96a07ec47e566edd50329397f54bbe854b7dd6e54bbb4da4fa1b6deb298564;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1dcf282c4bf4ed462c1e432efa2674a927f1e8f3188e3279b97b7c90a09928367e16cca91d93e1f86654e0ee3d4234689a33d370611f7e53720b361215370739114df58b80b7263ae32c430c0e827e583cb6aceb5a0799b332394ea72b29ccf6bea083234346cf987a7;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c40f7e563833a9bd86ddf09a65380c85fecc2f91dd016ecd8ad17e49ed65e32cc7ae05233a3da818c7dc58444e769a16686c891366ff34aadbe36ed4c6ef5b0b29626e7c81763891779be142ff96279161b73fe5cac128bc9cd6a223a36a51a823e41a0332e4ad3557;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h116565c86f0ceb17f024df727c8163be1ec685924e5eac92ddfeb8eca1ed33167d5c2a629ad316b7a93753a9ea25a51df45131c230503a299e341631cd4bd50ab294dd99f52e29c4c47c3a1e38d36507b3f5c6dd8396f475cb172cc475a0dfa6ff5c84687d37f267df;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h55b68cb4f75e0840d5da22ca87f734c868f18e5552bf130d92ccd595e43006bd02336287e01fb872eb8658a6dd56631de8509e25e9339d6cd7453a69bb66043f6f8387f1459843c9fd67a93cfc50574097705283754590b86ce77ee2f2d60d73f29d32b29d4d56ca4a;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c11830a44a8eb14bf85a7497d3c7ff6b69319dbb305d51e0b2827c478894963ad1c78c19ae6aef5ffd08154d696fea70fe44b506c4e55acc796a81435fd3f47d593232d0cd0f71e0ebf99832592a6ce417ff97b9e49127e78cea908c44b18f4c243faa80f4c0a06bb9;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h51cb4ce98d7b96e2555dd73627c4b8c91ece2d407f6b44cb6f5e98eab11c1197078b588e612aa3ec65d50410900ea820bf711e1f2e28a65287c809d1d5889849857a5a2e8df75cca56a430d368e23a62a3b4eb45e0aa36740a3034acd7d790fbeb7e75571cd830f25e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h89d4bf8a1d4a9408003c4dbcde0ee0448b5cbf74b1dcb22136dde313faaf2aa17bbe98ff8cc11e20b5db5c2d3593794857133294a6768f9a89e02bc166d0abac10e5ab1b8cbe2247b9eb5c62397c1cc00807cca29fbe87f9cc192f0e2f322e1a4a48643afaf76b1c3a;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b2ce909b3b1f5451eca6933a70262d488f407cf481c0dc066ae914d2374089c8c2eb10e38f78f90e6eabd9c87136de1f792de662a3a1ddd17c02e74e8d7ce4ec92ad0c9205ef23d9eb35617eb483ae90b6424f557bd7127228b3e9b2bca010167b8acd891a132fe766;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h11733d255e3c934cf4caea5dbe01e2867801952f343d043bd18957b2cff34191b526c184b4ed73a4785a855ea40bb7bb2d96acc9a8faf987482ac5122225d54a741ab119a484eb01a8d46ad7d22d00e7b5de86b564c81684bb159a4411fba2c650bc0d6ad22435183a0;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h18c4cadd5e1c8f3a5fc231d6d79d53c0cd140fe5f7182653be3ab8a1badc2d39bcf8255ae6bf184c08c043429efebceac82bab28aa66a51cb9d308fdb356a178c31aa0748bda83e32a14a2fcc1cd6f666672eab1b504c505d0a92801d77325a16a96eeb4bc8739b23a1;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha4c2507b8a843f13719d816084ae694957dea610eadffdb296f27b00fbe231c97d5c32ad8377413e65fccde2231e2b74c348481e2c613b9b940a1507b6b3cc7391f3de29ed3e25bcc1a1818f583597a7fde7b410124c1c26769e39f770d3d612a1a0afb57af1e615bf;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h86da36cd9ac01cacfb4d8ff2d53355719652b496e36afd3cf0048534a58881c6bf36614a35d51c5f5b350cdfc9adf3b2344ff4c33900ffae5834c83e7ca80038b52fac604f5658fc62e3b5570c9e456041685e04dd35b740af669d0497ad8422f57cf446b368c15071;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1298571630df0d75b01858d2e48f332303237cc3d70308deab8c263d15e5f6d4d5936e95b59b7e70140018cd281864bd94760d2b01b1dc9a9a07eea0937f9f25cef550e39b22b88277ab5715bd3772329104aa98fb85d48009a58fef7ee28e4ceffe762c31a20b04111;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha57c58606c40637b1c6cc16e6fb46756df239d4623eab6abeda497a1254a5f245b4b0ee89d8f619bcd4b117f751058e0473210799fe1c23e423f0354550f37941ea927d2aafa1ea0af1c7cf2042db90e2dd192ebe5faa7bc550b4c28bf3023a11bd45d13eb1ba959dc;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hba6d71b35eeceb403076b970611557f76c16e37741b09be4ae9b381ca2f928c9148336f1542599bfbc229a3700f1cbecdb5e6122c507e1e300afd221a1b018edc228f3ee1a5694b526a19cd90d224d1c68beba0e735f0ea0c8daaed8d54aa7dba379c9bc9a763f27d6;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h7c8aec4ff57a09d819ab1e49d9ce01cc14888559c9a2f91ae758f32f69b7a5984581146ddbf8778165d45a9b6f0717a8d06bba01882622a576c91f52644035254b6586c52c7d2a97ee7124c2a4dbc68628874ebaef27924c6076ae1d41a10b02404cae6dffe62cc399;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1908407e09dce169232bc8f4c22423b23b19d38a1fb21988517f08fcb62279796a27aa3296d696498d25e2ed296f172dc45d462fc04e87b79b29f1c78f5447c1d2db162748aabe19c2c26e1b475dccc58f1c6bd2b4e50a5d8af8aa510b605169ba4a6adee5656ac08c2;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h6bda09f00d9977c50b82bed610ad849c84f3f13c2822c08e1c7f47ffb9aaf7cbd7a6195d331ee98148d396c509e44798397039e1e96310bef43214125f93ba10131dc19b65fff487422285adfc1a1ca587f42dcbd71568ca02846603d45bea3b0d2a056e663f5d5f00;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h4d87720c2ce82813359bdf5bd234130da41e5e474ce5f69c1635ffac0ae7996b78932a33881130df4bb7b967da2dbcc6ebb941af0d18dec01f52962c81bdbb8f6c6d06752a3664a5e0eed8bf063cad8aef3372ea293929c160ca26250a616d409d35ce14491aeaa045;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1163f9c76133bc9698b22242a60e357a7432cc7803010d37618b4e9c6557ce54b270ec59aa3a0e704082e453595dcf004e0aada3987d147bfa1ac812a4177046faaf6cddaf3b85c2c8ca94b506bcb5f49c615c05e9dca3e21ddb27aef970245ffc6e152197f867bb155;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb4b7e27d4a63971e951173900e0192a8be8bd1de78c95e1e7f5845301da940eaf4dc0b0c4d0a787dfacbdf6549c6e168f0b1b117f7e91ee5d669ff622852e39ceba3974ec3bba6d8e6977a6edb4ba354379f3252ba3edfe916910e37840db048cb225a15b9edef2baf;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h8c64a7a15cae4795a69a8e9bee8ef046c094160b089769c41ff3c1efcf25ec35b04268e6eb12983e194912fb7d671e1cfa6552977ddf07e14d80dde6e892ba428210cd1d4a0f7d7c8346bd29c4fc2836f9e232fbd14f389d81343093600f448226b742843dede0cd01;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hebbb88de08717be13d22b1b17ff4c66cfaaaf0ebb4581e9e5f6c9df84e8bd63cf5402daa65da5680a9971a5008f980bbbc7ae3b0b9be92e286b86561d380dbef288e0fc435a15252f2a9a02b696010d86571f12ee42907793e3d0f840112600d75a2c05d11f6a6bafe;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h7f7c07ff057b4bc32b3cc32a082c07ebbcad97691616cacf3d5bddc6d8e8efa5c14a6a0c944a8bd0d582fb7d037772e16116c146a6985b47387b0b61a1e95f9dab25113abb0cd0a222a0911fdd755cd8b89c5eada0326265703246d49f4c52924384cd19cc049a927d;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10f266a06b1b4b3da4a14aba5817aa1094ad831ec0ebbcd4bbe799f4e8d81fbaa6ae8481f104a61a6bd9f81fb2ae6302f24e4f616c16f43812e647e5378cfae5df9c3501bd14679242c36f3f5d295448ff89ed32c59af624892f777d9c859bb2f0d8c85c1ea6065d144;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb7e697c8bd7c50ee22d5b2b7e22d38c97a495105043bd1cb3d3e4c75728dc6f85e6507a7285df167db8a4bd467f6b5002070c149d597b5587711ece9e0dc7b8ea356f7dfae01752ad6a5f37a03c6ffb615432fc612bcebc6a81b1b7da108235c211ad7c13e9929f079;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h27ebbce873805969fc1251b2b2a65dedeb596a0131079444b2f9d58fb9910291fbe89f11eddb0e827adfbd8d14c90150fa7724826cbd5aa26957f40e57b82248824e9cc19fa7e4d499a8fb37d47715369e01014f5202d597d5f93970a7855a34f5db63c8ea04c7b59f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h19fccc55841f1d8b2c76c7a411bb45d077ef93b01bd2911404febbb9c60d0bb0fe29bf7a6246964300b3bc9a01386ddee1bd0ac2705dee6c51ce641ef328f90cbfb02477025a4e289e9aacbb4ab0528ea9713df9ed368e4d5f34b5ed358c1a9caf063b0fd5878bb0f5;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h6efb3775df530a4395e478f1eec395b7281bf7823d9be39197da4cab02e4d395b2f1226f5d753b864a1d3b9ca662b73cd20c5766d142afd01e7869f62aa57589b32a1ef247265fc3790802622d4d21d5daa8ef427113110cf1f96c6680befe4f8f33ed9af66be2644a;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h750fa741f0102e2fc141669de57ff24209168ef2ac4aaba9442b9b6ef53000569c141665835dc45a7e5401bde0f71f368de0de27b4b5e3c642186b33a195e542fd3e7abb9e780ae7d6209217f7b49a6ba9fa27bb9299b8705d5650fa539e94ea3a6530660b3a4bec9;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h165171af5901fec4fce27e0f25ce0e30283eaafa374a417d518d1aef6ce50fd467f6893ef3842e19a7f1adfa17456cf5c4197245539c371c1e23afbe0fc4d7e68f5147f3824087156f988f73bab61badb5700dcdb001f560f03fcf27abc0535562a3e71a2164186ca66;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f45477bdc9d90da96d024b9c9f136142a3aad84d65d89025d78f25ddfa36c5f718723b7b3f51596e9e02a8c058772be783e5406119381a66617385e51bd8ff895f9ecb0225ce1df22428cc08307e304532d9a452634ed4f0c80da494e7e90c3b8388fe41ad01497303;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h16c066519e8ea4b8bdc957bbd64243074faf3026ba98f5de9c8fa665f3f00d6e774658d03040d037ab66418dd4302f91c44709be5815dd4c1b9ee75fac9051f27bf2fdd148e0c632822dbb442c00bdb44214cd420d3aa3bd70ec3a3188c06c791a0a0c4e7b9c4e5dd4;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1742c0e2156476b2bc6705e2d85e782f64e35ddc64cc3ecff44dbf5b18764c6397cc01ce7b8ed898fef3b5609cb689069762ad0dfb57d02e3e56118e55e85c2bf380f557bae282972a280aa47b61457ec85ea41cf6d02f886ed16822f8f6068fda2a128645a567f8431;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb1f2b4736a25e93d291e29650cade2b56f11e39e284754e55cfd2c199c64da7fef911f4d8ae34a5617b01ae9802f1046075cac24e68e44d19dd6435241149819e56a263ea0d843d57088eb26b2b9cf51c850e94996b4845668d68a814b769a5d76445be0f2117a2723;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h101216ec6643f6a556c436dbea707722663a358171869803d81e9fd1281a7dd8c21afb9fcca7464502c902af6ae76b40d5d1534a342710c106f2b1ae31f0ec84448906faff341d96e350b02a88d91bc24ede0e93594424a94392d6a06f0fc773663bd691b445aaed0ef;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h82baa5e1c8b73ce4813d3d31f1092990b87dc5aeef8bac740b93a3d0b5cb0e652cc9358710d5b3a774cd0ba39430bbd8f200d775601272fbb307f9a20149c5eb6b44898cb27665e473fbdc4e9648c9400d512759c791a5f40087ecd8c9e9fccacccfb525cae4c12634;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hdcd2720590a80c02be35e232823c4377d12660c7cc5c6f7a876ae55229fcc45b7c9f5ae194c830560d6184a3fdaed3f7252d2f5a5626ca1d0dba254fd61fb0fe32ce0ef47d7c16fb1385ae59f7a6c4a7e915f3dd2889fcec09d80f74c644328f423a0c185e910eac9b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d4a71699ff6d440287edb86bc9800236f8b40fe78566efe1e4620b2b6857f90d154c0592891578aece557700e9de2c3d5960159e90cf8fdacc03425ad9154b73788595067b54015605e48271cb2488a1a098701cf2b0386fdf8e84610371393aab287cd9f115cbd926;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1cfe7b0cdaa4ed8a6917f38f62fa64836fa9817df8b25f4be6c0bfae94e39d465bcce52fe113fe87effcf0bb9a90b5af9ce0a2ea35c1ef57d4730b1ef536a1fa3fd996dbebc6e91398a09e10d6ac3c02a628e446316d7343cf5feaba30d757764949b3f9840fa66151;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h67bcbdefddc56790324e2713e5ea43ff361fb011a72b0b0c616ec06153294a57110dc8c93d9bf801e40306b86a704845e10198b8aed4b02d3f00f76f2080e73a7377d230558143f53f598da1630934a5526f81f95367a8fd69ada0b8ffe1828875679465d8b0c7204b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h9e85dec66366b9a7c7528621353f98ce60d733441f08c7c94d18f60633f35553b96e6d2bdebd54f7a1bbd7e9ebc62b27b90d4a234183c5f49a8df77a99aeaf0585490849728a6fd2fcc87e4af194dd055106f1eedbb80bbbee352d142ffc2018c1e81f55c156984f23;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hbdd10b14cec001f70d9a88481415054fb47a97e75feab21e0240f1685c5c43ffa1d44c5723ccc1cbf1a8209f159ca0aa81a0562c89eeb8a4dc2b68ee85c83db357a7213a27ea7fb04dd56c1472d3a8e40c869b444dc29d4872b4bc23aac32dbeac3aa370964f7a9f10;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h267fb4ae53a05e65f71a68d35561274f476f5d3f995be60e635148c9e82287687dddbb977743db919aab46bb6f562cb5b209dbc1971366688196b94554f37d8148a428b8f1543b0c075932746ec74d2bd57a132b0cd3c669079f9841453159d9559dceb3d88800e43b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h198024292a2ff1114b1c3856af8dd979a913ba80749e813d50e990adf763decf4d3c7431fdd59b2b365a3d10e55d6d8d164c54b5a98e95e8766d9b9c7d0a9486d6f2f25e953399f99339c831c1a7c11a2077e562d1dd3a0a3c264e079a737967c05b5af31c785c91341;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h17e1ed72e6e1109589a2128b72bb049803feb3e74f48c035089410f805737b5e6f6034c2de24b33b1d412fd953ae65b53bd995ae55d484f0dd16089944f348c6bb40b5e47c67cdb871a661a1b49fcbe678590862476d362e86fa4ed1600314aa0a7ba799fe9135145d;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hbb708f32fef65fc4360f33d666bdaa49cd8e59432fbc8eb306bdc5a4b77d872b9c8721cb12a9ed1b74340f3d8bf735e374539260ac99d6af5beb2c61d18ed026ebb16a66594562d63a04312e96949d5f49d428f5463a3ae2e3b9511850ae8b6b3f635bb79916e58d47;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1329ef681d46fc6699abe99187ceb26fccf63278e6b1656aaf8f326f9f5e1729963ef7cf8aeaacf66245f8520a54a56ce4bde23a24dbc2df57c7f1857a8fb269267a6270d7eb6782721639dc34d9ce1474e8971faa88de7b363c556fc352b1248cf32038a02696095e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hbfadc6cec274426173863994fe5594dad2dc868c1d3d666cc7819809803b2c4acbc316fcc9be76b97d09b1173c681cd1eb1653e276b47f725cc9141b63961f90d90d8d6a6efb9bdaf35f48a004a5a6e5cac4c06d3cd31abe9089595f2fb799dd502b5c558e6041b291;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h150871376a942e6e93d71a5186e7970bc680d4f557c71678113c7ccf092537aca432a378a560898af35a0f99241c381ec1d2d2ed730bd310ccc9af7f93312bb89fefa8eeb7b016fb833f0f8d3ef3f5dc705a38db7b1181ac7a3ae2ebcf7546107e607369984286d281d;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h4d6d7f495bc67a864aab0eac1dc6ee468b3e938bbf13b5b56254af8c474d1c0bfa8e5dc9f61104289928fd8309eda11bc22aaa15f17b0f67bf8b5bf4a052da5f57fcacad691a38a9244efd8ee173fab43794201cb27b2e5011811eaee938873b0b52d01965346943b8;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h410798feccf2b0aad181126da9a5236ef432b23dcf10fcda89e9ef8894d904fd5a59938bd02740f87519352c2a237da38c57378d5d9cb9eebd3e625169254d3ce8a3c98b93ac06f20dd0ce667b8b2ce1a18006247a2475a4173e6fc2edf621841346abb7ac14f72af7;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h45bd2a9b1a204cb0a0f31c970e86393848f6d1d8dec4ff95417c4b22302a9c867817ac9da62378da021aab45306a06618bcfa4d0786b97009bc8c8503a91638c8e10be925af6490450d182f5a220f342203275f4921badb0a52afb8cedb9a0f64e620aac0959555885;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1cf921aed81dd33cbe6dea45e3c1283a29d0f1a3db745f437ba74f6754de7bd9afebdcea48267694128b89677ecba579ec2f028ef243983741853439fbb957861a97c27d965642bc2f715d6b8f4e43d93e0bb8b0265e468493ebe7471c4152993e7e5663832f97d01b2;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1cbda53dded7c6417707f8ee4f0b7b1a5b5d55f1cf0804616e7cf360e375add820fd00bd055d0d537d646e45adfc63382307856beb89338a91753f31a4875ae23c0ab74ac8b4aa744f77458a50da355ca092b498cf52354dfe045cda43ad2db9432edf21e0a6c0c79b0;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h985f85d5682a9707fb92c78d84a0e355e4b5ea130bc8254535eeeda2d4e5bb7f79d90b9fc6c53ff9a87c978877bb0f460955afa2becfefa4b5ebb98c882c353eac456a03662ead04a89cb4baf9a038fd5fce80f8fd7102cb6ca9f81efab74d93d9ab07bbf9a198ebf7;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1567ade15b88973001686e79c698a6d2e8a5964637823451a932054610cc231888b4134018936b5af0de7561e7d739b109a324e00a4a0f9ea1ecd8ec0db31901d3ef03ff980812061a11722e09f043e6d6e586b54dd6814ea6ca28340cd5ca56d4383eda55ffa9d2913;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e4e7c10626c38bbda4ad60d543334ddde7201b5c8dad04be43ef73f532701b78959c109f584c9bee2ecb53cfdcd6f80c2dcb12308a173ae399807033058424ae96223510b95fe66e6eceabb99ffa0ff9ac69617cb412be975776ff536ba6679197b0f981387114bfa8;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h190783c551513773ce225b37bca9bbd89f185d7c7a8f810ec8f3f7a97b473e573036f3552f4b9da2a87265cd634d8b7b35dcb48d7fe6a59d616bc187deb12ba8b25d954b41ba84b8c079e6a85775998d5cc76acc7d086cd3ec772233195c960c8c37028485933f4dd2d;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd25e833c013c2cfea0a955df9d1bd67a2431e7a7f9ef7d1b739f92e097b97a82a2a1a2bfc5350d5fe0921b76970f1249c67bc32daac2005810f23ca79f150d0a8de982f2924433eca89de86deabec1b887ad5e8761487f32654a607427ad627533c18afae87035577;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1840457282126b41ed77c33da1d972f7fc01f67bb089f6df6233f3a6e276ebfad9c668db4af45da39ae696c8547acb94762b866f5d638ad856864bf3d9ca9ba08adcb7965347585e0fa81721ace817dc729f7c949528f65045c921135ba528247ffa9ed687332f92f9b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c60aa3ed64b24f38bd8f0be869a0161a92c92f0b71b656cf483b4ececedfd56938678f58ef158ce9aba0c15894c05bf04371493896c138064f9f87a81a440fe746645b5609d80db14631ac46847436163b08a2f920a9271d0adfe6234755b3321f70aceac9c853d3fd;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h3ca92fb2147f56c36861f7c528c30f7d3eee9799562d2431d25f7efb9eef29efbd251fea558a599a3e4266ebaf64e046ee3dbefc1e1b6b2d9dcc157f511ecdb644515632c8aaf81cfc28412794b640fc8faa6b2466779dae71aac2bad84495ae4a2601f08412e67e24;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h12be6ee285636dcb4ef2a45311b160885aa5fcb5f731f68683acd660a6708101119c236355bda7a1f89eab740919e15412f57f1fcc1d17c0fb737a4d3f6d65ae6237725b248698e79b2cd029498b3681c12fa106596402a96354a128202f829d999abffa13fcbb22db8;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h14544e2f97519dbd0200ea7525c0526d20ef4b707c0a80eb46a62ae5217c367c81e3dc22e07ce936d2bd849f59d54354290ef35e666c9e1a672f876e99904c946c402a28e9a4199885789755875120a613b085e1323cf245198d7b7f7027ff6362670309b7014e4f23e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h2c5743dd5f4605e159fabe9694f9bbcd3713570e2eef0c0ca8c5e4d55a91375b6fc8137c9f7f17868e04080690a6d94cfdbf4e14b047bbb914d25bed85a364a957058925584e08c166b624301f93079357abb58e70876a15c6f59a6564240a797b92ffe82b4b619dda;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hed8572f840e0a7ec818374cbcf5c51be14946ab1220929ab099a7ab3798c3965993d1f78422eb991316512a25854e3c663876a79baaf0e1ffdb81b4c0d1cb4b3949e9aa316611bcb52f9ee11b925a855bbcdb9255b7c993f9c0791fa7f53cd9f59a581f457fb3c1354;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h4c8324253e897c9048baa928e7dfeabda81e40e0a3da8fa793dddf4267d687933db9cbda4294fc594cae2d71b83c9ecba0cfd9396c9e1f03ea3a5fbd5e1a4344e99eeab0ab201e7373762cc68d7892c10cd7a2802cd98361e0408f493f7731fcdc43de96e8258b50ce;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h6c4ca88286c8d2775ca7fbb07d06b11fff0c405110ac53af7dace5c110a88165f1a28ed3ab2d0cc7de56f84166ea6a8c78f0a27fe5dbd849c89c9502a5f6ef0632cdd789299f33ea1b505d7e813cbfbc1fb8fa4a064ac8378529dc5b4d057a627d27d5df51fd563e66;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1523950c1aa3200e90c58682963a6e27fef17a3579534137c208c07596850c1dd80696d85d5004170ed7193b96952a2284ddb913fb981da05d4c0b7d9741b2229fb9968a618ddc9cf442909a9669b84ab0abcbbc83d08bfc907dfdbce90065bdf1331190711d7e9fa27;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1bfbfab350050f1585e8601dbaae226ad7222df0cbc6be2c3012b3474828cf112b30e14cfc72268e2703205c60f5b49728914deb5dba77bb96791af086e3ae993b6c3090aad0b46daf786f415a2db93709e337dbb442d91e5f18649c0fcf58bf6362d1f857b90ee1858;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1796f024a42712c114498c6a7206ea3ba639371b35e081760aad650767c3604bd09e235960811f05e0d5cda3ac9e986ed429e213101df561de54f1ef7e9ec72db8e2590382253de9f41e0ed595f970d6c760925d15285f955bab96d2cbf42ba5e8f07697a5b2af941af;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10cf03051228e311a1771d97da6d38d8f52112798649eff171620a3dcacbde3f79aa435b8434c54cbaf843963fd424e2f60bcd27b1495a5fc380441ccd64815e192cacfb06f3409f2f78d9b475d100ad117dc1153a0ddb147a6b3709b356833e5fbd719cfd8dc06823a;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ed2521ca6ebd2c4bb0f8ed6da8c1df2015c533b27ac970df9c2a7c11d532b019ddf61adcd96b7cc05ad03f62a141f787baaea514263e89e56e357b5d9dd3b8a402388302f37bc1878405c3c90ebdd8e39f1fcea63d94b5d8c9b42a0c83487f4126a3de1de34607f086;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h70fa8b2b1bd8e57ecdc9b1868a341222e618e0ce6c5be6ebaeceb217c7ff613cef85ce71f14896c3be29720ebf61cb1cfb730af54ad37c2d955297e061aa53cbda405402571593a2312c2657272c869c229326c6ab2e6a80c3c4652391fb9a565b7d96a391888a45da;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h122a4804644c1c4b4e90ee7ec33370d7066650f5ec499548487fb33843531c55a70dc15b060026395e42f5ffcd8a9ff66786be85ae6b72c273d8d353fe5b92da24f3c5e836fb7885964736e3c71234fee8fce5b142d4365dc96270d61a5889d6bcd21e237bb1fbbc9ef;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'haa26d716e8d2699cc7777ec0439b5cb489775235ca0a382bb5c83c05d228798cd5148120ff563a416e676b05ccb4cfafa0081dc408c3dcee8e13adefe9944da8853c2737682ebc4a82271c9cda5c22ebf19081a55628db75b8f99028e05c3d1e8e86dfad0b47b27de0;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h7cc34262cdd711b481b526f209957be4c57205a075a93195fde48527309bd8aabd08769a7069b464f5a3ee542499ceb2770252bbb24dc05c9b5d3d17effde520f68a573c5d00f3321e130bd4e8c9e4a7d04d36ce75f898aa80508066274cd7d52212186d818d340ee8;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb14281075f76fe018bedfa462fc048676d5169b6d2d54d0e08907079cba7eee9c24459a15423e422c124f13561026307cce68e8c9bf23e37422109ffb0cf0d293d84888205e9a01f03ae0716d033dc16aa9e360c859c5ff2b117aa26ab84cd1e5833aa20b0906c3b95;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h3e7bd5cf5c5e6518564e1bb4a0069241dc6603492731a4fc51152ae69d63a9912b8de876355446649d53ad78babcf07abce18c613555caff9856fdac1d7863ee2f59c641efbd86a80fb3eb3d4c84b2657358cc5f162877c0dcdc12da178d0204840dde26e694efe3f5;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1478d25d27af0e7189b021b48b3092281f85ca3fe38f33cc32e7fafd5c5b3030b20496cf01699092aaec235c888c96a3f1e30286e75059f63e8f2aac5821e99726b28897c101f9d1d8073d8dfb68fdee3b42039738fd56598b43f410a2457a31adaf57d2e6475a42b9e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hdbdf56030f5e060f38b769be916674b30950bfc2fab28082806be818b86717850a6ba04eb4be7fca41d0874856120e84187cc10bda14091b86d2336410cb8c57e551ee6a89562c367d0666627196b5c0080d6832c626f025de2dd5391dafbbafd85062da46d0d37580;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf0b11cdf6c7049f69d2e8c5b1111d6804d020934cc01163d8aea352bfe23ac0f710ebc17dfd0a88a91e195d847a189245a8fe7b90312bdf0d470f51e50f48fdd07d325d2de24055381d4a9161d6baa963dde1d235ecb9caf54f9266f5b5c1f541a138d8b947be977b1;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd17eeafa8edc670e0d94df42c66ec2f8e6b61c2e2ce88dac680f7764e5cc0ce7f64902fa87d0abf5a08296a6cd9788f2ac4c447dc245101a8b0da9a25ccc3012b093c4426cd7b28462931fd0ec721795c74dd92d4f73a1fb17fff3527d8231672820275266d9af09a8;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1de37ebadbdf3163e12d7b689ac9d5c47770d5d68b646606324f3cbbcec3d8ff437cafc13dd6180af112a064795c173136169ff290bf93d7f97f70cd880d4a57fbb520ada7e40fa8b218b7620acee6a9f69c061a5760ad198b65418c07f5339c09601efcd0b0771c206;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h9825121b2b17696c253961cfb18d042857603c033e00d7db7bfd5c54ab120c4fc76505f9d8e6baa7ab5492bbe46bc53f000a9df9e9b761f63fb506b406975027ce3e4a7d782e7e7b7aa5a7ff8a42c99ac6cd77713a01da406cab3f6daa6774d6c1c77de94807288941;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc1137a39778f7c8edac04cba72d211e27239a6c83a5c92d55f69d6b17d5236b35c76aebf4986be86b1a96cc426e110130327ea94c1d661533ce837c8885d511a3c0fadde0a77e2178be68154053884efd90b5e7986c5a97b5438642600107317a9e33f581f584a1104;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h197b1209cc32ac9fabec7328cb5b5d0ba53689b24645a4508d95234794fa92b504ab50c27c2cf000d94d671250edf611aa36aeb22109ac0bfe8685f1f84c9f250501a4b6ef0afc05e9be7f91d5efbfe038675de5aaf2736c908e535b94bcdccf87e9f4f74073d901d65;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h243e5f54d0826368f97efc677174bd5c0a0b446eb729cee3fb2a524bc3bad47d15d712b32c2a72425d1511f52fdf4c684a9a57d343dbe5452983550785becd74acf80350d1af20c4cccf0254b3bbcdfc258d5669692150d562aa9d6bb5ec0fdc8f0bfef790ec5166;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h15cbd8d979d58f6b72301184b86fd413e828bdb74ed974a87e7b7ad922d78d42f250a5a73ca7214f3a6b5c8fd36f8b76eb7a7243e15b22411e2c51e1995678969220c51f5921f6e3ec5bed0c69484b5a58d97a1c1233057c90bf7beb34e3bbb43111cf63b3a95dfceaf;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ad03d492d7e058002e35ab95e400ca78ee0c72ca9c9972f153db2703948973c89682004283529d2b7b76b9e565675b9f8d42505b263da01cbb9eccf6156aa069c1680db203c5f48b4d2fde0cdcba105f212a5b80eb8919671ba27be37e0b4c172fbea24b9b036a28be;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h25b7b11136917a9a769a35c109f596f873ae9607634e6ed709ee04257f83a5b4a7d9a9a8c81dc76c8e0670297986cebb9d89d07dc2df73e7d53db5f7831db501d796b70741412a4e5e94363f04a6f2f6e48e9e91a55979188eab8aa7e70dce001fa43bf47969e99389;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1fcd80f3c320f2724031510108e02df12c30962445aca2e736a54231b90b2f032757d64a30e1a9bf0eb8f5c353414c5fbc494c2e4c077be8a4ed7027bed75e44ea9d7b29ae296d2007245614e2dfd8204d2a30e05e87c8da4040dd53d2c458666577f55d5e84f9bfe4c;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h12bdd0d3f576ba938dc25cd3838256ee55f550323415680688c4beafd440098897d9ac4552351dcb65270c7625d66d4111b7ae3ea865ffb20bea64312c2f0085161f3143fac807852a8e12d3e8cc8d53dc85dfd90670ac057000cdaa858c8677e4b10bbaeed1a42a29f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc27d25ec8ddcd9f0b1fb2dd5e1e271cef9933f32460fd2e9826c04b6e79c15592adec87b4d21f8b6883cd26c2619ba2aed39031357d980b1ebbe935a8dd249f40fbbafba93b34d41d89287a2a732a84ba599935583c9db338c6215bfe8dfe160b130176f5a52a48842;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h18d6ccbfe1a73c443975acf52ead98fde0b4ef365647fd4651f6f5be35294f16cfde51c9bd0d911b9f9fb0268173ee2341eea6ea2c197c50787c66926e9eab3e92cad0a0e2642f284b8483aa49ce196161f032bcb42463736245cee069252b56d7f22b983ace18615e1;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h286125350f3bcb31f3ffbc76982dcc7eb0d9768e699b8de43ee6f4378cd03b201a78269468063893d7473c33f7b46e5a424db5e2dd3f145351ccb245e0b1b9ef5996422161bb97fc85400520f6f83405824851d0fbfa62bca5f588601e80eb224a9fe0b695ce70d1e8;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h107dc0d21d999aa1342f568b9a232e5d19ef617dc692186290d44ed48415ce17c075e4fe6cb82bb939c9e364a55e668a98fd82863a6f4fdb84392fd7e97eef74b7e683e417529d2071da0c6aa0293bd1d0b1ead954be2f385b8459a65e119fee780c0064a9df99e9d9;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e475f553dd50e454a954473fa11366abadf86db8d04fb86d3d5e47afc2ccd0e141c47877f24e9c3020ff05598260e91a95822196d969b67fac9e961b4cd19ffb159d4ea72a9de782e28a7eae372ab2dc9718337ae0a4821e0bba0e9dbf281d8b687e10c9422484247d;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h36211e5a673df7e13dfb87245366e0247f680def2591bacdd35835d7ffdba9a92302c1527eb234d95e2a31e20d247606e59dc7d89c20bb74d24070835fe7c471a1c07f052903991ed5f571484a4fbed5c4b737c1bef15d8754d72f48f5b5ca028c63e6b1b446682714;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h114848d605d27598183c980d433d50bfc4ca55f747d762d2818cbd3abf3a069c05e097b223173c274e60379784a00fe1361ab9940cc5264a7025a698b8470f12896c20ecb2611e2fe744cb7ba955ac00b708782185ac2056f237e0b19b76bd1026334b7046b9ce17198;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h76edc2db1067f61bc2bcee9bc580cf1838f0d88f0cd5006c6b8f743b6bb73c15153aa1f6d98290eca3f65dd44499d608fb61c4aa4f4a5c0b1d2b86c7fbd0e7b64a2fdd78f115ba96c379e826d793a05ab748be0fefdf50cea5f780d8f28ee62052cb32814cc4443f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h6c674b08994673ced7adcd78d3b0a51facb93a4a78637e506834ab3017a2925d0355c707ea12e823602c777c362017d39086170577eea71225e3c3aee6231703bdf633198a958c7f9fa2eef164b63d248db3db301d8e824b4711b94e03118e51206b19805a30af220d;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf724e2be95984de93e968816611c53d8caef7c90c6297e49e0a283ccf0ed69f7a10a97be9f2ab2d599500a25b2b489334c1cc8febf7cdfe4b780571b2c8317fc3c244ba6c175cde9ea4d4c03af5f5ecde477b0898762b8aba7286d3192e6aba431afed2adc35589800;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'haa247935ebfc2139883c0b323e9c620ca050ae6aa6ef7d1421b035f423830dd20a5afafe6e8d4b754e1074a967f94422e2c7a58a4b4de648747b4bec6c589bff97200cd8c6cfb5921c9ea1144ac8676b123fe4bd22dc731a0105991fb9888ffd8ca162326e00703f6b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hee2d366d602898b7287c634692ed2f8a5d21751cfffcab6a5d94f68b76b25cddf5871056388148770d14cd8c93b643294ab75cb26ba5027a0946af60aa191465b379635e7ba28b6e0ceb94b4c1bcd887712b79a354d69a467c2f0f1b507dde85a3a6ab6f23b446679e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1db322656d0a642b9a6a6b22d89b971aabfd0f08fb8955269e5b2b343c986ebd71eb3d52526be0912a22dc78f313ae71426a9e507936bf513a6c25a896409bb3d9ebf64ddfdeba8f3448c1ba4b3da95aefc0e86f2d0c824bcaf8475dcbe740da3c21913f768f7970fb1;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1866b706e65e0625d991059db52af6cc57d5fb8bfdae569027845d6f52b4495d7d50064cfe3ebaec43a7c6f6b04dde67e84288451342cc7cc458d0ace2abfa6346b3e51e09e169b9478e5d3f83382f579d0df23bb604b24891d61b9efde75c951fabb7abc010cbb0359;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1511a6739b613015118ace7f42e443fe4512e1339b05b08f88c3d422543cdecbc97ba5d91565319634b74c69a9ca943f3ce35867e934e49336e133916bd456a693f58cf186d15b5039f9afda5e5dc4827b3cf41b921351a11677162b80394190f907e4a605bf879b09c;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hae923fd28480ccaebca659bc1fed93a28266ba0a410c719ca285cb88a2fc93578ae6ae45aefd3e53baeaabab75098f2703c04c64a162a357fe1c553efe79250d5ee7d03833ac7b31be971cb89b4fddd51a7c301ea63cadddfe37822a7e3fecb114f8cfc6c2f1fa1913;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h989a7b9b195e14c94e195edd0bd98543c468923717da4fc477be25e5b5b1bf80bc3cd0a960c826ba964cd149407a416657bef84c70c1c3ecbecf9e37f17fc97c269e51c402117e301f7d856b1501a3dd20dd39851b98c53b37e637a6302fce43e294d434b0600a2080;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1db0b79f50c2c9759e1ce64da0d34985ed455f3d6db94491942c3af7369d2ef49b7d2bfdaa2ba1bd9d8fb5c08e16ec0ec6f6ba523927548df18288d844abc084ef6df2032ae37ca391e9747b6782841471363d91de94b83bafe9c07593f109f2fdfc386c3742a74dc9;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h137b1b54715a9098c88218772fc1b0399b9a4d6f6878ef001487e7fc2fb0a6df73e9d4ed46d2d90019cac9478e73e3f27c78a501804cdff36d55d965363cb702d4b75db314e2166a6430ffd7bf1ac4f8a784fd2b6fc75e312e83bfa3731e2a3c8619ed365d620ee34d6;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hcc1e41595519045cb202ec993573f06477ae4389bd61c8ef72d8e80cbf9f4af3956a01a6d94a1f45ef0979dd074da882655b78a9853d4e85a98a05a23ec4512c44c1cf2439e60253a2e0088d37c773de2615ab74c93ba0461bd65cf960931620f1c7013f6505de388;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ba827658daa19514b4053692a28fe4dd5dfeab0effb78669520fb49df8e2bb95ddfad50f5d0e5b27d28a6a980de5901e418a593161c7be7e0e9f14ab152111ea9a830a7e39a9c2d16ddf2c2276552793e7b767a3bbe7e4bded3f011b31eed8c781f83cd28bfde99bb2;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hcf89d3fd84b0c8d9d84fabd202419470da8933ca035291074dfff6ddf3ca2340ede7ed0bff1474fc214e08d8c2326b23911c4116cb155674bc2d9d1036b3c3f7d8dd3cad786b9e101106551e332b75e2d5a4d63b9784b51f1dea3be1ac4ae7fb6cea00c761d00e629e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc671bfd3fbb491f89fb1704242b3e0dd028ba0c25081a1b9cbbee0b0ed764acee9fcd0b0a88e0c3bc12603f53f7d2cf35a52dadd2146463c35515442a722b22096108d93a0523dc058dde122baf44e903b35d5fb1a8d2b2f01bef18240f7285377c09517a7c9d1c567;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h775ebc79abc6286d5bb3a1878c07c13476a2ec2c4d6fe0bfbed9f8cab7bdd238133b0129ff59ffdbe3119bbdf4037b5ca6effae35c8cbee8de8a0a05631d5c5c452f7f1b4dc44ef42ca8114c2035c4f27443f0eb5aed10df704f29713127aa52cc2823772bfb1f7f03;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h7a7e7636410059bd580a2d982d43cb34958435cafb58aa6539adf2b4ab3df26b9d9621c7bd1e1217bf5b3d9dae55d457d8ae8716ab934cb4e309192df9fc59d323c7c97d8d9cfb02e3641f120ca5d5f1561c9f7994ea850d4c0cca9dbc6f430191121015be4b3cf154;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d8c6b98697b9ae87d04ce44366314d158740172dd2b24ca79b064142a70f71a80670fe778a2ffd26d667758c7ea8352a7f3cdefb69294525788278e8e476283ffdfbee8cc1f2d859887a58f9c34ff101f75cdd58c3366504bce47b67591d8d12a4e9a83be5020a6c6b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h191fc703bceed579387d0fc36f07c3a3334985731a5989ac27ec748f0495461e9cf59656cf55b3e1b977fda5229071653b3f1d996b3cc7c1a2a717e862b601a63ed853f604114e528ee3f08b06d85a9be4375c04bd9953aa684cfd01d37c8046d501633d5ca627e58a0;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h460ca9db5fc56edeee0db0c8edbf4dc87660a8d3b9f9a084e2b0416ce3f4bf56427b74f06cf7151c13a5d0f971d7ace6caee40a48313731f4964d45a1f6e94ee41474ace1bbb019a7e111db4da7c1623d56f79f199f10c824ba69b7e06204356a282b6c3e55ca2eec;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h5acbc83147e4e054e940028bc610fa54c900b02e9f1bd58bb0eb9ae09beea6a3febf5c4dfd62bf29b95c5af5fbbf306a5548e28d2b4f7b57ff1a09c32c9bed92984756e9ae763595146e40cce4f9454607196ecab34c964f0b1642926cc5d7e3deea7e9ac2975b688c;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h154c981056cf0d2c7dd739c94eaeaa88acd6f6f8157eb374a5f4310f2bb05c5549466c3dc1990419c261e011395feebf3b0314b376e262f1123025259a1604e8129a4e26098371794d45decac75522953afc88b512e092c131c9ea344bb8e368f77cbf8b1d37f7cac53;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h16635f02c022c0f4a02502ca1bff8d9f8ee8614a4a7a06a5281f65244937722892e41d45e46962bc7c9da5098f39e67e7851b8256d4dca89123293c7f0da4de90f35565678467d09938dbb0796f1b5c4389db0f8338e34add4a3d7f5da6d3b48adf6b175596441d46bc;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'haa4f5160c56e60c805646eab4323bba80359ec13ec58f16b6cc20ff8935f68bae46140284d7c23234e7bb5625c9d7f6e373166017d6e4aff4461dcba43d465340c81c38b95f7916102c329c9ed2951bf0bd015fb0c48d520fb96f0194dca59bc54357dacaef8c677d;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h6c40e4be399e3578f7bc959f2537e221654060c70ae91ea2f2afabfc36f4d84f32259ab6be984838870e05a64e4f56376e73a5da69281f11f78e38fd78a924bb15bb9bca142d1efa63dcb726efee0e063ea82b095432ddbd470008f36cb885b9b0c72e7a93c86d03b6;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h2320d1cdcb8a900856601082487a5cb531041555c6df323226eade054e2aa6e8293b1908b4b1081308ceeca1cb93016777984265057976cc6226c5e36944043f4bb627d84a8f4dac477c0caa0080e81cdfa9ea9f0f5a0527f0f4f12f3fdb8fdfb6dca31f80078205;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1005f5d5f13d543b51c859359929f477e5bb101c4731b4330d12468530ac347d3cf3e6abb72d227c55d6e29cec23779bd3d6083ab6a33ff14438f9dd25c66ff3db991fe20202362c792d3ff2647d91040e9f393ff4302e8d0c967efe5e2eb9eab227d090a81a7475e76;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h2fc69a446853ce1bafbe9bf38ffe71f7a3d37c2621392326ce287e3f4e34886615e0c8a5779322127c867757f4e234b5c96a4e6d01f2d817f552fa4cc0e78fa1adb23beae6c28a04019bc5da63790d0ce42d8119f9c60d52d4a7f69d7610234f1a5346fedbb0afc1b6;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h12af77e8518dbb74e274bf215a4b58a2338962d95688e062333027995496faa907db305830826f9477cbd7f934534cceb77c90575b8aa68acc4161cd6a465556e4c80253562dc5043969c49854391ba0f0b421dca0704822a30080712944214b6135013b1b260553c2;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f5c6ac0df5f31ab4bcdfe1c42a161a3e0f8ce83f4716bb48cc37af4d6ed0888dcc0f3cd3b1ab3cb8cc89b956d61b0a0156293bd993126953888c032b4e98271eaf80fc3ed1b8c179600d912064c9210271e36c2a3c3bb913a21ee7696daea941523d48e3d76fc2a0f2;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h18768df8719e2b0848c4b8fdd72e770d8dad429a4785278add7f597a082b96c4f3c4a8a437837c97570c20e15a03592e38e4203a2910d4fc31153b59a7d9c8b53beb1973bb1e1d4ee90c8591f8c806515753859588ab24af2c07596bd2aab5122ae6f99baf821cca820;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h111ed761494b22e8bf1f2fc628bf00d09bdc7c1381397e6a8e83fad1699aa8ad78567d4e28d1603a4ecb5ba32f97d89eb1eaa2db1e4466e4f16f039042b885880594469854e3ff60d5265078ad85ca929205c50cd39865eb88563b2944b9bdde24e17a5bda608b1ca9;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h16bc8a28fcb5f68a03ca0d6312dea0733338a1d76242ae8e948fe8b9cb4f86d6ebd93cfd6e5f966ac76e78c826ece0bee97fe6bf9de7da69530ef158533cfcd179d35a53c2a3c15f4ffe9ecdf49d2fbf371322e8e48c1dc838de2f6b3f6ca05f4b07f1e33369758a2f7;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h142f97023dc24692271fd8d1612df025ba672805ab1b15941af3d0a776f84238d199c7cc9e7982c3a281c97d0ca654d928e8ab30a1d37897b3f0517b42a84793be72b0ab5f751f22469c9afb998e51349292cf7b334b3d95536cd36af2f9dd237f08827066f0567184f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf2d2ef2afd61eb45a255875ffb77cc11194dd6a88255060769dd34b37b0561957d3263363fbb8230e56351e0237d84b71073a53a6db915a486eb5526bb398fb2ddb973e8f617a42a1532049eaa461345ebe753b9280b0ad88772a5a9cc0a64ece3846f6ba4ebdccc6d;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10c69b1a54ef522c18d861db0ed8789b550cc27edce4d4e54fe53ab647fba837d1e4c91c79109a61544106aea354425c4545810d8feb4c81b743949cd88de3f452a921efe52efb1a4c72ea4769d40e01d9bde222b37191f255eddb93054d6ade9900132655ad4e1a4fb;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a46acf626fba5615a4470fb647f8617330a1103d293bee315edd72d3ff65001a9bea7abb12f6e3f7d16508de3a9ce5b2dc4cd126ae45c0adf593f208a821347bdbb0854b0f6ded45b1e9bca4cf392f17db6f7d4c8a6b314cf3a94ca2324dcd79dbfb7532f066ebf94e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h14900a267cf4360adf23a4cd23a515f877f69962773a32832fe4461ce352ba7d6abd65a0b35733506e7c2cdccbeb97292a566390409b69e89beda47965e6d6ae1e575eb56aeff1d43672af70f71477a4a7d2f090f6bd030df5523645dabaa28a587e677a35383930863;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha428e8446bcea4da787fbc0975914c8f6e57fac2c6f4580e64004923cb6476d63974cd5c7c6907418361fd11cd5a26428bf8731b5116ff3ff967813c52b4fd745053823a3cdb1238b710266856197beca0a7d14a9b936b5fc91a56e3ae91dcc5d71d0715e46996217e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h614ae608ee333f9a9baa76f909ffbb7312132d27c1f78bb7d3786aef7dfef73aec5642007913b4fb27a538ebb0aeacad1c0acbabcb34cbd4dbb501dcdc1a266702b0d80ae905a15e6cd725af37b494f27c1983d21545724fee83ddb09a4d030395bbcd25a3192c5479;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc5150a56f3cd111a48600b90789290bd33029f1dd9158e3a16de2583e8040f7cb0fe9ca54308d3978ae5fa3008dded0f32ac6f700cfbce3a30a246335166b33b97313d0fb64884f7cf2ac94ded71aaba55955a560c29188f689fbe5a1f246456ece7c6171223b89aa5;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10699f597abf1ecbdb6d46634aa2735c66e8fc319576d02bb69afa8bef4bc08e83cfe18b7dbecb4062f7291ad7dbb13ae1b359057190c16b4e9d6a924679fa0a5e0292f057fec17319afbe908e47d45bdf358ee351becd171b1deb6bab88de9c72def8b73dd2b66f827;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h18fd162c42eeb9577d672bb517e96982d9762b93b5f49277de5f19fea47eb3ce9b982d450f445808ae092585225f01d898232c7ff2c80b2617b06c5782003aa3e2eb5a8b32ed6b636931881287a56785315363b6b21bfadf5c0127ca7a53e3a9b9ccd9d7bfb1da0e2c4;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h7c209886fd49eb0da396e60d005fb7e107732d0daa90fe5797a5aad23ed17fb4844bcb7f32faf54bd4923b2afba95ddc931ad8263e16c9490051b08058c9e41f4dd8599648b05f3a6e9ffc642c4a90fda1a4159e938d299f249b2c369d6437ba9f53f64b6869eea84d;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1fc00803673521c19fbdaf0c4ef49a1980fec49842dfb01576283023e9594ac3e8da576103c2ab533da8c9a139d2ab6b8b8405feb8f0b1d12cf60202f1bd5f155646a148ea2d8e8321b28265da616b35f44c876a3958bffb97dc1499700271af7af4a5b244f9e5b3858;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb906c2f2b3cf956d7b8fc69d34dc76ef970cefa4c7051c46b724a5912cb917779e1566d31a131e4a2969ff319b2a51249070c176796b25235dc281bef2f964c873606a8c990dd6195d92d1a15706ec38f44d75593d3e546c892d08207b8aa5ba41fcdaf87334fe7241;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h12d18847045f2902594d160dbcbeb32c9dca4bed519bb2e356d05e6971b3b35ee7cc827e3c17126d75dceb65a7d5f9de9408724a537d741a14ab22bae4032d607be33ae9bcd01bca594ae00b8ba8ad27913d0b2bee4c87415aca1a984554ec40dbdea38af53811981ba;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h5f2548870f51975cfbcd9f43617932e75393b320a2a49fbf54b505b244f8b53a973a358f770e4ad4415297d227162fe2388eb05edf88b5ee2a4784dbc6bf6a900eff4cb2e7ad0e292ca247c85f835bda3cd6e23a84e110533cbe8854e40c6afa8cdad1cbf81c5d184d;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e867d3eccd99cc9acdf50bf4b00940c4c41b39946fa76bc53d7dc80bad15fbe161a078d25d603d40e74ac24f125e2a1f6616156c09ec0a10daddff4ec67b5fd8c3faa290ca3d69cee0844cb2cab971ff9fb18816129417ac8bdba70dafa31d57b9dd0255b501f44678;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hffcae7107741bbe159c8fbdaafbafa49b4a7b0deb5e4855b4a71c881a7b841a49621aab893c96e36a0b318326fc9ffadf2c3b7e0829931910cd760994053d9f8f2a5a586dddd4b367cabc96667fbc723a4d5f7890c75cf16ea60b3a730299b3fff76feb7e95afcd1a5;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb438097fc9bbb3c8707fd825c43eff8403f1f6fd45091ca690dccce1fdceba93bc806611ea0608cf0ce1bebff33ed9f09c83f4532836f297d20509ccca8b61c0186f847c677a69b8458ab95d32d478b979551ba6ea58ec52e4e56abd27b010d756bccac191db1f984b;
        #1
        $finish();
    end
endmodule
