module testbench();
    reg [0:0] src0;
    reg [1:0] src1;
    reg [2:0] src2;
    reg [3:0] src3;
    reg [4:0] src4;
    reg [5:0] src5;
    reg [6:0] src6;
    reg [7:0] src7;
    reg [8:0] src8;
    reg [9:0] src9;
    reg [10:0] src10;
    reg [11:0] src11;
    reg [12:0] src12;
    reg [13:0] src13;
    reg [14:0] src14;
    reg [15:0] src15;
    reg [16:0] src16;
    reg [17:0] src17;
    reg [18:0] src18;
    reg [19:0] src19;
    reg [20:0] src20;
    reg [21:0] src21;
    reg [22:0] src22;
    reg [23:0] src23;
    reg [24:0] src24;
    reg [23:0] src25;
    reg [22:0] src26;
    reg [21:0] src27;
    reg [20:0] src28;
    reg [19:0] src29;
    reg [18:0] src30;
    reg [17:0] src31;
    reg [16:0] src32;
    reg [15:0] src33;
    reg [14:0] src34;
    reg [13:0] src35;
    reg [12:0] src36;
    reg [11:0] src37;
    reg [10:0] src38;
    reg [9:0] src39;
    reg [8:0] src40;
    reg [7:0] src41;
    reg [6:0] src42;
    reg [5:0] src43;
    reg [4:0] src44;
    reg [3:0] src45;
    reg [2:0] src46;
    reg [1:0] src47;
    reg [0:0] src48;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [0:0] dst26;
    wire [0:0] dst27;
    wire [0:0] dst28;
    wire [0:0] dst29;
    wire [0:0] dst30;
    wire [0:0] dst31;
    wire [0:0] dst32;
    wire [0:0] dst33;
    wire [0:0] dst34;
    wire [0:0] dst35;
    wire [0:0] dst36;
    wire [0:0] dst37;
    wire [0:0] dst38;
    wire [0:0] dst39;
    wire [0:0] dst40;
    wire [0:0] dst41;
    wire [0:0] dst42;
    wire [0:0] dst43;
    wire [0:0] dst44;
    wire [0:0] dst45;
    wire [0:0] dst46;
    wire [0:0] dst47;
    wire [0:0] dst48;
    wire [0:0] dst49;
    wire [0:0] dst50;
    wire [49:0] srcsum;
    wire [49:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .src31(src31),
        .src32(src32),
        .src33(src33),
        .src34(src34),
        .src35(src35),
        .src36(src36),
        .src37(src37),
        .src38(src38),
        .src39(src39),
        .src40(src40),
        .src41(src41),
        .src42(src42),
        .src43(src43),
        .src44(src44),
        .src45(src45),
        .src46(src46),
        .src47(src47),
        .src48(src48),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25),
        .dst26(dst26),
        .dst27(dst27),
        .dst28(dst28),
        .dst29(dst29),
        .dst30(dst30),
        .dst31(dst31),
        .dst32(dst32),
        .dst33(dst33),
        .dst34(dst34),
        .dst35(dst35),
        .dst36(dst36),
        .dst37(dst37),
        .dst38(dst38),
        .dst39(dst39),
        .dst40(dst40),
        .dst41(dst41),
        .dst42(dst42),
        .dst43(dst43),
        .dst44(dst44),
        .dst45(dst45),
        .dst46(dst46),
        .dst47(dst47),
        .dst48(dst48),
        .dst49(dst49),
        .dst50(dst50));
    assign srcsum = ((src0[0])<<0) + ((src1[0] + src1[1])<<1) + ((src2[0] + src2[1] + src2[2])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15] + src18[16] + src18[17] + src18[18])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13] + src19[14] + src19[15] + src19[16] + src19[17] + src19[18] + src19[19])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6] + src20[7] + src20[8] + src20[9] + src20[10] + src20[11] + src20[12] + src20[13] + src20[14] + src20[15] + src20[16] + src20[17] + src20[18] + src20[19] + src20[20])<<20) + ((src21[0] + src21[1] + src21[2] + src21[3] + src21[4] + src21[5] + src21[6] + src21[7] + src21[8] + src21[9] + src21[10] + src21[11] + src21[12] + src21[13] + src21[14] + src21[15] + src21[16] + src21[17] + src21[18] + src21[19] + src21[20] + src21[21])<<21) + ((src22[0] + src22[1] + src22[2] + src22[3] + src22[4] + src22[5] + src22[6] + src22[7] + src22[8] + src22[9] + src22[10] + src22[11] + src22[12] + src22[13] + src22[14] + src22[15] + src22[16] + src22[17] + src22[18] + src22[19] + src22[20] + src22[21] + src22[22])<<22) + ((src23[0] + src23[1] + src23[2] + src23[3] + src23[4] + src23[5] + src23[6] + src23[7] + src23[8] + src23[9] + src23[10] + src23[11] + src23[12] + src23[13] + src23[14] + src23[15] + src23[16] + src23[17] + src23[18] + src23[19] + src23[20] + src23[21] + src23[22] + src23[23])<<23) + ((src24[0] + src24[1] + src24[2] + src24[3] + src24[4] + src24[5] + src24[6] + src24[7] + src24[8] + src24[9] + src24[10] + src24[11] + src24[12] + src24[13] + src24[14] + src24[15] + src24[16] + src24[17] + src24[18] + src24[19] + src24[20] + src24[21] + src24[22] + src24[23] + src24[24])<<24) + ((src25[0] + src25[1] + src25[2] + src25[3] + src25[4] + src25[5] + src25[6] + src25[7] + src25[8] + src25[9] + src25[10] + src25[11] + src25[12] + src25[13] + src25[14] + src25[15] + src25[16] + src25[17] + src25[18] + src25[19] + src25[20] + src25[21] + src25[22] + src25[23])<<25) + ((src26[0] + src26[1] + src26[2] + src26[3] + src26[4] + src26[5] + src26[6] + src26[7] + src26[8] + src26[9] + src26[10] + src26[11] + src26[12] + src26[13] + src26[14] + src26[15] + src26[16] + src26[17] + src26[18] + src26[19] + src26[20] + src26[21] + src26[22])<<26) + ((src27[0] + src27[1] + src27[2] + src27[3] + src27[4] + src27[5] + src27[6] + src27[7] + src27[8] + src27[9] + src27[10] + src27[11] + src27[12] + src27[13] + src27[14] + src27[15] + src27[16] + src27[17] + src27[18] + src27[19] + src27[20] + src27[21])<<27) + ((src28[0] + src28[1] + src28[2] + src28[3] + src28[4] + src28[5] + src28[6] + src28[7] + src28[8] + src28[9] + src28[10] + src28[11] + src28[12] + src28[13] + src28[14] + src28[15] + src28[16] + src28[17] + src28[18] + src28[19] + src28[20])<<28) + ((src29[0] + src29[1] + src29[2] + src29[3] + src29[4] + src29[5] + src29[6] + src29[7] + src29[8] + src29[9] + src29[10] + src29[11] + src29[12] + src29[13] + src29[14] + src29[15] + src29[16] + src29[17] + src29[18] + src29[19])<<29) + ((src30[0] + src30[1] + src30[2] + src30[3] + src30[4] + src30[5] + src30[6] + src30[7] + src30[8] + src30[9] + src30[10] + src30[11] + src30[12] + src30[13] + src30[14] + src30[15] + src30[16] + src30[17] + src30[18])<<30) + ((src31[0] + src31[1] + src31[2] + src31[3] + src31[4] + src31[5] + src31[6] + src31[7] + src31[8] + src31[9] + src31[10] + src31[11] + src31[12] + src31[13] + src31[14] + src31[15] + src31[16] + src31[17])<<31) + ((src32[0] + src32[1] + src32[2] + src32[3] + src32[4] + src32[5] + src32[6] + src32[7] + src32[8] + src32[9] + src32[10] + src32[11] + src32[12] + src32[13] + src32[14] + src32[15] + src32[16])<<32) + ((src33[0] + src33[1] + src33[2] + src33[3] + src33[4] + src33[5] + src33[6] + src33[7] + src33[8] + src33[9] + src33[10] + src33[11] + src33[12] + src33[13] + src33[14] + src33[15])<<33) + ((src34[0] + src34[1] + src34[2] + src34[3] + src34[4] + src34[5] + src34[6] + src34[7] + src34[8] + src34[9] + src34[10] + src34[11] + src34[12] + src34[13] + src34[14])<<34) + ((src35[0] + src35[1] + src35[2] + src35[3] + src35[4] + src35[5] + src35[6] + src35[7] + src35[8] + src35[9] + src35[10] + src35[11] + src35[12] + src35[13])<<35) + ((src36[0] + src36[1] + src36[2] + src36[3] + src36[4] + src36[5] + src36[6] + src36[7] + src36[8] + src36[9] + src36[10] + src36[11] + src36[12])<<36) + ((src37[0] + src37[1] + src37[2] + src37[3] + src37[4] + src37[5] + src37[6] + src37[7] + src37[8] + src37[9] + src37[10] + src37[11])<<37) + ((src38[0] + src38[1] + src38[2] + src38[3] + src38[4] + src38[5] + src38[6] + src38[7] + src38[8] + src38[9] + src38[10])<<38) + ((src39[0] + src39[1] + src39[2] + src39[3] + src39[4] + src39[5] + src39[6] + src39[7] + src39[8] + src39[9])<<39) + ((src40[0] + src40[1] + src40[2] + src40[3] + src40[4] + src40[5] + src40[6] + src40[7] + src40[8])<<40) + ((src41[0] + src41[1] + src41[2] + src41[3] + src41[4] + src41[5] + src41[6] + src41[7])<<41) + ((src42[0] + src42[1] + src42[2] + src42[3] + src42[4] + src42[5] + src42[6])<<42) + ((src43[0] + src43[1] + src43[2] + src43[3] + src43[4] + src43[5])<<43) + ((src44[0] + src44[1] + src44[2] + src44[3] + src44[4])<<44) + ((src45[0] + src45[1] + src45[2] + src45[3])<<45) + ((src46[0] + src46[1] + src46[2])<<46) + ((src47[0] + src47[1])<<47) + ((src48[0])<<48);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25) + ((dst26[0])<<26) + ((dst27[0])<<27) + ((dst28[0])<<28) + ((dst29[0])<<29) + ((dst30[0])<<30) + ((dst31[0])<<31) + ((dst32[0])<<32) + ((dst33[0])<<33) + ((dst34[0])<<34) + ((dst35[0])<<35) + ((dst36[0])<<36) + ((dst37[0])<<37) + ((dst38[0])<<38) + ((dst39[0])<<39) + ((dst40[0])<<40) + ((dst41[0])<<41) + ((dst42[0])<<42) + ((dst43[0])<<43) + ((dst44[0])<<44) + ((dst45[0])<<45) + ((dst46[0])<<46) + ((dst47[0])<<47) + ((dst48[0])<<48) + ((dst49[0])<<49) + ((dst50[0])<<50);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h0;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h5390c1711ffda6c06038711f8750210d58d9695e8c32989499479924cda109878986fb36a2fcba65b8fb6a109656452dd8344df27a4ae940d2dd54ba74804c552439f11c5471ca4893ec324777e8;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h266df0d21c5284da2c4c6ec2b1c87830ee3a99667b1074457bfd4e350cc49d9200625f1f82a3a461094ae92901394507c5598bd69c76b3adfb919e1c331f2ab3acde770601eca87ea6c50a22bbe0;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h11043135d89aa1e17d5669f7ae2185c1922570a360c86b79d4369323c278691f8650bf0cf2060723ab8598d7c9d48f41de738b748ac7c9d8cd72ebe2f60c277ed307c5cea5b34bb678e6144770f93;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h15180c5baf2ec40686990fa8a895854e5263fdc039cc7b21c1ba99922a6b320315d980aaeb209256a8afb4d0c26d290989769cec882d13cf8f4e5dbed3f30517d0f86f6d755bb00c3cea936463319;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10baa263ec8a67c5b1514631353ea74de50d09d72f27de4012a99a42182213284e038074f92b31907c952facd54159b1221941f929263f9103c893de6e6bbee757116af4c78a263000230f192a01d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h2889801dbfcaf3a1bcf899a43d8c3b06d4ed00fd3a83fcfce9f65a4b8d37c15794c425b5e83e36ca4ba9a14cd3c60f6f0b313d481a25ed097138bd536b5d33925bef7b42679e2344c8b150e1c231;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he8903e97f5a0d65936af4c9e8c0982744da866d5f1f71c9de96a6e4c88415df4cc543234eb6d8c04fddb0bae4d5c2da09b3c510d4def5334416ef40d1de1a0ea26a7fc2eefe86929d31ca5199840;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1bfd2ac491626748fbce69025678884f0412aa5731b7abe783e1a9d9bd51ed77f894725339b4bba0b1ede015667ff3b3b1298fcb73404b3619722326ea374ec23966a52712dc97eda95d47fe91f72;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h6a50129ceb0a42a60c99ed2c5b8e87a1d00f79f5cd97ef5f021de8c82e862984990443d8ed0c27ac8926e9c32f08d1e4f0649826ebf81f0a5aa501bce69d04925d987f3ff2aa525c3258b6c03f37;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h33a100f6d20cd98231a62cf51bd015d1f12cd24ed72f63dd9eba51abacc42f5b5a6b71e02eb941bee0c747d5ce3b624e90807abb58dae881dd5f2af89f0cb4354e61c60369fdcdac9d86ff9b0845;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc00a77bca04bd76edb019db8b4e1d99c7f405f96952af03558fb34b1c2cb171851f1264de7dc32c32dbbe0dc671b962ffd672d21358965625776a3a3f3a7e73eb1005afd221e7d9303dbcaea87ad;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha983a70dff6a6955f181bbe30208a3da9345001cdffa67b108e66fa5d28758127b5c6ce3e896ca9450b2d002a062d94bbd75cc96ca5494de7bafbf19d05bf039d74b33607afcdf554a07e1d95e7b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb33174b7048e74937f55ab4b4811b54ace435ff9a393060c7d2ad6eee3f62440314bf02f8d737a9ab741d96dd479f5db0a696a06279444abc4ac64fb305c5070886d97caec13db5dcb8272e5effb;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a90c2217c0e64aa2e35a294b7230aa0e82de88379fa7da0f7b23df4f4e8284409aba7e12a7c2541ced731cac7fefeae427daa2a2161de65b08160342f7fdc65a2f2c1611ae7efd672faacb42fa82;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'haa34ca84dae78b50b68a5ac897855213389ba710749bd54694b54c855ee1e6173081fddf54c94bbbe7cc152f538aef74c29532a8bcba93848b5937e012a1396b8eae90ddc79dcc69fa4578946a61;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1480ed2897e75e8c5b6afe6d5281005337f185097d5d3896da29b0a7e308c3dfa7f9a0ff73ab5dbc8d557d348e94651dec665ebc95a92f508ab7e5a9b3c7003afebe9b6cfe4d1a8bcc0a82951bbf7;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf9257e8787a88e9f79aaf5fd0d03693c9d26de2ae928cb986caf05d2056f656d8c4de954006e159b689dc8b9ebb7ddd51fd6477a7f65f57ce939ab9b0396d2e0fe2307cd75bef272297a64bac8c1;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd4c13021f3bb4cbbcd57cb31194fe443f618e13d6721150d265c62ff11da3ce0d2e869a2f6054a09b77edb7aa3d0f2d89a0587b39f24da46f825aebf0f2eed3b3cce4ddb5186b72e3ae321cdeb6e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1885183a5de88b1f1eea39f76919ab96ab019fdcca92df5d56d9b049c6178219aff674c3a566eeece04982020a1c2a08fd43d30f405f5746a3cd29af1fbe6d384066cbe42d7fdc56afe11e44eda6d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf4839b29846799f407adca992d81b1b78e5abab4f6657a69f04f1b210dc224ce09a897b51732e0e5720bef17838648643ad14d029ee829df0cb0e74bf88db2f334a6fc6a147e48130697be21e8ea;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb775658b19759a3b95aaef2939cfa50136b554600307cb5e461ccdf4b9c2432571f8ed69d09a835648db2d53c06f1ff6730b8c0f4f9a1c43639169759815ac2dbc65a879ec5433d216d3e332b6b2;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h92b625438294cf1ac74f742f132bddcc978a44450eab3cccb786c67d8a2e6070e4411c5ebdda3e4740c0222876beee5d3f98aa018d4f80a195478104a2c1333566ba141ba52909fee16672eca719;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1503a918f0d03a4e96200c9770380b8d0fe549549be3a10e406014fc5833530cd540c9e5e55eafde98f03000f9f82947a18a3ce390d4996ca2126238644c9defaa23c36e1f0b9bb0a045ad58955af;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h188558708c14f70f2adaa7d98f8ebc0b916537fdd65570754fcdc4b979763be59e79fa4df0da088ec09f7d3d8962dc7171b2fc3b65834e89157a54fb338d679f9de2654b2f118db0d28a594b83463;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h4e2c0a6fe4eaa963e1f0daac0590297eea951421fe411f9dd68ff396b5fa4ce99839465ad6c9332e676cd35ebfd0815014adebdc8b7bd2218b06dfb091bdeaa2715a7b7b1ef30a1500ddf73339b8;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h470ed2ae81807fb7ecdc3916dfffbef9a20f0e3b53cc1f26b24d657c851df17ee45ab9acbc2d92032739a4da09a54a6f0e0a3f330326e9bddcbc34cdca454f66f1be2e1ffba6a9331b9553dec659;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h11113f68f25b90ea24ca055a00b7d25029b4ad68b40136307f493580ec0bdc9747fbaecd99525d3512d312b375886740ad9d23c084662016d24ba607f3ed6e04699e7e4bccf0b40dd448d71187a19;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb4bf4b621f0976e87e0f17a21dcd7a4afa6c82c612fae91a1276217dd2413ae1916fa551cc602d760048243134b238b51d6a25848d84351d46a1e70e1810f1786014c4d6071714bc73ce483049a4;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb22181b7456810bdc80e5a38648620eb1caaeed0671d2ef788b86d975623c7f316663f2d282cafeb5ffd92c9ec9a0f303e5c37d1f014942ca31336ce692ae935c788a7fefe228b83525709a6d700;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h845083d33934dff51bd6eb2f810d4e9a5c5fd959ee6043294bd2ea29753b578767eaac8a93f15f5119bdb77fa412845886989efc0d3bf9906c149ee4cba802f34340383cd7378bfe456f5bc835d2;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ef6cd953742d8dc9a1046c72e8e061db5d893a8ffc171f35d29c75a994fb6d3c4cfa478cdba659e119ad3a59326c9ba819f557a183f71a45032c0971b312eb1fb7e97aba8cd3b54e3693f0c8178f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h2915997e1137732f7f8ff4146f9a19bab78ef154d38213dac86b559716a54461824877652309640f54341ad86a11dbb2b20a49e92a16d760511c4fb96ffcc7b7aeb27e886240741ddc8e8120a4ee;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1026291d9086d5e80f4c8c4f028dbab9e4983fe29092f7ff04353fc81a4637682f605742ea0c4595625755c0462a87214d331b3fee6ede5df5409dc730b9208554e5482144afcdecf89e55ff72d72;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha0dab83e75967ad2fa03f37ad09de43aa08fa84c5c59854b877989bcd986eb953a15d96c848a6c27ece5ea671ae3c188862dd35e281f6645c0757a4b52fa348bef1821461d5c7ec916c168db2494;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d1da823a5ad60958c23462636a5f8f05266b49cfe461cd0ba849de676cf6183a339ab4f6c96a35865aee34063098ad4d8abfa714436887f9be7ec817e67bce6ad9a5a33f42888dcc23536cef24cb;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10c6639dd7cf9182a813dbdf45bbb5f3a4b392769d00d1d66c52212c6f752a9cde19e02bed7af21f5b4f5d3ff996cbbf230742d207f51113e12a2625a3c1fb2d82b6cd9d0d844649bb40df196f0c6;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b6549aeba5146e1a62d7435767db7ee10fccbbb5b6b00f244fb8cb32ba125e7992295283b437c964dfc3652190bbc215cde88e7dcf07cb8aeab7aa358876273a43fd2f39afa5a3becd09baf41118;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h9cd93774189d3e03931d7dac546aed0b28acb586ac238742cef5b3f76fd1143db2eaed588a4a632451c9650786c70845d5fec8620145d5e5759d744e3430c23ba322e703d0f8d95b81f41aea13f1;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1112899bfce08283674c4b610ab3eb05536b8f82babe128f47093cebae6c5598efa95f3c60e5ba672a11b57f8f7be34a085daf08436f32bbf378c9493e4a831a853393eedc6216c5df05a2b173689;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf593ba7e9353263cdd510e9e92e076696fe6566cce841b257c1ee17810e3706d5192c49a500eda6cf39b1b597fdf4141b47216fa34f17152826af829c8628700ec659afb580dfdc1a1a14776e00b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h14085cb7293a9a2455ecdfd07fa415a6dc829687672e23213cd1645702847551cce6b7ff958d07afb056a4319838e7eec9a90803ad65a7ebee5f54327fd0cf2e7a473709cb1f08711f07dc1102c7a;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hfdb85756e528ad7b9812dbb31d37da6d79c31b72009535c62ccbcfe43585224abbe391fc1572c85451ecc2ce60b6eb8612521a04ab85d5cdac7d888a9e5b78b5389373b4b9cac00f68456994733;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h13bfc88e589195062ed02b1c25fdd970d5db0960758058a21217dbe0153014f68be6251c48f2309208b7a953f7ecc52fa0b1a8f101d0235e53ddf427fc2487e12946b71c5e1a6265b2d743a9d015f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1849658b72c4c4beb76e3c77bd1f5eb0d0925af754598f324cdd7cbf208250e275d357936926b6a4d47efe5793da6b2389e86d75fd9c60c2d937098f10f03668492ad5930f288f9303940a39d4e2f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hda9d788ebd096a667ce3bc191be16eeb34201c0fa54d6b2affc6a6ca62d028126ba2b578ae9934b80d05506e46bb7380ab251f3d35229d2105cac90ec0ce0ef231f644b956d1be00a54dae795ef0;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1fadb4f47516fd494219b40b8386b237fc8f5f8ad41945e73d77d708bba821dcd2aeb0b06275aae98b185a26784d85253cb9d6336f35010061d2ab836c46779ec0e46cd42d7bb9883702fe1d24ed8;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hab61fe00129ea958087ad9d74d3d0809f1066777f9fba6834b5b42e12a655e4dd7671b70ae3e0696b0acffbabc1fda3b442697d823924b880456300e0e1dea206465e2efb4bdb8b26f7ab82c8405;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16def7ab1c03d448174ab839c6a302b3d24b8cbaeda217346ec58ef78f78937abeb8830426b50b0f56b860ddbd831680c64a3a0957c28f19323c4c7827109c21ee3f3d2c31f9b5e8dc8db9f83d542;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d6144af5b9b837cba3ff773f23bdc895127452b3ee45124496a188ed791b0cee1597ef131e72ebcf5b0146a115c62188016ab63a0542cab71ec2e42a06a5c9db306665bc5b7841972a799e38b6c6;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h15ffd49958d6b89ff4e561808397a6c20f6a8d3ae15fafd77b8e4bc6294ead86001cc12e853f26df2139675840e9f04fbff98224fb0583ebdfa2db21f7ab9962d3b28a270a2e12fddf34f792a0ff6;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h14834615d92c4a2c61732bdad4e211264f5f4098a7d8fa0334d07c2a49d056368e2b6f4c0c888f26ade496a22b83c4f620a71e2cff2563c6746beee2e4274f6bab4907637d83b96883d99c203d9d5;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h6ed9d520caa0cef4b19f80e13c74c7d5b33ad604edaa0a46431eb7b2515fe93cb794189ff13c00c9656b24cb32ed42d24d05d7712d32e124c9737b536538fbb02f4c096583b1b44658732405c867;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1969e66d78fd08db0485a843ded5098b1aea329f00a6ac56f7cb24106504ca3adc4f8f1c09c8b30311b8878adefdf83274b905ec811215bde40f1b3e7b0805959d6c664cb82c1ca632edb54c0da33;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h17a57a8498c0320a79607af697619b295860d1bea22085711944290f8fc9a32cb012b1237500f726430b7a4e7af2b1ed538aaccce3066c7d2d1f9e4de2570e6e45b9a86ad94aef720459cd6422f6b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e09b95efb7c1a8ce9db09c49877e6483da728f886111c72928d35c457efdb379a718cedd495e0380731eb69af1cb0b67c71e1e7fe493374d3488ef59a93a1406e11e6b28c83a02574d9e336578d7;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he314191c6f09e6a9b6c9b170c00d04efdaf9791a8acdd227fcca925e414e5add561d11f0c8334f9528aeb95fd784dfa17a60e96670375e73a7670e6e1c31fb116c025c7e299988e74348f9b3d8a;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1169e80038721435da4701cf523b7578d923f785479fbbec11d0231476db262b91e96f235bcf712f9b0d1fd211129a1e3c268105cfb994e970d88e17123bb42bf2167702c7b9ec41051101597cbcd;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb1f732fc019d7937369479fca79cca6e620db1e79e5d83fd21387e4533fb2fa9484e0fe1a1c3d99e996c67c5dd406470f198ce06f930c2a63a2862a6e639f263706daeb35c4db5d4cc75226c86c9;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h19b4518ba80da8293f8c54344553c81674a84f4290a783a806cb78bf765caa807b64f7b0c25c3ff03b9269104986ea70f3eb6d922e0e595d3abdae7ce2a8a6daa380eca4c6975ec5c7eacca894b20;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf5b03620995e02ca5f80dba57a1a508548be37efb9b0e63d4ff21b9ec842fa786b5ce1797646c1b4c3665a75714154fdf08ba05e4482b3f26c73993281d6892ab7c9a980a68a3be70c5383942d46;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h8386dd08cdfd5fc5187a9d4aba93bf813dce170d7f8e378f1fb413284430bf74477ba3054177ec77e89397ff44d63d7d9b28b2631e4e7a4f2ea93d3ed3e746101a6a1d56ec6cb46a6c2ecc7995cd;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1fc9a568571780a3a1872ef3a58840ebf10fbf55c5f9853cbe9794627a690a72239e207c58f9f0d8b753a5af8bd3d18bf239f66687ff827d18d7888821971352ea6284b30b22b8f511a223a702cb8;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h99501d9853eed3ca20ec264cfb9a8ec26c0379d1c7d63ae3d3a6a68be32071bffc2d839375d508b526be97e884fed7592f35ce2bdfd9c3131bbbb38885ce1ad234a966610094f6d36e27b56586f8;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h116d7e607f218843655fed5fb29a5290142711203d31b075832166f7e25a3d6d358a1bea3e8302373b174db3aa35a81100028a3e961989e0d4a5e1778ed00c8391e88f447b1d2fc49341cee18be5d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h618fdfd7045bf84a1eb5a99cf89ae40780803e81c381e2a1238d1735efeb018ca6b76d4de0bb251b3966b1369100a73fed7b6657051e3cc153bb4279508c54d156c360fb3de036b98829cb2ce2a3;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h4bb862bd0128705145dfcce670e6b59ba9dffdbb894f038818263844f25295276256ca41a8b390f8ea61d6eadb79fa181b0b77926bc42b2c4f9fd519273379914a3302d36c10fe4a5d7f6ab4fdb1;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d37d4e6cde949f0176ca119e7486371a9eedb00fb995d3915779f6c472c93347907cf5be31ce1e6755a455f0186704b17f46c302f93e2a985d2e2fba01706ef536eb880eae86f4db26f08c4e124b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e98784729500907a602c7f7a39992b8511c64642ac9dd69a3ff9a7552b6ccfbcb70e1c831e44da0fa131c5903ec76737b24f7423ba86d1767e5a2fb8f837e51bd40539f9374527cc39c0a7cd748c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h9e0557caaf44e000e90a78cf9c99c942d0d39f1c5f457f8aba013c2729ba900dff9f085f2ab0c27335386d564ae412ef66114a4b2070e3f0af481b2cdc174c0b923b3953e070e1c665fb78ce842b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hdaf0a9040923e7e65f0afe019f7202188d956ad6a18bd5c738c12c8cda8f8674f1f8d51ba726178abee4543ce269f61572322a8fabb61c15487b86373f8161586268184b40f263b79aa9c96fec82;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d01ff05741cec68926f8387e490355af54f0cca0c18d24dad9a00ebb51f874bca542fa24d3e321d856752ee0ff7cd6ca975c1ef4e00c823be53f93be5b5957d135f50c43d7b1f343e28630664ddf;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16b82a945f59b1ce3e87acc455f1e954057bfe9786c9603f2a1fbdf89de77330f2789746501d4377254cf3e6d7cd0d692d8027a0eec59d401a393b78f5c1ea8d412306a46f45e1ba81bc91ebca41b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1777b1d92f55203f1a766557233cfb57cdb233660493fc7c6e2e5b316f8a7d4ff703cfb640ce419c20f1bac2d74c2160112ea761a47d498d095aba23c1b2480e89c09b7fb706fc2da28c9d54218e3;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a35c0c5c681f63513972a0ae5363f154477e064d7d6665f42a31db2dcad4f89695d9161bbc216a0ed9d51081ef7b9f2a95e5f5cb14b5d7e986e95288c5f77c108caa5a9f5a607703768e50faf64d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h917d5d1df3bfbf8b1017067e125ca48e391ed3c8faaf381e62e3b13c70891ce33df5f185c353717893fc909bb5d511dc13719516272494d5cea1f3d68c4167ba612f75371710d00fb333f1aa2100;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16e61313a0b45912a4f00a9492ab462e39b6745d45013727f831f323c8ca8c8fb4e6c6342af858b6e026563ecb736c9e47f559acad209cc688f49f5496d6a13a8a142e5fb03604dca2a30635f3050;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f31f35d061bc33c8592c2f3d7617d055dd2e4f92b4614faa4862fb5e96f82f520985ed78f1209ec81ee85afbb4a4f797afad523a94565ae5d66b6eab9890f359cf8d616b5649bef0fa1b85b72a07;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1beff63b800ad2074224ed842a9914ede2928f7bd95ef75ef720359f4fc76924f2cf2935c2765a14b9ee5c1eed5b33f153bffeaac27bd015164c2433eba7fcbd67e69005df375892ab1dc57bde6dd;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h419783109e9066cefc42e08e3c648d86d84316385b8909254f6f16da6ca8cb317cb2e54fabef120d11900a46d3b68b9a5e70445af6847ac51d9f9d8a99edf141e0140d3e1e54e0ff61a97c391be8;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1699886bd19d883e205f11b1fc0fc6af0d7cf88b5469889fd533c09a85dbcbab335a872bed82b91bc8a12fc318aa53a122756e78a8b616cf59d464579dcd1efc674f516e1b8038a0cfccb49c29c5b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10beb9366dd3892eae0e3aba95a68b67411a4b179d97ba160dbaa1f8663d2cb08356867231ce138886f16a531da83fa282159d5e50b73d9db8b9efbe8e4c1097c8b1cc2a967ba5a5ffa770ff2b2c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc878ab1a9322e95d123472116ec03fbf3c63c6cf5776c06182278516a1ea0660610228373e6cc00ae89c411afd6853e6c2c37802275ee529028d97c7c786cd9b96cfa9e38d95a43fe0c9cd33e907;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he81f9258440a3288a85c1c61bf16a20d3f121a2c05de76359893182f85b7214705826bed9cee6a74104d72fbbc2ef725de4aeaa3d74168b37a10261a5d10a580486a33b96734db29293b4af0a80c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h4c90caa5cac53964244d587fa8b15c8062283b6f3b29219948a9f8deb1fc764aa49da78af7c576402063e3fcb19d3af706325f654b2ab0005a1a3e40ee4aa9353a313fa52fea7584a4839b0bf86f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hdcfb47e4756eb258f1a504f7a3e0d4a1a6f8a71c4c8d7624577472d87e9a721f7cb2636ee83d17d540c067ccd4de79fc73c3b1c770edca6ffd9d142f86ee1ea906c440ce3427dcc8700caa9e01e4;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h22cf5dc20e291e3de5d789795536a6fcf2ec5c7b3a47e9d0bbd22fe1568b377e3fbc4da1f294b8eb35dbce9854b02808daebad9c91d7116ce964aa0892d80101ab9898893adb71a999f394ea3534;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h5558ea2daa067763ae9e1ca6d0c555efe7b61f3c5dd340294f04c258f149234e7e9d0eab3949d26f7f4faacda6f67b45b1c08cd76832cc32c0fc8285237cd6322df8bcbce69c2623f35ea5c7f31d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h8d0474b4e18d06de7ec2baea34fd0821b27738da7012b010287eb4b50eedf656239782f46cf272b0ab303f517b0d9e5d48176deb6fc08147d6b051fa272f79c7603d1a4d2cbf1fa0b1959111883d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c0a17a148aa0ba12f34df686400497f1a3dd45cf45dc3ef757bd5537756c97d31f6182e661fcd3fc62da52acefb1aa2a4d70b0f3cd7852e88479a44101c8f5d1bd728ebae93e2b78d4be28fbc5f9;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h773ae2633280e1657adf19ae3c1c8623b14537795f3a5e680436c5ac2996d1e1787d8c69d2e8cbd406b3aa6e70a8016a494752a867845f988a0c45c3311a9aae2f4ad5bba6553c6e9b129df81575;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he4ae70d2b11cdb0113585898cb2875079ae891a72307976c2aa08c26bc3e6d69cd03e12b748b4cf56fc38101a3797bf4ae6d7f2c7f3120192542d1f3d331787e84fbef521f53355fc636c06a283b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hba512eb2852d81f9214a2748aed9e978986c0191a5ae8e57f5f865467b543ae52fd0b7a133842d777ec57b88a0760171e8da7e2144c2fefecb2f0f3a3311a9481098778ff30a5923705273b7d59;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1fe3d47cdf7c59b87bffb4f6be0c1023a547b0c1e1e5bfb6ec4d6336499405482a1f56bf21917268a3589439df161a1f1432a0c5ca970ed279e2016c12e7fc9ec9f32147f94e0beedc35cc9020240;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf8cecc9564c52e24b050d4b1c410e7092c0d6196eb9eb8c46a8ebeb718a60bf78f4eefe7ff87c78d7d8b3913403c4c60bd3e653694675600e67e638d80a7efb907f47ae0fa4873afc1f39059ea3c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hae431a823fbfc26bf39696e7695debf5817dc5001175c536f37ee699b8f271f8d8932d98bd6b2fc021e4f1e13a4b62c95dd488fbe7e9210c617ed75b55d06388f9ad3d9f759850adf733777be6e5;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc560dead31d966c03ed53886e69016fa152f31afbdaa3bdc713c694a46085896f237c8038d0992e10dac5a010fdee5c470e25d5458658fd9c49f6a060d4ae25d877fb0952c743868e49bc78c5a5c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e0bcfc083210a0f6b0da3929b209274e26f22a95d1b27dc0dc13cf042f5bdf6f0061bbbb80626cc2382d06ea64ccf0289ef656bbe8b88d684f1f312c2f2208617b07ddb7d12a77b93f72490f6480;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h22ef7b1d9d2c85725ec809b62fe7086c7a065d07df024b40d46d540ab89f1713dce7f80186fdc14cb130589ee5a84e4ea5051bd80b64dda5b030f639919dd1fdf8088daf2b80b2dd74e7cb961901;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1049f7c8ce602d9845c4af4f90610b14298a72f02496d21255b0edfab38f6d4a3088b24b4394225b8edce31fb58dc0ab3503e8f891fc6b132e5dbe9c2d723921e1c3b08b6f9f00a4c6216d6a95515;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h18cf989e4a14dffcd88a14e5d3e93d700d19f63041cb7c05e2735ca5831f529f613ad7792c9c7d45695abce392a249741377aae62ccf23ede485b23a84672195c807aac673c668200a8189fcbf0ca;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h17a7a37eb3d868ff8f689e3dbbb59ead108d9a5850255673e4521d17def02071536f131ceadb2f9ea949e0239137610b14bfcc9491aa9a31cf4a7ae2a69a13b84afdadd03dd0669e59ba1612837e7;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h3c9c4f337fbabeb1387c946a520f6c68885df358ee7b792f945a68cb46b90e624499b711e8692cb93e0949ea8dda48799335085f4268ae76fdb6cc369f1615787bd05703c8cdc6bf5cf4e3ff7256;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h117ff6197e2c727b2211f6a1d3e408ea69fb3bae70bce599fc9086169d7d55f513b0cdb8bdd4182f938993b0ccb6c9ba14eb41a5891b2869e272f7fb5a9e6af8c84d0e97fecd07818ee0b7d60a585;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb29229e40530297e65a274e13d58d0f3d58d8f2ff7e039e7d1b942c2d0c34f94c5c2e81f3bb9b75b694a94cb042eb0c206fb9e83adf7990727490a6be568c43aeddfd2ffe46c7fa7a8e6cc3e301c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb8ed6ee1f22d2bf7841214009ade8d6be47ce3af81fc6d76d461a37744030232d7fa1a6ec865a6b6b79b5971787511f742710b127cd8e4983836b1f5af40cb89d8beb3ce9103db87be3da188abc4;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h269f27ebd48bb0bbba82f2e5aeead267ec01b2082987ff5884d11c321c6daab9a603bdfb3f5655df8be5a6030a748359dc870803713d116fa38db540ce5a7d18b82dfbfccdffc2004bff5a663b3;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha73334bcf960311c24cff9f2a9d2e36d9252390f5734ad8c5917dd92243ebd619cfab7fccd0523408655e9648279ca737d3373588a6ee047f3c063ecc1f1c709b368154edf0d42cb96c2a901d548;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb3e365f58b39d5883b761a2908002ad531446ed9d6702bd28ef7b15c3d0dfc83092dedbac10bef02f50b0f9099971293517a891452b5bd5b10bdd11e16d5bdc9e5451eb3589a696f2d7f8981ac19;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1fa0ac50db84473b57f8f161ef6307a2ea396bc16b8538af7581746e990cba4688f80e8cfe8cb646581d5d85778757bc554e115a1b944078996a6297b1c71c221bc33ea637c8e25c7139328753eba;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h924b03ca70c9a006634b2632b5a48ac366d5b6bde3aeacd1e73773e9fc043826e618e2d7a6103bc16a472c0b19e48cfcadb173cd4c6aef864beb04d53bf149da89d928fb91fad2d564bcf852417a;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h19932d3b555af95c4f84cea74ba66fbfc867bd61eeaf4489f68e4aed0d580794ca697925fe8c396390e3deaad2676750178995a3341a3a746a81342162fb2567e4e3175f4cd8ee154c12aeb9dedb2;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h20c0674da62c4e6c3576ab562c730610fa078e85cbd2aa70fb8fec7f2a055d513bb0e82bfe2cb1f1f3ee3006dd03ba63c9f4949656c9884b58ad7914c434992d423f33c5d169fad2ec26216c0b7e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hfe266de56ef2d688000049c99cbe201b14947b8ae7ae7a338a7ba761362f60842e77a745ebae550385e89ee497fa3e4d0a6c01de4787118990b049ee5a1138ed3257e0b95615a5868773d2df10d0;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb6c9187a298da7cc61b15f7a82344f9aee598cc414a647617930f2c71223fd7e0141a2bfbc756668906ed00a8490823f41b91e01bf2e7b929b950e3a6fab53fa936f68583392a746ac3e2573db01;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc7e9e50971d49a2254a5be07043b42167d69340cb90a26e6d260195fb5f3535a544915fdf3b624af214d8c21d83eb30809dce751d6aee8375302a18873f793ececace0461d8ceb54e9c359ce5dd4;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h15bad38190834f9fc267546866e5458987c5be3dd08826d0fb57215df868b63dda94183151fba1ca2b675eb658ef54215767bc8928b0bf95b405ef406fc48e13fae5e7367749057d053b20916f705;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf93322f6ac4d5f8aca26b87328ec0798c8d47c97b77b1468d5723377e5d098808a1fb235b134eee7abfe8240d474872506e2b130029d2afc7adb384c52fe80f91da67213d04666c88a220cd91ee1;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1963b4f10c843cbdd244bb13dac1959574accc98fd693d82d6be7fc03902f4719b71009667c6e9afb503eb2abdab1597217c9e2bf6c66eb3309019258f22ace52fa078c5a2709745fdea88b1c420c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1261f14168d24887f415c0e33803117c3c902dd776972100df460791218c72a9d705e32ea5901db57b70c360b0ffd63d33cb96397b9c915141a056ad83270261ffbf7c7954738409e3af7fc40ddfc;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b0456bc47776808dffb06bfee8791a357b0dcc6a7b3e944e4fb06b38c846f4fa102a1aca310ccb2a2f391a8752040735fc9ab7e7b42e1c800ce566046a7be9e8a079b6faeac6d804fca8b4ced63e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h14a7b73fc4b03fe31476c2182dcd1f9892a58daf5491b055748fd551ce70be0a3bf29046e32865997cc349b279cf40f4a6f92f185ebc0af8dfcd17f0ca2bf5bbf56c5455018f96bdbbfc3c13c3764;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h14a55644abe5b72178991f8b253d1bc383017d151cf7ea475be8eb37adf50ac6f10af9a47e8f28d6954d9be296e08a4a6ec8858cadeb67cd66b7126d9e6a34668cfae72d01b91e2d0f7935bd87b22;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1032630dcccf0f2474ae96b01b7b3a728fe2e5accfaf5a58ce90d962e872236a135e550e8f00cbb258259c8c4d0a00db1ceebb2be4786b9234d8e7d8c77611e058b5535d7ca3b30fa9da64d738ce1;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e7d75e526883f0c391874eff273b51101306d6389b5d70da49384bd9f79cf8b8cc46c2c4ab7348cc23ad5db46e43ceaeedea46f248c2fe0c2c7f6ec5fe32368d25eda0e54748e319d46dea0adcf1;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h89851f40ce00bcdf575b1ed236e2c2f9f43439bc2b0171705ed645ad1346d3fe78114be2cd917aabadbe33f79b5d4ef81595b740541fece5d69c101199241470a9c73798389e54fe2a41f8c4d9d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d7f2fc470306f996221e1b3a612a665132ec3fccd5945a7cefb1fb21e8d04bed5ba3fbe73e5eddaff9da36a293ea37928ccfa94a5ecf193daa38046a2056bfbd3fefc8a1e4e4e9b921430dfa5d7c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h172bcc1969006e82c1e76f4d09cf8b60ec234d4f1c342be23663ef67d92a64a7f66803627a2b271a2f7bfb4b6e7bd3bf58daaed93e443045b2498985f4a41e0a639c7fb6382249e7019fabd9fd06b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb764cb0b16dd4ddb2c8d70d8fa9b32b93a20a38c75ebcc4aa1f7382301b6ba0bc30a68416f61e48174b577a38fcc551b1fef00877c65853c912f9e04c2138f39b608dc31a43596b1a2fd9e1d920e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h8798619044af41e5945900a0cc7390dfd5cb52eb10d85f9f1e0b9e9acbba582f6f8d0fd407d010969cffd448cdb95951233a68446c1e3c0e8a6027ad9ee05b508a9ae8b5346e0fc5cdb5e717db10;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h17d71f295339d45ff9e5bb35fb83453332d6dce91963ad6793b35128eeebcfbec980ae1d83e2495c49c614fe90b2aed17ea00b853d1f42c9451c799ec4da887272ef37f6a07279b72f7685a5f7379;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h9a9b1a5b1b402d72d2f3631dea87077b077d8773690a047bd59a1ae16e6920ac2a8dd92b54bd83475d07a9616ed00c752d72250b83d06fb700354bfb77d39ccc60720319a51e66ad045380f20dbb;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b6f9027edd4586245b9cfef372ffbf3732c795b08a1e25214ea22419356285412672ce09b06e382977259d1864e688e96fd0ac41d487316cc800f905a93b38c5aae278439c708e73da2101640062;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha03974976b135e334037f16fb139fc29c42033be4df43e5acacd85b6e5eb0deafdc73b2031e037d79a2015d241d96f97099a906ceff54a7aed30b43e463e886f1abc861dffe39b0160f15e029275;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h14fc815fdc48a2e2ac045d07d1558316e8d1a8c06c1de9e503d781f9da18ef5962e802f5491e491299da9a213f15587220d97c390e322452928f35035ddc3b12e648192c808ae7e0b464785746960;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a7b2b8a290483b6d3e2ee473c86c1a233f7400daeec99b2dde987b2f200c1eb18b2904dea7a9037818775710295ed41ab855ec3cd4f3bcb5538e5b8b2f92d45acb8698e65d4efc0e3f56dcefa73;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1595913aa6ae5c710c722f9f038f45590a76cdef40756e41b58904e01045aee905ff07c25c7ddff4007d32bfe6f75a21c9803579460dae11ee97adcd078b3c7c3af8401fdd4386de9c182e278de74;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d39e824be00b2114ec0af69e3d3f8e8f391795aac5e634df587272e82aa97ce42802e1d9eeef589ec9934894feb2df67d62a46d8e7dd88c2936850488dbcd22e6b611b689557bb4fc05e7894cf14;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h744d2f751026092a2f59ee3fa0e123a6d035ca1304b4c92cc5c785d6a961075edbc71c80252d43d2a52459820ab3baee809fd5ee4d394b9f31ec7069c76ff209026aa538a373ec10309c24093c9d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h70564f5abe0c73f41f40b9df4a5818e5785d2c7d8f7881ecbe2a6627444776ee83ff5c136d2f6466e9250fce64b209839645bb828c09e77b5b6bb81f23a0c816c0bb4e7a65e225dbe2a726f78912;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h267b5cde43a47b8d3a3f251914b00cc98b8cda4a5a2566deb7eae4c045cf2483b3360fa0d40b989e62a549e92b1c45d5f571206632c50912755a10b1cbba0436aa0dfece8319e4a80ec4056e3ed3;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1fb0e7d2fb5777223b87414c39c76ceb6147a32a134dcca7c4bcf3dc21799634cb5a0d7ba2fb58b1ede2146eddc72d6346d5f1ed1003aaf5a7c82924a11ee990b175ef7a010c10e526e53ad3789;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d617602ede768b053c9e634ec9f6144e03c3663739d2c6a6734d6048bfe6475983b21b12df1269bf218cac32f745f4bf37973acedb32c50b3c759aaa43a95a2360fe5f2d38d77eb8dea3adb7cdd4;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h143619dd51fa8705b068e2adca27fa99a5b8007b4d64622fe50cdeb53bfb68f46215a1e3cefb6815dd2fc915f26b5160f1648992b4a8917f3660beef6719ad3e60d92d887f3dc08c43d5d0c8918d7;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1728ef392fd9e09104aab2db5ad7013253dd110d55bcefe08cc2c831208e70b5ea8d94f71b3fbda0c2cc2e6a4ccae87f8ea2193f0ae350902aef00c652db13f84e55fa8eebbd984b0420fca755603;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h153e147f069d5d608dd8cb3c909c9b756b49f88a0179c98abd4a60cb07323cb2f238d5ba44d909a600b308bd84594684b6ce445d150a7986f2cdef61e154eb3f17ce5bed9aa8020c644d7fee8bb91;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h11e1b9fb318546376491b0d32f86f2bc62dfb96014820499ec03e2cd08d6eb0b4bc7377a8b9c895bca4855b63e1800177f9040e68b120daf8d6fd4f7be2d1ae023046503633fa2ec6012acc13b566;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hae0ce4a10d1dc61ee73f2737f133fb007b65016ec519717e7623f57477a80702e93145675a569da4710d8f63b8191bd9fe42acf8ac9d96d1028275edcb5b888368d5ef69b86648875904a7517041;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h131b2019f894f0a33052a6ed02e6b07a28fdafec82b529e4c9fad635cc0b74a99eb3c5ca26a62745a8801ea62ad783b597f52b96db5b5b293f3589b794684b8d3f4acccc79878987dc8f534fdf2ff;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hcf16ac6406e2ad5b9bb27c17a2e436ae768a9dcd1e722e908e1127539bd92b0ef4580a67818dab752649b0e0c24455f869153f5974fe4384f5e72c164f4b34c2c3af058ac7b36259f7ed9dbb7dc0;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h171f7a859b0f80fa7c7616780e29e13c5cfcb849aba4ba8f314e4c84bcfda8e6560d03ecac6e35df04bb4249d6fd14f24e230c7a576b148b639fe187a346d57fe61208db3ad568881bdfc9032f68d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h6cc2dcc8a413fe086115d0c290870539b92c54c1c2af050c36f8f791024a9d03c72f11718f61b434099539a75063e2502676b1ac0178431f70cd8fa551a43dc5f5a6ef5208c45ba921e2fd592d96;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h104e3b7528a21e1e22c74597dd544e4a4965f50e9015946978f82c2f1fb52e7a6b24771168cc8abafc09b97d1ee83f63f2292275a0a7e9534c43b0e0d65e907b9eb3ea96c4a2754e6309c6038369e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h19eded16272051e3677439063aea121578938818460a14767a91fc50ef11e2fc23a5d0322cc04e51b4362483e4c54eb223252cc247bdf70667580a8dc4f1748a5f589bcec5474a283d2247ea136bd;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h8a0cbe853d61717756cdfb1283de0ba0f6522413f212f0878f6009d0bebe432a51f9ef91cd68ce97eeefed0bb5e8c00105674f166103d6ea050745b2f8c545581f6c168be817692d3af0a64487fd;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he7e284642b3cf4b05f5b70da566e54a56ae6752f323deaecc1cb9a0655b2dd5c869dde9f45c1a1e9a371ba9020cf33b90613b469f0e39bffc142692458c67f933048151bee2170651dee8c19d0df;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h117605906b58e517d3f41f93aa7dd838cca5704e3249323e77bc83c92f29b680e2f84788c8882550cdb1a164c4408264a64d712206bf89ddf6bbee515817ebb7d5ddc6132d7f115b6bd0539f6887a;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h4ae1834072723ba18e15f56ae55fa2f150cbfdc9e460cc9b4ff234904db697735a37af79374a4224af28997733b70776498254d63a8dea8d37f17bd416ffbfbe618bebed392a7988694748b62308;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h18207f9adb800c202533005752e339d8ad0c42c7340865a93ecdf3020d01e78a1b648781ac4f92c9e3e7f4df94c8313af4066e4bd489526c6600061ee6d263cebd600ea84235f34b282dbe00ee5ad;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h401dac8e4b0513f57f4e897849dbc3c938627c8971be4dda78109fc69d6dfd75bc7df46d25cd63df34980e77426d4f2400365a91cbd3db53efeb21c7105f50f163ba08455cd09a43ae4c2ebf1dc7;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he3392aa74648f52796f328ba12cb9db6a927fadebc9f0b498da51ead5b380e0b897f4498627746a818a932d73052ea2bfee74fe93e0c6e663c469d804c7ff25b444367efc54af7bf527977db8fb5;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16fd64302e764646e52217da2297ea436a344761e27a89fd4055dde7d293d646bbd60f1b4771bf77692776b8b83399dbf0c99ae3c2bcd4c171daf82d6988137e19bf6dd8e74654c9379002357e5a3;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h134ac3f79711884878648b7f30b668436ac4765c1486635e9040c182f48f79dbae8d0b31380f6fea1899176a4e7cfde22022e7368673ebb2a49439a531feda3444d4da28f7da3bbb9e738d31e3e41;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1375bc8fd2d4989c4940705b2d27dd72f6880b563029f3b748adfbd3ec6700f210f1a4506f2ff8087c999895bc7f6be3c670bc49279f3eb8adbf67ffec23eecd02ba443aad271f86631da5f321bde;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1db967c1f59901dae79f1e4e0e854b4e6676fc9d3412f8586beecd94ac0e9177b59813a49e6c994a7569e97ea4d0ac49fdabd703ccd7a825bfda15e8a9c3a6c2513634aad0f15e866e40d853c1de6;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1210bf24e18657ce8b4e9dc9813af292c5ed0880559f7b4c17e749528fc7f1724b2021fb854b3c560cfdd35f900d7bfe5cce9e1b18b96ea5bdc4f8af94a7b8f9a8fb0e8eea1bbe4565e6a4e3d8cc1;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h49b16ccc5a12fb9eaab38a49375e05779a43a758947bb9cd02c967d926cace7863f23976af120ff740ca595f146cda99598ed5bfd358bf5b40444f8430f7e9c198b0989ee3d4259a33bc34a241da;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h329a1590286586383845381e8d98d88abea8d1016500f3faa2047d33baedafdbbc71a1c453aa39b904678e3c0fd72ef206a5292e8887492c098b0ada24c156d08e48ee3dad894e148e0cc13e9be4;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h4b2b0a711f1006c18fefe889ad22eb36233199608971a3267feddf965814f9079d98148eb3e035f35f918f1e396f60be5a80facd594a9197bc368a2610c2d2818e1793cb3552ca1fc1be5b599c82;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hcf7e6db957442672c8ec9fc5ed610a89436873ecb04d313e78a4d9043aa4b804f8ad1d8254c6bc72a7b6e7fe307ea1cacb29ab17a36ddd47ae264a9cc500b9ab564aedc68a0dd1221809ecb1c52a;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb6e7e0c55f001c8ef00a41e742765fbaff0e8e61e0678ca252ee1e4aaaa94d90a709d549704fac8f8421219bbda571df00594ca42043b393bfe1e60c878764aa679778b7a9cfd2258214cb8d0159;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h113d457d6b859e161f7a34dcb2a8ad5df7927b364a733f4f9255f03ea3f040d80e0f08517843a6e1e700e9436c5283ccefdcb9aebd82a1b555ce8333dc9bd829d653080e0f2ace365b299d10c727c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b66238adbdf82433d5be1f2bf8370f9e9f0709e6776a5278edb21b1c6df341bcc8ecd27e53eb8051c30b86c4beb12cf7a06fdd064625aa2ab2831a0d26cc117c9a33c655ad15bf0d9b9207e9dd2b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb2c1d2bb997834c7d762162a8e8714cdb61a847746ef5913c323a97aa47be787bdc09bfdb604b903dd807920b95140727d5e8efeee222f138e2e2976383198514fa526999417298a0dafd10cec0;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h44eb1c3910264a9491fe46310488be9bb31dabbcad11c823c3254239e6886d9988eccb74c212509649d70f705f60f12a72bb3bc3f3fba23a3abfce0bc51d46097966b3a45a601787b3977bcbb3c4;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f05b30b5238ab2f948145cbf9776e9e3d250e896a6e5452e8d35c8248e819c7b0cdc8ce997eee977defa97d84e83ef75ada6872ef1d04528da7dd153453c473a7ea4ddb5d2129b148cb4c8b2ffa9;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b081b699ecf15ae3703d503eb9571d8536578b1b4ee09410ca5fd0d6fe0b50b0e4b8747a82720579a6f1fcab50bf958b08026a6d310578ec3a8ce34f7895c303aed7a2a755ea4f43b83af52681b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b4b0773ffd235907f76805fca0a00e15f2a7c867fa78790124535d24d2ac12dfd5788ff9f93d7379b661584630647b70b38acda0adcd7a612ed605dfa88f25853a70c42072cac5ffcb137f2e9f14;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h11073a311f0eb83f53f80c69e52063288a5556bcd3d227219ff644d13075a77f410051eeb08fb70646ce428279226fca574b717b07ef94aefa164bbf59da378039b64af262084a9ce7a3c1fcf1645;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h33b00d031463435eae65a290f955b6dd06c115c1291372858272b8ae7ddcc727f7adf98e305a02f65f50a637ae4a1cae1a2f671407308b45f6a4db4adea299578143dc66b8d940acf34f78ee3f52;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1661873346af4cb28480cb7baaed1c481270422e4d0c8b30ee643bc8b1794a049c7bc5891c7895107bb43866cab61d25717a1ffd9b8c2e094f4dd067d0f3f7b945de1801016bbb0af62d0ec3e3483;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1640a2b158e6858fd61404012222197ed2f8520335d5f774604600169fd0abc2c663e27e49ffabaa9264a29b6c5387f5e5fb9f79d228a0cd41b75b2ba39b2e943a59bf1e6acb8eea353e856c60057;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hff1d611a149d81a1eb5bfc5a6f8c5b9f319d2091fbd0e397fa29638c6ada388dfd85b80fc9649bd857ebeb930e0c02942a24ac0109904f5d012d9e4d593aaeb2396f170444f1578c8f7fae5a97c9;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1fe110fb2487d0adc21611b174dc4e27848a755ecc1d4967e622ec11eef1c84824c1b6a8ee7f70eed45c5e3bc51c660bacb2f3b90c5ae272ce91b7437478011f42aa20cd7e188e4fdb0dc50c8ef37;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h590dd9e91901b75789ac18388f157d0eb92cf990a29e2f425db0b9e295d9503c05a520982b3ada98529874ee931a51026bb784740d9a6256ef66e46ac73dd61b345db8d7d103f6136727776c0a64;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h13ec84f065188a24848fe1dcbc2f5699415ec5c771881a0bfff2a4f236c0cabc756d73ad1a655e03752d23d2b28d59ac5490d9596f250b3b974c423b51f26d36fd8be467d4a39053ad75b60f55d40;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he6b79a5ddd8a6b9b64d92150618df22b44e9e90dbaaceb745f86aafe92325d978e6263a8c25dd98aa8a25a992bf17424b6d6f9bdf2cee74903a122b8a74877ee4552f6008daffb823949397e0242;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hca6e18a79bfc43836241b58bf14893e52d4a9ce4c70d2ea04ac086918c673855870b84c392f2991aa724938e00710327a7a04a97da03f0b28388fed873e818f0ce312bc7bb4adedc887bffa89d66;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hdf2c83fbc8efba99049600fc3e39b475fd0d7bb8043c429cee16801192e283401a496581bbbd6885b73788f6a725d87bde49d65df3b60e6ac521950dd653fcec5c43cc9e2bf2f2ca2949173f1c8d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc0eff47f240575cbfaf4a81b07e84b5a364c73cc7d6ec1bb71d33d65d97d642e2c766beac35b47f25cd567d65c351357fb29cd24f66c381e3748a5c89c6da2e4cd05cd23b4f5421cfc14500ab15c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h426a52d93c77933bdf6bcfd05d84a1654c5e965d5609df2903a322bbc3dbcde5c498cfee1182a198bf1c36604771f90aab6c5da3ead75c58678342faf5d3591dc65d141fab96851ed7845fe200a6;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d3b526dc2e37ab8477e78aedbdab4a8953233434ab016aca936df048b34ad7691e7d1fac22b25de1c9334c91a2fa260271a86c1fa4db93bc264c76475922490c72aaea7df1bdd7daa91f2ca34f9d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h67377f607372b5b7010ca702d4e77719c3e23cf3d2cc4afcf1699156b1c691992c532fe37f9c44c6befa0b2ee480bbad597c2b3008f4d3b5d43ce3228e69f01bfe923bdb9f781d3eef38c9df8c73;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c90a6472dedd0e7388f028a337e53a3df7628c8a72dc37bd03f13602d402f852778de977d3835f634ec50d49352ef9e4e991dec7a99c7514ab16b4b9069ba78ab8b9d7698a2937a9fe9b8ed32af3;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hddb1b2127e85c67fa43945c04f4df5714bd81368ea0d11be81b6a8ff972600d28ce89e5dbcd7ca0a29f1882493c1acec9f33c4ef5beaf0cc90cd54f295b398f23ecd060715a3f7c3df9d19195729;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hbe17c5df42d68669966594aa9d5eb79e70768f2eb127c22906ff236f4b3903b2de5592644c6479d1b4acdc7afac296c5931ded45c157b11ad767e37f0b574ed397bac705d3e04a9c6e6b5935711b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1893d87d092ec89e60c0040e48eeaaf1b30b08e1312766c9dcf3a53daaa259c33715544e59d2e3aa8337e8fbaa327567b1ea5b76b62fbbd1e709450773a30a0134b3463828589aefb5497ac2f63c8;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd0f3dadf9dcc8c52725c316b62c4dd279a4e82c36bb529502618c5fcc870806489c19250e2b72750b49e7e785f6641939de67ab5abda1b47b070a1f7e490f4d8cf4c379e272eb7bf40f562f9571e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h18f71b806a0c3c40bd03073e8a1c6401a7d67ac09b01cb332e9d4880a34c6ca7a7f7ea578552eb2b16ffa249ee028285785597200ee073d157f9d5b91e6f0e294101a1bcd1b8866979498f703d322;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h2a594ce493a8fedb6d0d2b3fd2077621f0a9c61610a72c6643d20dfd192b2c6ea36d8944140412f88124145a36a543516d700010fcfcb9341262fa2baf002d1028190dbde37377faa02742e700e5;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h187c16072a36825d5a6806f8af486417066dfa123c6d5f7425037804694ec054b1d29786ee7236689401eb4665d43cf32a093e71f1903260b88e469416cb304f9e74961cfb892f76d2a3c3f2efc6f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd38f64f252a203be7dcb60d94c141bd49bae7106ddb2b3a2edbe31a9e4cc3e581aa717a8445f16001218799496a7f6d07b60dc669b3b38c32b1d4bace76d2b354e13779ec3053a930cc3b28f4f49;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h69a3bcbbd9090fe198db3ecdb0d7bc320ce0191d64b36786d342c705b80d64eb8896d66313b1dd389f3e4fc912f38992a8b9d1b049d40fa73e18aada423679a7e98a2896eb98aba304cf5ca02aff;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h117499079ad174b136301ea0273447a40bad8468b404bb39ea4d7060e66854ed996d5a575bfb34ba6d58ca6e73f4d5baffe3a1c99b33cbb0e43760dc085830d4ee0693659190a8b745e7f8aade48;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc533f6e4ef11ac227ea8695661ec1746d81e5e4bb1ea7977e4ae884902a19e64e2df93d192a261d1be44b696263c082864ba03c0c0e90d31d4734800ee6be31d76b4a26d443b806343d24cd2edec;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hcd5369f87bbfef8855928f10e63af2ed2f2baede273ade042b97fb2a905acb531db9a96ca69cd01ed31d327d575791ca587d5083ee6c4268e2d6fd0cea95deb60c718541125d528d68d6459f57a5;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h13eff43372cc06efe04d5b5e33e71a2a21a20fef8d8f64fbd094342b4a4ca4411bb9ae64efcfe1d1ffab14cf57b5425899f8666bfc5f1699be81dbcdc75872c2684a7609118548c8826c444298c56;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h572089f7b34a6be61545c53712867a9418acced7571de1dd00a1198e7c0e32634ed7fa5d096867bb32a2198c016e335da103c129fcf97e715d3dea1558c3ea2a8ede48b6d5d4ab92e29333157811;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h22ae691ee544929a181b5f505aabb8a749800daae2cd0e24ed3d0b0bb4297d26d615174b4fa57ac7617268cd7292a7453b720e11135bccec7ee400e916bf887afd5ae7e989f6f8ff37c177864ef4;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1df8e77016c881d0559b16c5984399a290da8a9a9d4febd7261b30e4fb39b312bafc97e6e3898000273312b9058326e0d63a73284d930798ba549b47940a45ff1c382b86661b78f7e0f3deabd03b2;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h99fdcb44eda589473b9f1cd8798665d18fd249ad845c1a360bd59b09680e8f6e569ac7e6fa17be14e61419628be92365947edba0c354cf5d9820c9b9712c1490c2ecd07951cac627dbf05b08243d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h17d2a4575c6c43ab99df1fcb468927f847ca05589294b7164313282c709dc1b245d8b2690f21bb1fdd693b942d65f1d87f63404b85625906fbfb8f0120f79e0ee16cfa7f06ffae9cc61f15ba7e7f1;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16b699ee11c09891ab4ee1031eb117b417c4a456d06454c02c484ac5074c8e01d6e02f9186f28e320259f221ebbdb2af5c5485bbcb84789479547aac4117302cdbd27f25aaa18b8230345d3e9a34f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hdfab67255a306ae2368242df30ff902ba40697c79f06a0189cce5a9cc39c815b4aa563bbc680b505975ee508ea28209d70d38f0ab3a01e7da67d7439c2918c72ee061032fb4310a318126ab177a2;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1be0acc13d5f957acb7677e735da8a7db641f4c6b4399f011d05b474a170061eecbc6043faa9c650e0d99e22e74f8abf71aecab73b7fba81da2ee4583ed148fc4dddc5025db60463a38ecafe5d92a;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h195332d953e2f9c805ce062de56015df22d16c20ed037a283b05e8b076599d86ca84d4deaf2f189e9bca97d9ae8eb4111bc8144f9efb203b4cf359f33f3a41b7d3ae3fa44fd95ecec24f70f71c900;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1dc12108d88354a0da850c3504c7ed7e25f1caa2ec7ae660bb03b6d877d2199465190b36a5bafc6026c063103ea726af18077fc52def12064c925ba8190a19ab80e42852e13bc29b868a0ea0582ed;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb4d4bdf33d576d2eb2ac6ddc931137e03a8b89cf406efc644ebbb82163e5c817faad3a843a776d997207010b891951fe4f13d0ea8bb8854e7608ec2e7852d3ecaadc9764ef8c845b1bad722c379c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h145b15e5743a044ecb3dc54dce77e04e50b20f63bb96616005afd9f1bc168e6831dbea350567848cda4e3a41e78b8e8652c0e6081e00d93274bcc1b3f3f531991108c8f15b8f337daf3212657b97c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h14c6106bbe121bcba171d7c58cf038aa0bcc92a21b924032a552270f3dae312b6eb5f487a78e606da073a795141c633e5b6b01cf8e5edc43d4208a60f304cfe4dbb2c07bb352ca260aaba4dc42a9;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h87f8d31bc54baccd0fad75d13d87a76749b36ff1af0e8ea3a96f3ee5f255a83ab796879b7eb33abd6e41f995b08363bc4a887590904ddd5c4ab46a7e43ab243ab2f47d6c5ee67cef471e9698627a;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e92bc1f9712a2d145d84bb93f47edcc87d8aae23971c8a20ec6f3b0280b2d90ba1fe55faef5826c13ecdb2f62eb86804a6490fc4522178efbf6cbe85c2046cd93bdffcc24a510dc7f2071775d37f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h676acf1e550739e378b837ebd9500befea37ceb3a8cb4f8e6c50d34145a98a3acc730a800ffbfbb1ee84e4ec455107072b2d2bfeda46866be2851d3f030b832d760da5a547963fed4b6150bc01a3;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f313bfcb5743ad2b1fa51742a36259391a5560682fa724d7596add2bd29cf724ba03cb0fd45a5366aa408b2878aa23046c67f7dbbc4d4a9de52379d703eb5e512770cf6c1133140a751367e0c9f2;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h154e459d120b5ae598f99d62fe1370580576c582e430b2b7bfe306ed3f10d81cf5c3092d6e851a5fb90e6b1a64bfd7e4d262e6569605bfb6479321ee000540ad97863cf7f7c4709f316813e496fc7;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1fc00cf598f60db0fbfd676819435e5877f919b70cae094e048ee8ea9401f2a83c31a6ce3aa7cb873c90f7116fa1b4b9f7901b8ec9266286dcb90e234944ace97fb57f34976b3fa6ca537011fd2a0;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h24475c1e8a8f0cd8fd9cf486d9446033132ae74660c691b02a80c0280f5ceb57e72dc9802d869b389febbe86230ec58db36bc4a65a76ab00c485934a3177813c7c066595e4b452d4c00a07075e5;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h4e34b597a793cd85379f7db1f6d5c1d7ddeb7a278e855c896e4a0ef2aa8e819a8c52c263a3115c3efcabdf0151f39741d6f59f7d1b76b2334faab5e7772b014804ed3baa0c670b448cf14e4897b2;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1bcede49ec909c6b3873ded11d00f5e5abadbbf7894fb64eafd72d6d0261d57f7420aab5f5fe2702438e45146370c80f7f534990b66e139f83f963490cb689bfc480c0ab47169d1ea590579f5bb51;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d5defbb69ede9c264012e710803c8c28821934c3afb13544fdb5fb352fcda3e352596220134598772b28211cc0c5795b71551c03e53a0131769a1d2b647124d68dc9adbfb7abae087a0b8b459bd6;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h181f7f9a803114aa4acbd112bdd1da793d5c6f398c27261cf8d60197a3b7009dca13ab95fdde91147dd762d70850f37471c4f4b5c787e3eba831ee7f2f28b0f1644bde38dbfc940b96a17c2c845df;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h2d7be2dbd0b258588803b2b92cbec1efa52caa5e725eef07d22be0f32fdef332a1100dc6c8f1788d6ff502ba75901e6614acb17962a9f21ca82ff40ffdfa68702867263ef024fe8c9e81598e9cbe;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h13f7dbaaac34ab00b7f92013858e988019c5c35cd40a047551c9e8a0353ea44a6609f0c47b41a1a42949653b0659b717f9accab6d7ab4cd798ab952494e57145a3de701c60af3d7f82aac845040be;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h19e4ded6d1f3733339ba77b267cb3a2447c48b05dbad53f97b788eca92ff03df1825457e1f6a457b1b08da08e1e38c137e385609fbf6c384830602ee1896604e61a689e96c58e67af41d2f4b464ea;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h119f6a3afced3b44c81d0d06ae3c960e7b4592d8655adee62e30bf6fd8f34d5038dd512583740998e0baea801e24cf7603c0ce6f6ace78eb65f85288b7cd42671bbbf1dda520cab453a94da10596b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h9219a06e94dac4dadca88f96819d4b6001e4ffee3a78f12ecc713730eb219dfd1f7861d7d8791a17ca7be26d7c925cb6e13710ddb2b5fc0b016255db7dda03cd86dd1146e1dd1f3277c0fb5589c5;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h14ec7517beb5c75173f03d98ed1ebab80aa138d43118cb258a3bbf9719e15b0d940c673cc9b5a3762ba6675e1e4a4caabc860aea7690300d292861d4a766803e610f0f22d481943504a78952035d5;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd6a7fd411f37313ccf8a030b5f2670312f45c25550bb8d9af0a0a742b45b8ef10a9f56ec68216d6bb3e384847a1c8c93904168b81f247deec6fb11176e8ac6cbfc64fc9947c6b6df5c83b1d2973c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h14e2ef3d018eacdaaaa5fcc69b19b51709f0562f30ff711e469f64f5a03faadaf91b46e5213570b884f4772e3aa728bc95b0760c6f0f45924d2dd9e15bd144b27f7a2c309d359801dfeec61711f98;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h158ac9561ab78fed2a82693ac7968aa9721e1cdc84dfe099abbaa65a66f3d8ac51f57575a1d090a54e4907cdb694878f6431671c0c1d4c1eb029306f8d4a2240fee13464ef22b7936bd534c0ddcab;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h109714f3f79897d76d3d5e06ac6ec168048cc2efb93258b1df9df863d579c6f521e4e35d4687a80cc15e37bc68e6c1decd72eb6b037c0428db78ccf8bc3f40213125ac87040697337c2729e9b680;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hbf2dfab0fca879506f42bd2ea06e8bfa5b6f3f1a0882248fc168487212190a20e2d6557fcb222b1cee5bdb112ce5839880e951f7007c9329e1152b9078427a6cbbf44f5d98d37dea6724275a708f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10f94a46bb70e4ed9a9adfc8cf3accaa8ebdea5af544a66d60269b07865e23d3aa3933ca9f08b9ce19c23c5e4bd540c18bbe7227df946543c6b360259dee0f567f28801304d7a5ba1a2592236db45;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h3b5f85eedbb441faadd8fdf966620138200adba7b27c46306d352e5d71e418aba753ee4e49b771c3ebb8427e1c5b8db26329465e1d30d5842942ef3f7a372832a21f2ef37630f29b76238d593c7f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f2adb284be1700fc1eb0d5c051668430c3ddf82da7a6b016ab6a0e7aa59ec37b3aef7d3c8326f31d00ef204d045fdfd75a7d155fc67a19227c9ba2ac2d0fd60f9676b5a96696064c183e13765f4a;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a95b9374a04b3cf98a60e18e0b67a43415339a04cde6c00736fb3abedc1fe834b762159641ad67e4967291d732e62b2a195552933a7f8ee52b31cb61f5941f6edd0a3fe757693f9ad23cfc0c2dd7;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h26e24eae5bdbf44ad44ac0dacafe4634339a615042d358e429267317d367c023ce772df464d24f7458d7bfd191eb26007c622a21fa2125a5b4a505995c95ff4f2ee81648f7f4cde7cd93257fadea;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hacda4a063cd527c98a3fbba8f5f73f0aba5c4d573f4836d31dde1c30a766b0ced5f983b178ef63c7ed3715e41ee353915361897deacb7d9cc41b7f96ee54092fe8c025e0a9f84a4d744fea31880b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h5b53ba6130a6a1917af109474a1d8ead02c2ca294f4711a24d93533c763c75a16ed4df593d89bad2f018b1fde5396c8419bb42c98ec4cf2c06fe77bded6daa52d2b28f3f4622d59cc7ac2451c2c2;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h5fd979fcbfad9076eefb9a19282f9ff8a31d417ff89dce66fc2a92f0eb8d2a86eb3129d1aee6de2030aaa75f39af262667238a6ecb3de222e24e93c4289ffd90ee61583992e92f5ac39353ca301f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he18a9bed8caa7d5fb184e057a8032465afc017c1b07a57ffa3188239f62d8a814196f2c193af725a91f4a01c86e4c15228b2b32868908c02413e504651b7ec8807616dca682b02fb6c11719a240a;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h14fc75fb571e7c0e08f11bd94459882605dafc3f0adf7e4c9660e799a69576f6d36136be28c84d3c71a4df6f0e3dfa421cf33b2286ecff8a7a91611abf908402b949059f81b26b7cfd9ed8e0a3702;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f5892b18d5acdaf341c409efe8c96bd140252665ee808a9ed09efb69f74f23caa225c2ce90843ba4eb7a1f7c3d1f372efe2d724231ef1d8a6ef52a44335140f594b1b07605b2c23ce38eeebf6d64;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10f23cf8db093bb922fed57251e71cc514895c9d77ddc51fa292265a21cef16b1523c81291aa1639cc1cf773908a57a445bed4d4e25687cc7d95b8bf9356f6dc0161d704051589592f40cf49396f4;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h170c26ffbe5cb1e571c70e3392efb0b17dffd3f605281f140f3e07629f66025b8ded9c7e5bac4047f067dd04ae6c967681bcab7f7438f2c16e494b2c20122209c3e47ac9decbad7a3d489ec4c5efa;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h5371981d43ff7c2cf65f2010df66fdc007561438e196fc531b97e9ef43786d6bd25f4d71d37cf15b02a66f57d934989813379097f3fc792829c26f36676ce9c334d8a6fd6e98cf0b8a84afaf76c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f313a4fec23dfabdc0f8d162a4408f483fa713a7140a14ac93bbb9f09db3a40b5d1a5d0a7a745ab054a3ae26e1d197cde055df4253897b7e45519b9f6278aa61492b08751dc49afb05b02443d656;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h4282ea88debd0687023ae114f3d7c2dd99670bb618992a5e2d4e21643920793027e627148557f6e70f387a6053a20df4de963e9338c8eb9c0b871792a4f98874a9ea26ab691351f913aa5db576a4;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha5ff02c9c31c4b86576a78b645c5d05d1120d91c40b2cbe391ff33af3ac4ca54e8cbeb6fcb2d4cb3e76ce341a0ba54fde1d79567f80de66a4a99dcbe4603fe46dc6a0e78d6717284f463d9e44de5;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h81840aa17075c7e26da1ef4f760cf104f09dff4da445b126016ab563c59160130601a0393da3f2449378cb948f241dd290af05c9aa38a7ed7b9e97a4835d1e59bc617a1d38d3f971bdaeba8b5e83;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h62fc7cab4fc72b2612f0c7b3b63eb4045a9755bb2bd5e7fb1628e910106d1893e63114123cce6d078d8cf1dee78f72555959773b26022dd40299d55b47e824d2e63dec31c6da1f09e068f977a040;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hcb596aace5a83ed9f0fdef22aea1f020f1c6583e5b235b51adb9ba0d1eb67e5a8215903d5468199bf034e140b37dde74afa08bdaefec7197ba8be73b780e15bb4509c95d3f2652645f1e53d2b64b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h15b379abc7ae306720b665ec8016c199f1c9cfee6f8fc41a44e4a7ca1033c503be79a8fadca84b3fa3c3a16b59e795c541ff1dbfe82cf3e72b92fad02021dcc3e0794d583342f072b2be82f3bec5c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h489d66a6c09f552b4bfe7f596dc3ef98574b2d44686620930e9176901606d98631744245ff60251c107c1e055678396ee9e1588de6d6490c44f526b452aa2bafd0e0a91144fcaa96efd5a93e6bd5;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he1eb5da9ff95c57ce6722d46932b383d9232a8be3110a25dcd58f5458ac8820b3ac2aa6d1cda3fd00a295dfd224c19518db3b7ca2cb2153201cf06e96147aa2af49cd24ac0d52a24736385543e83;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1268fd6891bafb01e5dad9816d974c462c55cda8287f36993a8f92dac2dd112157fb6870987bb3adfec30a3fb9ed7a4d8fc6e4ecc2f2ffb1406b9a7a5f9c90f5c9b6945976f233a99d9447b7d1f32;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h4628d5b99ed5cf4c4f5745f5269dda8b78dbfb6926e827741bdcd960e45bd3348d9e5daf328980eafffad093044a7881e2915d1853b919894524695fd760a52bce41b12880a570d0ef5ca7db233b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h706b3d1e68ed7ebf875084d398e03f78f2bf3d4d11eba63c968b824e29ad16d336530ee04605dc7bd0627b58c855386b20078169799010fd7b87b2cd2fbe07d8cc1e0951e9266681b5e9fbb00bee;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd2b6fd19e511dea94abee843bc6edbcfc79d7465de1cc8276eff1cae0afa55b8f2d239e1abfd3b8a089acb09afe59a21026c5236ab48599fa17123ca3497b944401663a7adf40d354ad9bb305372;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h9a76f3f9e86d9e8ad2e385f2fa909a1ec08a7d8c036d3bfe2b54c7043ae0adc493148fffb702df3b75231e0d0bac3407847d5a70fcc27f9dea46bc355be925cc4821e873cd558967419aa0b23c01;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hcd6c2e44ac059bed96a92778a81dade902535c3e873ccba5e3afc4ceb7ff55699134f3ca12a8c1707179fdd9cb6514a0eda721358b556d44ff15ee95eb6fa571ec5b269846f6a8431548240b0f61;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h15155e3fa5612202323e5c9e06464e353706886f15e8f207035159b481b5b6086f9c2a28dca747e387bcc8baf9643e9a2324d269a18ff6fde78c6dd1a0588de684c644125b4f311ec6cf509785b90;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h4a3c7da8da642c7e38c832aae5d647e47db2384beb37b8163455fc95bd2cd1fdb00e04b05bfdd23c3e2fa4034251f7a07792658198bc08493cd1dd2971412c81c5c1c79e6342d15cfa8173a3be42;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d95c78851e668b8be6a699dfa4514fc404a23486e0f89d0e11e8186037615a3bb05903ebd5a9b6e07ede6fa179a1dfbd50ceefde6f70b2770aab43887149b7121616f5670b69f064699f282c664c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hef92d96337c3006c4a52d0ca01d9e75550ea659b3fe4eb0bfd910761b8096534463e8cf6d327f39d8d5c43bacff060cbeeca89928128fa7e7a6b6353b78375ada3d15324efb3fbccc2943c71fca6;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h708f99699607ac00392e9e5a30455cb732250ebede96f2bfa5c9d8154fff83e3fec5e7d853892d6f1602b0fa2e943c40253e5e356303a53870c922c349650719ced71fc34c09e37c350b3353e69a;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h175141c9f8cd2428d3b7cff08a0a1b715c0aed810a161d4920bd7ef8a7c423db0bbbc7790254a2bd6783be1844e0891f8cf734e72704698eb4bc4ebdae143780f3c421e6bf0d027fda7da9eb5ffc2;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d0fc96d6743c17c82da8a426a5737f3df6d5869ce1c4a3ad2b19a28bf0b0b3ee3bcf1aaa5023679b03adbfbff310e519c8576b25880b78b69a4919bfcf1372a264615422b85539563e4e30036d94;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h329aa89ec3e94d1b05d1307ff0632eb30a3c28178524bb9b787d4dfb8e4c1b84aade5e562e846b8849d51d19e38a604736071f6bdb214c4f74cc46e2ddccfed897cfc6d880baa9c51d40c93472d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h34aa784ac6f18b02c787fe9e35e70fcf3f91d5870c5d0ae09d25d3ce782d3594d57cfd22e2dc9cf54f64b6f6b0e2caedf362b3df094c3ba15d675b1aac59a0cb99c260391425550a9a300e3c88e5;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h17fa95bfc810171ee133a6d50da38309339d50ffdc54d65afdaa0e8dcc886605f913e9016a44e7e826a8354dcedb4d833141d2cae49135a755c5f90eb470fc8262615037a63573d6ade18e32622d2;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf72be975dbcbb8ad3cc0a037a3f73201ade1e8b8b3915976467e86aa31efd80de68ca925903748e63d638920543c9ad27d2ebc74e135b8c9c051c3c94118934f04b5e1d845475fc8fe14114ee356;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf736b18911e189afefee60f03482f3b3d1494284db611d81648cf6fd4f0fa80a226c71ef4ff68b06e5c221d03ed1477748a187991661f4a77751b014223940888aeb0b93adb75bc88aa696bbcec4;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h14028d88110625efecb34eccd0fb9abfce44d752e4716d3954c8e0b4d869b4510af804f65e019326fb7247d7802a567c0cf9fd86742bd655e8b0acfd7030bea3d73ac2d9fcee8efe15087fec723cb;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h17d08345969b019fc0126ff9a3b2cd8b4dcc6abc781db9b6188e638dd02ae710a24499e5c1f5c5262842ffdac04610a3a5d5c12b06b6c85bb69f0b062bcc8165d5d8ae24e6feed5972201c06ce763;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h4012825f63f211d8597b5857570c9c2ef3950701e87056670f1af8c9a7147292278ca90abce341c023e4a39f57b666ebccc2739a3b9bf772342b731e7cbffb329a709c2b18efa7cbe9442fc052de;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h151d5a982d718fa7c0226f1f2ecf44058a6e52df9f53bd1ca771f4e64f474a54318e99cc1a9cef2954d9febb4543cab0bf845234777614d192a271e47b8a327bf3fe0fb5fd0493b8a7b8a0bfa5768;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1be4936bd1ee827abda71a924facdb379bf526eb0620f9e0266ccc244c8062e6a6502ff0693f38505096b17f9b9d61361e1b80036ae4d917cb3d935fd5209f70c5cc1536dcc71482177d9ebd64f3;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc1888c03ac187f9546b338b143170ed64d0fb697f9d93d27189b15af8cb0cde7638e9a8adc5e8750d54e0cb714cf7c5367d84c45c6eff54bfa45cc25d3e70140deebc72d7e6f870552058bf21392;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha043546dbd21c89c9d35683e58a143f15b83d8ba27a0d8c7d7f37b5fb0cf3aad10011ec7da02c9ce11ebeb5b89c13215e69d8aae81694d2bb5c84e988eeff40dfd904e7442de667be62b17b2d75b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d6e8711666d220b51f6350d7ff0bb4cbc4cf4f74efa0b77431ba1fb9a1c6aa1efbf84d3f304bf446a00368fe67434e4c6c266dbbe84084482b27e5908b14887481309f649f6e419589bd6e7927b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h210e0f03c5306f11ae29542056755c27af57d53cb4411b65d8a2bff332ae6f033fc289118af4c0c6acbff2c727dc5481d5271b73879c7aa63c4339e0cb2ad6e1a208cfccc64168b35d8e244ec2df;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h19ee520f59a793614ea28cd760c3d98f48a6d2974a9c3edd3c7ec06d1f27dafbab72e4681b72ced60667b1c9af4229f05b89882b9aa7e990f658985f0cf67505dd7aba6abd302fad8438e65f726cb;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf4fbc294825afd5a3b1d0fae1f4953c12b9aedea6e55b41bce26189d6f423aea000bba990bca7056c539761810a1627c2ce1b7f599808df12a70bb6e80d8d48e70f625f0208d627582728ab692e2;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'haea6164d954ca06912120ef6f6d5c2a11d26464e40aaad1dbd528e218ded10cd4f47a84d2b0f5aa10286267ee81cd7c8c7dfc2b0deaad3d91d29996b59723d38a66ea90fb8a245410d6b039f8064;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'heae68ab4c8f3ff353f3a4a7ad41e041e36661cb32d3da321a63b1b0a458f69c734a50ab87cb0995b6239e30c6c4f5375fe77d9cb0351de763ed1143254a2ac85c6647de2c82f71586905dad2f293;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd2a7fe2e9d3836c2a1d765b18f6c7858c3dd5b659e928465ab938d4d549ce1f31308f514cb10c658cf701612aa2129934c6eb3a20383335fe5ab99ffb17b21e6b2b6cd78ed39c94dbd19b98171ed;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1877c85577b2d12336dd93567e15fcb7f618aa40fcfc7b8dd014be019fcd4b7c4bf6b484fb1ae2668de2eb51f10d7430ff3afecd59674cf9951db27c35175206d62abfcee0fab72c3e90f94922d75;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1919920852ab15301fc34a9af2c529d2ae2924f41c8e9ca7b124ef5933296830e2ad334549f3e6c2a930a50a472e4583bde25d611e5d639330791914d85268f5e3d73015068a0e8dfafd615295b7b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h101c4af9daa62a046eadefb0ba99fd476cb23cd18980d78613743e98900abf7f9f48e35a590d3dfcce0e30e7b7135abd12d9affe75f6124a318be4b994d878e9e47796ac5258c6615d9e1f2254e1c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h750981c8c222ce75ef875efd4dac2ca6358efe5a4929871e9502311800d419e6dd9dabe7c683db3807bf943a34070c7abbd066d75e98360370f201f7d97a227d9da720b76f98a1baf48d5f57128d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd0dce9eaef9ecd552a27a229b851c367d637a65bb5d9120263666329a10a4bb13ff987b1da3b5895179629536a01e6811cdc127c963b3b4d54ca288597fbae9975ec956d85cf8451ce4b9b83987d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd52061a9e1e2196a508e85762026c7308a8813d60337becf0398cd9ab97a26a6f64a65d58984b7e73bb9e45da1fb2f1e1f0c676b044c7d19daf7fd07c697992705ca52afc214ea46e80917b8fd7e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h116a2f858a83e20b1eb2708849cd13a4cd813a722ffa753872d67cb1dab59f931e7ae4676a7b1159095d3376af9464a77aad2200b07046154be874c6a5c858a361ae58e03ce9f891cf1ba1061b98b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1faa97be941d5f927969ef894885d91d1cf1c2c7f666f5af5110fb82ab567eb6434101b0d9562dbf6ebf5f13c1b596925615a0220cb0cd9dcac23e1dc2ab79c9bde5e8ffa26c5af6a77f53c3edef;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h2d82e93b3a24a50791d727048683daa3f4c74095f29c507596ea4c878501eab8944af539bf7ded740d5c775d0c98255f921f953097f964d9bc03d897f8f656a1cce3e5ae2ffeb3c37c49521d0482;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hcb5ef9a47bac7940ba7fc5d5b07f231bc4c6ecc2b42feb0e1e7908eed16eec22311c7008140d4afae6380975e04957cc3bb01ec4b8c668064c3ceb78baac422c0823526d8c1e38e71f08c8cd0f53;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1358fdd2fb503184196d775b6c5ac0d4bfc97ce928a6895784785db9a13f4a55f7767eba404ff91d1c7b682e3e62d41fc6418b6980441a730c58ec935c712e708ab85923c7ef2d0d68ddfc56fe61e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h8fa300d9c470969e0413066f56eaea7a9b39e1f598c60652c315a8f84e6484c9c218f6357d16a6d5e2a0e4cfdfdffd5b7327ca0a0613b33707a488b7698d1029b96c00ec85e00d1239a4c454c30e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16a7142ef92095746c1bde15cffb312f4ff3f1e308c8ba0af761c722471df0a0baac5f9e4b1339072e06a342e4561369d8705799c67d003d6e1b28004f35e5f9c7d300af74ea3bb9a3d73d5ba236c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b00eacce2ca53135914ebb6fb210d76bf4f9462f45c3ac61d5e105c3c58a38eb421f5206af159fca878cb77e72158a6e5a0bcf93ef90e05d4ad288a73ce9bfc9bbed858c51109bc5ed51ca7b24c1;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h14f05d624c9d629499474294a3931c715cac54585c4241b887f0c26989b4521b7fa55338b7952770295f4a5ddb33a58a7ec9ea99eafb83ad01b92f054213cfe1fa526e4814b7371509a67fe8a9e3c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1fb1e547ebcd841078a7fb79a4cff473a4319df88bfa567ae61386ae70b5ed81480e94ff50effc1b53502d335221b10053971c5367719f7c2b2aa0d46e08d074039b7b78bd3586f4b95f7e099d5d7;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h4294230832cf3fcca405d7f0a7e35f20dd27920649615da998dc9d8f0c751d5c35a420e5331f58fb7dbaae06fb043d9d2998e6c4506b8e99000d25039ad403286503846aa57a28abacdd0176178c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h13bba9bb4f96d55b2abba86dc54bae509574f9df32121ed1c071235fb71153b598dc1135467841a5053accd7676b5ef036cd38d5050765492f0bb4d0429ffcfd1cf18af5fbc1df00ed72c3fdebf8b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h668d249ec5e5276b11893df8e0426eec0b13da50477780a031fe32cca55c501cd71487c423f7071b7d630e4fdc705d07b9ab66a7349c087d45e619e1c3e21af21a56f9ad740109057552de53de77;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hce03149f9f6c2304092f3ff007d0261060656720080475f78b767af64b83ee683dd5b771335d5a07428d8cd6588f6b19b0c0e0bfc5360bf619a1039299b19f0817f936a72cbf0ebc719e1fb18b43;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hba1045a49a8768d4b79eec21d4f6b9af22c5ebcb980f51540288463bb62746f5087789f8250f292a8f91acbc9b578c8014039a635c10682a0ca4ab58075eb662632f1874bdedcf6b3462531090fd;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c4ff51902586efccad95210ccb55282fb28f96401e9c799371064dc7b7e6a54e89f7066e2394b16b94df6318a985260df017f386c7551520fc4490ad1ad0d0d7ab1b48e4866722e0dd725a044d96;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha1c6624962afab146542d75270c9dfd4b4c794e3713d9a059db857c7800dabda6d4a4c358d8bbf490483869927631020d2e644df53913468ffe8d4317c078d2b8b14d1d04bf39556826c8852d67b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc3007d8f2f58c7defba50f7d30f35714e5f9d0a1ff245ada8909bdca482e00829e8ff11b085920be6cce742dc82ca23f21f3522c4819ff81103305a15f1fb4f11c41eff09c3358acf4057757029f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h11f6d517a6dedd40a899a8bc3b437bcd756ff2c47b99f23c9e677561c73b7653bd5940f775eba893bb564df55f6cb93bc513180c159ca299030ecad9485e516e4fea99829d061333d1865beaca3e5;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c0835956beb862a32bcfff509b3c49d73fc639280754a3b51a36375e97eaaae980acb8bf1de7e61780e9f2c9fd6bb5d1fbfd98c9f709348fd19f544dfc7cf6ee486592e71387cbbb30afe77153dd;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10cec890b3e40b7cad9cfa95013000d5c9039ad45e2753b9b973fe55a55b7a0e4957a2aa7a2cad2137beac3dd417b4ee304e353c60ceaaff5c211ec9b2da53a20b665d8a0f66871fe12f4d0189a1;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha56849ff34f726732db2906167c77a036c62afd4ce5262bcd70024acc4785f4599d72877109af48f94d71c2893c52e49d4f75a52551b9ae025aab4500138d31e94ff39cbd3c2d9877836d92f9f7f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h259653c72053a69deb5e7cd0e913b4a6d31b6ee5e5e058829a51457c4d65c4e9755b8614779730fcad07c441d3b412b26031956ee3b5dc3e3d19f4a609732e3b77f34ca0d9ac0ddc5cbdd69092b3;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h160831921395501d61c58c28669202539a7e73e81e7c97ec271a0aa4ec05e2f8b97a5cfb909b2b588224990a1729a3aa627d5a332c4c2c1c5c03c8a777e238357643bb86cefd88eba4cfb595d8acd;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf28a247f8585ab89de6a42009f802677840030f1ea446d2c64f52c3d74cde567c8ec2c24af742fb662a6fdf039198845ea0668a05d81041ac2fcbe31c0f3abce41beda10384c20a93b5754767e13;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h15105651a486ce270e191a2a2f16ea1e63f173c1c4ed16dd5b7f36b95b1bfcbab834363eea5dba50665a925b7926c7aa16e5a09f637501093194264ed6ae0baf8104a85de2122d25eaa12b61d4882;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h35b9d28fab256d765325dc212fd3185c424fde6c134047550266b0961f607b0796ec992cf3c50f4ae12b2e96c086c08ceacfff569f503263e5899adc3f830f4b1279c6be77584026f2388526ea11;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h12ef7230769c4fa9a587c000c3550831874b66190484a7adcc27ed0fb1971e11c99d1be56f2b12b28dbd3848ea6b93af2c4d27ea3dd272334a06c2d0098c97b7c0cc472fef43ce1dd07384923a881;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h3973eb36dc66b3cc17a5d61480f269d9a2861dabcd5f26c1e695fa571bfcedec1b7a2d2c50a8d836734d0ef1d10b46170b42ca718b78d3f3ee18ce398178c11458b5054c700bd8ae6b7a6cdaf2dc;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h9ec7abba4317ef160da74332edf824c925cd18e9381679b7c58300be29e8bd80ce99413ea905b658a510d82eed77a84f8b538047a30037ecff62d996fd3183c0ec074f0490b5c2f19442f7201170;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h6e4123ba117dfe11e067c3e3532118f6447d68bfb63f7836fdbec97cf77ea6c45a623fc6954ac8caaba811799937cb45d3efbd2cabae0d3c850b525fb50d26c30f53474801c7bba82a2b26bb1662;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha476b677d5bf0ede5c0ef954e0d15662dfa9d263e034f6e98953a657f9729f1271583dbe5fb65a102361db4271a141db487cc6b99e898fb63911ab40113d36f37cb681eb11b1fb08977608c098f1;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a9c734f3070f81dffae3eb60b735f1e4940ac978f70eb400735eb7c317d744f2fc6d81cf58bf72b90cd7252129e36da0b925dfa611a16780141fc2c676d2db72f7189679180120d72ff92863e89e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h5e89a2c6c0519f962df16c63aa03918c54ccbf577fd250e1d3df2f6ad436c2a768eecbe78286f4dc81ea7beb2f9a23a6ffbc5c0adcc684e97cebfb026b0fb849aec94844d59842f00fe8ce599efb;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h8c1e09432b4d0c4efcef77b7235d056e8535722ebb1412e8311110da8f43d3dace7db04c6f9abcf9b34ce765eddf0b6ce107779b231ce46944f11b4e1828e3946ee7d1ffdf8ee0b01255916f1317;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hfef52156403ea8da4072d32173f46060cecf2b07733276cc7cc7a33176259d5d2686e41596886d440b1a7a8f758a0bb1d70757f0b5f229bb4a91ded3c931adf9bc2e6dd5d07a1cc5cc991f1f973d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h3327e0c6067206224ca79b064cd3efbe2825ffe0b8b6c4dfea6e3276a10fed132c019aa191244f2a76b4d770e22d54321644aae963aa7dc2d073a100f2db2c67f1e5fcbdde3d2c7e11df3887f866;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h6388eba6effb5a657c3545e176c2693e925fb26214412e091e92a9a774f0cfa132774e21760016835fffa8564b95a7bf3951cfca705ceb14dd6d484c583bf6ad790e0354392a698ad78dd361c721;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1354456577fba8833dae2b29f1e54091a768937fd3f2614f335e47ea90c2176a7f60a9ed9b7c26e1b55cf3fc22a46d2f6ee5f4bc17b04ad0de60b637a0965a7c4f1fef2fee0b53b15eded14b2bec8;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hca8bf17f1014b6b0a64af8ba0836517c86d8481b73f41b5c1fa9314c7ec3601f4b423c75d4f08f6e2376c588dde25cc632b55223da7f9545c742dad21cadc82b020cb480511e4c25b64c1d8481b0;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'haf40a3f8ca4a75d8611f531514debfcaf970b58915dfc5b04f6cc31dc84dbb72dd0806b4c28b2560461c90cdaa1a627ec9ffb9dd82e425e91edc4f6664343005d654e18f9681785b807ccdb4e25e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1039865ec26b9ccdfb6f56110402886e70c2dd8c1310786c851989ef56660a9ba63e5003b370d0e91d50aafda2ac3ccc8370e314b3c9ddc2f1af02f19c4dbcefc6db05a91378d769bca16cde16a30;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h8297cb9668108ff8950eaca0fb49a48fa0a1b764f394f384c52676340fcac782e069e7ad838477d66a64df85b2d78ff243e9f4d00852f7307969eb8a00a0910f90b3cf092b421c226df8c2bb4f17;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h11f2f7f6a97a0e2c7c5ea8c6f628062b7f9d4942be5193b4e60de865b123b240320a4f810ccfd968ec43feff4c0b57893a1db857f06d625f9d14377da409ef6f400d5c9664cfcbf4af6e3a037554;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h814d45cb66048e7344678361f5850dae2045716a130562c32ecfcf99b831cec8542744096ed5f6fe234b8fdf8ef6eaf6495bced03d2b3e6e2d358e449f896a7a1fd2edc40aeca5cca26b9561f834;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b5bdb3a5607f7e06d00712ff26efca2d25854a6d6d6008f0a2518db4089ab4f8c3aadefcf0ef032d119f990aafd273e7a4f4042c8f7e5bab5550345d424363a6c1fe7411134502a91917b53657e5;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h18db1f3c8b806b9493e182f751c15bbb80b77ad26b188cf29452f6fac28d74dcae773b9f0932cf9e83af7f41c954cd4391306bb3807335b8ad1d9324f46f506177c05f58a2b0b867dcd12400be855;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h9835b2495aceb39ba1bca96bf80fc6727f9fc56b336742ce9e4231f42c5e6ab23804c4a10dfadaecf7ffd82ec6c59dfe212f9cb0e00d699c7fee0eb0f9839f8a55e720cd3fc7374fdd98b4af399d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h4261e40f765f526d65a1d0d56bb2eb0b654622b6ebf570a469820bf14dfe35f29506ec576f6dd54b9ed29fd0c65e1e1385976615e0975ce5c9262649e9f73295bc16b3b6a34abdd092fd4dc4d24;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he19ae147e695b92bd30516e4a761155fc2435c186b9e7aeaa4ea5666e8f3fd540a8c2bf95b960f613d13dcee8e29a5f5137ae14a85a7ffc06c629b15b7b4d2b553fb06c607b8852c1c49f63f9d3;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h63d700506a75f4d7194192dbd104a4d3f82732a8ac9fb7c675466933cf4d7091de12d11c3e88cb8cd57dbe8d6971e83e64bc894ffaea78374fe1c6b20d31677272dc57125503c402d6c5b50751e4;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h6bd43f8a2483787d5a0aa3ebc33b785b95575061d15f4818cd73217e639d84e7d346cf6314fecfca85d6a605503d04af3029f8ed5e78cb4cdd1efe265219d9de8aca2772571bceed882a9c08b81;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h50358466d3cd199e719cc3fee0832025db4dfa4b887b7a77178fede8813b67cff52b13c7712b3fc0763a00d945b3f455cd6d51404e4e4d34a8a417bbfe0ab18f260252e719283ad7bae79a4d6d66;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h61f41eaa6e6185868501c90167f2f79688e6272822695c198a4d260b12e69b813ac681cd2e316fdb226d83bb19aa8d633f0a01b3e880492db80bc7ba88c3873954b6621b1863501a226348227792;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f1eaffb4b61aad6865c2ccd93ee116499f8541024219f96ccef1039427aba5712fdcc76abf2387bab3a0b08729b71c92cc7e83a3b8818a09989f3d557334be47a0ac126e84b23d573e9d20f9942a;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hce61c410657f6a7d0f7b1b8c541b5d99279541d38e5e53f9e8a558c191dc7bb2b6dfaedacf187479211bca95986e47bec0216142bd57b26d7249dc18b50eb3adb7c40317c38aa45894d16feaa45f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h30f7411c910ff84a5d8c927410c7ea8e5ecf8e1f7561fed54347a4e3cc3cd915f97c0b35bb1613713d6d77a00be99e7d64212330b68030d87ef161f86f052085b26351db5f8029714b12e81831a8;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h25479bcd942933b62f649f3e5717e2019a3370d1c4eaa2090f6b402e350070aa102a243be60746ced87bead28db60831d72589e1b973ea210aeea1175efc370571395a4b6aa2adaf471707935bf9;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h13fedb766c36992ec132fc18a5c943b3c36fd0db407625512d00751c1ee334a40929b27ef5d1b792a9a01a3fc63f31a57214bc02d2a5396fe8e2f4cd8782a9f1f35fe7f40309b4714f02dff1c2be;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a81fab16940632a206c5a0c7381f6ce6e161f4c528e3f0b483e91ee2b0d4c05d3b29de1610d484c73ea937ff5989116fcaf0f49e4e4f5548f9889af425a177928bf72c7cc6650779cdf4dc60d71a;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e8ff7e0ac2f67969fdf18629d3eb551b1134bd2e5024d0ffd44056856e216497fddee6b799de6777444256b48647335df3d04563b2f054cab83592e8c11f9c43491044af3ef05facfcc60ac6a72f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h15e3006dc13d01fa2c8b344007954644d44d483bc5afc4481e3ec67393b2886548fd61cc2a3f3921026f61652be891b698536a980784e4c6a9009ddd82b3413742778065dde9087afed78a2d267fd;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a3e1c42022e1f755d3b843871c97f8a94916791dd599fe57b541a4ba9ffd8e3618b3c5a9d5b5dfa26f2d9df6f2dda21cf8cb6a46afd370aeed9e1993955c8b57581a38d4a3d7d74b2055fabd1c5;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb07f25018c186c731d67d9756a1f8065b54a1f6ba2ce5278e8c7b2f41f06765606669a8c76e384a3f2602caafc9053ac3e0e83a5ae415b4d844b00d500f514f35f46df0e5321f922257eb09299f8;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h92ffc0bf211e809c6ccd73c49827b761bb033bdf772db0b846809830690a2929523a1f7e0d2c8abb0c75800ef78885fbcc3e4fd697374fe99f10c5131725a8f24068b635c2e993734c7122743e3d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b39c30f1551f730dd1e2eded3ab2eecf068a2910f8c8cff2ab6cb9dabd020e7f06992f9634ac946d4cf60f7b19106c2637ff87d19c3bcd09e3ad2db2dfd737119d2ac53064d9ed6dcfc66fad82dc;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h137e3abf2f3b145bde55552c69e517418e0b1388d8a512572b14ee1745c1eb20b3da0df4bae29bfcf823727fa2140ffd8f97aa811b8ac4e654d398b05d9d0469a51df836a33816ce266b906eb7676;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h94d10474456bfbd7f029870eacaf0631b834763f21154059d4df3fac26c421e57bbd122248a0c1a4fd49697dea12d64e4ec3564687f3451b830853a8588cb68b8639495b0e69088bba227f6b75d5;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b55f9485591ffe7e9779dfb34a5f4cdf99858b89afe7b7e791f8f2320f634a9fe57e9a973a55e044ca6eda5c3c26db386149f0bc93039d385e2b7887ba2f749752f92f812e5f1f3c07f3aa663105;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h191c28689b87c3a8ba4fd23a60b00cac2b9c2958951745c45ac84b7e3f29a5ac0ccfb158f565bfc6f368e07084f3d4e1d01b0da68e8e645a8e8caf038acf4989881b4828ae1b1027b691ca23b0bb;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h108728c0f32ed83ac41b0a433e706ccd25af87c2905734a51929ab7ec419ad0f904dcb57594d35977a1204de412b6f6bca350856f599d1dfd0cf466dd0ec00bef65e270979d44cbc3e2cd7794c027;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1501c05acec16bf762582af362b12a8150788e4d1acd9da7e9d4d435f69963e3da7d5b9d9cee7847284f7678243ea349189f0bf0672d1223ef633d43bf8edc8d12c445e5d202c071be1f3aa220ff9;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1362576b82cf2c2cbc32d4498048fdb5e2b6a47a64bba63f94f37d14491fea123ca4fc23453831c4457db03e83e3eb17463b76fad08186f7837ef776f995134c8991ceac143e7ce12e9edbf22875d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hcc2c17c3a20409c82e3b1ba6edd9f87b85f800fff5128fb98171bf9d69cabcbd5f54e27b1b2e40ebbd19d291ffaf724766b3f5534c788d57046187e0bede9cc7d82f15d1366ab9a65d894bb1115c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ec0a6c43605f01e2ff80a50f7ade9707b9bad6eac13ad899603877a06c8a5ce4b19f807ba665ca9c5a8c6666317aad6883b9db129633ab6b6bb410fdff090e1f6e5a342e50bf48bc10668ebb5f34;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1543329bf84e43cfaf4738cf20b6404658082a779e618153145aae41c8b28e7dbec95cc8d8d41625f76a26471246d7ece721176bfc65bd0b0e9523638d1fa2de8682816311bb029772ced952ce4f0;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h187bf80959a2c12ce4b0a3e65cb0120eb417c9f896277b4d2935a32f7ed939379a2f248ac92fde48b410c31fe8f6e89ed585bd0a55e5bed1a05f46f41c5b8438a376460dc46aac185bcb461bc279c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1fcea5386c0f58cdcf84f3a872698ee9dd91f9a8f3521adbbc10de3db4ba51f851b83384b99ccc45ecae081cec7111dcd2e3cd5bb58e62c2c13957fb97ab5c6527e724dc20248935e1af9585359fd;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1efc5b359e6d72b146d788f5c15331fa19b2475c1e78e574732fba2653aa34f0e36db1e0722d82ab7a79d8d21779f8c5f8431a40daee8272066ef6d3ba91349ca163d30386fbd7e4875dcecffd606;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc0aed42b2d9fd0b22376db19c7780d1c622ae17a29545360d5ec69f6f60a8b1fb0b7ce69fea429dbb743388bb6b5a0fd3e236ea84cfb794a144f734d109157e039807f14bfbc514ff1cbd135ec83;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h183b06aa6229d9eb626ccd7b124205bf5ade9c1bcee26a5d906c01f79675cf498ac4832bf31cf199a33d6d22156d3fc5f80d39380b1bc7cda960d76babbbbefde05a9c08174ade44baab4a705a6f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h11b8cfee8788f057d2fd772e8c58db1326d51a50ed265088184bfab91a0b444d0cf483bf1e1ce6bbba089a249987d65537ba97a5eb61039c7398a9442f72d104354c01a5bfcef366e24ccc52609e6;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h46b6f79c74195365e393e1707cd929242e55a562ecf5d0a7236125794f0f160896f7f2fb11daaf4708db61823bcd59966a7270ca8461d54b7ab49b97c91736a5ac221a37dd96e37c8ef9bc3c2040;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd717ef1b8afe33f6e5b67d7fcb6ab884e18df84ff2b9e02f3fc355d091680dac532d2ab56bf0cea52c86f9e595cacb88a328089c54af042d85b101cb83647d9c6375cbd5479d5432baa88456446c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb8bfbed7299cf407356942579556f7494c04c869751d23ad466ac0595ba42404f7a7791ed7006f9c2a8e9b53314e67b924f8678fa55be4c7b9f78e0ef4282f42bd1446fd9b0f386f2c22d90f8832;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hfea02efb49b5422a2c09fbdc1f1be6dd721160541e5a14cd5b2281acc6cc3e2f5a18b04d680b05835e955064ce8da45bfc0575241bf5dab959637491c7e35750084b321e32c6671b2cf21c6d570b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h82a7a9aa31d100607aae4364614e3348d6bd2a826976b7d5ce0d76342eb6685a6e8889401156c256c2d12544b311bc26e796c78e079198cdac9ca6a964f4c5d178fe20c61d77d866f629b0967c0d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c153170014ec8030d3c3b872d29bd4fe0db25da44052b61cf6b10f6168fe86b7fa8a8e6df206b1f3416b6c3cc290d225350cd292b476669efd18115840cb644fbee44d882bc1bf7268f2c89cc600;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hfbf708d09fd640e4e6e29de0b3f25e3d693e97b4429a6715c145698d357daa1a0390090cd8af90e90b7aa05bee507c41c57a1782326c6ebea014b84324d6d7a586fa173cf3eb11ac27d1d0bc9419;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h9789c9d990cd99481d4ff5b48ccd7265d71beaa3d1b1135dada2fc29a765301a83a16e622b3b3699357512c1876a2057dd778d82ba320d24096dc3bc238828cbd47a4af962648a1e49d0f8ceda56;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h12ac8bc57b81eff4336b7fb3aad87b112de20f544053e6e62e80559ee8d468819519c317839f502d5b4ba8f24fc8933c3c680f13faef7b13c5c2ce39a485cd71c2f4fd8352d52163ad00a2ccfda4e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1deee99a0ff001906eee5e9b18e053a3b8b8d82039c446229a93180d183ad7898e7bd3ef64feec26b4c1467ec71c77b509aa7a21870cd8957732bad009c706e95b27b6d4064f4f7bedf1b62ccb155;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1873b190283893e84f97bb8aaced81dfbda76458de25b28709b3b640f1aa7e4f05c99aa52ca2767f67c67ce10e281092ad3c7fe08631aa829a77bd7634ad282f9130bd7cfba9e2f2cf0c0ee140e08;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h7ed61a2c5f2a4a33eb838cb864b4a24dd8d37a27b0a7cee4e95deadfae1f2b1d608234d626582aaafc2f30e044b5b6def19c3cc81d95bc4f040589e213aa546c3ea70f7e47486c54933d1041f36a;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hddf7d9e9ba08b7b07166b81149f152c5c79ba372902addbcb5c948741dc5b5803239dd5770ed3b12b311bc678f6ec2cb2f8696f524260e08c672c772dddd3f79a22df5a900931f09c8c2e50db06d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10d89155f57c32c5d28f19d1d4098e951d5a4aa3790bb0e98e764ad8f6a8f65dcbb0ac14b9ad1a134fd4b65c8454a502e79e342a47241589da55c44fb61157fdf363541d40b14655efa3d89cd774e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h3ff1cfe7d99ffb770c23784170c3e1f30c839a4a4bf5a7b5cf6520beef8266458e89c5c7c3fa9ff63c3e8b52303cffee0c50114633246a3fad31bf08b46203b897f659a009998d021eea92f43fa8;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ed27fa51b16292fb8af18c2913475edbf93452b388f10c530a6425986ca1678906c7a22210e266d7f0f8b699d0bb8ae860ef60a1ea54a1b7fe93a51623758fcba7db40fc39f42828883378c7f5d4;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1de667b43aba39afc72e3a7ef2759bb78e58e8988ae394a5abfcccd69846d0f9b2b5b8bdb10ff18d8b0f70887ea7120c8d67694675467a11c2d78a3f8f3aecd5c22c5bcf5c8177a03e8acaaafca00;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h41710222b8779b435c0a6ad5967eab740e112b10acdba966b23782c4e4bbcff1fdbf4af9b56d8e006dbd0782b5b74cc9d3395965a641ea3a5fe7bdd73241bbba07cd2517a966fe9edceefbc5a45f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16613069c680ffd658d72ea654a62b37a2e5038fddab473cbad5e8cfe9229a098ed528dd1d130b36aa29c0a209d923b06e303d11df6588ab2e8f55a821553b645465a4ecb5cb754a88d642c7dbdc2;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h5b0a2f8c5190c7ba01267285752b2e8f155ba5af4c13572a37dc457e135c1355703865bc8035b3f1c151b2b8e0e7372b35cae3fc54118c818ae093cf9803f0552ef54b5b2c65b53276f9ba76b7dc;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h19684f0698cf36fe450acb9c2f4a03cd30c543d927af061ee86e1f4dd1896bb97a892226ea9bbc85410e24391472760739d466c778b391994c62051926b19027235017127eb6f3933d0e22b9b9de0;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h12da4b76f149ae2c43fba7115562ac5b2692d33b2fde9f342614e25f7d414b4b6deb2e5ab4213c063e9612d9cb6f04d341d3cb43965bd5eb846018fb8bedf84c7bf18dade131e911b262b66d79a45;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc639b23fb221e2f2770ab3c588cb7c87c513eadc738540bd6535124e8ea73f0f65047b0d6c321cc65cd7b2a6515feba817b40378b3de6afee75b5ac610ea6f1276120a25dc5a47e4dd752c55f244;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ee44f816a04e410e265c4f06214fb7e56c595f900cb5dc2b42cad8870ea85fe3bfa17cfe516434a7606a84901b364fd52c616b4e5250895b1bc86b340efa1a29435ab3ab12faf7557169fc1a6185;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h8931eca89e6c9cbf25d5c7595657a9ff40f2eaf1df7a9c56625615a934f49dbdce75a61abb75585f6907e1e1758eaecb5cfbaee84611c76f714b0a40a6c1141f1c32dcfcd673be278142e14a0dbb;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd8d379fe607957476aba4aacde81be65913513d5ff72ee0aa15d795f3d051297a3ce3369da939ea98e8be5b00d71dc58ff63f6672ba058aacd7cc118665634e18c6eaf762008bfd973734df36de6;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f1619a3fe8792dcc7bd445854923da6b69594eb999bd275ef8db03742b7003f3b8cbe6dd3402f844ce62b7f3ff9ac6d2de2db3176141097889b1fb9a6851d3e22d0af562ad53c851ccaa8759580e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h98ceb2a3b2352137c85565987871781bb8238aa1fca2f53d6f6c13e735ae301151dac2ceffbb356352e6b1934486f338effbb85d9ae78cc1926e97c76a9e5e468b0229d43e4665862f37b1201579;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1378463215ef231e742e4cb58856ec60cb407849b5698620e30647b00648d8888ca60a517a74c96edc19e6731fb43efbecfb7993665c43c5af5552c9049d3ac4caa59b59eaa40d37e862f4fc7634b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1cf461660ff37ae8fffc2d5ea5e343c5e0f93b64c48c269ea7e35ac424faf632d3d88f5a1fce40c955bcf04082ea850846f72f2746bedebea5326025c4f93cde81f74ed045ea8abde52809799e68a;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb1d98e1dc3adc7e4fcaeae0e01809aa5dc27aa852a9d38fac7fb3d477abeb3e7182980b43abf47043d13c2b72768a6719edd08737125bb91e6400ecb49a03b12802460c2d780be98d844276dd8e4;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h187b853e557e9f506d7473e12f26f2e51b8c922344ec575f20e27376743bac9bdb71059785890a6cea760eaf050db07289dafc88d806c220b6c7df00d50a680ab68ba284965ca95da5e62964ff82a;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h9429a06b9da5d7968fc79533de53f6e4361a1a92725842557e12a464dca2ec4c84130f5d581528111034d3839feb0d7d8e0128a75ac717c0374231fb210cc37c53748ac57f18a23aae6b5932054d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ebb949c3a8cf833bd61503eb28318746909412050dca1c539b6c652fc20b5af9dbc79e932a3c160771b4e8d8c73eefc39e79e46126043ee2359bbef8e8c0445c718f0e721108144f8b2e907d2d69;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1388bd781ac2e68a614713157482d4ec7258fdcf2b513462c0c09ba6cd8520269eecd8ce45f4ce4e984d31c572b32eecdff37f0f70dd9ebfdacf8aaf9e79aab989c44a6a26cb10583cd01a422d512;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hbf3fe59247dca6a44527783b14074a1ecda96335c95047f2f76c5fc6acf12a6cff563f4a5384a3dd15815f8cbe08194cfcf8c22af5d4d54c8c0f340b553393c68f1a7b89321510fbffd77604e512;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h8b4452c4dc3493a6952c049954d5a03c02c285cfea91e370463e7e0cb363f379a06d550d9268f3e2aa59c889d1be1a6a2b19c8634cb64cda9e203d9747938f3c59bf16db4f6da7e0630416e50b3e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf1aaadd4bd4a91ea0b4aebc57690f5673332338001cc11539e404801c44a4122092821606d1fb30e9394dc84ebb6e07fcc423cf3a95dcf6ae679f656c6db564e4b8262c1c54e2aff21d500c4d903;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h227f97c3ac76518bd02f6f702b8bc3215576ed898cb55a8569373ddbb27bbfbdb86b71e9178eb14c57d0fea6c09608099d45be7dd2e10b7750e45fbe1c6fdf2a97ca85579f19b848c0b0de4c2c47;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h69bc5021bdb064acd6bceebbdaac82c3d25d56e041c7a4e9938c89962321eaa45af53ebd71371b0e448aa57d2f67a53caf4cbf8b8d7e1d0239ef3f576ea8120b3ed11b6e93bae7976ad09298b25e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e951517a62556b282e59bc8a2c45645fd277bf3afadaefcbaad23c87ff5e3eddbcb69f042af6d303b35ae1fcc757bd82f2f224c248c1250a2159b87ada8a2e0da3e0312a220e5f2ac4ed0aeb590;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb393c52ce042cf8673df06bec59b9919dacff8e76e4878720d4b9cc0bf8128197e6c4a05a553f10dc6b296ffcf365f002c899190d25cddcb21b20f129f33f31be59d2786f176863363d28a6a6ba8;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1608dc2b60db0fd9c1ad953f7362216f2e51a9e9ce8290b04013bbfd550c8c19aa497a284acc918d40e438436f6e27e5415949585d74eff45e85e3cb45f62f43783bdafae0cab87103d3d9aa1d3c2;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1172410745c1347da43d38e92060f5db47a1c1cf11de038aec5e5a57cbc031f4f99bdda69b3f3c5c798c719e604bfcb949dbdd9111b942c27a8727a5ae13414d5798d846c69cb91f2ecbdcd4c2505;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1259b4a9feaaff301051e4f80d896c5c158e8716fdb9daf62af4c2beb2c7886e16b5662292c2111fcaad7837b0e6ad0d9c1929128a5b45bc1479e09086027e7c9ba40fb95dffe75cb04fe4a579bd4;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h11c96c61a72c54d0cd1d8485bddb9d28122f8f418c539eb17433dbb64aca6fe0db4f94d97a505b2c11e8d4ea2adff2408b0f2521596a52ed7d2999f544c9aabf8542da8d29ce717c7b526a3f96922;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a0a1dcef7bdab2eae79d14c2686da0f78608ce1efbb69192ea9f9f89a13a72222f51c469a34ca931d0cb1dcbefb7edd8b15d271676d2b9747a720ac18420f641db0b55dc63650897c696df70f4b8;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h5ed98c86b922689626af1e3306e0c13ec8859dbee1e8117b2bbfe6be9111c81896c6b4a91b3e260fd7784e0770ab158ca9fcde301e7239c6edfd7e07ec076424be89de3052bacdff88667d741b9e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h166761bf10103d252d208a8ad3200d58af8821addec93947bacc8b25029ab0833d52cd810269959b8b3cbb45f014265645a218dd928c09240ec7dec649d2004a7e0246f106760894abe85b576fbfa;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h62c4725a336cc96a10f262a3bb5f32da4f14e675ac2822b202aee9a858f761c8a15313630a850eca37b691eed488fe40013ec4f174628424c75f67d781e73fed4f80ef9824777200991076d419f9;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a805020287d19f4f12bc6ab5adb77db7fe81545bfd831f007763177186b23c0af987c5588a3ce9d628b25af09cd8de81745c392fa09f459e7e6e2a03f70cba2a381e241f60166323ec1945f26e6c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h19870f91293cdb5be25b026a28847f61729ce6db8ec5ccd65b1adc13a5a759d16b4203f851611fbfd2d7c64ac9bed88f8480dfcf496aab130f9bc31de2fbd1c5602724c19e323356fc88f35440579;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc4a7f51b4d49fde1c5f9ba55ba53aa7a7c36d71ca84ed9fc9f5b2902d8db64a6f523162e20524c1684e5ac1805766f3f773904785e907fb5b90c300177831b233eccb951e63d97aca2117c71d710;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h14958f81d257c6dd112034c0031dba0b7c00e5eefd6fc5b2d5352850cb45a06705694e22124988ca433d9b47ff76913a36dc50209410988d3302748057c925909d6dfd2b856959f8d52b514d80da8;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc4685d3452ebed6f565d1a114b3f03ad73100e10119560a2b3836ae68b6f34bb276086d9925a073cf9feb7d925426be68787c74e40bf7729d91d3b877710c86a300848323d7fcbd0dd577cfb07e0;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h4eeb64c54ef38e5a4707339962a9d5379588826409ce541c86244625de97c1f4f80245bb7323b6f071f59be11dd12825a0bb0d018f44a1dd4e737c6ccfcf4899d8cf6a944361d2926f5287b8dcd6;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f8ea7ccf2671012d3cbd27ce65424d492f881be1e5876c081c83345a0db258ba4f25c358decc16624373047de8dc1b6fa121eeebf4738b5d22a7a9ba8db0ec254de7adbf92b02b0dbfa75caaff7b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1989fef9b64a84850804b8b4df6e0d8022e55796617617dac5fc6c515b3f67d96c1531e8b3682d43ca64bb4cf2f6331d0795392c62b43b721b4992cc1be46df7b0cdd5ddcea78f7fe5e6bae0d4cf8;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d942780401c8d1ab3870fff14b4b045dbef54a9c40d2fb23092b8cda896c4338f870fd1c043fe2bb6deb04ecde9edca7ff4845bf1f7f49776815794603f3ea591a9db0a038d9083deece2cd60e7e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e7821ea7c0eea5d998d708fae9b5e57e5737a863e45baeb10e02fdbaadfe60e496bed2b1614c6ea5a4dcb1f910e49ea06956617faebfdc99366d697aa62e0441e8e6f5adba8e814b1cd0699cc63f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h109fdc552813fc84ee05dbd350fd82176a172e10daf217b738f94a959188ab35f4428e92d7b6d0d8f08b617319d12dec734aa619d8d90bb1759edd495776edbcf026af5d88adb162bbf03e509d6cd;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1645862aa4faa219462302f405bde9ec82f1513e0b98aa2541cb45f68630344bae4d4a3f81f787a8d5f12b77c2d1f232637e2bcea42e0548c36a80888454deba37cb78b3cac5f81711fcac5ce9a8a;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h995257ab7ef280b16a70baca83889419a3c90a49c3d95cf796f726f5f785a7faf0ffb3d013e9d8f557a4d1e9e1673977b6fc8202722f59fc00b92a9b56b890972bc329b85497b7722ff732191429;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha9137e4732631408878feb651279b0c25b920ddeeee4c1650a745497d72c5c01fc624e5cfd989fd36dbe6e493a5a3c2ab2277aad19261d8a370d9bf7c73cb41fb573f7c5f867f8b3597b4ada70ba;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf890c9a335a738e70c4aab883c09e89f2b39923ffb583f4ab62015b37f2f10143e7db580683b1bf34db084665bd6ea7e6fd30972e13c52b31eda21a66949dde70178d4fed59edd3a36aff9581544;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h2707520a3098602b3baf2490cd41fbb1dfed924c90a175cc168edb5167088946990f36d1bfebeebfe57d3241a6df8b5c8052e5101b32008571e129f27cae86805e8cd33220209ea00ea44c2b9cbc;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc7e5e0bdffdef68dfeac458814d9399cb4254dd608443f2f506a49291f1e1ebc2d9234aeaa3832bc6f44a041570ddc1f50f4d973720fd8097650eafe0b411ebde07bd783c4f2ce92a4863bd5082c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h132d0e299bcc2e59f3da2e9919a63243c2df3799d86813f589e618fdd5b528bfe0e0c3af497f8017454f6c0bb7c4e1b5a00e2b3ee1e65a9dedfae313ab593e33e539a174b98721443cf2d6e53cc10;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h2685becc986e7dee007e18237cd3a00f44b5eab6fd822e6b0922d81fcb82a9ac97984ce582fa7bcd390fa1f618ee3158f19c519b41d6927f3270d43664e00f20fe57b1d84f8e50d4418f24853c8c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha91fb4732458982c1d24d6d597d1db052afdb74539631a00038a692d77d52918eb0b9394847e9052702ce8ec7bb7edc1b3497732c43f3de40040742681022cbf041866b38ef34dc1da332693f356;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h8ecfb4796f1f313755fee586048a780c5ded19196e54194459f28042c6f5121780e687c79910617cecd970b970449870b4521762f925868b1390bfe6281eb10014724763fd086c94ed01016266be;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h28a58731f7a43b33aa335cc59840840baa85579fe04a0c97ecd3bf16003c9077905a15629441c47263980e2c0e0eac894c69a3b551bb5577755d8c2449888e924570156beda03078a016b27517c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1537bf65c47ebbf2329b55d563d9f5cb3ca25985608262ad37dedeb608035268f5fec8ac4a4442a060c267bc050b7ed10e99818e56464869d07748814b43e49046961954333dd449b1801d84d7049;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ec6a8cd2d0d7a5a56977f2b8dfc1c0ba68be2db0b25a8ef1abcc9d1a381343247a840f8e717603656eacb8a091a92ddf66f0d5c57c85ec2ee326017747702a467e5f330656ee87de0521c41947b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1585d2a03cb7ff48b92ec3a4a9136ae50b865d3210d7f65be8c0122140d460c604f605961e5a4e8bd5b6028d90519a1a921e312b6d33aa1374609de6c69735b327c5c40093dcb66c4c1e594999ec3;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h7f5c7c85d8f1c292cda99f29f17e728f9ce52282f7b92ad3145467c264ee821c400a8bff7504ae86951cd8736d189f70037339baa631b09c85975242e2b309dcd0ddd12d4c790cf232c37453030;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h419688041fcf45ab9da66342d7af9df8b55101e05efe568214458e7dc725c92b17ff1453024014781f850bd4c0d1fdfce93d429f4cf0dfb6950d0eb3177b0a5716279b513f4f9ab48eb6b0c66d0;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h9a00b435ba4a8ae750a9a457985f7c2dc0afd2ca4876afaf7de81a5e5b161bf52ae7a377eee5175bc63b3ec15a00edc7ad0ba66e00d39021b801b34a037aa8a6503d9012192a5d9b52d5ac1e5c34;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f03df34e71e9f473de72424b910080774872257cd05d3f1ef5d35d7547780785d96a3b1efdbde04cbef9116c69a8c5055922f0736523a2ffe8382f46f138103aeddb8f3fe9bd0785e80bda7128c8;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h19c2d2ce114112358c923ab832ab028ad110906447060046c5502a60cf2620e78bd92af9476a3cf7edc90954709bb166dcb97af8eaf1b2462896d0a5959b52b407da9288c257a3b41779091664f35;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h81171ecc33000ac055d4c8a5f4897ff6e0c9415a41d5861ad047bcc5d668611fa325396cbf3b632e48c6fcee3de81266159b2774cdb2277b657826b6fed37fa8d147cb872998f66b3b1db8b3fb44;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e0919b84cf5e2a5538dc02daca769b9fc271bd59f5a3bca3ee73a2ea64727f941a4270884ac8a9f4aee3920d7905ec968cd7cd17b494233ccd30d6f7ee0cbfb94afd0839eb9ed4c956f3178c5a14;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1134eb5b921042690235581df5ddb9b455eafefe1a8b54593e1ffa853a061fddc62cfa15f162096065ea1d2910f2ef582f7ab67b5855b9edcd88c8743c9800d79ca2b688d0f5a8f69529c73cc59a6;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hebb6ad9c7d1f5e7841918ec2116019b0c817e5dbbd5545b0c4f5723b539a56e24e2203f0ed8acbf23eccf7639bf07f28ae7d4396da2475be101fba32a5847b18b12bc5b25c5df6e910c69a19ebfa;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b9037f79c939d689c55b13ca4699a8f2708cef1e2150f2ce8f82f2231f454f51594e17ffa364f77ff4173e6b5bc91b82e7fde8483df3998c9e337c51509bea3b77a7460d132b8fc1ef9e434bac3;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h6d6dbd310df0dd8b31eb25325ff40cb1dbcd0614635f69adabff88a21573a816bb95b18d1ee55c35e1b09f6135d74ef4d10ee7906f27a29dcc793af661bae1ff03f7feea54280988c11e5c171408;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10464a75d67bc5ed3b626594efedb0176041153229246aacb97d5f8d6c2c6121606d32e5b8889a9fc2dbea933e07f37647e8bf954edd5bf1bb929d964bcb5f3eb51cee1f9199741b0ba7a3097e3b7;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h499a8a95e28f45b336a14a9a73f7348ec1b7abe914dadfe990bb186b1f846612e1c5ae6fd20290753101dce86f021505ca1c2f1d55bf00653c8bc6c8391205c03c5a37fe1e71f4d7335c6fdec397;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h7ce734f951e49ed74f63e76b8d286cd5ca2ff044c8b919f457088b58bc5fadfa28638c6544b438c0cc09384f6b4c962f7b9b88acb4e53fbf8d76df4844b3165d0eaecb126f6bee04699e66cdf88c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h15794932cf44d0a1a59312ed61784babeaa5ecdeed60820dc50b1f3239830d5d2a6d824b74db671ab6a2d84e8c5e5b941e47f7fe3eb737c293cbe834796bab982c5e518689f21d5411e04a882177d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h5cf6f345b8fc87e1ed3a850a50a2a47913d704ff0bf872d1cb909dea6d467840c8d7adfcacc0463c251d5368fd797d89120b1db634b63ed95d5b3b89d173aa646ae662e67245f7dd2ffa0569c491;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1150ce13fe02a332c9f3eccd9350c14e44802cfc335d4de0f298ace852ab7e2222eecd7cab101305bc7b6242bc400516e58bd65bfc4f43509d2caa6fb418e061520f89b05a3c55552064fa7c444de;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h11be8e6ad8b1ea052a6428586d902e00eced6602cc4aecf4db6d5f0a16a7292578d20b31b65916ad7eeb1aadd21e01c50c9bd063e0491f844920a3d0ee547899d033af40ef2958c97da3a37ced582;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h282b84cf953f01522d8a64805490945f19343d278c509d213d0b93ed157ecd69c34439a5994ed28f40389ec13359bbb23fb61400d799afc72a66725f48aed18a548626b5f5e7ea1794dc0f888b43;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1bb14a6b64b622d6a883303497be0f837079a89318c1e0caa54c8c5c04a335cd01963a3c48547b73cb6680ca0e737de95bc65410518dcc4463f4766f65d554a66b05d9155a44d5a2633c152cf1acc;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf07a9fd9064c5f057e7ee58ba2cdb97b56c20479c4eca6ddccb3c9185b9aa33a1dd7c95a3d024096cc65738fcbfe775583de4403fbd29a0c590ca8a01135f9df79342431076a5e4c93fe6981a1d3;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h161c165d8b5ed1985d0cf24a6594980782c802aca81a773ddb872a58578cc55f3ace53ae931613bdb64ed18c9b1b793ed0ed9a6fe90e41028f7cbfedb193fc75efd3785463ef8127368c2b68ff777;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1434768c2b10730a0b54575fda85fdf9dff9dd0f3b1860f8dc041aeebe06e946b005d369ddecaad09737c335ccaf72e2b72639c44359dcc2d7ba6d5e79265d5ff9437ad127dd1335ec923cde18a8a;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h44c2707131514571c20671453d712dfd435fcc18d5dfe4bdcc7f4f85fd42245e0335f71a0fb1b9215da8d64c16e59775f2485d06a8eea602be39982837bef4632742624d9d9498463a02ab88bb94;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h178f5e646188de8e0292304aaa2ef1f044c68dd197b4c74ce187c0ef1d5fb5303ba8280dc9e3852ed14c73561f26645ccc4e88bd808db3a9bc5d71b49723e87bdc70f6920da0aaffc293dcad8c297;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h11a92239324e736ec793d0f48eef6613ab250d3ce33d5a23a5b26cfe8b7184ad75aece4332d09256018be3c5cbba298d24f97c2a7be92eb2092be8b61390c31bf32e1b4f67776cad5cf5787916087;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h606a51da52508628a2889a9308e8481fed11c0dfb85d0c3aa9a6408d85cc8453a67de70073a166c078c13ffa34e427cf4355a190fc6e0aef0e7068ff34f9a8af65496d4df4948f02af042d2a2bd8;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h18aca56e701d9f6abe25a31cab8b1ac9d461e68557d9f3b2b8992ba0ba713b441becaf566c2ca5d8922a531d89abde2a60010091713831ebae16192939b73f74c736e1d7952079602ed2b6458ffe0;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h9ceacd5a5de900ae0b909ad78a7ccf2608f144a44e924ea60a1e7955899e0f010cac4fc1a1d4b968064cab03e29a426fc0294e1a8fcf8e9b92c00ca550451623c6a1b777138130efc005f7a94c43;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h106d50eab65a77c635b65b4cdd6ede309c2e44e88262bb0ed863b0a8550cbfb8db9e3e0520bb2591d26a74585bb15d52075a36dea4a6048685ea3226e5b1d6e9b8c96c92e1f219def7159b503916b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h6788f1cef02d7cca1c4169cfcd3f1ab07156914e7d918f5600fb4b6a5b9e67684d86c8496c538c2c9433b17dd9a085db4ce4527efe79d3272da0ed785bb528f62242e501f29447c17cdf9cfd263b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd39ce28d6cb9b601118ec3b39b8680de38749c05d04249a10b4ab481e533319eaf35903727c938f3a4f7e6f80c3e3ed37d3753af3cd7e24ea919702b5c354468ea6a1e6ab447f3e5e601c6747161;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h27c5215db87eea4555df71fc385fe532078a21fdc885eac8911604272d743a788bc53583f6c624f647badb66916fbc16368d4c4f95786a3aeaf42a8671bd76365bc1ce82420d7a5864c5fad07eb6;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h13508e86d1b19840c9d16554d1aaa7c94d317c0837ec5b9c02b302acc1f98d3dee816563ccf0496fb76d8d7c10f8dab71fdc8e80c44b7340087736bef85fbeb9900bb31eb37ba1cf634e446b25c58;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h447ef44378a83e6d6808f84594bf23272e16e943b96993374181109838c6d5e43ba3f0dea989da4e37814b1880900c719f727e73a94b4320fff992595f2be8c8d0aabbe1a77d435af9ead0b38699;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h6ad78abda5fdede2346b6d5920f2fedc5511ff7a3560e7db903ff0e310df820d15781fbb44b3d5313921fc4dbebd6a762dd42c4c82e7671f54daa4588cf339a7a034ef332d249af7012951547dc2;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb8243ee887498c2260f399fbfde51406a924d3a2dd6c132d41991f2873735ab2a4cc2ae2e2f7534f36b49de2f01cc08be3fee885d420205f1ad91f6c805911c7a611fec05a8e6af67ee88029e17c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1452a5f819b746ce86db2c22542a8f2e0ff2c4d3f0540b3dbb2e74dae6c6c66d5b9c587f6077f5b500e5570c951deecf4ed3ea9e86c7c0c74335a0d9ffdd6dd6a5715f925db2380148232ca5cd66d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1776b8a88ced372773f606a731fc930e542fbddf71355e706f710f0635ee56b06e227132c04c46596b5dc5fd3dd537171cc79d374b27533de2e331cbbb81c4c25fcba14b7ede3a6702ce88ad03dd6;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb19916b0ac730926ceba4bb5e8de0dec1175eb3d89064dfa2dcbdbccfd61f958d3e7026c54465c41d3f88478777650d90b3448cc568d633cd778eb1b07e7850ba18e44a9ec801402bff26ae1b4e1;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c2ec007e72061045bdc4aa3e61e481b91e8d33f0244827cbd84ccb6f792ddb033981719dc2339189a2a87082824b7b77aa786e21c260e2b049ae7a71f5c434d43ae4fc12c4b64080189d504675b1;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b02b253c9b65bf9a806c81138d0cd945812ee4b0a834ca56e426b04b5cd65949d86a4e54bfe87a57b0b972d7d16cfbd7085779b61f7914c7efa0e9ce76172461f98edbcd9d072f2c771ef5421426;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h169f000e0b005bd0af345111b8cb6d7e9cea5fa0c4cef2253ff6b9dd61b1b4de434cf8a34f0c14f9eeed2149fbe41834464e54eb3244d8ed9fad7d095d92122606191009965b7876369e19eaa452f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he73fca53e3627807dffadfd5e8f66e00b656e8358fb2eeeb948dacb8761ae1acdd97f1af39f17f88f0cbb99707c13b67cf1cfddbb25aba397cf69face8bfe644054bfedb95ea2de0ec2174ef091c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hdbe5dc3509cf78c46e5c98902b9d1c388e60e70f2b2e76105ef97f2d5be0af48cf02f37e6c3199355f57aa61ce695d61be0de6e119bd130f7858014b29b16d930aface38ed363bb46dca10ba5581;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h19982db7a32c705990b93e344ed618956b4f4a9fa305587f140e9ff8f35f1b05f6bf63a05e2855c66a6e441fd82c8bba6d826dc33a1d93eea6cbed95f6781d395302dc845d41835c2c26e35cd3906;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c70e49ea63925b39d1c8202021cd15e9aaf60caa43b86d6da2834ffcdc142aa633fa6f7b908ba3e491573c520a38741fbbf1036089b607a64b5940053131a4c039a1de6c9f367d66c7b9b7ba1a77;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h125aafbf598d5b643230ed65f6fcb659c749dbb601f07316f938e02e5d2ddddcfcfe0edb6e3f236a5f0f9c1b5cf73fbe8f084cbbdfb2ae97d6adfc3cb411b5f63616b97fa4dfa5559810686678c60;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h15a41185c134eceaa556fc16dc70a6bd2bdb7de1d462f2031491156e56e68a97ee0e6b040c07c141f9a21ec6601b260995e739e28f92f748ded74c4f1b0d7f8058bff8debdb0388ffe7e590d2c278;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h128d0cbb2fe553738a7cd71ffd574d9eb5ae698644b0bb8db235f27eaf152e66329de64577c207d5637f1f6e7e0dbe763f94eda226e9182d42efc9e2f030cb0ce170831686c27e8a86d3bbc2cb511;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h2ac0c527d449da1591071c3eecbd8424fbf2b7c981def65eb611493e48dc219ff0fb614ec9248aeb46ee24e2e92c2806df4d1819c016c1349339373a4103ec7bbb632a7a743a81653e7dc3540645;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf5aa5e37007004021ac6b7b889868c83055698d6f77a18e00e5995039dbd7397b9576a504488c50a04e1bd9f2c2b458aa2a330e0bb16f68d700d5c56312e6048b16f621ceb4bf34619338e3a64a3;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10cc1e38524789eb0812f97a2a10bdffbd44d736f1681432b45bdfccb580dd7ac8cefcfb957f14d50d8f98e2ffd01ae9c8127f90c4fc38fc441d56757e5ea3599a9ddf6e9f341093b148a2c54ed57;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h101a296bad9f7b56f8a4a0661c2c91ba1a7b5e731eec305b6fb6943ff4c7f791b6510ea7907ec3bc0913ec4328cbf32a1870018b7acb2c300eb1d68d974a2534273e83735edb3d8902e0f8688e547;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b1f04df757899f03d93be6c92056e735f5ee9456458427f6ae55608c842069cd9878040f04e1941b9b68e13dddc5798d76b3f4e859545a336013d08c49d0c231fc7cd4294fa07b7d378de33b31d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd6c1e7e1a324af2365c28f566b098b083007f73d654c162988c18920dd2215e90e327a0f8a0e71ed3198aff9c85e1a81e2ccf7f0d394bee57c008ebe292a6f937374c696f8dcec52c2545927274c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b138d8e464d7eab310c47edc917225fcad6a522391ed2f72a74b170e84df2615c1910c57f97c1aca0d9b36f67ace2500d50acb3499612c9f6e380cef4c9eb702800a9a7cb8566fbe708c33f190be;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ba00d1a7124928a1894753421502969bd0299892989391b9ef9c3b58a1587fba1c45d4a969920936780a8813d83b740c9c096aac7f96f915aaac121987c77456f60aa6d827b38e0604ebdfd2236a;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hbadd1fbf7f93afc6fc492a502d2ddaa0e1e48230a9d51574581403a597332fedcbbdfd6e5927101ff8149e10fd341025b5f4ed3339000d31701947cad789c1efedec941e8843c5e558e43db8f6d9;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1af4220a0ec0ae0ae7c02d5338d975107cd7ce513ed9fa627202f90ac55d5b16c811e0fb95d062110050f5bea418786baa527e31d2d0055dc4f5e5fd42a524ffbe5e518efbc5ddfa9dd42a832743f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c5bd13a855beb73edebaa5e36fc4c60fdc65a6cba4b344e17f6f79f649eb6843389014ad265b4dcc382244ecf6601b423dafe71c81188b4cfb7ea0e82802e642e0fe09bdd73420fa49e987229ef5;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f1678c2b1217be2d35707b447245aba37e6c775820fc6230cc6a0ee87ba9105804078d1e1814ecc22abae88e09d55e15760641711c405bc42ddd203cbaaded7fb27a8ff77ea18435fa990ab92645;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf684275ac203398fc2edf1accf9b1d52a2f773a4db8b89fa56b4764ea43ee9aa825a174e9a6f8db19c2bf2e874143e95d70ad5e5023dbff63e4f32bfabdd5170fb8e55787a66ca2796721ba487fb;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h140ed051620b81d6b6953de226a11b8e88938b2dbdcfd69d15a0fb189d6418eed1929ee5908922827bcece9efff12af22e60a1ed749e39a5fb0dd4bf944f18b1a084a3f926dd24f2186a69d2d0f0;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h959310295c39cb6f8fb05e945f1a8d901aab46b91c86489915e3b5c39a37d3d04565d95e151c338f3a06c3cfbcf7720f07fbeacfdde3de1accbcd9c9eb215710e1c980c9c7093a11a19136081db8;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1135521c07e27e29178a6a7aaab346d74d3dc9a724d380999ca8f84c6578bd814f3d1854e637e5d5f82d7e9af454352ca5f2c213067e5313fd11a8f17f2ac45256fa6180df96de4a60328860c946c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc05364ccfe0b8df3e5f29320b329ed36494b728360a06e8eb2a2802705c1fcee6ddafc78b3baedbde1e2be3f4d6700f86bf0da31a2628a7c66b37cc821efe1ee60898ba7a8f9a206a0cf56a69119;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h362d4c75f0c75fa679395b94ef023f7d9f6e25db4ee099d80e01a578c7d5783d9baf97656ed5f9401a42ff9658437fe24830db10dbb55864e70e981df443e67c362b83b753cd3c5ed59141666e79;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hbf6c6875aef8e8dd5214222e5bd38811f7c6c70a53b256b8001ab9c248495ac8f1c95ef550bcc4b5e15f23434d57b3134c4b5e514e1333470a79a1a794d3ee0bee7d7fa1e966059285d70dc16db0;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16c52fb8c424d1be7ea30097dcb79a3472907aa81716711fcc4b9364eb68e4bf3f78bb2ff72abc03754da4fead0b1fafe9a457a4fe908c42f6a2142b0ffb0da31fd2b31a115ddc94826246b2213b9;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1505092d4aa1faf9c09d3453fe9fc0a172504609d12b4b0460a0343a179d5107a661a7b3a9e4b10719e1e5e1803457c460427977ba639e6b912cbd28f23f79164a3d6137a556a3ddd57b28baf3f33;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1834b786e07dab92f9cadd44001c7526746c28b6df168aec18e664aa9c5061f1c1551da44b7dc6bf0704ecc7d7151b4db3b9a848b6ebdf57390fee36dc11014279a38a6bafd7bb36a38877cc323ee;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h15cf7057644585c7857509fc89bdb722322419be4cb8b81bb7b957395724ff9152ba642bf502cd7a46625fec76803d01b8681389cae33dfabbc6c8fcd4c28dd901b8ff15c3a15dcc2655d1b8152a4;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb4ee2c942963c61ee22d4f426016f1f5059cb5357be1de4b6145c7509ed69f88de6f0eacf68d22a4877f110e61ea8572e2ef7e7fdf652e279061ce83577728fff3d3e67a7beca06a95b751d9c35d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h15355125ef9c2f7841a3de151eae641972152ca0843dc13c1386d18b39337a9445c9d444031814c636599da9112074441c92a57b493627698b1bf7d4e5bd09bb3593fc2618fd17bf76c3b46b567e7;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c494c43443e608a18382044057887b6c320a79fc7ff8c72702289a1a682e0a6f98227ed6f8696838f1ad74493e1bc47604aff447973dbbb80d641cfaa6860fef147c78bc1bbb6ff16d1c2c20b902;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h66060208689a0dd840190e4b7f6a7a52b00026b1337ed52488baba15a715875a809553d8b41f253212ca15e9b0012e87389aa8a80e9313c074808603b4d3ecf1282e301a421bdbb6ae77113cb48b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h139a740388346a11957a68e10a465dad9e4ce20c1ec378d75fbb649a1c9afe31d97f284fafc0b6e5514636011dc44ff42541d1e3169e63afbad2a5bb8111d690f5686c9f98e9e7160d67bb1ff8295;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h109c4c51ed50ec9294b904f635d8181de47de36d8b1325098b82400fd94891719e291e469d782cc09fd2dfac8ce83e3471cce7c3fe055b0f77ce6fd3b7b6eea34cb3199ce69f193f6c5c5f7950;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h18fadb52c75f5aa6c0f75433adf60e1bcfdc57375f68868aa31469b7b35153622aa30a9159f86646acde0afd979809ce066b0df92c3cdcb6bd6f486e75cc8b40b2f076d1004afa91594f8eac6798f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1303e6777c1a0345954ecb2e289a00a9cafd9e7d68d0dc02a729d5b0276a73fbc627e389a6c0f5ac9ec5dc3884d5aec8589bfc8c283e81f0b60be4f806a90e77376fd7743de36a4ed9623f55f8613;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf0c7ca57a523dcbe815333a837dcae2dd866a41aa6b29f81f39137a99731fe9864686187c58ac32faa950ed837cac9bc96ab0b075f7dfbea42a32bafc96a0e1bc46f29e4ed73321438bc7034017f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h7d9a3a882ad99e74676e39f06e02660734d87d4943de1ed48d5efbc4f36ed85b9bab890f55f3457f0c6ee9ae2131ef165b66f0d06432cd2c5166929260f9e50b99ce7d8b7b6af2475819959661bf;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1fbfd5f74d4d7532aa78cf77b798422c7f31921c2fba9035a46752360c3a222f5bd0afd89277ecf1da4228308a3c2e1f958d252e2dee5dc0d9293abd6266deb822a2c08700b1a3d3d380f52ac382f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h12ecad6eff1cabe851a12520867c78428daba266ed90eac974687a726b91ea8fc262992fcb46542d52909e0b7de2a33cdf103ee6e9bb8a5397890c5f775d8f981bfd5f201cdb2ce1a05e0cdddc68;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1939524101b0b4ccd88adc231ea5c95ece8548e50b4f8da1f6a863f1204ab34db6a7b48caa556654dd8f318c7dc3a5859b1d360aa0af27ab7b9fa72717a08b6e3f6060fc5bf9c382c60a0e8ce1c37;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h18551138f2abeaa83c78824ce08f81c380e7841064cf86fcdb5716d757fcdd15d59a913dc7d6c6e13804209f1dbd807a8af84a55b1195aac0233ae69458a650db656d72103f79771192d360d11859;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1dd6e3d213e47dd47dd46c9e57cb578df0497e4e4ff011a455b612b8512d4ca90735060536dae2873b9fcc161c348e15b0ea9c189b0c7f554593dabf50a85175015198ca80784e04247f454688fe7;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf2e59395e2a86982bddb85cb7b9662258a5f1ba0cc4277c37af55cf0b6e5027b207cf74bf005695757b92e7c28f71007b1fccaa0a09e428a69ef4ba7bf987e66c23ad3968c398c42c24938770c39;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1912d3d44eb62b1ab9ab3ee71a9dc4bba4899a68951e016f4037a1e661f5e2e923bc4e044e961c11e22e08969b8a33c224c27514e6111af9ebbc058337671d40945761d492047052d7643b1ffdfe1;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc94ebbc033d557c1c64335ce6558eed96d19ead53e1cea7330bd0517645a297a9eeb7ef846f2988296f8560583927884d2d9fc1005aa65e4cf7093ed376d42302393675643edede7b005f41182e2;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h108482e1c4cbf54cb71953aad3bbe6ddba817c7e82ce579e7da321f7d8fbada49a2263df1b064a810ec95cdcce912fb7647e088d242b6b81172b72cb9344c34e5f9b966895e242717eff96c1c145c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h5d11130524b99dff8debd4af85ac928636254992af1a9516cfb2a72b26efe7eb00d5ad084b305764a81e793d5c71c1a5e11b4c290194be08483c30050b8e449cb31b3ce237338364ae112db9909f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha31716e6d1dd507b5b5793501c4b933017ace6338b414e8879c65c9d70de676512a959b868367856cbe8d985fe22a465cd47e6061a97f55900a53f9e071f30e09f26cdcd2230577968df57c7fd65;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h819b7405766444b1f8370b90049953e049c17ae04917100d4c4ccfd132b9cd46d2f42d331b6505a22aa5bc044d45f3f383b4f2a093f69057a8d89e96f95288251c4eb6154b564eb759592188f913;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hdf9deef31e0aca055e5e84930cbddf08302acf68293e85d257663fe502307ca979c51f72c0288b2cded99ce63c8068aac1fcc35f2f2e23faa4df1b99ec994befaa665d91553010b355c7d08244f5;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h5fc5d52eade38c88fa7d2780131c96ed160e35a51c3116f7e0d4c1369431a06de723aa04bcb3682b5a978ba7bf7bd48c4b2d994e769f977ec0ff5d8c13cc265d846278051416ed67b1395381ecb3;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h112c91ecdf9274634ba260dbf6a082ba3f53add782562f1fa62553dbd9295464dee3e6eeeef9e126390a8b45a22f1163eb25a1df7aeadb841876c30177d9ec7e9f39466b8b4e1908a0f23a47f66cc;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c885792107f3ddbb8bd59796e704c2a5031f8e900ab336557cb043f9278df8323f29a370565f202395679c71ee2b940a5f0d71f60540bd64abe7827cee24d3ab93fead8a21345d23d9d5eb1658f4;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h19cb2b2d6c8ffb7e0e6a8eed6c342062ec5cdb6ccbb5ecb5c8730d9ad9880d0d9cdf847083d58d9339cb6639e59e8f27e6a311cba15c0de07e713a40f1c4121fb6fb44b6b355556173f1147cc235b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h14e85140505087bac427b84ae578da7de116d36a96eec96da25cbf6f53fac5598a60e618e2d205791a6053fbbf541a8b24c9bf33598673d081ae0c7e8b0c5ff4b0f1ee1e16e3725369a6502b48d44;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h471df7406972ae12baa36fd17472085a909670a48b389198ef1377aef3f06a0fbb83df5444eb290a2c3b077b9846184eb730b17fa8e308d1aa50df1aeaa2e0b2c30378983cfbe91de2c983c42303;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h5f5e116bb0d28585efa2f34a145b4cc196e99456f327fc92ec3423144ead1dc683b808e2218a450d6415369d92e0570d14ecbb8f2b9f9a088be7fe40cf5b1b903f43c38cd29687d6617b3011251e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h595d3605d77d13ed2befb63219522d178c2622cc11b3be2b30e2e86f2d321298c1a6359d012e922f1136e594a185888a35f73d17e5640a269474b68878921d32a7ee1b9af1abb5015a7d2172713;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd9a7879fc1573bccb5ebe5c2e6728b0154e4d3f25c67f12a469330f046afebba336b4a62db51a45e5fc132d7160283bd1b61dc353778949301305a446b5f467a9fa52328163eb9eb5f05d68c23ac;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h8987fe84454e68eb443b6f9a00cfa4268a4a7a2ba476960a9183271ffb9307669d3846d4cd16a2b7482ac9c002a0f402d0c35a3c236da4fb971cdfb7327af37c865afbf10dde168fcd89be267502;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hab76819185264f4eaa5cdb092c4b7bf9a809fc9736c339135367fc40f1085aa8dfeb77152308504237f3a5bf7dc3c47f4914ed589b75c96ddb3456837b91e4b4acce0ac50ebb5570bdf89a2f40a7;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hff4bc2479fe65162c877aeb344825a39333b772c87b7ea37a2a0975dcdc19d806122253c1fc0f58a42df689d375726cb8a0641e4f9454fc0b25af35789f4924e8d88267f27c6d64df957b76697fb;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c6b8c87ecc1a299233bb1b72d9cdb32296c21cca229fee7d3fae95c9e45d87e2aef3f611fbe2aa83a2e0859ea007e6a0785622a7404982da4137cc03627a1b6bfd67ac73c4c9fbf370e2435d04b6;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1735f950c37c4199852ffee432d414ae57a5450ed65c4c454ed96aba87d00dc75a5757d1db81292d9d0b845b48b378df4302ad2600718f5a4521409ff628166b47d4865749449f0fee34801ec4b0a;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf588fbfb83ea9618564146389da26d3095c6c7aa49509374bca553573bb61ba9bf1fd06e5a904306d6538e135edced2003bc819f09e38e089c3198d1cb8951678dd65d46b89d6bc84516009f85a6;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h12b55289d49c6e66c436250dbe136e619729db92f109b9d8562fdf27f98090856aa7269ce9c24eac4edbe54748665a501921773317f847a616e84704fa5f221a18fe533730989b24f3b333c66eb0d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h34931360ed2607fb4c59c5a94318c2210d87eb3c4583fcc1f96ac214a16271ae3551b10acb03f7cbf589588275bcf666e42b29c11186d43af865f3e63e3314b5643c7f7bafadfe693721db436a4d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h17f6f5026be2c9ee4198506e6d77b66214a4359bf4d2c12b0b86ce5b22d732cb38cac8bfe58cefe5791bd844b9777b3834f5b76427ddee4d7d59b42f2dd8176221ee1478155d9501c809a016369fe;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ab4969fad04806bc78247c052fe160521a28a65812a7411132c394b6c89c7ef8e4a32364de8cd41b59123f29091967d68c19f6e0815c4d6f5c05ef81aad90456c02dc6b2e9a4c677b6fcd27f9e82;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d106bc1b529e61ffe72e8cba5bed7d0d4f9b4258c4091b62930ee9f1b00168cb5a457f8b84c766a90fbed23acdd945718fc7bfbb88d43e5ef23cbb7e6ba5c748f1fd46a6d788736206f1502a6abd;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e93e8a26bc64dfbbcc8f76e5e15727b6ab48911542142acbef1ceee49e0b7b238fbb3e88e1b21090c9fb0851dc183a92864402704a4bdfc3ec743ec387689421a8f4cb1fe6ff6100d0f841c90ff5;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h12eea10e37f89e7f47200c9fd7014e0c2d30e23ab13739b6df23a55313146ec391371a56203833dd641cd3fd3e79ccc3b3c9cc5d025a15cb2c869570f6b2207a4769a75298f5c198607994e15d64f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h148ba85aad5ccdef7bad25da2d37a12b76b995916909953d1358194a53fe4d5ccefeb2f738dfff5ced886f6777a1d73374e55a91f94f0c670bb681c44dbfcd036a827d36fd902c6f614dcd002fbdf;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h14ca946ab8d2a3258ad9fcdd0ff61a8cf7cb1258a2a16d5169ce14eb19f08ce4c0a826f00204547936170d4386aff7a5cb85c50b888097ff2570f9c19acb61be5b0d90a9cb7af7418e724d85294b9;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f3505bcf2c2eed521f58e938fbd8395eaea8aaf999284081cd1d864f3fe8bd8a8122a555711c65fcdd71cc4e2d1a6b1f104436f1c22ad14e25a751eeca94189e3095d4285e95c56f8633871578e6;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h183e45f91b672dbb9d4674bc36a73a129c8f225e5d03009b537ccd5a79681f67ec9b1467f7bf416117530f20344a2c673bf6339e5077d7beae03054a220b72877b1fa70654a86132892e93d0ca3a0;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h76dcd871eb45c2b3acd6d09c83a9b6a00188105479132dc045acf831acb695f162af31ec28c056411b3e98a08235543183638677ac9a8937abb68a87d890087b779fa9c88cbdc5c1433aa3c0c2e7;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h523f131903ffcccaea16cfd7a62ba118f85ecfcffd61929e6714eb9302f342ce70cb3b1611de87d618c57f99fca723f94aca9ceb428c29e272018f020a54f0c65b2ae3f6927c5cf4cdf9731e945f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h134532e1e068c926293920c531dc0fb90bc405a25eeffce03fe95df631606c03ee7e2584250ea340aaf73001f9cbac64543e540e83b994ebc0d21846f7bccd7d4e71768ef14a62309c461cb839a67;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h285d2c95c08d9d9148f9864a7bdb0c17d5085381bd37163746d22fba92d58dc48738b49a4906d8891730ca6646434c9816579dc558f3c60a3e35d6a31b0f0f2f3df6e292c2eed50a25e3a2f45beb;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h18fb3d231c5cd9bce44f6472d347623cb30ec981908ee98bcb1ae941523114d5ed27a18cc0d55753bcf480ec5297402ed20eaa1fe82c6133e13dcc964fa01b69fe67bb6b8546394dc1c10ce5fd5b9;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h3de31839ab5016a5e8fde9e05a5480a0aaae4d043fe0f760bf056f5ed77dd2b2ec1f1aa6f7d56660b6d3fd5a8f07c70fd606f426e9d6c93c1e703601b5bb5bed83a4276dfc82da1b83970c2e9826;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hccfdd51f5b928870b026b233900a987535e4efcd35efc4222b7302e44592d920716ab5698f46b65e5815264dea52cbd03e32b8af7c846814661799d79cd63fef66c0039fa3d05cb3fabe699c5644;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1102d7e79318832496e1f908a2c30f4874d8dcf92995b4277888e9d7a58d2f156c698034052d5bb622eadcbd8efd0bc4b314b10cc36d913c9e0317640ae8d1dcdfd9d48ac96b67c561312bf7bedf5;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h149cfb03805c983b29659ea5029f5b0029f74fcc6ae1f889b0b75c094becf24954a2fdf97f8a99034a95f6ee389a41cd90db5a69106a9114855f7f4b6d0e5a83c568e8d59ca9f2dbfdc65b1d77ae5;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16bd8a298dac7cd0b15f7fc3c62546a85d81c502bb71f7aa15965a772441687d4588f8f85c6143972575f6627b2af0446252ea152b58880a44ae1426db26da29b3374677d0418a9e22396c0ce8598;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h9cb40f38872c00343958f3d9f8e06ad76f1814801926fa8ed16177959a8a8cfcce1842bdafbb3e3e8f4ea43323cc82622919f904e862f02c3795c24622ec3af0e89a79cb9bc2a82faa4ca59e7570;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h559e57dc766debbe5d1cd6aa4fb978a91afbcc7db60e293a1ddd2a99c1793d8b98af0b86f8e35a4a4b5b32c1cb209e4e011fc3999de14e98f4a2d5ef7e293602e3da82e9e1832b918882c2473225;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h14dee59e1e118162757d23f9d4d5696b4dc9304707adc356f3255bad1f878fc9a44dddc45fa4b55b2e7e74aa30a8a1b17eadeb08271ee0a18516b0f2d0b3e7f64dd02e899e8e5f0a4286767fa4712;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha2aa39ddd1a3ca482cc5e039ce52062b84ff6c2085a71b981d64e204f25d54fd5591e21d0174113ff07a59a18e00deb80d3a5fee08dc39a2c98b5cde7f82b1c8481f6e0adb81678337f8a578f1af;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf9e238c7eff1bf1b5b8b82baaf84c03385fb96a03af1fe9d8964829c30c63c92d2021326811e7c71b16f4241e9a99396ad7aa8c6ed1c94e7abad81ed9b75b8b8787868673235058d8751d19de853;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h6b7430e2a894ad0a057fb7773461420c4617fe101a7825b6f53ece6a312c27b1a92c621e5eede0970aa6471171bd6f5b67af9920a8681f6a9a696b2b3875c99560525b3b7385b799504a6a232f3c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h155639702206361796c2bb99d95a872ae9c7e7b17d0842ba29832e1aed5eb0f193aa2ff028c921da286d7703b3e5d6c4b5cc4bbeaae4eec3eb31c78bcf6a0ed84ab728b95677abea1d97bfd61fc29;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ee1270650b289e5f3b05a62c1eaffa88fec03bc68ebfdabbc261db7d19dede921d3d3f03ca5486443f4adb5126bb6e4e324d5eff78641a38e5aed2da94b4d2057637f40bb23b8d1c3d3cec760bd3;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c8be1d9c5e05b37393b59810100ffe60af7540fc43ee23cbf1ea282a607f1c261c0eec795e2f14fb5e5c1aa7e0f5636a99ff0e90a07f90afa1d46406591b27590da72885be3bb2fce60b78120e63;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a267f346716a2454bc853871d7813b7f21a35fe557f04136cdbfca87df40a825e84b3e79ed076294e65e70a7ab15973a8e938cdadc37cd17508b51525bc1c027bfe9a7c3d89cd78d694d35437028;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h4258612c3e205f12f0f412eb8423431012cafa911b16bd3f95eba8367617cd63d53a9b4b1d70818a6ff510dc6db6374c857810d5acd5adc63731512f3a667dcfbfad1d382ffcaa78ae7c133915a4;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha8b03e41d518814a22e72d9c991d0736e0f81a6aebe32356e210367f9a9cb300caedfd7b3c4a31555835c8846b8389dae9b509811a035678e563cd954f67cf7437faf88202fa922fc609949a47e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h883c1d63d3c770669be711c460c190045ddf773b801a874ec6e80ce9f3a27ed65f87c9c965ebc862476da46c4fa3025fff1238c6214fd86ab17dbca44a67bbba933623033eff2975a4061d2a2d4c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb88658b2fe6ec9d4eb46d8d66d8dc7778115cbf88b937b37e7881df3adb61d8f4a184183a8244866dc180af67686ce11627abc818aee0931323cb2ec019b789c26fd7fd6bc03e57587d7eb6acce6;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h18d326afc0f3cdb8a60d744727d48210b5c7e36bb9a132af9015dee001324687abb2540d947d524b871fb352f15a8d0cf3d8a462a26f62c9399bce0c1259e8c413dd105740fbd90f36f4c1426d824;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ec5ef479152259966ed8e1b916ff64bce6ed1924722ecdf2b54b0b5c33d96157701eedc697af881fd2b2796e8700fe4f5796a2aa50ba5495e0604d09d443bb5396c5f4d28d7bbe706646c31ac352;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h175d1a2ccce23060303dd75673b0dfd99a0c6c57a11bf32655700860ad19a0c655ade4e370445b1b65b63b55d541274530db71a199ae83f93455a6905ed51b40b5e0f4973b137c809d8f54c5911d7;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'heb698ab005649d470ccbb0d08f7434fb296b300ed42a8776916322943ac66881367d48f712addc6d27f7d37cb1649fb2e8ca7fe223e5c219719177bedc541e6e131329d4afa57bbe6e1d272dbe39;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h3da0d0555ae7aa63ada59b8864364db01902adb8f3fbdf600271f9a5a5629ee26773b813614d8bfa072eaeee41bfe9bcd04d6828baa7730a6996087e14b51eb06a470e0d44d6178ef32d3fdb1911;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hcf1c338556366281875a35b5ef374a67d7628352dc9822652636a0747340eaebc7c3f28bd5177947735ec8aee034fe4e02e9bf5f7394da93428c364088c553f9bb25141dd3d309a4101b14af5a98;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h14a34a05debc88155a82a9789fda964dff62b0efebc1d1b9524728055a0d45619ffadaeef82f74bbe8345c0bebd7c541046331f74a773e7d981b383eddef7e71f3f9f209aaa6199b5ac9a08fd396b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h145387bb0fd1066c9790266c94c3fca2af4ae63f7f9ac560a5b93fabb4f9694056f74ffcb34fc747130907cc58ad7438d7ddff1bcee347247a2ce105261dc30b0499f46a6fd6f30b14162320c7fa0;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ca6fe9f9d64a481b1639b34464e83af49f9cd68731e73e92a96cb5322d3856ef34947e578e5644dea4550cead5df67c5cee8dda4d5e4d09798f54e0ea5ea22e85c1a8935a48d3d00e9ec43755d27;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h12421c591b8099336ea7e0340cdaf290e47edc7060db01e8c5b13d09cfafbe434361361a21f5b498e98c05dcb850011387ec6993b0ead98e5c987905118ddb34facfc487d0d30972ff0d4da6ec211;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h5ee5abfa96dce9bc530400b127bc03eb22ed6fb046b74e4c7002c5c637b49e4da06212bd4ca45f364271c591807ad82fadbbe476614b62128a5418f165fed2a8ecf79492ee1a80fcfcc4367d8da5;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h9fd51236b66f33f284fa52386883d6a59e9c5b337b8c5d7d59412a4dfe31591807b32a57fa8a78bc8e01541d55db9fdfd29e9bae291debede6a41fe0aa5c37533e1a40c69cc03031d0af532ec3b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h17fd23fb0ac810f668e6893cede5b2aa8340835e863e95a9d5d7ea1a3e5d12a489463492edef2d23c5be874d470fe906d0ccf8426bc603ad41d67677d300ec278886fdd08627eb1044bf4adc8c365;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h214f84d316f31d796eaf331273b2b5e0849eb724e112c3e04cfe1618c75aa4b63ae6b8dba103c1452c0cb1512b088fb11ed515e18219dc922d2902ce0059a7b78985200cc5b3b2cc6ab93ffeb7b3;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c8ee72d8f61a114c860f0bba67167fec6d6c8ace4f7cc3bcb059bc74201af5b1b7e039fb44b3d07daf61d5d4a1a2e9f9bf7cde77960eb1df190dc3bdcfb360af6597ec7c86bf80dcf0254405b8f2;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b864a6a2f78335b562c7eb24b6f01f9f3816bd75eda82630f99461ebb8aa8a7b654bb648a3b1936e53d4885b8f4d5c906cbd93db7aa8de1c3cfbab5c936b16d5e230d23d800500af41358ca83e25;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h93d0ff8257a03e5d25bead9d815811920ecda7e50730b0ebf4725623fea2c21499b01f54edf72491c5dbadc4f7ae2976248042f88d4d8f4c2960360e26069d7ea7abf41955c42d957d260a75e4f3;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1588d5cb168a6c34a9510238aedd9c433357d85e2cb25fa6159af5662beb299b1128ce11ab1f5816a0fec841936a9e696bbf9973f647d6cd511128f3b223ec9ceb81743ea469e803aad97a69fa007;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h455a6bb2b566cb4fd08f5a1323dd1a416c5593b1f0318ff7968f7e99cd44c382ab038e8d3c3ca654579554584b2aab40c9ffcffecfec7290d32b964a18ef59739e30fe25a685c20a799a97e84e3b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a3e14c5ab24f2f8ba282f010462febd8a2c1b2b612602fdd4d93a1d8c55da8824f1717051cf35100b5f16b5f6ce57ede1bcb399daba029823c31ef0d830da38a6f3dd029fd7d58bf301e2dc5e44e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h392448dde9664bfd0c8bbdb01f039594698747e38925b5f485d271578c880af312ad05a3cf129944b6a7245b2c573d73e8cc1595da5f6cce04df896ae6cc8aa4a8a73f4fbe9ea5787617ec12ed5;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hfe5297b374b6c13b82d22693dcc24c6e39fccb808b042e3718f8af9bc9091b240283db6d9ced55c60218e414591df4ae5cd00b763b3e963ce0a1366df63fae5046f7a10cf978dedd13999a707887;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf4241819977d018302e9d831aa9c719179e14fb1e96a58977a85541830a394f5ac27ebe3cfce0d6d7cb678f691611e36b98b90912b34cf3284002e7ce1119abb6314813df9cdf6b3a67ecd8a8a47;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc8dce4f2c9abc99742dc380dee9453f2c7678004949be7b3a92c596fdbda5e6fb360d39afeb793d7f65172dbe7ba76fd41945f91c295e7254d608cd4934ef3bcef8408a91e53c73185219eedee52;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h29adb1fb0702a4436335a748ac744dc82d0ebe42065dad37fc76268b8fe0959694a97650f9db8715ee769ac8b7b962ed6231b0d562f6198b98a8215158adc50f5383b89412bb3c93b61b84e92735;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1792122d8b33c33d7b820843bd72368193f432571a14075f4eb62105ec5575db1efb0184d4815712a9e28a24d010ea69288a0d3f3cbb9e0792ced4181b4f24661a3196f70e99ccc5516805b270e72;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1bc22de1dbd400259be73bb12ed65eaab71d03cac183d9213066ea6a077acef5d7a69d3c2de1ebdeb5aa3fc90d4f170c20c315c24a17ce575d3fc3bfad5ca72719ffcfe909886449f9b42bd491b83;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h7f9d11e9d64dd10ebefa0f5cdfc095c31066a8f586f67390f736a140462e986fa18457ada25daa48ca60b79eefaff6fc1567e911023828d6244f267f91f7abef3b0cd6a8f9fd6dc27b23c777bef0;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd8af3cbfa6e5896144cd7d2bd68a2ae298decd9074357ee55dc1642279bc080f4ff6cd75f92b63feb17b886e5ba192a22bb09c08590fe04334d1f36f7d3973578aba565a4a3ff2727ac49aac2d87;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h664bd6b661f5a0901756684668bc7a9943a2ed509ee4f4090c32cf5a047ea259511d2fdbe3250bfadc6c9b87636057e958d8b05fe015f5e39f1d826e781429c6cc24ad16c181707a1d8241d00642;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h185bb58f9141ddc77262890180f9141f28d9ab87ad753bbed709b5cdebd9df673339b1fbb337643129f9c5ad87d878c9cf7037006f567ce9fd947bfaf953c7181843c6ea93461a39002ceacdc0719;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h22c1c7ad20f56ed13295f93604bd32b3963b0c59465491b56f0e71289886dcb9195e3e6aea53d11887461ae9305b37516a8897938d959748ed3719cef5964f93cb32f3aa67c0fd8e4e31d711df30;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h11a1bb6b4c9ae2691439423aee3d544895e605f0a15f96e4737777cf08bc6330d436f3ccf39380c4303339a53ffa43c176ad42651bc29cd0b8c9aa309a31c96d8c6d9af2400b2fb1f6e0463abe555;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h5d0f6d638da5b81960458216ea94e5a5d006392e504553608131848573d1f81e037ceaf0097f465c33d097b5ba8bc37b0b77c0d9da9327a5ec7ad489a8d5853e9d70a79f5802abdfff4fd32eed5e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf2522c77b188ebdcd500677af9fd5cc1b71dde8f6995275df5e1de1bc1feb94bf655eaf46896412ebca34d52c35f8e09e24bccfb93c8d9aca8272cc11236a0b31159c24a83a1a95edbbeec33328a;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h448a88116d9daa6b367d8f59907491940ee280347afe99470519fa441590523e8c3d010afc5aea4a3bd0e2ad556dd65de0c2225166377103a342d4e22e3e760d115662b98e4f37c2062c7b857f06;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h17a40be650d5a2ab9ca95d701a7738cf5fd6b72836959a44a59f8c13b8b5f35d0ca9dd3388025d2fb2ba506e95bff0cbba8412a1db4f8976a228db5a583cbc11672bf24d3c12a6b08764706ec29b7;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc3cb2410b5691a6d568f746548fc48ee13f344f68f98ef924fd0c56a8ea3b451001c33ae1b4d02017fb4c0e577e672a5539a98d3a39930b0cf2ec097297ed113d8acb891e85497832ad0fffa157e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e6aad5552b77dc98710aa560a9323e9a540d3824f1ef441d2749eef853a48972427b32136fcaa8ff22cc9a7eca3ed892a143cde80ee6daf11e0ed8bad9a2a2053058b6e74f459b66b5876c9c600f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h575a5ea4d2968831ba4b958a2a0ccd980a80d4171558f0b287e1fbcf1b3241573124039def444cec216f947542b183389da6a437b211334f0ecd689cb435c59498aeca712a8e26fcf5cc4315642b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha7bbcba0e8d1157e12d29fc6d90d90ff27950cc43e5772b2ffbd04efe12794dd1474f2304d75065a0504fd49315e19306ebf0cf392192c5ea625cca7cc35d3335c1a24f8df7fe915cc89b9170fb0;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h409e61463b000dce5b6a097dd6f07cb939caf61f0a6366b456f8ff77050b98d4a25e61d8045e37caf7ff1ad2e58bfa07f5c1d208a0c56723d9e94e3773996e749826b18dceb4eb94f702c4e0e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b66753d2087e4becf8fff70c680c91a343178166729b68e7cdceab8c1166ab3bd52e2bf1a03e6ec8d46e34d050cbbe910106a2a952d6f221b1d2abe5ca7ca095e824c02924d744dd25bc947082b6;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h2422d53da5bc4ab40790f0206e5a4cbee5c97f01a91156c15d85a5f548cbea0cc7f1df9f478234f56354ecadb0562bea8a9f1eb82f7675fce5330ddc8c71e6987407dee56543a88e6b9a67d8ad5a;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hbf260e914cc06b7b9546e73c1348c41c31c21fccd1a95c481b37a956908cafc7df020a745df37943ee0367ebc218c29b76c64544372d70a859a513682b9a174b934dbf3530cc5cd477e8e44b2dae;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c60715ac648682e8595717438f3cd781fe8bc55ab0f0997035121ce843e93baf646cdd0f764f8ef3c7f0e1f49b244acc1f8a6f8cc3550f9dd04a1583fac2f7774250e074f4164008463559bbc5fa;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h191ec0ddfa8563b8df678266765f974c91276ccd864d7f864ea28caf7f7d1a6efc5a3664acb30504194a55fd10a366124b0f0126a871a7602d1c2f2a20d17b21b569dd72af8dcc108ae3fb5656d0e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc665b37108a7426ed57fc85c88f3b521ef3e4d29d576ca74d2371e5b7589ff2990075279716fb6c8e761832a629215800e3ca4c9d50d23d8b910b99ed58815530c6db0ff6ccde8c11fccaa9536ae;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h12a9cb8d075ee4955c63fc5199a546a6cfbbf2afcdd32ce30b39076ac0770e1117a286606d07a5dae24b621e47750ed4e87f898551a12825716540224d2828f8e95112b6e04495c10c2f0e38436b8;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb7ffa3760f054ca4281d4e49ef4a430f8cfa0429ef419566e83b57dbaf5986832b02676893037d7c4156e20ee90f43c9a89c1266611f8c34112a79155a37a83a456e3810056b1126f063c81de5cf;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h477becfacee702a6f1954955482c972f5762c680437aec5abc99fd45a4fc79d666460db28012de8fc03960c56e7a4f156c53e4a1dc01feef916d8a102bc092abf2ee469ea3bba5263fa255ca338c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h7ddfbaf8f7a68e5cd2f9f8c7bd1d0deafd44003fbdeab3f87eb556378128a5146ed3ee9c91a4f2d9883c954926799cbad8a005b72bfe12be301f747d006e96b95de1ba6148da525b287124af7589;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h8c0dc8d91fe4d2b902fc56f581e56076a55658e5de59f6c61174c37879f4619feebb7618f877997854d96cf4cf08acd727616c37b2b57af0ac618921fe020df860a1892fcfadff0197c6c19e5e36;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10801cd8703f1ebf4e66dbfdca51b16a03b61cc2ca27b5051e30ba2f3549df27da346cb08a13c1c8df6f5f2c104b066c0619baadcb0601143c8a27e201dca31c2e64328137445001e2e8701a65d26;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'haf927044ee7643da055f053482f58cd0c8dbfd9597d1725a6528130da3b0e911f96750441ed658265a256e0048e195e1fc4dbba8415336a6a310cab2dcbf60738fdfe938679ae3209004633162a0;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h19c349439cc9de082041d42a77ce00e48d95d6a42adbff1ff578468939bd9f311aae8c6928f857e6fbb85ecdcd359ce7c426877698cf995d6d5051877675ede4ab3662d239b1767690776193677fc;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a0e8346ada3fe4948affc31d0d4eef4d07beedc327f4da7f8123eac6b2dbf4c4ff5b40d65d73a2d3419a0965a00686170ef6a0899add7657de986a5bb041a6a24684ff6bd2d0853e57851829024f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb23ad991fc1f6dd35e2c5f4f7fef102336e0930ef0dacba7e8cf2e2264193a0b0876fa4281456dc268f430d0c98b66576404b9f5454df6b69213fb6dad875eb4a614a0c4d0e1228443158840b43d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h83a4ecafcd2656595084683d02685a0a648ec650bb697e509a9be934fd0add1d762fa105407004b6f94b6405a5a7e35a4c6935ab73ff546782ddfad4a923ea176a45b679fa522b7b34ff64660fa6;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h146d71f9be7a97d97c82abbb184baa11d959e10b9c1ea67d244c6229179a3b49400bc31a61e38db75bf09dc2973b80639b12d4d4883e759af797c877470d8ca68a46d44943e110fa8c78c6e95f163;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h3fab0b1f541c4fd27f3a03487e23a1cf7e1def30fda3e03e7e23f2a091b01fba5fb15e42ae324ea4ef21a226411ca47d69ed18917cb8628f9aa698b88c2f368dec96b866a4770da842be2750f44c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h81d72d1f3e7bba6c98be1b778c3947eb9fe2306d19dbe74b6b860584362afd8cc663da34b1d6c0562c6d0e70b0c5f698e1184a9257d7b7b90f2e71d98864eedd5386d74167530c69bea78fae6e23;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h143704b9ea0084dca2d0c90ed60cf2437592a33cee72d63ecee4e5797679239632511b0663670e450617a212b3b2418738df95d311d3a1600028a3aaca62cba2f03e4aa9ac511f957fe785a5542ef;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d0c431fc66e8f33b6cf1c115cc8e6c346facbd740d45d2f69e6f17e48420447e4570c01a311589b7b4a414d43aea9cb5a7e28712a4123d8c468c5aba3bea068965a4205fc7809ec8265d03d1349a;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h9444b450b4255eed5f3e8985087ce7d2cb1249aad1430d94e35fbe4d92f110953a4ee627b95d6a853c66a607ada360b2e61f2d6ed226abc36465a336c4b1615ac541b86f1ddc8ac55a7b5ff060e8;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h9e6f5e9dfeec02f961b861d733b37d8ff260e8cfbf5133ad6a485993de656a923b40f9680524cf81f613889f5451b1c4510240513aeeb27190dd73e4d80316a98103bdb6c8aea3be8ac75510cda5;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16ef04bf826bec3c7988a6cd7949ca99cbf362d3f16e8e783f15e0b1a6dda08991be0073ddcd4b5b431ef045f90f7a06bfb493982933cb338a423e0a4ac5b934ee892add61eb21446389b1bd87544;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h6c2b29e7f18eb1d96b7e9859815da584233f0240e3b71da0bb7c7a58cd21ea138ce94d6a803000a9520eee1f9d65f5114fad3b6273c9cee0706cd0a205be03c21cc5c82b1398f114546077fc38ae;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc4382e514e360d6c4b6957b67e0bd7343a6cb290af8c24e619d966273d6ffd8b71754aa9e57236169bd8114aeea57912a55293e7d2a2ad9e7b0cd3e797b43f2052f9c28c77403252c34f88b13040;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h99e6816c748dd1a1ec0c1d7bc3c3c45d5e79aca8fadf323e398bf2b2e9d8f833ee3755c7dc6b57559c093c023bd611ebc625830e83c7af76f0f74772a591b23372076f9c3066eb75c74b0e39e03b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ac963eb497ee3b039f4500ef23f24f40130f36c6bea633d8f85ea619126edce217479892fb607240d276d5f880ca8251ec44f41d641cd4671a218460c4b6e6da31fdcf062709bacc7daa4309f4a3;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c0ae89791c930980e36e7e8f0b8554c910517547663e63a5422e20ecd4d92edb43442e5fba57f2e54c1ce352835e7229de968733aeb12a838976ee670cf5cfc72959fc1eb02e34a243a149ae8db1;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h12fffcdbd40e8a46f38f1bb67fa9bed2da2a7063bdb2a04f40ba6d2473ce4d5c44b49ad65292d44609585239cecb5bcd2cc163cc84fee10a042d966057091fe74c8c270064a432e7fae8d0325370b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1266fd2f54d9ee8c4dec143a9ddff763b7e708f07842f3820521997331f1f65b1997a769a215900164b194a96a11f387e9302dc50294a8245599819a3589614e86fdb55128e965148724b29448584;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h13e8784944249d9909a8048bbfbf3619f15cf2e4f5b98f2c811e4f9167600164f0d3990f61b55d6204c84ae6fda02b8333268d73a33e70f24fed78ff5cccf4e50e04771e5f1e76877bcb9233898a8;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h17516bbf0cb65b7dbe8e18b28626f661e5d614c76e8f2d3dfa990062a8ea09820fd1e996a8f25c1a6ab20e7993e15ed32772f8e985c00e3124d123720c8fe5799b793672dcb0a63c3166cfcbc379f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd84b4b726ff5b48162fc66e97d6d0be6e86901c5c1f67a2e79d0d10d7d570c3cbb48d83faa2fd3e3cedcf0418d9e88e37c2355142df36724588090c06f72fdb67ea24d64893dd2772070ddebe227;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a56b2df77aa62475fe18a3e2a6150bbdbf1ba80c15caff959c3da321bdee14ce5eccb155182d302dee6caf8984bebb51d0096410148698593ef1dfa55b946e1163ea89fcd6587e50e51abd72517b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1782d82963a6a8cfa1655dfd54c99d4e3f838d77c2a0920974cde6b64c8f706d937f3bb118967dc0d633c23d8ab53b4060232900b7a7930e88287d2ab9748ddeba96ad430767f2f3c6543c74b8d2d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h63076bc8ce6a5dd3cf72d91574c04b926be8ef9ad3bb794e362eb7b7fce15e30eee1fdd4b8fd631770e3108e45dc882a201b135788b4d97daf73388cc112bf56b605cdc49459ae4f462c3cc87bba;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h103763c8702a7ad2289a2cfc0c6c04031738833a89c4708f1aeb748247e89b1078a905e72fd858887b35ad7524268ab8f647709a107fa2ef034ddd7512658fe869657ee4a4468ce5f52a6deb9dfd2;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h15726ef92e1c273eeb2cb29c12334d5db912bf7a52e6e92b61e1f5120faec2d21e605a8597ebba842eb74953f4aa9be2b21e5b53dbd3b5cebc2499effa80be4bf2eb1a19c5dc18d96185da4c1cd0c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1867bc91816d347fe95a73c6b5da5a26e40197929d9710d262bd671685eb338fc04a4172e7c404feab188c0f0d26a481e4629e0a3cabfe5d674a3963dfcb414b1bcca98fc4c395f1f148a51ccd138;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h6071d0a606e85150d3f0e72790370846f45a720ba1818aa2ac9a2ed3f02dca3b28723d942beb1c257258b2f029677861e876bf70ce7ed67b914c2f09ab287e2a5db1098a1af7c429488e17120eed;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h144b03141cd2a01e6fe5a91649191f779c3b406c4b039b0bc1ea96f66e7f2b0d39949d8b2cd95535da27cd753ee59f58240cea1b55880f5d866706b8025a80ad1aab5f499f5afe71e8cd59869104a;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ccc1b70ab686a35538cb7bb5074497222e0196d99c615878f56aeca8ea78400355a469b1b39618208344c251b1b9f741f408d9f224029273acdb1b3680e4a1d4c1b67988aa93016d75d43102afd6;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he259681dae8809dbc04e5f7944578131b9063f12ccb886100970b6d558df5e500d87b751243e5f29843d5c6578e6b02476adb84cd99e616b3f2fd0dd1f33695c62fcaf1d34796e90059bebf00a8e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1928723b42947dd65306332b0a3d2996ddc457f356a05a53f0cb53256b297c27e099af30d40fb013fb6ed346fa4269bb369d32892a6fa87748e9a1a09de2a3c1e0f031af879fb6e2430f658848f80;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h129e50226abc7f478fcb8c2e4fe41426a100939943e3accbe440caf81fb63053f6913dc1e2e733018528198a092ef051f7906e2e7f8dbc5453a0c926a2b6b11f25389cc6fd3d174ec48ecc0875aa9;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c27f6a5419ef12186591dcdcadd1d2d36ce8eb41252b3c283f73e6c98866aa9c5fb1e5affa1a0fba66cafbd720d890c9ab6865a1e2314ff49eb2da48da7aa2c9611810a84783f533d5e2454df300;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a4a1aea6e1d4f5b078ac090ef26565c61ed333b2753dadc6330df92af82694d4cbd4b00892c5d1b4962608a2daf96cb5c531c6e96e66a83e1f04cc8cd0dfa2fa1ec3e5e814bde87e367399c23cb9;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h6d416e9fcf8120eabb593c8055f6ce803f6ec0737577475029edd207802b5e0d8c01f9d5dbda5f115be7e63370d0ed9bf64dfb0f07d210dcd7b30eff0ab0798349ed0f1d6c5760edbbb494280697;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h11ecb79561ede582429e25649a2b4987891a0107e4aadd4950cbb6a7ad3df2b32532d04d7456c33d8d111237a82f4efe2286983436c4cf37535bd051c85a36f528c0256de817963f4da53b232f039;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h188bb7c371c28389c78f39637bc32b8851d3e44918e0b2d712a27a868b8a835ddc6677c4b993e9d7a224f3e27183b69c6b8fc2c7e472a205daa3a46f516ef41181b45a39d70f6303fae1e500c7b99;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha111fe02def7cea787b68e128a98eeba91c874a4a2de5fe3a22e704eafa46e549a29daf295588b3a2198394ca2048b696100dcbb005dcb3084f0e14fa800e95e35a62bd8ffb9670feefd8f1958af;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h182fb19cf32968bf359978df6d158c4ab2347afb09c0d1c787def0710934f0e8f2e719aee8349668b00a46014dcc1736edd2c639ab05fbb04c3890fda38029911b90febac0384cc375a98437d8306;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d8904a7c1f08accabaddfd44ebd8e47fd04eb915fb489b1cc4efa6acda9ebad9f5a332e7de9567db86efc593a33598f19e311777e2f870f054cfc5ca7550e392ab3a88d1859dda365630f4a0964f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha03ece6682ae8978f2f6e4cc714bc05dac099391e2d0d46b8914e9937143635d2eeaf73cabd5b17f1f8a616078268d0ea86663214089b8fb40f412dfd4a8566de8868c6fe9bfafc9b1e696ceba84;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd422defbcda55f6cc96f0099ad6492832d99987245b2f3722335809d34fd4c60c01ba6ed544391acd6e4a4b37e3148ef45f0c29c10e661009fb5bf161528556d8c1722c9aa9eb7d7eb033737e71a;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb2e0dda05530a197dcd6752aaa37dd6e9249ce0474f0ac28ddad2653929aad225c488f8c430201c8aa38b8f17c3d5551001b07d1816eae9ad8ddc71e7324513ffe08089d7e60172c1017bb687683;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h7072da50de344c749fa5bcf4c8a0822a234d7c2e87c6344b0fba1e846cb912eb06151675d8846350cbf9e4896d782aec97f36e97d3630b488dcb871840b34811e8f83ef46cf49719852d59b4eff9;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10ce51e9bd62e1a4ea84dcac7ecee25aeea8926d2256f5f71ab4825826176cbe54e60c0479a5b588c7db13476fb0a3b9b0b3cda4af8e5d264258f3b8b8a1b1c989d3656b02a98d0b61e535c9dbe1f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d8bf74e107df853fbd07b77574e34b70e60abb0ae5295c12c32e7c62138d2250739754306db27e9caa4941b0949022886faa28869c548c1b42b64d21a583a246540a0a7427a8f43585248ab40511;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c96e4f7535d2356aa0d28c1f3d940eb0acdf6481001313939b16f98a08500a55c4fdc7763e4663a34016478c6285fa472627ae4afe65cee99ecff889bd4e6c2435e1f9185d56d814463bc5d36204;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h14677aacdcdbde5565b6e5df4c63d34e7c194b27d576ef69067f610a1e9c5ce6d5a5bef3e1b253de9fbcbc8d0a0110378688873212c71b0c427fd95c50c1556e0672ca1c4d961be12b1c10f237ef5;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1bfd0465bf0d1a9372b70da44e24b1f809261657d65eb2497527bae124adc867e1d4ed166b06776b47b54ee519ab5c26e07e2954d7538849b00d77ff56b2c5adc391c92d5f5489a2b6ac2aee7ea97;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h19f3a8698889389b5113809ec506422a6200d8087e6f584e91cc9b4379d510ec6cf1d2700394f07131715840bc35aa3f832a836c664df5f0061428dcc3c14fcda0e06a148ddd41cde906cddec404;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h13960ee8c716564016ddacbb9a033d07603a3fd279b6a92a57cb230d32a113adcc7dbb1522e85bb2147fb1306f20fbd952866fe67a062a45125d338edd02193f677ea8838fd1aaf334df3bd500d7b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d249eadbc362cb6f0992db85977f219f45b2df8aa83fb15ec1d5673f82db519e954db383a65815142242ab58bba372fc6c51c1276343d3ea8c17c0bc900c4a1ee67283249f866a0eacc84eadd16e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h24b0d391f1d38063c427d47dae9c2b45c812ae66cda486526d79996665aa6a97966f81fa4655daa4c5c799d6814a68eac4feca4521d1998adc1dfdb68619ae8de2102116ee3def1bad162c2dd955;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h168645f70bd96b008655e9b95dad1351f362f20c104b45928aa73a4a879b6da00f47696514e37519719556fb3ef2d916c9c077d9e40fdacf2adfe21ae1d3625836eda095c7a319220ac043eba3859;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a31e66305f93b0a70a7ec5fb6b21c3454bb83a4153c507411fbcb004789c12f310e3e345516c1de5bb5df1491399781a70593462ccb965a787716dd29c49df7660eaa3d0e74d9733430e4a16c90;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ce6583126648811f772bfc72621c436d19fc0258e117862783db3addff7304fb06106e727b98e965bd84733e229b3d13465aaae4a29f0d30d31978566950514008fc19819958f7a3d6d25a6756ea;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b5895303357082827a262e3a350973a38182bdcd213166a891e460d66c7565a6dcf471e6610294f90f03e3b6406889e7d12995e941cc1ebba8623abd8f61a345f8125ada97184519962ab1a4ef4d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c177e019a4538eaae1ec257e0cca904841fa6b325a6f80020aeeeb514b86266e293698f666d0c7d78e7a4eea9385dcb725787f1ab967aeb17a025446b98e50c4f29a2734222cb89b6d9bcefae9e4;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h178ae8cd875f70dbd55c6e3bc7d38d5a7d8e4c32e442858b2b3326350fb6706d932f2a20257d0f6c6b609a63370e9ad4def2809700db084d123e3d28834cbab2d3e1bacc2dce7082fcf1e6708f40e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h545dee05d60db9376f9fea87821745525e9e201cd5c7942fc4d91e1f0985c0e2d5cd962d3c032477728a31a93a13a574ee9f40c63a6d117065f848ab43b39c995a6720ffbb8c19052fe9063f4b2f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h3ed31be741d084fca9a5a20c7bd7c53d10cf2cfea3261c4a2f8040f29dffcecf55aaaa1641780b5ed69458f3958ed7367128abcff9fa889b1c9b41e366c7b2199df421b9f159be01c8487bf10fca;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h57e27adb4fd0a33ffa3b5e4bd50491d7264ce18ae75947cd466c86db7c81ffcdad2df5ab62bd51bde577567ee1766fb7d6e603df2feec020613e71e6b20ce69192f316b4047130c6062e37fe37d6;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c06c3e361729f41f6519f69d3b2df1abbc88010e2ffaa6284633fdf96e831dc513b9dae8195a007ab8d7a81da68554241679e5c127c4dfab1da524e9574e4839d7c91745a71336e0fd2b1583efa3;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h50326187b9844a7154c38bd4a8d516ec6fd903fced0f8b26631f04299e050479241d1a4dc198099037c8df19a4b04ff30f55c1b223897e535eacbaa72cfc9f53f19a738384cc3ccdc917960a6311;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd653b30f405a3e1822689e55deb07c66f80756a75b64ad06629eb3f53d7cccfbfd5167b2cf62255f60954ee838caafa841bd55132b8827ed8480942f07b4e592fd8c98b3e9182194b2eb6e40e79f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h47d3a6599c6076a44047018558aaff6565bd8f84f3d70e11ba1039c3655e5a88729251d0f6e14ee141533d4f9defef727f39855af22d65ca53c64f8503308726a4b3a4972270ad3a0234d2d324b1;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h153c45f2225e3713dfc489c885ce383baf1af9c032c65e896cdcd42ef9dfe4d7078d2272ecdfbc10e7b84dd9682c0c23a77d5936c8df96437c8c8f7cb6e8943ab1eee504256b2367397eb7db07c3c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h152a02a4b4c7aa1d912e20eb40b33bcd07b58acad0fae88a6e37b60753dc41bc80e23aab10912d82ab28429eaaed94e55dee3b9462067a016918a7915bdb3ef6f59816d117d37d736c46089a5532;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1511ad8ae11fc4120e1a3b4af3abee98c4af954527c8b8c5dec9b83dd2dda58ee4f1fcf81c24936e03498f914af8ffc5ada2187f82a33f228dfa9cb14037f6172dc6ef6c9d8450440681ce45be582;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h17f69436884a6013776f417c64b35ee9f98a67855b8548f01a2269a42a81a92d4ed7ca63c3fcacacbc9705f22e87246d92a408eadcbf563f3a161aa5b5a8184469a4bbc72e74904f1c3ac91327630;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h13d88f4741c671447e9b093fc43cff2fdb07ae73bb2ca7b395b932c1744c703433e749af2419bb3473563bed5a1dc985416cae641f650ed97c53c071eee6fe06bea542551db33854c97fbcffc68bd;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1bab03c63fd5a98cc1ab9aa369dca75f54f6759177379259cdb659e6bac970d03a48da6340d55c6c588690fe131001259bebfe0cc62e94301d989818543ac0d077f66a6c60575e330c8c3313a8b05;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1af30d3a69ed3f61a46831ca61ffd8a9b1cb48d23c6feef197ed9fa90f8d944db834fb12335b0072f6068a9aa2838ec76cd640d87ae42c8f8c467d9ca554c44103101a9bf1795ae0937a36864ed18;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h12a076502cad6e95b99d436bef6198a0d5a731eacb75865412f6f6b87e5b8d1e806ea25070d0832b92facd37e078e8d5a78555b59bf4d796eee0913d6a5e707f51bc875f836120ffe0a242ef4e3e0;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h9fdefb0db7d8252e7e59f954158f941442e5e9503f57d88670dd341f9ed3c4ee8d6662060771db1aa11b82e494bbb05704d9b3a29acbfbf8b5431818b91bd4b82a32a40cc2a8182f4948db94d9b3;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h13ccbd24777945f8f2eb2bcecdbbbd6578d16c1d401db7502494daaf24f569b78f27f509d5ed6f19e123b66baa8684849ad6b02ca2aa037825a829912da62272d94aeb571503126648e5af43c7f99;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf961bad4a866a6577730b354f23651a03ea0404144478f7220535fec9575f4dc139765852b5ad5471c8fbf86b9aa034e529705ea3d15b05a1076894aaf41780ffebb23b57402851fd2f7bf3074a1;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h278fcc4ed762638a80720976574a627cc7d2820ba1103c7c5df8e74ccc6a280f9cd5c350d636333ab388adf74d0aca59d2d05e033a26165cc3a13c9b570d8123073535cd1ee53368a75deb48833c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c99481056b3713855f4992654433fdd5ac9689815b5fdc8e1ada922078722d33b1f9e111f95e5cb5a42ba907fdc9a3fc739cc30496dec1e6af5cdce1e4d2def9f32122766f85f3fdbfec5c46ea31;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha5628bf79d357c4cd95a13c6e5708bcd8ee6101a003e62c136d64b964223da23c18de74b9fc3b1cf413b4e2b367e443d872dd46313807b9efcfa7d0c1c9261c788bf15987505806831317d20e28e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e97acadcb5ec4ac7a68331f1e97f4997af166a8b6990569b4f1febba7fe01150fc0e3e22e3a0f923c9a45ea89545df67554d796610b3d0a73636b07b0f95eddbf8a7072aa609fd73fda4add6bf3a;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1cab5afe57086e2c222a09d6e4ea048a416f5ae154acd9e286434e6b75ef1ebd1714de3659d80c4193e812ae2189dfd6953c9a691015104158e079c0e5c14bf9094af9058ae19cfaaa9a41a539c49;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h53bf0a966d335b5b6ba144e2783de7836406572b07af1e8f0261568fcaa246db5ab044f47c09c359ac361d4e8ec5ae54972324a470349f7f735d0e70b348ffae047691ffea461ed562bb25145f28;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d745d0dba501ab215a9c0a1f45cbde8086aeddbcb9ac2208306fc08137aa75338f7a5a57f416bcf47d4c11dfa1880d46acc9dd3b6f4ccd5489e30935dbb14b4c40d2fab8972e4638346f5fe7c1fc;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hae3a4b2e35e6c133049f893cd6ee9a8a43e7e656a431ab048eda6ba0fa6e00faf58e0f16985dd224a447f89c11d0da8454c31ae1e2e8330200d9e57bd28637bd5664924bbce663ecd6bb04d6cd51;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h8d0698d6b441be20e4013a9b6fffe458ba33a136b1ed265ad0836026e67c3b6237cce7d7f2f966a2f5c6ec1594ad56098be2b153f3ea2dba6d43b9afb1a79acdd10d940b1233bec3afcc4e35492f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c041645ad9f15e036d0f55bc771ed02aad313bcf0a28c1d2923d8e555a2850c2aa61333d2bdcc5a4f05c5f9c80a7060934a6a02b410d9b79b891bfa4c079bec87d3b76dd7966bf022eead57b07f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1757d7f9e6d9eccfdc49c86be03ec918f401b726a0066415a56be232b5213869aaa7ae8d47e43f39518aee8d468bf8c17147e8e7e78d9c5734dbf3a2d66ecf2d8b9e2534014595faac1cc30e19ce7;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf0489974f00b4124b5bbe0196310291d624f674c0c3cd1e8c402fcda3257a2bd7b0dcd7dfc48d1c4b74f65d549b00683b576286e0a71b9676afbe5b82c91bdcb80bc47c93774053aa6ba458b99d4;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h4246ffb616547986d33c5cd9af3e71578738ff62cf25eef9a38a3c7085b30f487bf4048762c760221b63fcfc7e589a8bc8ba8db0cc8a71f13140cbaaac10a111279b21f1c4fda68f8fb965e3f8c3;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1fb0b1ca49bb289c4d6e3be1722a5140bc0464bec1d73852153eec1df8a6526c95898894841ff64edd19de8cf6b11f456b81cf9059c10501d43af8679e6f8ba55b6b77840b0b70f336077ad45701b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hac9cda3357b6251b082cca30f766aa313bccd61343c8bb318af825d2bd835a3c62f1415a3337386cffc98e110985f2cc97ead28e8b5afabc28b471a06ba7c96da780f1c579fe40cc3ab591c7d4d7;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h7e6ca4edfe5fdfa090ce9fc585ed6768aadb955b1d5db6e5ef589a685c1966e9af69b561fac5ebced137c8e9791986ba185edaec092b5cfa97f53ac503507b7fae0405a3ac4e3dc6369c4f11b5d8;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h8a738c2f1dac91068d81232773e10c650dbe2315524389eb030637224bf3b32e8d8acc91ee5b82a6c8d8e165f3f37367e70c154b516215a805edd961816aa5255ffce0cc1fb1d62283c138d2f962;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h176b1803fb8024633af9bae1c4d4394f8962e73ce83871b864d7a7f868029728687a564098226133bdd1b77f601db8d042f228661329046f768e805178745b2f1b64305d57b9346ac46ac03dd449b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1366eb4ee156c32bbbd13ac6376a8bf5f96999895addcab70c16154c27e7fe472d8887e86aef521886eba6e80b42a66aea24de4c8e0fe64f9ff44a78edb1cdd3ccd4d2b4bcd545ed96ef60addc12b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1022380db7e1e69f98a809a9d83f957d2e23a98089d8bea6f91ccad8f295d171a47ec5529383988046893caae48396593a19964ba6bf336ca12ae43c668d236621fe3d39beed4727c6cb64b31b9d7;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h105bf9b59e2d1fd63d3ea42c607e1a2bef2e434dd303ad3a7655be597e9b67620765b03e9b24f0431135ea878f74f364dba32c532d5eb65e18c4af153306739cf818f14a30e5233421bd8321320a3;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hfc28f4e5cbe13a78fc2c222537cc1253c4a435e36b0c53ca1be4eab3a2093a199810ff3a6a6f1616ec1f400099010a00c62bcaa56509375e471a891346352964e505b5214f1601b54894d3f01d4f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1169c1d1c1043fba9d4367eb9578153b5ceacf265a85476c146bd0c6d54b11949f2ebc562fa4cc942fe15dc90e672f096c97f6743d63d35f98b661b9f9ebe1e00a67b6b2f8e3ab5ecb7397b615c4b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h4667e76f7b737b43ad1f4f0dc813144a61200777132f2fdedee523a371b44f39e54dcfc5af5010f47fa628c0d4aac571614b92700a81f41fe37004e78ec425d2bf315aa5518546a6a8a938b953f7;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ef44d1075eb9f52834e98211b6952c1233ecc5a5d01eb6e2fbe3a9ff8f9d8edee440acd33b36c362bdfc07bfbed9ae753e60bcb033812ce011fe0ee8ba704f1bcba7236bcd736f0c3fa5db0553d5;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h79ac86637216a1cdba9f2edd1c7525e74cd73e16c4797505a974ee0b050ad9f3f8700e30717544ca35319cc92e9dd628e00e4bc90a8564d15e33854fa9247ddc3f3c99100d3b755127aeabfa7164;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h7e3c287bcff18cf477bf3d34066b0dccb2478d97a42a46921ff1e6ecdb25d7593020a78f942bbb4f598a4401a0b97b4ebf07e15fe8573c60ef29b2eefdfc8b791c0bd93ff1fc169781d32cb0812c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha2d2f37155fe15e9feeedb01c222c28bf5709f7639ffcc955ce7ddd016aa2e5f54bfba7392a59102afde1e34001eea781f923da362741d78434570ef153a5737c3535649cc3d40afac19bc4649c6;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h118654f39b06078053680b490ef6de40bcc87967d8d028e9f67f6280fbca1b9a6c06e744bdaf5d75be6b4eb0b4890ac8b8591e20e5762301e9220f8fbe1e31579eceeb7ff65213383ca09dcbefcc;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b6eb835fd96b53c2c4ec9b75f6cd83058cc41b63441f3ce62d14687f4d4028e01214c2ac8fbc09037b30eb8174412ef1f2a96a512a03d4823321a752234a78c2e9a43dcad27c6951606f1841ed3d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h122eb52513a910933baafb88494453e2adf04dd3da83b2ff4e7395553c26227bfc5e003fbc80273bac8f87620eff485ef2db8a6f5e162228c4724ec3047d6a7dbd237251cebd3b1e8d1d6b9601480;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1056c527fe35366d802c37a3716f70887360f1d8fc8079efb440e5d2a81e63ee69fd64b3f527c24c78ccf6e7ba48898baa304fe3d35f086a2010aca687e8f6eb45bb298355ac4e1d096dc20c67b8c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he51c9a35e35f5938fd17629f3afafa0a30a1393959ab6c515f2919d3c3e55b387564f28fc53a64a3a2a939bce2d4dc5542af462883ebf76d8b759acacc1d7b3fec8b631359f6af1d37730d9eb6cc;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he3899f24d52d672398d3a329fcc98b2cb2b16e2d29d2296523dd02023721070403f599d73d092c40d2161af1d5122bf4cedeb09bf37932baef89c67d220079e9ffc9f80dd244dedac4d2e27bad97;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h14b3e429921c8e09f0f3ba5c0f7720fa5f42079025a94e83e5db4130771ee40705b90c0f62e49e33f22d51ad15483e027761a0857d8fcd4f52fe8fa0d9634736a17f3833909b96b0279168b245b93;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he73e17db7c4ad9f16be0cbb5514002c77081aa26997f75249ffffc482cd1854e883fcc1dce9cfa39a4109eef33b804a9dbe15e1521bf84c5f17666a29f8721ed7f1a94c803db0afe1287483f7465;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he66408bae9e047b6d3b8ea8cb94d2333fab15fc4647496c6c858d886b9ad2066c093c87c0685a9c5aeac0295e9574a87588398d5d8720832cdebad3d4424d71336e34c9bddb0f6aac63f7e22a6e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb456b4fcf26bd473200f8fbce366eaa72a5240d3f742b595d2b0612f794750403aa43556c2cbf53f6fbeab95cbc4a00a45674d2ce983488b53f3b9afdd4950f35b2656005e0440656dc61a38e789;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1649f470058e4ae33d288b55c7b310611462e3ccf6ae128ddd325f65e8072892d3726ca575712c003195f0635f30c7b3d5faedf4915031cdfdccc8b296376fa3eaceaacc2ed2e0f5819829d1f274c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h15cf9ddf1ee8a5e81bdd4f1dd56d0316733176079706d8605e102410b646235ca8409d033379591da2730d423bede35f119fd66084a5830d770e454b543a085100e4b9b720aa840f451f206da348a;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb6b4f026e048556684f6cd5e62f29e33da05f2da817a00981cd5fbd8c0ad9a3552ac4735ab634eba432449af68a36b27e330a995ac5f0681e518b16bab129934850212e96ddc613c600d9dca9bac;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd8ea0027d8a6188cc432233d974c5f4472b56d722073581a11e354f8f3502a04d32211f94c6d1df7500f73193cf643fb381e332c9363b3743848adb3c737a1e3cc589f2eff0a3e85abf45f975074;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h134d600df41e785c23cd2c6153851ff949ef479b25317e82dc864e98ccc9bb310ed2fa8a4f29d0e685feb5073c35222d311f97f97ed93ae707c886e6537cae5ba75285814e513eb8b5cccf4ecb5ed;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb51e283ac3cbef656f13fcc736c4d5b08de5a9357c0c1214454358d7a4f6230bbdabefc4c4e7d49b14f0ca11a413d2b34060904fb6f81f0218620e6d826d112fce839c47a16a9e7db2cbe852a0eb;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha92abffff07a4f866b6c50513b83c2724c4a05ab691c536180d8ca4f8aeffe4e3c00bfe90f7ccf58af84c769d1b24014a0093c0b303ab9e56dce1643845ef89c688a4456c1403ad3c749a0eca48f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h43f8e99a8a982e83db8e1a567e471e03a19a66f3a6e9211bceb67186de25d08a4ae3fe06c6e99b81db107793b8429d35d01e07fa5d1d6e5143cc0802d3760327c8cfdbc89073605482b9a9a70c14;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha12adcaf627dd6af966d8e22001a1a7d2057f95bc8086c643e69195be47a3a106f4e443c12bb7f88a19063728a5a57c32c3795d2946fe72ac3e7febbf50759194c9f90323d742772a4d7111f527d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h2b2eaffa467ec698c7d0897713a5a8eaff5999546ac46717480a932eaae5fe8066507b66fd2921676242503e745f48f8ff88d60f46d48a267724bf72cf9a4d8c16c295ee919809fb75afb6c83194;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h41abb37c4ecde01cec45e3be4719ac5c8daec1df48e3c7acdadb6abcb10a16dc371db7d5a7b88028470324b7cf0843a88cbb954fcbecddb639770b170f466b8950b78da0ebf0b9f9f06548ab46d5;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h71af094e6c63d2cfeb8ca2581f14bdcf34788ecd68449616be9b2f35fdeea13824f7babba5b86c920193b65c6650e6decb17725b256306bc72d05038e80bd65e724bba8b18c947b47787bceec5eb;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1568fac0272d1167375485b14d02658af81e7166ef0ead7aac83f15b98a2b2eca0ecc0c3f11414e484ffcfc3cb36b562eb0cffb1059dbe34600a52f394786ab03935ff6c6f27e2a19f54bfb8d7360;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h6b8e306d19d4df13009ffe13d28d4d90f2576b1675a92c488600696866e55aa01bd284932314c32e58e7edf5058bed262d314407b165b1b587487069d7926b65f622dad97f7ca7660f2d334133be;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h53a686b20b5b9cdf59108c05028c8f6fc2dd02efd49a1f172c02a1586a68454f0fe6e84ab6929c6220b203aad369d0d4c0a8205385236a87894b5f19c1ad9a0ebf359c0ab5fa3d78c96441f600cc;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d809f75cac182b0b2d758fa79fbc75c6c1b46bd1155808fd6b5a8e01df5466882f34a19b406820e7441a05411a8ad6530b6d98693b46f3c6e781e38a001479a9270dfed14558cc0d69391faf1a70;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d2edcdfc7826e8b3a7a17643e45b7e8585389a47add62b917a6eeba1b88b62ce908520ba8b2c64b54b957cd903d0e038f71f023a074a39756b877e6fd5d853aa76ab8ad7ccbb8c3ec58049ac9efd;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1594a4c943413eedcb6d6d57b90c2b5d5b569106641594be58762dec5d8f6298e7d7ef6f10e75d93d90e6644b82191faef29ca998e5e58323124d8dc1d17746a2792569cb7e35944ee2cc30b624ab;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h145894e95d85899857bbdbdfc7b5d1db00b8b2356e4f744d25c150a0fee84f2aea289ee7031ff0ef11adc3cf49ab2af213071f63109f71960edd70af6ad9f05d64c592582e9d4db8266103b0a8f1a;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb4c602b464f688659739c013f4cfda22b58357d8f0d0d32e571ff1fe5dd44d823d511f9d22673a645cd74440cb41b9d027081a829f6155e23033630a5d22c980eb2c90f28310b75f5bff5e1c6e0;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h149513cd9f4247b83a515a1333a99515bb06c420b252cd8116b4efdc986a7b3d099ce9b72e365ec2b804bab065562ff37c9171e5034abd3b9a7823f21dd97611de4c0db535238c6494458bd69dd7d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h113a69d67bd3bfe5bfca9a33e50b47d1eaeaaf82654d9354671c672fe07e6f6c3b912f8826e8320cb02fa043c7bcbfe34f84bb043179b1db3c2788f05954972dc5273473bd2dee902036977461ae;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h12ce37bdfbfec5efafac4d8a8c06155864434e389f7a0f4faa24606762c6a5220e380e900aa4894324707b98d1a9e399f422a622f1904add1eecd61c9cf0805ee21d4266b81d90ea577ba1e1b4291;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f19eb40680e4ba1c0f076aaf85152db4634f92d9ddd2f3f446a1cf6c85a182766ee8496d03c54bf5bdebf91a58e74039dffc4a37bcdbdfabb99c04eb6c4abb123f85bdd37dc9150add748c78a67c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb54ca66dc8801dca10df8079660c603b73f60533c5dc284fe6b29d007ec8580d40ef78c87d7526d645e8373befd8255b21f6c2841b7ac5ee666d20bc37977ae5d560d6cc7d0e11eee8cdf67a63e0;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb34c2dc82020217db0bb5d14de0cc752006da2cf728e6986a436fd48cc78cd0791c1dfa8988879c2cc332508bb9b88fc96f4ea270200af543fef7edfdb0c97f43e3536aa408ef05e830d8a4daa61;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf308131b61aa686d0bda444f4e9dd6a8357fcfc8967da5afeb10e2c14eb17442cb3fe3069e5e0f967e80b1e4883015699936a75d221a3a5cd2366065bf75be6cd1c3e33dd4280bcd769f4d8816c2;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h6cded01320732aa74cc96986efd08f3e7f9b6a3730e14e7706c95ceb7a387593ad5d2b3c3d8bf0fa26154c00953434fc9faf3a9104264842756a8ad9b1537cdb0d15b02c517f02a6c660f8dccd17;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h6ba2a3bc8e8fed255c98dbf50ea92a5e7fd53a9f867719f6d2517898ae9eb93885656640bdcaa2107a60f78693c7435df8d5da2b8fcd0ad75f343296311f17075cf85d7e910c7f44a69bbb2d9fe0;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10e92e62c90c589a79cbbaaf5751e0242774fc98fd91df23af59925c06c62531faf84bb0db6244beee929fa319f72844a2fcc0ce2c5b4588414fef7f435d407d8a66b9201797b6cabd82b82e6f360;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h92b13c7997b94393861462ef8453d862b407efa8fdd168f9831600aef225ad6376590d5020595e391ccba9895f4be90a1c38139fe05d2f6e5c5af465d6c57b10ee0b85a110ebb93963fa45919cfe;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1942adb47727c7477bf0f6934e81ddb734c1359fd75ff28de0a6c28ec8eefa6d0f2bd80bde7c09cb99b9e04c6c0451aeddde895bedd409b8939656c70d3271abcc21035164ab66a015dca5959d337;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he78717a3d0d68f22e1cd6ee9aaf71ff5fb456137c3b0d5badc7e4c2dd69feb2f04cdeb962da870d4441ffca8fc2190d614e7bdb5a37bd823a3b38a16632c065039f3878553c1d07ad17d9def69b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd13041bca858c2a0a63c147acfbcab9fb56522d62e7542fadc24a779a9fd530f4dbc9ed0577006401164d1e05ec557a5c3780e1a5886fc243df4977aa372115dc72165de7e7fc03adcd5a3e620f2;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h45e25b851b9a66dfc584c4f9c4b4dcbe518a6201284868cf000b66e48a373c01739d819af7217e40baf2192aaabc417cb4f684e3ed84fcd0f936262461df6ee148b9ac35e98a6ff87bd004dc724e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h18c637a73b3826be6ffc3f6fb74a50e3bc840b08fa938584a2fb15855baa3a57ff1f8329b1c9927fe31e3ad878428b7dfe80229baac5e1b132003e27120d1ff43c06682f18d577370be4b9ac5a949;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f08091b2065201c109504d312ca6b8ea4a0faacf353a316acb1c3403cc9642cdef3d29f4754f79ad7cbae6c5797a5a385099c2369f937f0f58d4460db1ee8537af31ff64ca3c13393146aef4876;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c6c69f6317813b24188e991aebf9477b55e5baf49eb7499d07e9cbb089a8686d6e6e45c98c2fef51fb9ee02be2deeaa982ad8072c6357b9cd259ad8d4840b3b23f19025fda6516f238279d15cca7;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h956e61e4a683ad4ab418eba2cfbdee7dd84234461dcf409f23d66c30684a18348aac614e66aeecc97a25bb4e2820021426e870d3c4b501feb2b2a2de669d34f82469955f540af5efc1b80add862e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ff9489cae75f2d5bbfb4eff8a00dd8d80839bdd9aa29ec23b5aafafa17222cfa77278d99b16b6a13cfe34988c727c06a4d4d1ddb462350466f273418778865b28077316d98a76709c9743d8af400;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1851cd5d8c14871b3a9437c93a9fa7af6f970575c8afaf74bb96a959e27e96ecff4dbeda5ff0e2fc308703293175f67db08fb6f0445aa136fd553785cd0f59a254feef4b6f9e8571621f4d3a8543b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h17374136835a558c4a3bc5b1306f664c2248d00fc0af9eb7171a3c48685edd24417cc301968c91b92bcededd59610bb264b89dcfe0405a846563dc73a592f843a1bfc1c72489c67129d41e5440954;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c2e3e7e88d3d458661edb1a90b68e334785fa1a81ed9154f5d44c6e8067b8ad58bee6ccf7bfcc07b3d73bda9f6eb10b578ca5d95a6ac9d42bfa827d50a6a31343203f73d9b7f01f659c8b0cd3f98;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h9136749bccfac2bfbc90ab3bfa3ce59779e6e1844f3a5657b4d11737e8482c6813f7f847a4d75d2fa4f38bac205ef335a1b88a6a02c3da6bcb93e9e8c8ac851fe54a052034274aa3756c0df6e50;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h8d254454ae46823737a3c0b557b8eb98cd20a97c6d58af28ba19eebc83da8934d3c423a42c682b13d61ce51a3f51f47425523872943d12aeceaa2247a0278863412ef5d06638e6b7eb1587568f6b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h14f40752f6861c47ce8553ed09696c43daafa115af04985b8397ee3dd3fca43fc0ee92b2df4cf87a5c37b4bdc7c7fcd84c947195e5e1516afccb861828b0fa6dbb9ff98a8619a561419ec1b2ecf82;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h12885fd945185cdaba288ffe32f1d6b778fdbfcfbf82d6927a085bef7900aa6cc27298401303dc57ef46402c064f003dde793294c4ef15225b175a9c73cc0c1f29469655674d995e8ca13ecc7638d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16d1e6393cd95f1ab93be7c2281d08bcb3bead4a1e2b97c1e21c22c979b6af644ba7a22c93b4fbc6fa6eee5b680b7f9157f402f9bea895423f7515739f5a56888693456e1390bc57bda0b5772fce2;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h130f077fe267965f0b742936336d5824d1775b648a4e40353e5bf373762ef0f9560cf0f27186e77f688563423cb0e83481fedcc4ebc476918e57491272712dfd235c27c13f39af89eab2619460803;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h2701b96ec4e955f73802dc03db018b6bae0afa9fa31ee164da5ea1b627806b81b17d971e4af1deaa75ffb3bac7fd8da66f0361a71c864b9b337b8b55ad95a98eb00b215c7905f9d0f3a276aaf23d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h955aade4b112164839d376539dc76174bec3516d5eb33ea43a373142d24cfcada7c5e0dd05c08a97456555d5dfd0f8f112e39ec1591698f4870c11d65a7eac961ae61e8a2362223ed4ed867d2e6b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10d5a7e3d8d87c0905cfe406c8dcbdc97de4536497dcb374dff04b337065cf4178add0521fe349ba2a67865d953401213485a7e0d1747a6bc3031186ba6d03a0b989b7be8c95265153a2b7d4649db;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1970c412224c0d8ae5a3b20974c0213e348ffef7db2fc6bff9177e1f242f8728d61e997db0ebe4d3760d6916f7dfa1715a99b86a0d9f9a264bd304446248558b2caf29af27953fc793b1188257561;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hfbd39c328192fb3c42e9910cb42882a75d54828fdf60c56df02016ad2740fef0d0458c306949ea2dabce51d4532a97ff6007cf08e1ed83b785b3369627dd6f73e86b27d9c471977f61415f8ec272;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h67fa9c17f5b8cb1bbd705ca36d21606311d79773dd4d40f1b9b38e814c8b2c75e4441e82992a7bbbbb777b49fb7c14466c63aaaec90000a2f4d6f3628708c686aca5945f13d99eb541b192cd22d7;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h9fcaabecc70c36a29bc3d9d69dd0cc472cfcb67b95db2a0aeb712957d08baab5f19ce3fdc70a778aaa284217ce5bc857305f575912129f34b1577d92bd57d736536b92dcc383e11ebc51fcea548e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a6343abf52f962b850bdbe6940db4e8cfd12b077afc60767341215cb5ad6be1141e5436e18e05988142067e14a8def2171852b438862e5071bdad79b2da33790f24cdcfda2f444bfacc34f19ca21;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f076241437dc9632ac9fcd4cca4886825ae758cd0a6534af9a6e6693c7e5763bdf977430f2f28c959d4fe41dfa2e59dd0155dfba3d15422f9c048d703ee0519d905061511bcc47d4bd7d08989aed;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h25c9b0027708409d7b07a125ad50a02a67d87d17180739c67e03409070fe3b033a810ba3e16d11713629e797ce2f4877f1e4f4e470f3fbf9ac68495640940c983a95dbdad7419a5940ed92044101;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1662c4b6776d369693726838d21dbc84488af38c2210bf53303c541fe712ca83d1447eb93e3904be4b44063e764ecb74ce256847cddc411fe77e7921b1aea2941bccce2ed09e2d9df46a32d1c0311;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h701006dc319c59ff990d7e80f184125dc5f947aead2270c1ae15e55415932874e53169d89a2559338956232fcf90e6c1b2060987739c67684affea9a378754d2e78c42a1e5212ed1c77aa0e368da;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h13b059fad4acf22b422070d5c65530e49e14a5625dcf22231256e83075723cb6add971c6fd64c71ee1071d0275fa3275b044ca39c6f4458a9d0e59b353b7d792f4815005d93760c9f8f8c65fd498c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1deb428b210abf370295aae97467dd2901136ecf4716b4e4cf07f59b320f71e509f09d4daa5fb213bcffd94671907f4fa7b77bd1bdcebd57308ce702f4403934e6a10a8c30f4f02155a355d2c0750;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c90ce76425dd1d8619d05d212a1405fdfd84627025b42d7df54d18716abbf124f4dca4408a778cb19322f5db9f75c795b0cea003a22f958b19d8b97503ce8cf5d9b53f428b7d286bc4c5daecbe91;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hccce4dbf000f39f5ba2deca2599eb27050a9bd2789773b2bec52b2be7f1a2d6d48d3ef06e98e35e8777a4639a27bef8cc9c35de72b2ea971ade52f0a44f36151060d3dae4b687156a9091e30ca56;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h24094af0dc77df6f3f45bb036f1ee8cfee18ba9124bf9e02a18622b05c90962ee646ccdce754ac5ee0200b0728fb248cc07ee8d9150b936888fb35efc5a3f6b397066a7bc8f901f98bac5c7d595b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc7411273253c2e862d3d292012fe457e27d79c959df1968db7b27791aa3ed0d7e0fe69f868e8cb3bee3fe255d114e9063feb4309f57c895e29b2b0036445942c9dc840483f0582107340fe976ac1;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1878d88180b8f62e803b08c081e09874266aef73404fa356e26cf1b6feca5d7712f996bcdff3a079f1f8726c8a95df3c15eafe8a6d3dbbba8d93dacec7201a26c985427b72e6a117831684d250e01;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h11dbdf66671b76d56696c013b02ebf00a7bdbf50ae96fecf186d44454ec3330ec71af35654ce7b7fe5238f12615016d3cfb2696c014171c122ffc0496f4a4b9665a2fa808038047eed4f7fa6b8387;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h19ed7d92a500d6b3af4ee790f8a7192aa756441c18f900ed776f60a4daf9b59051f5f49cb90a8239015a7e7c121c5da516cbf00779825cdac019c76b6038afdc2ef3401687691bd7663f24c283320;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf0119f3c565b61167baf9d245be624a4311891c82e05e0d32648ad74095fad6db6c2c73374f0bdcc25bdc616d8cf30ac58f351b7e5d9518dc6ed16f3660c3f9cd7a41ef65c09a63fb750c28f32a9;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1dbb567e37e48270a69561d1dd85247dc04e7f6ea587a3aff28a8a0b6c9c5d87b6e74594c54d8049d932cf6868c45c3128f3eb1686363a506fae41addc5c2a8b7a7a193fcd36a2f486b5b9df9ffcf;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h2adbfc8f072c5d13fc6c2760495b032dade85b2f187e61568d1286e47962911809f5d221ca49cf9602fc546cd60877964c903a083c855e489d39107067561951568415f81557d0654da1830151a2;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h15e784a5b8f90cf38e93822ff74c5ac7a8cc27a9b72f3d0b2e67e8e33f6ac992c386be57b83d6e742a554084d903da65513fc4b65e31108977c361ee58e08d66d9e72091a3938c5aa1fe520b96254;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hac1ab6c55fc8f8dbe045d5b4e500621972c6bc3ab52417a7bc28a4b47f197fe1b58663c022014745924f0865d1d1804114af028153430ba4aeb9aa1c36f4ca181556395df6813339e8392e414c9b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc9ca941b6d4812adb529bf0246a84ae9989fbe760fe7b6d6db2a5202e34ecca097c397a7233f4ca7a6c9a7ada8e7a5a71b97d4e86f98785aa023b348e10c4fe9984e1ead903926d4140459a076c4;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h17fd2f80b0da69a7a9c56eda4a26935ccd53b15dba9af2ba29c2ba119ac890543305f55d57a66ba38e689c882f7f3b6bc59e57e0699f86f4567e71a74748ce82e3f7e2d937988dad40c229adb34f1;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h12773b72308ac7f264d2b91a780ecfc4ed7196a790f1be1fcd57c1e0b5ee093dd19c66a890e5779446f39e9ae48562533f6540a4e5bf7e106954c5d370fad1c568422df7cfee60a73b4c3613176b8;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he72a538fa51952933071d34dc14a5506672f098b5b49a76d2603b624b7d83a08960e7f875d7fd022c2e331d11a8c1c8848faba4cd6ef0a0aa6e5fc48a64521db6449b0ea46557b99ce9142ea0c59;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'heec5784a3ee8fd19d79a395c0ff7f8ff35c02bb1b55e13cf597d196236996f49489c393e10bd59dacb0269f0ae5151c072081866be992fecb0ef0436e7883108155ef817ca57f86439e2c9edd03c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha3fc8e3537a3ccf8010cced0de3c83b083a330a275521e8bc2c29cc411a65e85e1fa6542e5c13464d1af51e81d450a162539c1d2980cb489aa52ed9b985dc0c749afa47f2378f2aba76d34b4d8f3;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hea558ac61faab4d8dd0c9b21807b320a4c6edd624c13ae308c9bd6d1e15dc78e4c37f005a27aeda1d1a13b4771b5dba7e60bf9a24ef3872f298e10f97782278c83151cc4965e2452a1ed9e224d2b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h14628f961386a0d5e84ba90de655dd524fecc14761c7803dfaaf304e48b7927dd843335fe6f035eece1d24fb8244035f43b3cea0a7a6fa1c4fdebd0644618a8ba137da16b26f3ab49a9c071b41857;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d49534aef2f0d85618edf33eb667b0070ff1645e6a3faf9fb17238ad3afed0d05882b4b5a242174eb0f83512a016eeb152c669ece8ff995b499c0e7c9c413a271a9d85cb2af8ed23b20a76b019a5;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he131048b15a8267b5b825ae5644abaa04fa98caa250074a7d95e498e00f620bbf403ebc89590eb11efc2a891b59828ee2fd3904cefc3e9879d1f033c8d557429e87be0d518e21a448dad4e287085;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a81e76ca9f51e6ab26686c36f76feac0022263082ae6f5b52df8d124b0ab2ca61672df1e496263cfc076718e699dd5d061d0f7f9c64f5bd72a122a4e384f406299bf25399c19d3c1e2917f92816b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10d179d99872217b3a08edd1ba6961e6fbf0ec89b6ec20b030ec44ca59bef8ab5e321a340a8050cc521c9c024e4565af0e6e5f0a1eb86101bac6bf6790e6a67bcc3a8fbda6a15965faf52f99ff65c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h8f386353d83d2f3432dc20fcc80b97b52ab54a0778c27a964fb6f2ad411e4439ad042bc2e895e0c0ea71c76b597f4508738c460d8c32c58e3ebf79a5358969873423ae11d47009d4fdb949c0769;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd998ca3d71a0728dafdad7a9d66db7fefd2549887091b9a7ec3a558221fa11bd3613bf6d81ea8bfdd0d5b5577996e07a62d5322f09a0d94e5822b2ca7e66f19bf60d074248c41227895203066612;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he10ce5937fe169092b52dff40cd0424efc5c10c99dc775cac74e8f81652fa7b2b7204ce5fef8a2b9b0ab14d9ea5c04c749ecdea19889902ac5b81b558e45497d731f69d5b03edf4259484a34db7c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1990ddbd5b96fa08e80b784d83147eae0b44fe2a11fdfcffe1d19248cb5e905f4e799991ff748629790791796fbb81bb30e41b07ea68c631e733b097a39e493d3720a5b3b1ecba8e286ac77524219;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h19bfd01cee5b0e2a1c52e2528c8207dbdb29d11bc200b050770742392eb15efa5aef07e2381c378cf12be33aaf431d5e380b00f564a1556456c16eaa4fcef8a07f4d3b202ba314023cd50c4aca3d8;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h29d91b117768f9873f56f85414a70fd5f0a809d9dd4b21a86893dd20b73a712af2e5f9f5e493564dd04c0e4b3a4fff774c433f176e9e4854d06ca6af5871b9d1e87ae4f0b63d66eb7f7e3a3ea7f0;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1fd2d7f727ea3d57d89d6e8d6b9113a43a8c9e8a097cbcdc2cec155a86c4e60d31cc14f6cb0d92c1134666a3c7f75bba4ad2ea5fa87a1ba358c0980bfb0aa7660afd6d44ef592e2c6336350991c0a;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h9a90dde08903baea072e26aeb70bc3f5a6ff49d037ef9d10d9e3fde3bd7f8c891cceeb17086971ccd7062029d82831f029af16d35fd46c1c8196adb398a77d36ea7b4bdb3d3634cb9e8c964a63c2;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h34a613c4961d0c3bf80e7c65e37e85f8e636dd725983b099f1fabe3991c07ec4278928d88b5bb61844bd8914a7a8839f0a03385f8da88c6c8b3743c0ab943c63f4d67ed47692f345d4104e2e4e9d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h152b23af42e6842d4ca4bf64e95af23e886c813c81e32aed0d73ae910719e81516bb3ca33f779bb3d636a0008dce7887d238afd22ccada056c2913543c1423f712c9a7663279225f2ad9c4f51fde2;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb9191d77161f8603aa7416105bb5f5aa544d6173a5071bd5ee67fd48d7aa3a586718e0bc1536a49c8eabd4e336ccd44816de5309ad88cf059263b4b0ee503c3bdcd53d5e80ce0ffb73c7cc27f224;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1730c1dc5ede5921d9cf7a9dc1cc62deeee5c21a53c01b0bce0440044fc0150cea1ec477e150bf32bf6574c61df4402346eec48870ea86c89bdbd30d63873ce77b5353933a7e1ce57aa9f75ce7497;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16b6c47a8bdd554c0c02fcc837ea336f58a6d5d55dc9723445edd547a33d1a1adb667a0e1ff2d064a2f1d34dcf930c56b87e51756ba7cb88264d72714004b25d33a864581d12d7d6ae7ce6079745e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h72555fdfc4d21ce211ece83f99d81cb07aacee7d9e6f7980f7e59989425cb12696a62b0a3a13a6398291ae94181b206590f604e9baae6e8f39764c1d6ece7a9c88ebd43a2b4b21f53b44fe7ede9;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he633fd75118452eed25bd6ac67e2db941d59ed9794fffc14aa083b10d99b7d8b7e09c9846c222a7480f5b163435e3fb9e153a1fa3aef82cafa8ad9854814de47ecd13928dc968e6d0aedd7598908;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1cbf1964ce968303580145c903a5c4db9f5829800d0900430ec5acabf88a57e63ced0eb2a0a239ed19c6f31b6f82e6b53a5d47084ae14873ea3c7869e6c77791854fa06deb1e0cde20b10c982cb8d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb22a6798d7f3b6021ab2ae39f92c882f541837afa2012379c0cfb9b66d1d7cff5bafe10aea0a44b718b769005748ebffa862c5b1c3573d0dbb402adacd7e10597fd9ecd1c11035e9cd72e9cc3e93;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h4b7e4cb0d5514a29db0a54ba24d802c8d7e7b1a9e5df8fd17e113ca406587e92cabcab18c98fe2df32b5aafcc504d66652e97b6a975a1f8e35126eb1d588867f2655781d9ba4b2e94c62278c9ccc;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h33e28638173659ccc81a063f75d326ce1d17382490fdc28f8ec66d93908dd652ac946a3d5932e2bc85eefcbd39b9fe13e7148ffa0b360dd0ea46069f79be37166cae722011e8c1af2375d76d9750;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h18897a3699051e2a7cca971db5033273ad230f853ddc4ec8cc7aaf36d4305296a032add4dfc39936cd1442edeb59379855fc966363e9cd643944d68bc092f52dba1695105808d8721a775c4f8b936;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h132d0980f7c8a28bfdb356411c4c9a8e0ddbfc62075ee7d00b3c0df38964e2d67f6b14c8ff3c6b00ec507191840f1f152c0458dabdd8adde9c5b1392b69fadfd39e071118e298757f104f2b53570c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h29e669382deb176c179de8921a111056ebb88f378cd199d9adb5627cc2cab81d7861ac6ccdd582a3c9a912f761c3d941cb0fefe9867552c3b273bf5e0d173dfbe3755b13be34eb8e23cdb2411d1e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he876311117db53083a870ed823e842897a9d1fc5bfba11fd25f9e8bf82704912851a6294f98f0def6645a74eea046ae48a878859cbe99d0413d1d9e05d190e6ba9b04a5a1681ddf3b19a010885dd;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h165c17dcf6d62deac16a744eb7fe35f9df2bc79f62bf21879ad1032e950c521d6a911f1a8995ff9a29c632a20f8792c3476523f31232a0f93efd2fde6a223f0c8d4ec8a55555455610c8e0b63da8b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d806905c131e379d1c054b4aef23c113fcb7f93d3d0334883b29aba36282f68dc96ef1b8a90af1c976a0fb49ee6f39fa59ad746d1c90133e7e57067a20f1746941c2afa4d9507400d18b0b0b99fc;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h86c21acde0603ac1bcfa10efe9ed483bc784ee144f2900b1ccc5b76e190d9292a8a9d8814a0e03a57a8a7db33fec2e935fe4fc20e491af2fd2d7154402c085dffc640992ef16ec5a7a730abfbb5e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf6f476c4d5db93c7bd22001d832cdabb53a3f738e5888f62d4462fa213493310e5e02e9f8f485a7f3f87d9542f41232920cb90f4e7deb88c3db87268c9a0db76f99dfb7f401203c650cacb635e3c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1839c81ade126c040a0bdca04a37d13f8a4fe383aee0186af1d33728f3a48bfd1c932b3e521e7d05a3762683329248f4d6f4a12a068ec2385c123408d93b1aef3c23ded30f9ec417e6a0e9299d1bd;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h5373f3886f01b30e7a297d16b4042aa266d34d317d4e9f7b590760ec083dc6be003d780e68f46270f82065eb6dc5ccba44f904317b259be13ae41d308bc2e363fc21b1f33045fe07fad12cc3ecc8;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a668307d7f6d96c0969586097414825d5fa0db04f1a4dce51db75acef4b6d856814d4c7d49ef272db4c6fa3b58529ea774db8465501a0559bf84e55a3b92a163d8e7ea3a7b8ab4e4718c1038f41b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16dceae52dd8f100c0aed9187fb1b4b760305cd3776a1f2c9ff6553a28e5e87cc6b611575559db297f37b02f911812482372c9f138066ce57b8ad8cb29552aa2a37a3dded98e11380f360b446ba88;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h9c16ab07ef55f5e8421eb3aec9ed5eef6c6ed3ce74ea018b80b836e9ea989539d55e907c05d656e026356ee059f0ca585fc14b4826cef94c776f198cc319665c4ff7e589b80ff93faa6c59cc62e5;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h7cc9ebf3692c00637844ed684751cb4722a827d9392f2ffddf32ae53252f5bf6792ef33c1be30c9f5385e266262e0622ec497bf22badd9b40ece8f4208d3e0d02174cbd47a299b4bf13ba65e6184;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h19ea9458ab56e0d2b3aab05309f451f88e0fcc9b6fde4047c64d81068ebbe2434156a88f7516a9c2f6ee6eb7692c4de37f8b66ad9e622ae92fcb4277492d2641164d2d262b1ffdf15822169f8d685;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16fe52e00e406133f1da75ef8d143038392795f418c154ed0d762df2221e6207145e0244b209f135965b88e696a60e52bb42104a45be89baaf73af024c814e44ee1663fc333398782369e5ea91997;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h12b864c14efe1757d381dd5aecfeeab971cfe05344ed76bc480225109b39177ec1eb9c1f838addf6ffd0f20af84cc98d4274c8a4c8540cfe04a24d98ecd01abf41ce5ec4380c633ceaef637f7c9d3;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h100a97004bf35b8f981b9a4bf8ea5014c04ad538da54fa73ef740f6fad00eca8092e201091d4d296224c61996bc945ad1780fb5d39b981ad035088b201e6302b1034ef75a370ce701b5f5fe4b7b16;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h11972b7c78ab3274569f2b4e716a47230e17679bb583649fe05a45e1d600eb6cd5567ae68e185a5817502deb42cfb6d18cc947980d88036c1bd38f525f1e1ec5b8b46c176037e26a5d4f840dcc16b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he2bc3dab59fa31a762d777365c9887a6b599d9d8dd9d49ca7f52ba741101350cb838ac831a514247d8322913b43ce4111d8cea6cfc9c73c05c858c4cf46eca7d04f7cf934785688b788f0c257a4a;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h493e9f7e64b4894b971aa8fa48aeb734aa3f97cd8d8ea455b75f3b0a5c233b8af0e4a9c8ed8476fb641cc9a2eb4b3ee9518027e42eacd0c4c2a1414e50b60132768e274bdacc102a04468d38887c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1faab493adafb99208b4b8bb0f9ce23c6cabe2e824428ee11a24a379d55c469b53fe4f2de46ce5d17d9e77e029c9fb5245374fb02f8e5ba7bc683df78fcf81d86069a1d8c52a64bbfbb3b5c3c8bb0;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a4f63729aef7b6712f4c589a148c5625a912e23d074afeff3fccba61243326fa3779d53b5c27f148c78d31af3e04e4fc718ae6a0ecbea43c8ea33ac5121ede39f26454761ef1b0fb629d0570481d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hfe0bc3cbbeb2329c47b66005ef5f1bda21f6dfe40e0007c582215096ad416a44a2167d8c40695aa21aaeed505700e3105444fbaa4a90e7c436eb05d249d873c23546a6c9254462ee9e7d1dbfd1be;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e9af93cd208bfa872e821c8b292c342edeae11d320d7f731d64c5d0a87077e25c7eaefe034853489aeda39967a90f15f03c3a1c8f720a6410cff101c7fc62ccab367712aae4cd9b1a5f114f18407;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e5948b9427c62aade5aac72fd49b64f84792ef22527af4d872d3f5607f8a15d4e12ae95ce47dc485f926ef6caac56b007178b1711b1e09e511b5be63f8ae5f20897657c29808abaac8a05468a1ba;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ef46e998b06ec1822ec4cf52caa3d3755d79b50f1eb6245841169d5078e04e0b1bbf20255b59bbe5c577628cb4129156584b6fdac013752c39c640b36ee3718d905dbee563df7d8cb4461cedf674;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h56cdf075f13e9bbd58da7e99f0a0b391c1a3a584ab542b8b592a00bd65fd9b8709aa67728e0519ba99ec900ee449ae8e89217229b01434727263d7eb8be7465a8622fb490b230f14d78084f3f0e2;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1cfeb02cbf1fcc85d99ddf49c15b5b9a191c1cde9784aa7b8f124116e92001337e08ee908787cfa13ec04ae22507ff6e5c9b1e11cc3210ac1a712f12a14c44c499e22f6d0bf10a21b358df3fec383;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he084a4c70299d7b611a176d1c75e787ea8767c002fc30857a87dcc54e39df39ad6ab663cd678b1f9bbeef90d5c607dd43f90f3b10bbe8c73b803398d0ef4c954f21a31ae598101bb977181453f3f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ddb4c3900637b4dda31be1e8f9d7bfe19f680af0cf28838bd1bb45ec03fe6ff6aca2575a37d49da200bc4e3a430fff57c18bdda25bd3cd458108939a0946bdf54343dc80b7433bfe44df3a5d723;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h62f698378d981d9306b4249a2b5be4c040bef77c3ab4640dadc38832f8e32b0789945fbe1bc2010960290cc13b13c4f0e24ca04d9f926f571bca8f3b57f64b2c2a242bc59b015617aa9685a540e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h19ae90c61e526c849c7000e975b41ad1cab34013ba86548d87cd67bc4d8ab0ca8a6c62e164c95fe8f333e3263e9d74e6e22b30bad70aa291eb635b0c9c8ef0e5d04760055ced530ab92855cbcd2e4;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a9fb6176adb1467176fcf50c8d1968b6b7a62771d9d5e0c6608c5e21a66e7b8d86dd38da3c489c75d4d07f7db42152243ec1696d858f06349ae10f7ca96dae7ff1b748764e6e795f65c12281b630;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f3397d148e28c437f3e43bee65cdc95bfbda3510fda65623c86b0301676f9eb494c5ccedf5542b5fda979e8dd8f4d05a8bb573a18bb2501bc9848290a8bef06025c9affc83b9ec05e202c74b777b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e398846b8b3255bc4994de2487eda931429658f029b7d5ba8bdbe7edada614589475aa14047ec778d015e433483c84bd63736e6e57792e4bb29987bd7d386444bcf4e4eb34c5f85996f3c7c00947;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h179783677136af40e4fc1708b5a07c902494569456d9a186e238390396da83ec38628d2d5f8dda07f52d139fb36e5885c4498c1b3be1420eabf53bbe86b9a9389ac4a029f7db796963e999d1eadf2;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e7676b84bd27690bd7be55a8cba20995ea866a3a5c2159afb02aacbe746bae16d6c14ae7031184e2d85395a1c3612369710b12fa12f265299148924aade671fbd20b04815b2eb1f398985569d83f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h71bc184b366b9d3d08526b353f85cac7ef7e21dd42c291fb4f1552c9533c3cfa1a93cdd0a130b31531f94ce1047e25f0e9a5cde2d43c862861894f48a2633736a05659435581756322899c297e17;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h17a07204f1bde8abd24b91eb2988d6cdd7e920c9b0df203d58c2062fa3687fdd1d9fe39f52b845f5cc6a24ab76861171a758eaa44436eecb4e74a17a28adc2289afd312201c9d3aba4b685a883419;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a9f93a022cc3e748991263ab8fff4989a5c26726a5e9e45f6461781c1ba7adf4f6dd2b8c2cd569c4e8a66fc79b51f261fc56e4d73196925015cb02dd07e18e1cc073193071ad001f16c7088b6d86;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hdbf55647a947abbdd38a122f66e49c2c59519d78d9a41fb43e00c1578613de242e7ba2d727d454097644a5bcadfaa9734ab78fa2aa780570b2d69891b91e5b962e966c863114815829c6545daf4;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h6660f3bea0e14acfd4728e2576956f4ca5afe0b3729efbab56c6d3a8a944a507eeab0aac0c2ad95705279483ff16e51a34b62943e0453b9de86e908d0a676113e580465611ad6fa4bd2ffdf41878;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h15ab6bdb6d9b49359e81fff125d9933f07181837662326e15e8f83c79f4843073e2e6d99e25ce0bd386e98d8cac3f01d985d3f7ca3f74d8aefaff907ec5110dc96d0c2f61a42ec7b2646a460c7b39;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'habb153863a3954d83d37bad8ad31ebe3094c3b06367a502729403823c0c8900caac50e4fd0414e7738707c976772532ff3f58e743cf9593037bc012c877602fb38e8a15a2e2bcf830519210014d3;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h4d76197297a4588f3bee1d91c9890c9e5c972180e1f41e8f920f983a6ac263c38af82eea93a97d5b58610289ab96e5420e52d4f7bae352d0de66a74def3bf1e908ad23864475c45c3db33e4e22a4;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h28e44f32ec71c3bffbd733e11cb3fa4fa4cc5fe1a152086521f839f7c3df2b40217c770b0d4ce2d6e5f599b7ed73def33917452c1d637fa022f59572ed87519acd575e0c20f5ab4ab54516d06d5e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h12bb32d88d43e210f8e74261314d018cd017f743abc211822685c27a98ee2d89e81c8ac45d8c8cf2dae9d4c01d3173b1ab1bd99b6e502ca9136d0f1dba3d8397f4216f922ece2183b8dd100a8fdb0;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hbb35cfd2c67fa49abbd856cd54fc7c2a1d719d040bfb392981c2f847d6332231343d6c7bae26af48441867b0bca1b49bf21028d75a97b8652ddba25bd3d7e283eaab648f1306231940a451aed0c5;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a49a61502c84cd78f5b7fc720e53efdd73ab5f72f63b8b4d5d16082419326ea71653c0338d6c56a5cdd4bef94eedf7437508b19f45b708309aaff18ccba54b76d31f341b5ccbc69fd3db1d8ea28;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he6cba615656ac3da70dd94353e589b43bfbe29a920c9a2ec6844d9474a5d9a1d718232cd41f52e97966538d2cae64103e8b39ae44566fc21c2dca79ac048c73d2e84423b28cd5d3ed5a6bd10fa4a;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h76271aba5e15968f2177f243050697cc62b85830b06cb025c791fc026181046504b82b9baf120c8f265e9f86a18fecefe3368f73497fb8f0f724850a785c598de96d805bd57aa29d30ddf374053f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f3787a6d27fa5334a8fcef137df0a1c7b56fcc9b5852706f09bfda81e855a34208ee5b16cd38c98fe224bab0713a7e11d53bc694a290df4bbaa617a8d232a96ea67de831b86202fceb35a1dbb711;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hafb2314ab705d5bf2059105ebf3c25cf489f9b3fcab7856148a3dc44d8261c9d6b5fc08afb6699179913472a8c9a1d3f7c6e83a007fd5f09b916a96faf11c6ccbab71dcbff5ed2b0e0644e560a90;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c8ed862e29432e9450669d8da209920c26d37c5136b0dbe878fe8e833103137d941b860cdcafc1fd153e37f853a9719f202cfab472beeb7f18116328bd5af7ae693f8dd0c8edd76dfe11363ca282;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h177c4c85656d4e20ad906fbda97e605a7516e0fdaf817cfcb917a0c5a90cc03b0392ef934e954bd43b55681c2645c573054aaab3971bb5a60eed5cde54f0652a0438552bfc6bd48967eb24dab3cfa;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h5bfd3ab78ce345628c1519a2b88c1291a743bd7c4344b52e07d8699f0c706ee735e660210e30ee8feec4fb840ab27651e3888ea7b6284159e26e8f3196d8df5bca38e289b47b7bbff97eac891149;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1fdc61f2dc2c0d604fd43009d572651a35e634a5b608e07b625e7fb3aaea5fe522f628acb95f72cfdf86a79ff6502bda771714d1d9424a0a048881b5e8d8558889a0f37d880b569e45fd2cfa89d9e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c1ab16820b45c0e459ae066a02f7ebc48b7299b13f16c0d5b8f5ddc0affef15867e8b37b88dcc86cd94a28c5b648713a5cfad06e842516b5745c1bac8415006b24112069ad9990f2c5ee995468a8;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc6ce3cde05d68124685447ef5d9630832ee90558a9ee592b2fc44421063e991c4b5de6bd634ced4a4fefaecd921408ea185da642ebe396c57f60f014ee1d42f5885be88027d04a8a7439b474be32;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hfb2e76836f31c323bf0437e1c54f3c244a685ac000fc2f11d002e4d46b5f59d6ae51c58f46dc0010cc2449c275480280ba6d46d4b3c2dd54b993a5b9f0542b7acc2e56d6f8b6787106cc70d515ae;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h15e8eb9eace2e77ba00d89990640041fcbb28dfa83b92b040b68e7d9bf5bb96174bf2b6d3417cf956a77860b96eecff477a09defed4b8ff9cd84993f7d2c994a2736494168b054d202c8281cf0bd0;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16b0506d8aec3d8e90cdd06fbca0f5f2f1fe3e1586784315616b40c3c1c0c589badbe88da2bc0ababd83bac4614ec95f2eea2a6c987ff85679699e9fa3a6471b99604c4bb5713b3a89e4dba739514;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hfa21251eed6b76316f1d237c156e6c6cb706eff2130735f617772438a51835da0fcf4fe221cacce1e8c9cfd7cfef579c4004844dec41f58f8153f50f273262db7992f5cc1486d017290901b36f1d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10b3685cc58cf8ef478c21fcf3279f8e8dbebf98d72e7ac35d48863939180d70788e5423694e8d3966b41c4b97cc2436bf4e4bf77d7c90841c4510e8e317a9bfadfeddf04ebdef42e6c7f8c5fe614;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16da0a91f5c5fd5db62a111e9f3d2fc6bd87bb03ec524c48dfd938d6c6c0a9a17d13dadf880e07d62618643358ad10d333d1c3531f3d6b47b253409d5700ead42707e4e54e0af980501f759659fdf;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1dbde4addd18a5be3190e76899a23f80f9b31b7119fca57774e4dc97cec02fb4b7e861a55864c66ebc1f09d59ef2665badf18483d949e63b367d6a600661ddde91f295105fe1a2a28f4276c23ef1d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f3fc994b9d8da56de5337c6f1e5e467178312005c75daf9e0684e93bf1b46b16700f4e164658a3dab94eeab48d3aba533dd26e679c1454a6c0bed29186fca52bb5224f198250459530bb2e63e809;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h6d742c877c8510027f9b1ec5d37dd94d788b48671a91ccc466263a84d62319dd5964b540a25593c95c9da3a0799b3db322a89369ff0f3145ea5c496ed8f19dfbf584ae778bde6f6fa540b40f9890;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h3adeb84c9b86eda5b27b6eca17c8396bcd4e7c8a4e9ef5828698166dce4930c054f675b2ccded2191da64bc56ebe58485eda4d14f7f4a7891cfdbc5e6562f4ff2b7b5391ce73fea022216033a035;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hfbfcd97ab52b44722c12020399530d91c0f67ecd73c4ce95eb8022da981ba7b5399305ae8368568755aff8063ec7cf763cc00d9d94343fd8a485813c3a27013246bea3c3712cf5b6becbdb08fdee;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h14d31da1ba1dbae5dbdf5f5ed6aee61906bc86b768d429a6c65e9a69afdfbcc2b1d4f62fc9224501fb0a344fb38c54d1a22120e28dd24ad527070455e0152b0a6849deb45e393e9b1d2f20bc84fdb;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1308a6bf3e8c89e4d74b63896f0e64a62e517cf9c11c33cd80192a4aea2d9d2d939c81ce12594edff08526dd3a73512b0ec46f1eb15c91fdbde7cfa76418e65ac63e23155088b83b615c111731668;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hcb094deac81a0a727e8176f3df8d317efac2567946cbcce0796363ebd1509305276a71375364f24cbaf841da7b1dff492294adf40dd8b82ca6dd410b3e8e4a27f52c8f0186b943ec5f2e1822bd7;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hab45b9414a822288b3b2e5588ecf78639ce660a483625a160f7a1ab29f8f782ae3326bef36388a5e5d0b0ab5b1b35897944a2bc54b5221481968aef6d6014853b72e402e14bf9a493fd0165a6dc4;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1764ad6d938d0201e6a95d569a6737fb1fba67f2e0d0bcd804912933bc1ac2f7894215e91435effc14d2d15bce3520b6b96f911bbdc75ef214f2a2c350d4a569c7e322b618eb6848abb467272157;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h104855cf74810d0279c13dee4ef2392b967ab745a2c7f29a9af1bf3c7792a086893694fd570c587e3ae6b89907679500664b11fa963b051c2705092899ed8116d4a3ae861b51eb88e27b81cd2c984;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1814eb4ce913415b186ed869b80c8b7953e7025bf5a09838c6f2379ca452a5bff551b696871d202f3ce41346a4be5c07b48120b9d3705c2b39392f68c6518b1c612707f6e4f9c14ca39decf6bcea5;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h8a464c385ffa75d9bac53ef2bef611f739d63dd46c097bbc5339729a7b56f8dbda0150f32bfd8b58abf02032138544228c9228790a59c6ef69a7bd8640b131a1f3da86a6dc44b6c3a4f5ca824250;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ef62b7228bbe0b9b4ff968f97a5a497e4026d721733af93c67fd1b631bc6c35fdb7203b152565f9644277ebed764a075fabe9d0645284eaf97bbd439bf88561529a3ea0b6fb1f1c1a76eeb8e264d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h8dbc134cd7e5bc5ff8c88a38e750644585e0f4a9ae0e9828645a5fcdf1825955da423adc575d5e91f435b3733d3118151bbb3b3b129c44126571d6401caeab81e2064acc0a6afac47989f8f197e1;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h18e719d72111a5d1fc9679337978355fe0be014fee16f5f2178567357a4c25121c6f948b565fb14a17995f42e2f07bf1a620ce1e80e7a845786cfe911ec75ba5c590348b8a2c3b661abe3cd8b2bd3;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hdee7ffce3b854751c71adf57641a3f84c617c0f1c869df830c7198dacf4800f1dca11876c0e39aba9698b4e757d22b60f2a9ddf1329697ebb3c4d6ced1b77d318993de9700d410074025a1d2b535;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d1c80d5cf37d3fa3bc82a38337ec1ce42c2258dccadec74ea5f3563a6f4285adf387094de33c5d4d3e2152d27a421554c19c49cdbd1d300e79cfd5949c5f10fabef298fc07effc4680c837a5cf81;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h15e7012877b0c0fbd5600901dacf89a4e960cf05798773b7539650ba5e90bdbc34c5260e18c4991e1b4bf3e4df90104f69bb8db59aacf820ff465f643ec9832a76a955d2b2a6fdfc35335714eb30b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h119c72c59b67c65aea88a5f518bc2c67e4557d2f110eabd74832895ae905f48023f6efb000454fd66f19b97e8075fd12c957faa7ab8e2b381dbf0122cd7990fafca087a645327b57c54cdce505c57;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10dfb7e05bda86933ff6b44c09f38df3a5acf526b62d18bb83c8471a1ce3fe2f61011b6a50778fbd221457a012c7cc15802156b395a3325f92fd445126dd104e933269b3d72137710810bd4abfc4f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha956c8cb582249cb432597a8cbfe1697928a3bcbcb19bc91f3a6197cc3927c5dcca4ab37901aa09c82d736324de54ee00b1d18bb98da2fe3e4343e84587159a6bdf56a024f0cec033c26415607de;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h7e6692e409996ec78b17124d3e8dbd7b9cd6e17f58426ae0aa75ea9dee1b332c72fc3dccf0a7e79faced9c037739a3572876bbebf453eda9a393fbdd9c92ebff7d60f59e3e0f7e97f7972f04f499;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf60d8430d7bab98bb265ba616b54d813194975c3784de92b1999242f0ee00d84c3151104628e8b0cfe39be825fba6d6bf5334dafaea752e148271e82fd79cde8c0362add1c7ae7b3b6221d9a79a6;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hcbe5482a3d2d9d173774e7b42b216e7590ec8f736bf3aa5e6339f02ebf0d2506c17ba72b5334e19ddf4579efb70b21e7dde428f1da5d1a8d02bdf3e28d080d0ae158c17ccd415493bcd196ef2bd2;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h136e40be698410360b72b9d9dd81a6fef2dd13f57e9a408f5f45c26d3cf3487cd44c7d65b44aba83ca5d404849743ae302e51f0a5b619dfb9e149e56e3cf6b2fc01f89a4af71a3e9c63d8c0a5a183;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h179989dea83e0fa105b7a3cc3b4c599a69d15e3ecfb3fa88bd65a1663b8ac47e82f0eb1cff676ca4ff2bd73528182b08347330ef279ee277178e58a742408e2dcb3c32466144d0878cddbcdac022b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h19671c73936ae4fc9bcf87e640069fd055c130f1c7cd045cee2387a9790b7120144a3bb8b5010fca5679796c79dd9340a79e6d3337d9c4c76279ef0b29dd9bc29acdb0c0d58376fb3fd186e1d678b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h18212cc46e6ee98b9201587738697830273be1123de5839ce9b6ef2d6e323b5d80da890d8166b7455ad757b557e426e2771bdf8dadbf7b61591af92ce33cb078dff2bacfc21543ff0cbcab34cd81a;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h987820cd6c53ce47ea6560fd239ccf2539a58c66432fded1182d3428ce80cfe3950d0d5e1dc2004029cd4938719fc5445350f55fe546b998ad3d352148842458a05d03071a704ae9a85fabc2eade;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h66686be0817dfa298a361a601e038f3dfa973026d1c778a39a094706910faee7f81865af820b1cc33cd9f844856d428a0c403ce372e93be26ff93e1e294f1f7d6d514c69c4d77a2dc127c0373721;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h295bfc4c33d6dba41f99a47d3975b9844c824d174a55269eff4a62ded3a84f32356dda95f4108a2509c426b0d6cdac35eefa672244e12fde3ae28e1ffda176bbcc3eaa736cbba0c5cdf5e6b0941;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a2c88de2dca323dbfa7a9abb4df3b69cf5d78c5733d893da3d1f6c11fd694ddc63913e7e95fbdf897b05f72a8e39f75e21f1a1bbd6064a6defac33a35954a6d3b20d42e98aa71a82efcb6eebaa5;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he0204cc939256d7a6a801d53213c76d0f882c32ed19ad1cf2304367e5a5d2784b29aca1985d5295e7a3dc11560e3266578ce6ab38d2db6a7fa956f2060bd43b949a72ac69ae9a0f5f7ed3ac5dec7;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h177dbf69e1394dc0a366f33c6d2f0eaa0d4080bd8206f1f1329ad85beaede3543975564a0fc6186020434beb093f309ccbf90e209566aa818bd58d0c8a5fe571245b6b4aa2bd164c72efdadb3eeef;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'haebc1a2645808a51cc8d4fbf7ea6b20028828559808d706163d7b479d65adb9ac72f67c4e2e5e17c2411913dfd5070c6b58384e71a89048626eeb406c12a21968bbb318405c00fbd30733b8f6eae;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf03915d5a65011d797705f56ac4742270b2b2c1f7039967b671f61497d918f6de9b507c9bc33bc4fc167e258e851c9f6cf56055aeba16b197fbe6278df2752343d85cb29a9491980072c9881a800;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h87caffbffaad36ab8080043d0c6c14b244b64fccc03ab8dbee7a7c2b67e5aef99e4a98e118d2567ec8406016c3f233a74172669f2ef9145e5bb0843f6d88250e3923c05668b3d8bb31e432280eb4;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h131110ee7f7a8f18398e1ec2608671c9e13877b616689c4e15a8aa2b6db185b714175039da310198cd28f84766373abe57534c457850a87bc6387c6def7db93cfdb1eef4f56839748ca7d5b1335a7;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hec4ede082d51e442e575a8d6093b7d596c11ffb91d2e6976dcadfa880518afe2ec09268e24b1df676e9b4b59a6a76f3312773d3c3df7a94285c7cc95133ccc42c452781fcaa382ba1581b547441f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h13756e5cf2c1a68336152b28b20b55c6b09bb3b68bc01c37f5d2c69c1cc0ea057a8d4aebc2a5ba3fde470c943cfc02c9cb06083fd3358dd059d6d773e49efb39277896db25803713b958dc811cffb;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h15b970d6c7521f0663308feac591a7bfb7f22078a793b31cc883ece5bc0bf27331bb85d30d188a3a60a6d5c2db353b26b44ed326b857620f18bd590d363df93a2ba214a325bb63659077a47cba3a9;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h17f89d24c20739a0587de23731df7d007fbde1111f06e1cccbf7abdb3897ceec713ae43ad450ed9141a059cf9db6a775b7021c2b81fef6f7e74c6a21e4b5c2594478b5ee189ec90dc824af69ce1b3;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1348b45f602bfd2e1f104e7f080b7d5e10926c6683c3cddc0d21b1722a0e0438706fdeb66375445e1b6754262b06cc9bc6214b37503cf14bd404964724c811f2b0a93bb1e41920a7e9bd7e3e400ec;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h3429410b687bab0e82de3fecb68a12add3e12463a43cbaafed5f6ec24865986945aed53cc2219da5ab866079df6648706e9510b2bf22febdca128a07acf5130fbe4a29d4d78b12774ba49ee2a83b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'haa43a886a58248e0a76a37859418968410d67894aea255963dfe38f456daa91ff85923045461e94d089ef8c4d17a1c5c41ec1c7f14218707cde5a76941be979cda6e466390a47a7a69da806d6425;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1457e47591d401bb2965e5f4c16b127817b5a7d5dbf6d8946e215d5061ad87d6381ac5d807ce0896e03df6ec5c20ce23e1415156d4c2e2c1c867ba8dfe2ca7cc677970e6987fc0520af3cc7b87d11;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ba6db667377891b7022af39a5a3787532a0e8fe47513ab626716267e034c4cdb186a26058000a596674ae2b19adda6c6c1f6ad90e54e85f53ac3dfac33f2f83a927109fb9c37c09dbce8ca6f65d7;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h102746f61c1171338b15d29bacb71e22caba5f40b55a18e345042f0654ef8a3351e2597e2a57b5d99d9d4953b4d05b2ff6ccf1b2166a2c9aaa74e11cf38070cc21b604fd64936074928c3403f8402;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hbfa50303a8a974d930ddfc9230a9b2de38a463315fe2ab31c67a862e7d2c810eb84f7093955213c83f6f231ec14228701ab57c53eac76987a740a4e2e93e40b8d1b52ffbbfaa5d39e6ac97e24dc9;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h96c235020f7b5892d146a4280fc2e3d2bb0b80d3b59560f2a1aa488f53cf5a789ad8e622fb735c1e4f744b43fb621fec2fee9d8b82de9574c4bd287a8b840e35eed3c864752e536a715284f8b3f7;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'heedcd77b42a24175b63e7799f8e2700e0b32b3c7c814c5c0ccae05ec16efd545b711a2802f33bec0d055e008275f57b66d876a0197b09ef38f41a1ef136a01d14c6fc1d6ce1aeb9bf514434997e4;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h746130b3ca8f95fc493520fc51038be5594e6f3012351c6859d5b588b9293fc36a1bbc5510ccbf432bac2d77aad44aefb14c155736bf8c944036e8bf4ab963192e73150b87d4ec5b0a78b6d85fed;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1cea1525b06178d0827320b9b5e11778eb2ec13e7576da63d2b7e825775d78a53de495bb55553ab48cf2401287c9fdb9e5d72645b4b542ea73f2c63ecd0a0b032565cc7ac823aaaf2a1938e465dfe;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hada93af85e0adb3b180d99adec9d01613110910c2b099966d3a27459a5f492a01ad1c4d8dba165e08ae0e21682622f1d1a895fb2d38b753adc12f3cbe41141bf174fe0c54189957d433e274db428;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h95f42086b77cb00e1bde641f63d5c3d85c62239322886da520913a2226ad81e50f62805222b54c243ce1236bf1a5cd2d49f6f55d2240048d7088c1d5e466345c44bb237200e7663681edf697d3f9;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd29f3e1e55f012dc3a40d828f936501b054ef294aa57a91601bd1833d62aa9d24e69aed7881e44e61aa7f382e67b6f5075322851e28811bbf5680d499b70807d6e0a063cad16d9b099ffe36a188e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc4ff0ddc78eb9efde0d63c3ee6908bb1b9b0a06c6f159f135e14ecc33db2f37b4b13537a8f018f157b4619fa15e8b46bab94c326493d7922c2d50d941b6df567fd5f0dc1dfcb7d0109210b49e89d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d45bb0625d59103d7a4c2d8538b3b85d9a51dcc80aa1f4bee682d8d40ade122debcfc94f0ab159ffea491195a8a80c068977fda947a691cea7cc54aeb98453440fd6bb9518cb86775d2d2c9f5b53;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h594ea7d6467a1e070cf4bfa1a46b88d95d8cc6946c2bf2b7767a2b830a8981a055e5d8b54d4c79541adda5807ff7bd6f383972edfa061c570f5656def813c95d99c7d46948ca1c82546b76929100;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h19007ccd166f00f54e4cdeff3008198e34ea2430acf3feaa4a2aead38cfe4538515425bf74fbaf493e8af68d695aaddbc772eb40c18b070f661552f90fc8c219c1b5bbca89a2a5052a839e837bf2;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h3cc8d7fc5c744deb371ecfa9751310d60a1d88182c92ee7d12b775c9512d6fec9690e28c6c0b2b804bc93e8f9b88fccc34229d080ae9e782c157e87cf3979f5551c95b4100666337d00303ce84f7;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h46a8cdd3a376115417eb1d21f72603ae3127355bd3afa6106263acbf43061270700159fee1ea86a381464a36a1e31beb3252ed2aef8d9ee28501175fa446e7a6dd7ab73d4d5ab902eb47e607d91d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h50b31cdbc15cd7902b57a8e924a777f009389345059612982dbbd37827ebb2e69a6a5bc2d7ee869cf5ee828368fe794176bed63dee2a0e4799c40179a0d7842a4c49cd95f87a923ce42aad97649a;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h11419a491c1f3f024bdd249e275d9ad9a3b03105e46ada08bc4cf2b5ee66641c78fb31dfd0827d810a5dcc1246ab076d08151ef32bcf1aa53da716a32562f2c46af1b03de4e4887dd3e555e542863;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1887a128e92f715341738b42ba677d6c6805c2381309f68b75cf361b78266cca0f878e8c1cacea89eef7d372dca27ca303d402143516c33046ee6431ae2ad43de48cacc68739a9c15911a3f1b63b4;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h17fcdd5192278f42af39dbf1bb2f2230ceedf2eeb941011e301d24bcb17eafa711b0c9f2af115f90992c66bc26813d42b11338584b6f96bff1c19eef8c96ab1a702e003ac1f48a043843dd22efb62;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h142f263fdbedca236f05a7268abe09473a5ce4c0d451e40434d9f79bbcd75cc178b157ab34435feb5a498a9d19ef6aaed447e2683604c1a94ae8fed4f70b5b2142e1d4b0e2e6178479187c41d620;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h9ae42ba86848c55e6bbc3df8476c49a076b105f9fe027c0b868fab65a1c8f164303369d0b219fbed6b7d19ea67a8b0d1a78eb82fa67f84e29b21b9c013aa05cd199f878449460ee5b6b5f5d3ecfb;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h3c19c4c1972da15b84dea305e5d46d9238d26ac994c7db36b8738359e95632ed300e661f6e2f249eb933991b8c7988664d56c3fb15f8c12d687088b4b646b020268a58ac4d5920d7bdcd0fe1ded2;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h4ed4cf699b3642b33632e6ae44d38bdf3d1a33c2ab3656a79161c22faf0e650ba4390d324a7aab8ff4f56f7d9097405ed1fafa95f5ae449a948f9728ac4cf0c9143c9327d333c8e00dfbfc1b39e4;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h2c5041c333a405e2f16a7cb5f0404bde639c903f6110c4e5dd405e357a6a096c8dda869df03d76034ea6aa416f70a940757926b6333435650015557ff9c1a9a49a0a589655fb58f6f778942fc225;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h17dd557491d5b91e965de5cd929bbc0f247e2cd86314c013ab1677e9d08e679c96fe525c7ecbc81299717a883be88ede031ca4d1c33b800dea4d1b06dbb9a8b422bf041bd90aa7f57a5c475c8cedb;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hbd3f7e6946e4f0fed9e2c3ad86f006a1d9e89aa47c4ebea455ded9b37711dd68d11befa4b9b3601ab9373614731c79f553e058efc842225942718ad3a71dbd9f8687fbd2e4c6c3f0597379801a56;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h17b23b3c765a5b86e67f384d851427c550e45f9e259868dadc8bd86fa9073526af0088e219c7dd7eba18b4b6353bb39b13001e8156873d394a16214198cc6552d808fb80f7a273ba25c561852d593;
        #1
        $finish();
    end
endmodule
