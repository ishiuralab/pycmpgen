module testbench();
    reg [14:0] src0;
    reg [14:0] src1;
    reg [14:0] src2;
    reg [14:0] src3;
    reg [14:0] src4;
    reg [14:0] src5;
    reg [14:0] src6;
    reg [14:0] src7;
    reg [14:0] src8;
    reg [14:0] src9;
    reg [14:0] src10;
    reg [14:0] src11;
    reg [14:0] src12;
    reg [14:0] src13;
    reg [14:0] src14;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [18:0] srcsum;
    wire [18:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13] + src0[14])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13] + src1[14])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13] + src2[14])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13] + src3[14])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13] + src4[14])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13] + src5[14])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13] + src6[14])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13] + src7[14])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13] + src8[14])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13] + src9[14])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13] + src10[14])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13] + src11[14])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12] + src12[13] + src12[14])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13] + src13[14])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14])<<14);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1ffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hab768f03ff24785a52f18ae930385bbc98d1146a1f3bc3618634c43d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h17d101fc30318363d0f8b0ef8063d992107e481172459d81037af73ea;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hd9597d80fe23f000f97f87502b2e043cba42d194e5d1e8aab868609d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h2465e1313cccc406786ca0f01f3e846af5431f1191f6a835ff26621f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h6467ba249dc469ac252d1d24bb742552887d184fde88b9ea1f41cd02;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1c22ef3c0d3005608276910696c255417e136b4724657d06ddb92792;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h19af16a0173a73b917d96b5922547043b4daa8aa0a0acd32a0605d2ee;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h4cbe142d221d089410b0b0b5798c1905635b38a2f53b2d8fffd900bf;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hcb2bbefcb12de8f102746f511c57d14cfd12ba7a84e10a5c0336d05c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1b43320d40bc743dccdec138453b192053e630548ecb262f64725ebaf;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h38c60851b721bca3e773b9e772379a9f5174b49c1295372673862343;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h37bbc27f804ef2e5cd50eaa5effe846b82c73e413d0c7d5f4d8b2659;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h90ae7655dbaacc2d666788ff1f0b92c503daa3e3cd1725664ff61326;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h14aebfcc35b1cd34623c4a6c683d873c7b6a39fa062f5b1b93ae05302;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h5ca2e0abe49b08ea1917b262baf5e2ec0a218021bc702ae113a623e3;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1e1e219c83dc4cb3dfd220b89988cdc41278624883e8ba1cbebb9ebed;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hfaf13072b9a2b0ab765d6783059597b039c3362132806d2c7d42ca27;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1ca259d711650b0dc335a7c022f17ca974000a199777ebd12934ac88d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h9088e5304f29dded0adb69ddc593daf7cc206b293c9c067150069d68;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h10edbf38a115d7ffe0983902810310f09d9455e36d918afbf9e99dda1;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1ec1f462bb617e5437b29668f8b5173b171f8ffabac9b493c8522b8aa;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1108688e6f2bf177cfd7b3173728356c7ecd0a5a7a6ecf0515d58995;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h116d71a7f9d7d7fcc7b1827b5b1c2cd6067053b528c7411bfceb607;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h13963eaf9ff418825f03714aff4d487d742e10a32b1e274122c92518c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h65dfb265a2bd86d1684f9e15a6569ee4d2b14d44c9c47a8c7ecb22a2;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1c3aec4bb98086eb91e8d518aa28e9cd7bf6d068b8cd9a3aab7cd3bb1;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h2ead3154c985c5444de5448629917251d5bac363a34cc18bf7562021;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h18809c1b099ae17949cad0aea0b8a8fe5861eeec46dffdfbbd18f711c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hb0299c98c21c41100e7c77a706ad231f9582603a6f60b0bf59accddc;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'he731756e8b2506a3a8c5d1314cba64b9f689b34ccd8884e988b301d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h18d8f0b692854429b6dff961f218689bee8b885fafc9bfef34660aa9c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h98f09df0a1e75cb053920542a1b41dc12d477aa3770b7a4bf1750b9f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1fd3b1c8cebaa3249197e3fa10b0301f5f15f091a1fef41da0bd6cb4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1aebbf385e2f9311b940a40a16c5efe39249058a3be8a2b59d275cc75;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1e2c6193869c4dc5cd3200cf123d80e9d8dca4a303821d827ce4d7ad8;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h18c76766967fccc7405e3a42e0b5d6a8020a2b125c223abb0f27ebcf8;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h127c282174ae6ae8802cc3a69a0377695bb9e54a82c4e5bbc54f87fc6;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h22232e7bfee93c9b47839ccf2e6195c57b139c8b29c737a1afb040a8;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1135f6f299ff814e701585405b0e3fe405b757be3b1a0e79245fd8cab;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h198cf0715b408742814643e635a8e859092f09e7a2ae87659349606a1;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hf9b4ab903c5c235702634740abd38195f15cc6f65f958d74b645defe;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h13ce57fe74b9980c2fb0b4261c8ac0ff38f838693f74bab05a639080d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h62a5ff84771857055f3fd77aaa0380a2dad21d53b646a5f34baf052d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h4f91c53b562b18d48c8b98bf8355d6a511e218a38e4933eb0a832c0b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h4f1757d840c9035bdf9d54c19bd135d1747b476ccd6ff17982d3d2fa;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'ha29a36f683ae509a27e369ccece91bbc04fc8a37802c71f6249e3de3;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h98a08ccf48aa2d710814391c255facb5d598cc9fae6aaed42e42e236;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h526a1b876d1e9f1aa749b9dded9abceb6d201a54c1f4bf2bbad52850;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'had69538d119b5fecf023d24406e5239c9a4573db509f9cf3c857b702;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1e86ff94d16956f8e0939d24c7cabb8903644232718fa13b6dd4fc7fa;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h2cca34f2fa0907cc068b208d81a4149d867b509d9fa2236474c02832;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1bfc76c7731e2b5af1cf5a09afdbd6ef2117d196cc338f8df34c93820;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h36c07a48660c4a0f5cfd10b7b7c98bff8fa250d4ef1e9c3e507ec918;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'he48df94a8e96cfd697f28a57cf723f59e9f84778576955183a7231b3;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h15623e616ce16b5f3ab696be54bb31a90c50de66ae4fd136cfbf1bb04;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h23b8b918509e09c5174079e025d5c3cf821b6dfc22203921e30cd268;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h5d6f5430841fe7da4ac70e8ed300ad49e8bdf78fa5d454a25ee2c8c2;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h13906d9ad158438d18c109476335299c25162c52d11b7e7107f86d140;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h63c8ac214fa09bd09c8843b068410cab18d743fb837d58f2e4823b19;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1ff7ce45eea998d66566a995d807910120a6843997dd2d4173681d961;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h18d225225fb17837c7edf695052d9ca372080cfb05e484f88344e2173;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'ha17d7fcdc32c4fa34c436a3c5c44318f562904628372dfb43978d25e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h16e8d9d6312ea9e44702be592b6b92683de34819b5c546aeabf3bd900;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h916b4c888d129a198eaef77518ffc068346bbf74b479b322403ec361;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h141c53296353d811742b389e2c385368afe9f8ff8584131f8704bfe17;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hda55381f6bf3950ee447e749cd987e074dfe5ae420f393200646a9d9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h192961d1c1213fd46d4a4896907bccfb55701ee7fdd3a71e93fba4c3b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1adca4d3c70277265054b441ee1518580afd05cda1b959280f8148e1;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1851cdd9514f774c802ff9fb19dc4b30b7ed33d5e86f7f14ffc4ea0b5;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h60ced89854984137db686cdf3f4800fe0d2c2df68def44abce1d0ff1;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h164e3ac74ee843860566ae71de05494ab1dc8285ec7cd653075d59f6d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h14d1250459ee38c98a8b42a1e31dbe4517b26b7662198a4ebb7ba4bfb;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h24f03498891d4217a47f4a1ecfe00e9edb9e3e519e3118e654eca974;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hadf1503bed69fe4f740227acdd48a9ace555722f1c15562a4ece2065;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1345b6bba1062d10af6754bcb782a689b32843cb48fc64cd0f6d80342;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h664b0b153b7531cf23094bc7cd92573a1135e4d14a0cef84eedf767a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'he2741a65bee89876a6240392f6fd416f769a1d45d3970f2018a81b15;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h136cd93d97506ff19433dc6d362dc02a1d9c82ff9b01e4e0b54144411;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h14e3e8a3d45dee54539d034e4d2ec9a76827df213ef0130cec7d0cbb8;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h88666d0f0347035999fc2e73967a44b60c1f46cad521131eb013072;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h10b38edd3cf369d140d9ebf6459bc6e010459a8bb4f7b050b66c31118;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h533cad323fbb7ce8b638df4397485cc9b02d4a49bd3d277f3243c562;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'heff7dce57e6e46d164eba1c548252f688bb6917f1d6b8bb6c65118bc;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h102afedc43c529da49d2c1483b5d3d7eb4921dba7e1d4ee53d82385ad;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h2bf31796c6fc27bb20587f1bc40fa70d5443e168da3f6bf3aa10cd0b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1e62629329a4fb4ad24cb76e6ac111c9c18429a327d4cd51c5b5885f6;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h989be5a31fe8b1e05f097244c3b92d8ddf0228bdec93f409c449359d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1a50461ac7a4ba5da4aa835f40a7003521fea2ef07bb4f68a5d707038;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1661510a6a8de9c869f1dd3ea6f60783f0bfb9e0ca7b6b8351fda7008;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h3a2e6e6d763d34ffb7a3868907a7449886c05a7a014e5a9a6cb08723;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hc2a9c80db6c2a0701783a3037566ce2ef93e778dbf46058195faea55;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1c3805fa08713ee65cc5a7ab4fbd0acba059294c1808ef98c0fe6a449;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1956b0c748e5859863cd7014242bdd70b67f67fea3c898dd3aea9eb90;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1a6710de7441a8f14a2a0daeda2af5620176a02eab040d5ac1027bf37;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h8ce093b4051b7273a0ac3e0097fb008bc3202105b33ea719b8824c6f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'he92c25f0eef33d1a49cf76a896916397bb0b8193b580a464d423a2e8;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1f915fd98828af2f3a502d18a788b6161562064c8e4d88ad2210ff9cc;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1e5b26fcc49770d7417f966d5b62bae1ae30b83f5ab20d46ef991a147;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1448c6bd339eaa8188e021aeba1ba039ab93524e29ddc07edd4a9b1c7;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1e3d53e510668b3f0aa163fc1ffc3a627e224cef38c003996fe2ae356;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h55f75468e114edb826aceae24931beddaf6552c9027858cd4a2ed34;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hcf96cf20f3b4a39c7f536bfbe076a92f1b3e079a2691641eb6c90637;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h838fb56c557a7bf027cd54714faf36f898d0e124bc4e6c3c3e806b86;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h773d80d806f6754d1293eba66c55341f8afddee89bbeddccd4f068d2;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h151926c69d3cc931810edfab644f95c1cbad3e56320d24635e9d2461;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h194b1999d1d4b12919e46e6f91891b4d5de175110f9116a64899061c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h61fd35d712c05a94cbf3d410a3eb282ea660cd13e1c81cadbf25e1c9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1ccc4215085fd88fd4998b6c814c6d7ce73da179754b2f5b57d0b7c00;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'ha8bb7fdcc2e4d0dc29c8fff22cb0fee9a532f893096a30741779dd42;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h5465e62b893ec8156648cfbf8a90b1a814824513f0bb6f70c36f050;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h5ff13719f867713b7954c423f1f1f3f90c3cdd01449f9bbc8badcfac;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1e908df2c3ab6eb64d00b1a76ca9e3ab8d276106191ebf39f5eab9343;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1d8ae92e662df011bfaba6420442e5fe8dcef0de80625eb8f574fd5fe;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h13bafda50e42934ec61405f32b3a318de78c20cb82461633210745108;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h13a1262130e32bb5ffc5f255c4aee3354e6b99ee79dad1953b6213589;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h5d3d9fe82200177a6c5ca9433b6c07d4c56dffa1b396d0276ad19a86;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hf61ed7eb725b1742468e92b97898ac4f94b584a0002eebcd3060f328;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hfaad1cbb1fdbf1b3ab4a9868b1109c854d20a9a9b364ae844653dfab;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h9b9cab21674ea6a33a909eb9c333b26d00d4548f71ef85555f4f307c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1e0a016d15e5e13a388038fb3d96dae2c49def25269be9cc1bc7d6ff4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h51e97cf47e488ef46419b580531d0282f2c894a12c9c8e8d67da7520;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h6ff84d45f99207b9648da34cd8e757768e592928edc38db670290aa0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h37ca2efba3f770cb42e5c219c5555418fc9f2ddb8b79140247af6732;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h4609e1134e6689582efd35220b6adf546af8a9d4d1f825bd77a3937f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h4012a90f9b935a9652f71ad4b92fda1862d93cd10e90831a8b9062f1;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h12aebf7f1210e916645e6dca12374a4ed589816b57901c2198122e5dd;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h7e0f8823a85be51ce5f19050226bc6e3f2fb49e4629f988cb0ccba6b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hd15e840ab8b47e40288558fbfbe2ace5bf79342da661450bbcdf8d56;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h8d19cb63a4ab670fffd68928c44935f54619c35242c3593156d29e2c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1f183aad2046df528e709ae38ef978e967b95ee33646ba7177f761521;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h15ca93eac990638885062115f1d8a0d51855ae000d2979b5ed6345fc1;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h129d629f7540d85436019f9e9b4f20c18ae3241ff758d00bf8801445a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1d3cdb5f880bfb94ced21bc7590e4924e38b41140c12de42bc20ebf98;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h558affaa0ebc52a72b73f19214ee80bbfb961364309dc279767cd374;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1ba159f55d76b6d0a0f77235e564e17bd6cfa782338ce0d92657d3d89;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1ec018a32b1911d3a1bdda189ef4b6c4a7b4bfadfc2916b0efa23917e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hb04201a4c1e8929d963a07a86baf32cc2f48d9d116c207e03088deb4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1bfdb6d9ad2b310b69e774432a62febeaae0a3c66087ce54316afd5a9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h824a62e2c90411e4a77921c99b56ebc4522ec27b98125a80c3ec5c72;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hb2fd266b9e6e242ed8064cc361f9ab1204c059a049f98a0a6c6eea79;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hf9877d06654ae01bceb05c3f60aa59c4b87f39f365a10ef973a29e63;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h12d639dec07b6fd7bdcd1cd5bb7ae57f949bceaa3b6ddf7e4197ce7e3;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1c6b11d74ae9e6081d46e1c8d8e8cc7f253d95ecd2c41a48cb2933a54;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hbb80106a6acc759c8000bb151ab8a8e9c7a768204b6b2cd1a1a0a857;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h18730f32c501b6ccbf67a9098bb91f187a401cd28bb222f8be23f1915;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hd1f6ab64a6c50c07152cd4d03ea5d8855c217437c748b5edb9122981;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h7ec4b1b9cc0382a28834eeefe6f2f5f121a34413f569a779ef149b65;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h127a21fe2fe1fa28215f1f56a9f6784b144c4e7f3ea5bf91a16dee92a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h8027249332a91f4a4d390af7a1071b4a9fe252d6bd7955592f443de1;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h17837c7d811baa65a6daeb3c6be047b8cd3d44e5cb9342d6e9c0bcd1f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hcef8ac0f54c6b4f0d30942535d92e49b4c6e9b8264056f12537755c1;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h174d1f85e3707877727966783ebb8d995386dac693e90c0b31793e3df;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hdb2be4b4492a7ff2ae93bdf4fa94773917dfc6d7566f17482226262b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h3a1c7481031ff5125a4864411ad87bf375a2308811df23ad276783d0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h12935e903020d6f0cb61f74a084474895e3f7f62c0d88d088b06f0c62;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h8a6745f8c09129ead42be5f459a765025c6d3c3b07effa9feb88826c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1afa4677aa4445449eb4896f61079aae99c85e182d5b8c178ff66f56b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h12641a14e409b4443260e3316ed8bef87a697b001f82650b996d55550;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hb5509181c8e9ba3c944338972b0044ede293f1c0d27b46088235fb47;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hbf1f5ef0a019baf3e0a2bc9025a9c302f36ea9e7f417c2ffc49477c1;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hbb7eaf2717b036ef9908f50eba644a91e4e979161b01f1fcfc7e5233;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hd20d4268aa498acc8dc2ece954892da7dd55a3f398d77e6eb39fca50;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1ff9b06604e9140f6e578682df4fb3d511a3c1bbff3c142d0a3be1fda;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h274d491ccb3835f9cd0e0377345267f1e65a2b604a15c6c0a830eba;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'ha25e4fbb9cd406b08b0804333fe122400529d24fbc0f2f10d60ffc0f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1ec4bed67767cf8681ac9b49eb5ce24cb7a19cca643c3c8f35ff18110;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h4470dedbca42227225e9baae2bb1c594107c70d9af2dd02716144105;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h137464d3f1ab496386a7ec93ed1d50f1221c9f9b7894b71cdb42f79ce;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h14d5d3d787208672b19f7772f3c43740811e023b26510b437fca77fc;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h10952a812e1efd4e63e9bbd7d34500e38b0b7a19c08487c923ed120e5;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1da05fa2c907a0cbd1e55230b6b80138a3e664fbbe6a0f29995665052;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hc4f9913c30908f3522b882e5a4b3cd88faacea8495b0b8a123c178e2;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1e9530b510d05636920fc005139a8b6f2da609f8b5a53a049b47b26eb;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h153ef29caad4851d2fd0265e14759984994f91b710571a1d1f7c98b5c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h10022790e9a2c00c9e3130ffc5000c81d63c25b06e6663935cb8845bb;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h5a72ab277a486b2908ebe751a71f203a4e494f9ee61e9583278969c7;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1f0f409a1611aceecb62e6f3daa4bca10167122adf239b1d4f02cbd49;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h15469523086526e1c6f0cc38250da6eebee3e0e55e012e74acf58b97b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1f192ab9e9f2ad7e153c4cca5fe7f36e6667128edb4d99b034a458f62;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1e536adcadd1f869e767fe2028471f1b517730de9f6693ab940bff1bd;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1b890001127559aaaeae860befd1fce56336aecc7a5235bb202eb4e5c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h194577efe15072cb83de5a26c03d8403a4c4a458a0ac4c8d1ca610e15;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1953587af18cff80611bb5e57d6f40f3911eccd778c6253a4aa48c4a2;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h193ea8d26970089f7c4e98fce23ef8366e4b641bfd82a03264b249a9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h160a36df69ac5dac20e418c1cf94ea6489577f5c9135e9e693b075987;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hd3c9fb2fba3373fa5671a0968de8609d234b0f5439f9300d2906f9b8;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h196f76a7a37417adeadd7ff57bbab394624c06c3279bc92ce85a3434b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h16afb0b177697382874c1ee4697142bfe3e27a66a1039d8d5a8dce9c6;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1aeb98240ea657f6cd813e2d3aa5a622fcdb1be1a8151cc25a4797dec;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h5be17618e5cfe38fe5749347724e7147791a3f6b7a394a9ab18f5d6f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hc0c06a07b94afea30105e7b718a3d878342bf078d36062f24ee11988;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1428629eea70692151ab4ce59533eddc44f57d3a9856ad0fbe80536ee;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1062a6adcdbd30059f492e7d9ff64d18e7f12afd0e54f998c591b770e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h6cd966fde810f7e6f651b498896aa6c20464335984de576ae4ba15b0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h7a3dea7f515219d9ebce20cebbf88bab0ac776a5eec4f34ecaee35d6;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h109453511da93339874bfa8d660ba8c2e2b81bdc232b90ff8eded3db2;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h19ce89fd50ef65defbf196c8cace3669f766e49463449d94d4e4980ef;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1ef8f1b2c62567abf347a3b49da836769f777432ffe22e7fc2db8df89;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1885cfd7a4c1d837d214a3b0201dde283e0e6af70799a16bcc8f2d400;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h17995b71f7325859958f27308bc437c54f83a659e2b28af4d51135640;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'ha6d88c2ab08ff0731af2be788af7db4eb86a0884f7c1d7766a6f58e7;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hb753707e15df3757b9aca3f0f523f053027da321da47f46a865633cc;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h17e75a95421e4769db20f4e9a82380678f13e279f0be59e83c5f132cb;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1c0ada25a7a837eab32b46802419e877caf5d70fd92fd2a0f2f0f9089;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1e46e1832eebf26c8846523934bc51e11bae7466ba61eeb562e3a421d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hda8331ccdff252218cc0b8430c1464a097c4fe70becbf5423ac99fcc;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1cc5806cd552e63a82db68e3eac33ca3f8545f4efee73ae1e4d6b33c0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h15ed5d7aea298a0244f90ea5290835b5c35827046b478b28144021852;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hb659f4483b0f83beb76e321c6cb2aa2a95b7f01f720fe2a8fa739cc4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1389ad7f035fc76457ac93647b29e8da5696448d48d400d21c4b2a591;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1d30c907021edc97fb10fcaa6634b82d89b1cbbe9aa67c1a01ce6c0a1;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1b9bf3c9b99d6aa38f0954a2162f4955c76695efa2e5943cd26925f74;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hcec64253f953b66090e4b914ffadbf7eeec4a69f60636a1475b10bd;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'had80335a5632c9fc17955182a03be3c557e0d463d1fc6e3b5b6a8dee;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1e7f6a61143f3b2e39b94435fbf843bff51db038405010cad558980e8;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h10dabf6ad80b7c1c33c7e6eb19c50b55a04a009726f564d5a8e4950a7;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h7408502c02e6b205bb4575249e9c78acd6cbf4e99038ab6b5e229be6;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'ha5a9e56c829bc17d971c4b480aa6bfd5a0cae1a13137c0b22037ee77;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1561a40bf2610e082d02ca69ad53894881f7fb9bfb4b626260bfbd313;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h14dafa05ca897db184dc041fca4a6cbe893de5bc3b6fe53292d441d75;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1d710a7c7c99d3e5736758f84adecd13f7cbe8eecebdcba590d295794;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1b8318b04a8223fbadd934019962fceb468b6bc8d2b9159dfdeb9709f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hcbd383c0d07c5f1b621f946935f9fca7b2dc30c04c02bfa849561fd0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hb47553c069f265421815afb1eacef625d99edaf4524ad68bcc417ed0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h7fc7a7b18db1e87cfba673850b4e058e645ffd3f46f585bc96667949;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h10692e67f9e9e539e0eefcb81946b0c0378af1240fa8f966e4c4ae21a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1bf09d443e6bd332da6fc19db4611139cc1b2c6cf8465a3c7cbb08686;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1890ec4afdfc6ca94e6c3d14a782d329fb2efdef7bde4e235655d01e5;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h3d21e60afa47412a2e66ef65dc420116252af59bf66ba72cd8a27380;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hc4fbe65ae5240e30a1104af92b1ffbc8b8ff35b983b013553f35613f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h193c09695742217a5361b3536f1b7d7307ec04a3fbc3518b7336b0df5;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h135e59ed3ae88bc083f1f85c140d5a059cbc50a857300d596ed6e5356;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h19fc4397cf921dbcbf065927ae40bd5c678d6769d61d2b2f87d19febc;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1187be2ee2b30a045afacd0d75e40a7bc614c7d371f9460e08afbdc87;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1dcbf4e19db8dfa54c4fffc703752f3d9210be5adf2d56a3218d5e3c7;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h194f0ab07f2ab5ac9aa6286df376906cf1409c051fd48e5b1190ef755;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h10c039a15c5ad0b553f9fffbeb408bcf4f0828c6e532eb3c63baa93fb;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h10122afee2508007d20ef203fb416e6eb0d416a55db396f601d6c1ebd;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'habee6d3499c2b756989a5c9f6d2a7efb33a26e9e35f5adc8cff90e82;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1e17a3eb6413cdd2717057d576f785968cab0e8f57dcfd5fd4b920d69;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hf54056fbf0c6e936e313342c7ca3ea11012a7e7ef47cc9d5d91a4d69;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h146f6aea01fe131793bf2a77129d2039dda658c6d6af75fb0f6270e4c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h174043f9b55478405daf3a6ef853781408e9fff0bd8a3376ed23caf57;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hcae11b2a80f82d3c99a5f6ae7d0d2b7e985a41cfa50696f817f8e84;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1d421220f7da317e591f8b33f75411bf537b7ac0a6e3873df65401f4c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h4765155dd3b3d63768d7f437ae61e3c5994d5f6277b67e1baefb4ad0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h93b9de0d1b8008679884e1d7bafb76c6f73151fa9a8a639912546a0b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'ha4c696c13e223a5d3f4320e0f78fd4a1d9e1e356ca60e383d285ce4a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h10de40048709519408e23e39e9593a5edfb64a1d1f5189ab5845e6a53;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1e70a653745d0e81be53378136d6caea330cc4f0b036757edee355691;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h11c8f664725b9d2b7b55f5d56bd73dd9663a1361a18db2b55d4ff3abb;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h98701439588ae5201dbfb1e27eb614f6c6fb33ff0a7d9c740c4ad41a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h10cbd1cf85d7a87c3a8223c33993581d8d8372851a451daf46e25a824;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h3a736a283f2ab27408da43e727fd9a616e1fb280820ca2bcdcb76332;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h80468d81ccc195230958ae968ff0072c9f3940705876ad15e0953dc2;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h4ed66e7e33aa463f5a3a752b0d7f74a72ff78b38be0f592b631f94aa;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h127880875c00faf15e272445a225914c9364a533612191c2500585322;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h7dd9f50e1cb50bd42622ed63e2a485c52c478b308652bcec50190f04;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hd071ec0f2020a9ea9990b2300c2c8d0496dd8517d245a4a07266426a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1aaaa07527abe601eff7b525088cd4b2342726b88720f4ebd9f7b3cc2;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hf285a1bf120bc8d73a7d2f9102af2347d8bf47afbb19135ab69ec68e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h553b88d3ca1511706cc477269f2e6757ef158c5796f0fb0077aa8b08;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h194d6a89c39818aea1e08459761d1dbfbf761ac98083969c1c3b33253;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h11edbefc5509ff2dc76904f78dd9eae2e6d9dfc381f9924f17a256a2b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h115f54510581651e7777aa065a3ef39ebc90788e722c4a36be91e350f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1ace262e37a7adc3c50d533059032ebbabf13075db05d73d024322479;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h199db1fff817b1b18bd4570a6654377df9a38ccafc2a7a9328fec1f44;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h123ab3b3316c4d62e41fe40d20a7a2a8882c45b96eaa5933379181f6a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h3d04cf917749c85b9b555eae8f45fc380d24a21f6440fb74372a8e38;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h6cb30f6bf2dc632dda06e8ffd741752aba463b0e6f270eea751de187;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1d908d850ffaf4d5c5f432506d11402b9445dd977aacca46753067e51;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1cdde911ca29d97ae3eda0a4a49d6b01239199564eb9d89f8a4ea3e5a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h37df9f93a6d68eb416c4358fc8605cbff92ca11b55e3c3b29b9f1775;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h5e5aab0583e0846fab0962b85414db46dd381d4c8a8ff54d9c45fec8;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h14dc069e9c083e01db6c2baf7859a7a1ef8ab401402213e63525c2bf3;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1d7ed5ce811fcf31143174db0b7a467f8eea21e9abfd50378aceeda07;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h86844e85d372a6a31372ae7a52fe09c5e357c106b2fb37c5e97c6418;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1447832122813bec853fce85bfd5c5b329388fd421a48611aa505acc9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h24b9bca4c55b7f85c85ea3f3b368c97e36e72c1936542b3e38bf3399;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h172039608f7573a1bf81cae559fabcb178826483fea9d142bad79ae1f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1e0ce6b165c0b63317543009b0824200bf21070db2b8958066cf5e394;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h2cafb7d72935664d1f0568b050b70f50e37001324788d053f868f1a5;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1e86c6f30d3ba3d17d0a0c15b11b58d19de5c6fa50e32f914eecfd83e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h14274879d3e6b0a3c39e8d9a83e96269cf08f9c087d5063bc6f801a84;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h2d14230d7c574238dd989f102a77fb2f9907ad96367ec5652541629;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h9094de25f023cbdaf1a4e25ead2a6a9fabc91915e204938f4fba0ad2;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1b709dde68a6fe45cb722bc5221a86f0113f3bb353af4d494e94213f9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1c349d8a6a3fb4662e4957ee192b37053f36200ab81d36b543b81c0d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h443dec93e9e2ac562b0c59b4802395a7f2019a2adcf708e627e9c9bd;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h94a1db524bde1c4ef832145ad6a89f64109a7ee553564b00db819b00;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h9c9181167f496d574130f12b2cba27326cd6d604b8899e688b700e1b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'haa45d770ce220fadfe649e0bdebc85ad3079b23abd6aaeb3f113e3f4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1df1cc335581d3b9661652b15db872c9ce8b95f03bffeedff3e6cbff;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h19b2ac389ded1a20f42e81fe46bdb24d9dff877081cb36d99b3d327b9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h160e36d042e42d7a77cccdeb62b8eaed112d317bad11629a83073f33a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h13f381f76cdb7b230444ca056db77fc980fb4c27a8c9fbe66db66c4cc;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1fced3cad20160e331b1eb0fe027b4246cd203843a45c24481dea7a7a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h177c4f96f828e7530aed30eb09e456c7e4b42d0ff7b73d27f52842f29;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hb38ceff4ba5c0791144ef48b78bbf0ec85e300d8e377d4152c2a8984;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h17c69da743cf96b04961d364d951ccb3d49cb85715089463e530589d4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h164d857a864a68950ade56e90bddef415cce2adc7f1b3a1e0b1b5ae54;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1057dca57915199e5453e9f55fe004b7849fd625a197fde38184b8244;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'heacb600e836af13610093b486cee4a004c38eed6b079d275df1b8609;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hf9b2f8ea2fc30b6b6dcd51117d7f530a4a7ee13c15291f3346d8ee4e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1be728b1842b79bfedf5cf45c3670fd1d78e739fef6d67a60519905d4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1996ef0527796bdfda7c202baaec14bf0062b92a2103fdab7929bf2bc;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h10139a0192de4563f762898823b21cca29c348d31a5c5b118888fc5f8;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'he4fb08b6cf476b3071e30f014c15f30dec4f7f155cb396c366e131ab;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1606929a0e7c6c68e1548a61bbac8da3ead50dc10df0dc1331f7ff78e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'he8da2b9a819681a5bc7b3ec575158a50eb2c98de1aca5a5aa63c1f31;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1267039fce7c58bf3528e91d179752f04c952dbc5475d5704404be807;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1672b0c20066365bc5a754381afb0e70f4d228be084eecbcda4802964;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h19ae3024ed884f6545b4320df66a4bf952eab1be269521fbde0605e4c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h11a9764e5e906991bc9205eb918e163c588a87acf128ed91e46d9c3ff;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1a0cd4de02f3ef2757a3da06d55ca39b9bd33c3ab622f8014bd0ab8df;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h14da1ccce26a13c886fd823f3b8a246d260580a8b54bcb57b34bbd5b9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hb72554087db587bbc0b76041e4b4f8b57483c1818f5ca784e372c471;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h94cd9d44f290a8d4616644a9b1664c715ac3e4f48fd019af215b5846;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h81e7865e81d481374be16170118b70d86a8b67bd017eabe6668be0ae;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'ha45090e9bab6993b175bb0b60f3c2dbb2af5429047b4338a2e3d1655;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h590074abde2eee0ee5de3adf8bc1f5d9d19ccfe8d4676cbf3d3d2b86;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h19713529db2593f388b98aff304017257d3b395a613ecf7e057194ced;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h8f0f41d013b73410dc3665908e343433169f4be06c5806eab7d84cc9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h23753dbd8f570e295fe328c5c403ed3bb16ce6be7aef52150fbc6387;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h361511aedc8c957f8019909ac163f6a716f8faa475ce6ee50b35a318;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h4c7fa28a77757593969726d4bc3573c894e26f6aee46ebdacc0452ce;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hfca4c169235002d4d32e855816beea08f049251b75e0316ca7689749;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hb1fbc32433684c5580b090621ba8451e24bc9ace6afdb90e0ade93ad;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1dc87c8c76d2efbb0220236e2e13811a0a96cf354c00ca1c834313ea9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h111e5b6c00cf8b747be26a69157de6dbac25f6090fbec058d0dfeac76;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h3364b0f44e8494dd8b8492172ebf05dc7dd3fbf072b1e7cbc1a038b8;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hec6757b3a009c15cc7a026566477b62aff59e49904beba65fbff9095;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1d77066a537fa4049afd17eda150e80125c92b68ead29a95ef48ccf7c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h7ca054a75b54092e0f52c8be4dfc9a96999f5545a9a3e5ada9213066;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h7b57f1fe7f9bf5bcb5a8661668c6c81633b5390981890013cf14fe0d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h2847c786b1e27f10a850fe93d2bdfb8460bc56984819532be0189cbd;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h3b7d934ae282211927f6406af6ce9ee10dde26d14621f302a4757f36;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h134ca4e486e499367ab384b163ac53bea98938b640a3e4db3038b664d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h2895d5b390e04b59dd49e9649252d2389d08416960f0eb7deb740a9a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1227ee1f34dd8ca4007ddf74690e4af1cb86fd98312200dcf743d7f1a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h282f7e38eb1476dbcbd40f17f5b99991b02ebdc38c65986017b47f1f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h143628cb89aa09d24267eaba54621f61b2725861996bd182843559194;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'he4853a52467bd92d13f52889258e62f4cb22dfcefc8d523640c2bdf9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h17a87892f6907cf554ea20cd7bd595dbfbe63fe82cbf8e3280d2e7b2b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h18f209e33174e30e3675226a32d15ef777f1a26f917d1384d071545e5;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h264120959a9205ea02af69e4797688392e75b1da238907c6466e21bf;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h68c41b6a201eb8cae30a2fe67d791f2c8154bcb3326cd58a356ed814;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hc41d219ebc80660b56375b108b315cf0f1fca83498fa126454b3bc51;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1f66898adfaab1ded8f9194c51e6663f528695227da3d1d3d90a91baf;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h18aa26185e0389e55fbb6fde02b8a0ef5fc0bf5e4d1bbcc918c518ed2;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h140511bfc335be3c458bbac8209437a5968192d142d2a1f157ae5f291;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1adfec03589a0eca5cc9a789b4fa395478bf43c0586c9069c8466345e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h9d73c6fdccd81b66ac2875eaf305f7970ea2c60308d8e878c1a0174a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h7705f9c28cf2fae6e8b426bc49a7de8f2285156301aefa5700429a26;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h2332a9348b1e467c1e48a4547334bb0682b4b4cfaf465e05a0b92205;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hfb5dd56e38a8b29aacec06e128116cb4dde14702d9d1f06d7a740630;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'heecda24fe4eb61bee5329e42664317dd95d58930c43ad9a285ecf04f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h183a13b63b9f87937b0a82f6cdd4ea7385c5a7c2eeaaf856d4c4ee686;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h26d137938250edff554f9073fd7fae3bbfca001fbc39a2777ddbe0a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'ha2b8f516270f5e9b29e41bad471f11ec4d31f2f03d833350093f4e26;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h16f8b7e8b56a620fa675e4b347e40a61e1748819016997fd8c2e4dbaa;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hf4a22512ef6652513e7e5cbca6b422317ea152832715772210eb5fc;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h68721af9c4e7e904424d1b9d33b5cb24eb0e4432cfb43b82694bd34;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1cbadaaefe6fca03d604cd9be1d1ba090da0d884321fc21b416bb5262;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1e126cfc2d97bec950ad17a74daf8c45a6341aaf6d2bca1219d5a3d5c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h141da3865d94c72267eeeb3c506650b22adce1b9d06920598af09fba4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h64a86e9d6e5de1be596b77b83a4bc549101cb8999f26f20744b411c1;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h10b2cac92e193ec0b9c85aee8295c8028e0f213d06a664456db869846;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h59891a3b457489d636824633aa32ed33b19631e84b13c1226b1dedf0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h19f10a9b2b2c3e94e9b98aad4478ae3050afd67264d1071cdc411bff2;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h30ec6cb8a43c73a9376ba17fb5cf829c25a5452e0f205ed7269a2bf9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h18f6f5106cb603d3cdf5bfd69308606081cb9f2ccc1abf13d62b3510;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h19c6cb4978ba019d10dfa341db04573676ad48b2ef8abd75955257b3d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1fb1663e752da916da5a2f665f69d846977dbeef82ed14441186ff00d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h832cbab837d196c8d72fa358e996bc15c47def1cb44d74fbdbab52c2;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1e61fb494898d96231581524b05117b735200994486f15b4cfc5e87b6;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hcc5a191d0a61df21f873bf3882794d85a3e19b2b91fe61fc20652811;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h10fbefcb73b3c5401a3d547ff3f521f9cd6faf7670f853cb468413600;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h12754ed6d65c660018ba2e5259a3a26189812ceaf767dd197ddf5c06a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h158e1d7fd92da9df35c8a680c730c74b37f8eaf5592ae5f515553eef6;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h4a324ca8172e143f1b3e9ae89d3dbcce11bf0ddc200f2f85cea1ddd1;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1e5185743d83c690f7f66c1150a0ee18c4c18e83b49f3ab573c0dfcca;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hfae5e32f956412dc39314c8f3a68e39fee6afbe1b4c31dfce69b0c86;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h18b457cb8dc6b228f01a4f0a7b1b5bb7eaa0426485487f574ae510759;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1972ea28d498d59de7850f134985959f5f3cee1c4f3e8f8961db8991b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1bf33d466af7466747df3956c1dec02b7cfef3f89ff7cd1cc433d5b8e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h19813bc005e01e8c704fb89be95a97887e23658026d6476eb31641ac7;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h93a9d6f60e3e8f4de8d3fcdfe3a567f6d6365c34b9a33577bb264395;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1f1f5b4fd43f96ffc02db0316ca5cb3c6451395fc3ce2e6512e8eeb7e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1b12795c1cd5e2c954bec4e777d91b9a9a234506491ba2d5b85b25dee;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h41f202a63c8bdd387384aed319773393a8c8d2b37dc63f24fca2e40;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h6a38575ce12e61894d3155ca5c968ea3b9b9cea39f6bec29a1ddee64;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h46b2cfe9740ced3b936b020622968b92a29dd918ff9cc91fd8f4df72;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'he6307023d67731dce17c2b3da1474336ce9d57f684d0302bbf525c11;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h14d30d62aa585992943b8b8e2da21e5a9bc084ccff719e723a591a828;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h10ffbd65206a6974d7a99a7a5e133dcf5c2ea1dd9eebb4f9fd531401f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h11e08fb7b7217db76b0e3d1d0b878c47f52b5361db1ef74c9660df048;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1f6d0481a349ef85bdbfce837832c2c656f4f39d4f2d7b392f76245b7;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hbb0f5741317e68f436aabb9e502f3d5a275113b41876298077afcf32;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1cb1501d1c034bebcd1d2728dc223c1250a8f67d2043ca733ff4a5453;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1256a85e442d8148eb42d18b2ae1c2f1ef806eb185f7dde5ec1e22087;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h3e363d8da08dbf67054243734d980488edae16425ca8f4b21f8556c5;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1dbfd6458ac51954b191e3fd141e2d7427f65c389f088a0896ce39309;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h169f2ab46cd75a8b0cfd22349c98fd8c84f8345dad67d72d36025946b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1090e0454c7c4258c16919d13c853bee10b2c6fe2a64b31f731e9badb;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h12eb639396c924420aa82dc6f416b488810adf8ad6a0fb5dd5f2b880;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h19d370dcae5e6a2ba1a679194756adc372a5477e68c3b75e6fac26557;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h10af0f236be580fe261a8a705515347c50904976f8ec0c7439308fc11;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1bbd33108461a43d7388bb1199a215da42ce4706f1cb208494d85586b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h17898fc04d67130bace77babac82e009c77d2e2633447059e6f0597b2;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1b2294b30be928d358a1fc9c9210ce2c070babbab093c89508b0a3f50;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hcd8775905f81b257b7f5ac4e436015a97c46494b50cd5ade26bb9df;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hc890d6ff65cac4c9e0ee1778f399f6514ab3c4a8934e3269e20ee922;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'he27259b3e412ecf41926737712828708407101da02ec77daf9cb5482;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h5e4ca84a0389050db766bf9d2ba838bf11a394100adb574c8d6baf1b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h9efd402dc7ac36d53939988653a83304c4ed88fa4e952a2f91db01b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h151d42117094c8ff6d1658ea085e6cb03ca1b08da22d1e1ee48ed3e9e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h14629470656ef4febccff573afc660ce64bfb756c789ab439716146ca;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h14a6e5a630300046a319bddc7915608c3b9afe97f9baaf11a92a46099;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h19c7dc1baf5c51ddc3bcbb090ec22d96a51a5bd223022d14d595e1e0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h176a401e0f5d20505764156052fc6e950abd74625df0703f1dc239c51;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1a0eac255741836088a4524da02e4c7c59cfd86ef465c55222e574ccb;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1ac09f2578d3b9df90a3eeef32c8510488e57104767599983dc37b4a1;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hb8353cedccb5e1a25ee60534489a75cc6582e64dca46f689c15a7c61;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h107b6acff034a6ca4931e07dc5c4db5aef0aabcaf1a40ca6a98141bba;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hd1e9fcc2ebd761715a13b6cb6b079eefe005650897c6a13d41cdcc21;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h59395d25fffe527a8ee25147c914d0f6be9093c15a0cf5470fdd998f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1f448e307ce0d34db7366993b0a3594c8b5c3c281128f5acc076f8222;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'ha22012d26b88cffe6443de58caad7805bca1b6f2abd0b60387e49372;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1f8f721cd28d0ba26bad115817984a2e81ac568da2614c1ef870fb8c6;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h5f8f603d2a25ad07d8609554010246ded85e466c75e6b0e9d97a8845;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1efabe5c4916ed5198357a23a05ab69ae9bedabd1964e53c1f3a3644b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hd45552263db06f58317b4f11dea484ab0df84099ac36915f5d3297c3;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1334c47ab9b0d73b4e39ec3c80b08ca9d7b6d0911885d31e9ae4975dc;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1c3d45c6ddeba873f61dfc39bcfd3ceb745150af0e8f589e26279f7ba;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hbc1ce6b60e4745999b919917aa47d076a33bd3059366349e2081b0f2;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h14d1e8202d92202bdf078bc3eef8d38522b8d73a0f4612dd0bd0f978b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h155eb383c54082b7b05f751d3db89aa8284402c4e3a439c5b0d2fddc9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h219e35c8d4efdefbf5874b4168877fcbbe77765284a16d1cba9c9c13;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1c86b70e000f086e1729664915a0d512e95a302cd63b1ba1a5f92d4e1;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h16a573f185a3465b54a654abbe60e64603f7307fbea882a02fa6e3d84;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1824e905c7f5e44235e0fc689da608aa8dc2458d191aae41cea404de;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h7124d09ee054cdc71dd5283c91a54718bea1889f5eab45b7f74601e1;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h5545bd0fd9a82e0ab33df14844c3329814ab9eab2af0c1acba973516;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h110c894ad530293fed38b17b8ffc8163f9d5e99869d5b420acfccb432;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1c906750fd9e5d6ad1e988a6192951d4fa4c25c9697276134fc16dea0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h19cf93c8ed871477bca66037a1273e8fa06576c571a7e71742a49a7aa;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hc4db899ad8c0afe57ec704b5415ae8c38d10864b20a9467280fe4ac8;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h15d0e15dc0585b9bd1c00ebe8f8029f765db1ac2994134875c5a8ae41;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1bb12403c4b02881acd5217786c0bfa4d7c79c6fea62a749be33aaa40;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1a87a90e04e7bef275ca26c78d646a383e8c5c523cdb2682dd22c497;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h95eed4a9f73dac0163567075db0d6dbb46815a5831a8f49ffe13745b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hbe9a653ecc13e9261092d016b4d2b949dfd71a6ae4297dc80fef3b8b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hcb2b46716935e687877ff50d44741baffb82e61498a757ad2fb4ddaf;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1e1361e9222317819608e359a8b3d9d0067a3acda8a1da9537a00db22;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h15e1d30a93aa764abf6cc90320d139fe488c51325ecaac2fd88627b2b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'ha4ff97142fb615c2a449aca9fdf3ed4300bb3f561b868ba3d5e35c60;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hf80641c2aeec4da0e1630bf0e121acf5d4355d48b95b0edca8a73f7b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h612f61e960e3bddd39103065b280d7992ae64a44ad8f88329afea75d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h5e0847dea35391cdba6f0cd05832cdf665f3e357d76584eb376a0cba;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1daabcc72ef7ccff73fbb7fd7c67e22d0cb39f4e4830dc1ec71501f0f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1a243a244276136b5ac4de0bdd88f1c15edebbc949eac7e76742cdc6a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h10770a9d9e604e6fd341088f292e566ddc44297aa4ab1bcd681c00ae0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h64c94dd16c2844f48f10155102e41a2bc3f9fa71ddcafc05347b15a4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h136217fad19261594792d0c8f855e83e23a10a99295ce0a89a4f33c52;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h36cdc70cbae1605c410c207ccb4df5a2ed53b06e8088288e19dfdbfc;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hce7bd2751257921834ec824cd4008f29b6e31deaa44d15c74e55c611;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h4a72ffba066203b09bbfb8295664b06ce40d420fc0a18da0c7950bca;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h33a2dfcbcc635a0ff45201262eab76ea3d2814a1769fe7a61a486796;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1b8e219a9959403d732350693dc6fe3d5b0e610ae6c7213b6f39c0f2e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1b8f07e5f76f30715d79c1c67dbc2cb8ee880d14a608c760596ff3031;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h6b1c04348f4e6c2068ca761041c1a2781366578e57b788135a11df73;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h110cf8a182755a4f891e378087fbd8f5211f88b7cc338ae7cf89e1d09;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1e89bc09076df7c3fd692efa0b93887c71bfef00c37c921fee8ce49f7;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1ff5d6d41249f1e821e397799508a68829cb79388b4d7cb86bb7893f9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1606b6169f306189f485af85ab265906e3a535b23f6fe1e6cd45db894;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h174b2e50c176bee907fc345a329865d2e6e417031bee843f32abe0bb5;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1ef5698c4b76d3b19d248519efdf9c7d9bfed3ac20b57c8d97a34143;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h9f30a4fa5df19a149ee6cf014230fe86ed9b87e7436266b0a6d23b53;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h6baf0ed1eeb5bc55dc56c84c2f0dcb9ef7c91106178ff9c172d841e2;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h9bb353004808ee48537eabc2e745f34c3d80b73dbbd0053f7dca5868;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hf4b7bf8d6394fc402c78fc3ef87a7ac39c5a8684025276592ca8aed9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h159bdee45ed29834d83896b87c83af8950440061d4181b23b56d71699;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hba93bd3dee542ff7d6a5be6a13cfe20cd1ed90a68d24038022708e12;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h17267e0672fb3932faf91e43a0fc6d01faccd18fee3b022705521f606;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h10ff2a5bea95cbe1b8f1bf48635bccdda6549b6cf0d297af18e77904d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h52beda2138bc945aad142d86f6f33cd8b2739c433e18b7b78a2c129b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h91297096212ba7a33e71e22c3d6a9dd676fea72d74886b77572af624;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h4095121dddeff42e7a90119cacabe85f2d220a5114e235174a3df144;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1cafb930951065f9ce193f6fc8e3e8529a0b9026610d50dd48396a58;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'ha2a6c8c38a2ecccf01bc7f027c7ef5dd79f23da6ef48afd07c638b25;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1c759190165a8158192e8c132fb30af1a47ce88dc4a5e77af6b24f1c4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h7c2cac349182605bb5900fa0fea9abc71e4dbe7ee2448049d132794c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h5321b935e0af8b0a828f72857e7596d869718c278efaed74ee35bc34;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hc2f55ee61789ae9d827f7a084fea96af9aa99e02fe5e84616ae29530;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h678cb87ae0a8ff899748ccf1d5a260702fc478e0f7a8a8a75aa13a45;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h686ffe6aec298a9ab651412acaa4ef6c4175630fdb3d20cf0f2f4791;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1c3e4995101db7b87ae57af6df63fe7ff7688e1f57e9398a7e668fc0d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h7893f9387793bf969009b9c1930e2d98ccc3801ec92a0d158ddb8ce1;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h16b88a19731346685c506e9b8db401040466cd9e14c0abd83464979bc;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h184aafe16c5eca975668049225cddaf8d1b8b8e92ccf2eb47630a41df;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'he73a6beb14bf086f8245f78a0d312f5d9d23ef569067295f71726370;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h180b8b9a072f9f0dd287f7b74b80a8eaf2acfe781e2b603d4064df1eb;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hefd88a1e69b434ed967a713a074b00af68656f82c451fa91a0d6df40;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h19d7d88d0db03bc4eb7208df4c7ca1b18c61d36c0c33cb7b32ddbc558;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h10c50f0335c32ca648510eeab4ab2161c77f6287144f6e0bc655d6e42;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h9b2b26af280750b631cadbcfe79b03559081c40c277a7f001f5c9e3a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h95496fbf6c270200a5b15942f2bae1cee7a7983afdafdf6634f974d9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1cd46754028de52dd90bafe6af2e00abd69c85ad9647ab96e91ac8a85;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h56fb566a67e7a5f55362425f32debea4547998cf6c2829e4e2b01c5b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h36a737508eb27d9abccfd9268504624736fe6a19be3dfff3c1d2849b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h148e73c47250645431d8e4e734ba5c0e7434914fef77f7a4b89cb37c9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1daa0c7bd192588ed7c0dc86811ba6bf645bd2e3b5936a383a2f24324;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h100d1b52e26b0e50a05400347779cacb0f63e3fbb476b6f24e16625df;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hafb7be5c380f5eee6bf8f2a13d362eae4cd522ef439d6399ea892497;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h7cc68c2a2eaf4f1aa9e4466aa9870acdb5947965dc3396167ab1316f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h12cc7717a30e79179b3b4f339059c3c5cf2060975bec3a697d138cee6;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1a8fd81f619d96f0138cd93b7745c31fde25ed02ec8018eb2154b73ce;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h823031e7e5191a750e1f49eacdc2abe22d105892478ad7032681c60b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1f8bbea26f4fba0f407749ac2326a93a45797098779d22a58c00895da;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1670854a92e047aaf4bd826f2a2dc1568b9ed3abb51ca06ebcd3722bc;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h301c50aa16fbbbceb9198d036710dec948e41fcef0f66c27e9e1f58e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1a0539f247615070f5fa351dd0fe6d21e89fcc2e34c70b522e6d9f891;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h182b2ca69fc748d0524d1e3d02d7e1577866edbf8613ef1c619ba06d0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hede14917a6851e6dc65c465cabf44ab667c4635881680dc65cd0f1fe;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1508b4c0f9322365205f34f00704c9bc717ccfbc48119f427133ce955;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1841dddc232cea3d74ffdbc753878af5dd721153a124cb863b17b4508;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h45dfe8639270abb44431fb1846bf92fcf5f97446913264dc0e8dbcd0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'haa4ea783c1601188e827e2d4d06eb7e8f81c2338eddaa977d35959bf;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h11f6a33919d0bb1c585cabd9b6d1790b49606e963a7e9069ebb7bc1d3;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h625c6e9186fbcd8e8aa060118029f6aefbdfb489be2a13b0a9197d83;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h184492677dcffe977a0ae8af40e1a6c0ee9323451a7df5a1ef1128ce9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1ef9d94014dfce8b725dbecc25595aa9e3ea7663547fc567a57c22692;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h190f6801dcaaa3b052f9b6cc025258afed37b8f0942f8aed7d7dd7bd4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h15b3665be6d6c3437d839b5b3291f72190aac956796f0f7485888d5a9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'heec68b25a522e22220f3543810ea4951f80be7c754024b4572e351b8;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1c4218a2c5e558e37006a52f4d9b13234e22a8c0e721cc701962ebd1d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h196873ac217bb96da3033c0288367386fbc55a7dc6a99bb88d952f244;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hc34af1f0a55e65e88b4bad222307579ceaea48acb324b97f674c468d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hecc8dfa2bab874b2dd1a8e0f27eda0a67e285e7b285d8e6ff1d61158;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h2e9c592ea2d743c4f1023218165efaaf1b7802e4ff3a59fd3d68f7b1;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hcdde54dfaa7ab6bd4b7051a56bc32ace32c5c8b7af491b43086ba04a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1518d90dc6201f92521603c840d842c1906691d5f15df327e97a565c5;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h8e7cac24a9d4f18e9a2051812b671695a5fb94acf7d7ace85de24cde;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h5876db0acabf9767225b1171377908b34d237c5b772d72033e7ef181;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h7e4836c4df2b34dbca3cacdca4faf403d217ec2c726baa7ed385f7d7;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h93340bfe142e3bed8083e7a744333fd23b755619de59b304d5bdd3e0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h6aec1ae605eb8bfc97aa0b3f1dc9883b20f2d268e7506ba16cda5b06;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h7ad9063ef299d5484d3ee8bdabe8f653f19c0094e830bf59e5b9cb27;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1fa9a3a7b09c07e77289d3ff3ecd7e59f9d9ca12f103d7440dab2e666;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h16eb4d23f4ebde721e59a1de6ac48e0ea69282d1ad559032469155443;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1337419d3344e51859debdfe9c8bdd02ef9d33cf818e95019e8b5182b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1005957cfe19823d7758030c9960b34552e3e4849b39bec2be406acb3;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1de0328761b2192f5774c49602107a7b6a4a5e8bce63da7802392ebce;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1d280e94641acfe98fa22edec1c2e9e52505f41608edaa1d0a0ab05b6;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h17862f065b5c2d343b67cd3e952246f54bcd012b46d3fea5e5db8807e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'heec39cf8ec81af6d66780230d1861df0ec82f6d2897e863090fb7500;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1c283316b4520f8e742d01c63ae49d426a595490abd158f24b32aaba7;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1fe40c1bbf590a98f4e7b88e7503333ab57e0c82353f2933365d094cb;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h20762de3f6ad6479a35c33a48dd9fd391a00e3464f4fa10580271591;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h14e3cb2cb298e6e89a2234bf76587d2f2ad1ad2387e5760ce7d2b028b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hb34d3b7bf75364da47a1a9429420ce5f9881aee4e670d5dd7962b35e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hc726c6c53504cfae1a7c042bf03a2ca0c11be4cc054d087b5a50fc6d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h901a10c9928fb56bc65320aee4c7cc9fc564bbda8cbc320267f92aa4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h118edda575d7d10afe52b14a4b7b151c88066a1e9c57a061eab86428a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h15855ffe975626cd53f7c035d61a483709c15ed6eab94f00ba16e636b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1f20e7d95409ea3674246c27649cb5177ee2774e27b307e1129474a0c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'he1c61566673544942f654695a2c3f5d20a0b5da47dcad6a158794fb7;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h16d9019fa437d4fc6c427c1d6dbd44daa6a0ed924579cc0c133245f4a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h90032ffbf49ff860896fee8b7bb2bfeeee5aa06bd9dbc62f4e5cd3d0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h196bb3ca1a7b7abe015d5bfe50fa27aca2e7bd593f77993300cf47c6f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h121edc356c2e72735f0e0c380d22affa06a4b59520f32ddb428268dc8;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h14a4b3a502dc5a526993b592f00de8d510f97651b1410953920784b66;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1df28c9ac17fc4196d69cab1af30f9ef94278e06e95abf085590d66fb;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h9efc44daedf86981b553f303ae72d9f933e558da120816be8ce6c009;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hf3b4dba2a114a9dba30808d2af76960a971764c118802734122a1a42;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h117f28038d2f839be4a26509b8a54d0c0df304885a9aec3b9fe0c8523;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h8d9f7c2177d7d3035468fc2da93974ce19e8a2e04687e67ac78c6cac;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1b931eaa861a5d5b436f50891b0cf1981de3e400aab6b00e0a2a8df71;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1af033a9a44600f15c854cb4733192e86742e210c640869497b3a4ffc;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h38d54e1415c7d718398c918727afaf288841e1aa2d054891dfef1475;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'ha09856e9ee1793c04dc4c20e36a536b916eb3b43cadb5dd97512a099;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1dffafc44d823d1da29dec2813bdab0bd141106448b7d43fade12a1f3;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h12e12e710f2c0469bfcb2bfdb1f3fce9e55ba99e16416f0a465da544a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1d84487234c5e0ce409171f0fa6216b89ed8f7f147edcd4229fa93239;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hdecc352bfd9b14e9f0145995876724eb63295799a88ba801f3c335e2;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1148e9878a9c62e524f871e7816f8f4f761ddeb4d453a86ae3c8f1407;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hc74d7ce2b246e5b0aeff32d8372a8c3a04372cee5f9f6d5163448a7c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1cef1798e7e021dc2170c9265a2286f671ee05a62d23be8d066f7fe56;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h13ffde708bc0fc47bb6460d397c4074db2a53715b118303083e5c3fc8;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h207a0d7f446ffbc9e465f503b1292d186e67dc992202f3c8af69358c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1d813f506f58854771cce3051877b585a0013fdd44d6438fb113570f5;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h189ff0acb55bdbaa0871fb046b172d28458eff5c3efdbdc82de31279;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h105c4147d831c9b95ee4f3b6d935a123a200792d40861bb95c931c40c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1ab65beac4a55690cf1bcaad412d8934ede919cb8407b52fa31b1818d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h8fad18ca9deb94931e984e8d02246d7418e3f86e80289693eac3a36a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h137e255dd4d88f747a5e0042b6eb74080879d7d6dad7dab037f688f9b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1d50c59bd802462ce8fa60d26ce0e9f456cb895002ee35cf646549ece;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h103c750cc087868f4e3e6669dd4ead5163603f6bda2b6f630f1e39a52;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1969e59d5d4e826a51b51ad5a71e82c5ff95c47937e217800966fda3a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h170464d5f4d937f036098e5ad21750eae457a5d5478f41eea8a921869;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hff73a04882d583b6d9353fef041642dfeb95974bc854c382268c291f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h8ae10648d2db45509f7ec907c8e8db26346c42a5361ceedd29cb4c23;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hbca18d37b6dbd27d601dbc5d1546ee9e6fb79d6040a9556e2c2c0adc;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h882147670bc7ba1e26ccbad89a0765ff75ed7b2acff09c76faae5679;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h12957096299f0183a624f92f8a80db157f0ca0d7cc787ebe3af991f79;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1a6491a6538f7c781d5e1da2f728c2bddce6e9e9f41160d51ce37d496;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h195a66661a6052841bede94432b1ee354342b0a931f8733fac8a5b336;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h303f3fe3c954b961fb1285132f86b71a9a15d9a04286318ce83574c2;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h106d561fa54ac29fc06f562dc77901c02e7c6222a94dee0e67660db4d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1976158861293f686bf11df7748658ce24df5a52730cf88f8e11c8fb2;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h173bc34653e2b14fd2cca45ffe2aecce147d6f1a2e09d4ed7ecbb64c5;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h12c801b19873642a447167384fe3f9cd5b5dbdeebdae375920cf8dca5;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h19a6e931ecb8f4d76b109bd859f248c09347a7cdd58a93e8a4eacf0d2;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1fe968ad97949bcf0e57c0d04cd0253ff06bacc8826471796ff8f7124;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1638360f21df9500f7f89fbe4a2238b17cb5301a4969aa062cef388e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1bbb7f5c56b051e392deaea5ba74b1cbd0211a8922c3deca5c380aef2;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1ee8a5562ce4fdb9315b852256713dff3f1994329f5551dfe294d0a96;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h9cf2f72a5c7a7554407e694a094bd965fbb92fc44280cd8a78e8150c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h30bc9587e143e25f0db6bb69fd7179669319ac3d698c66d1737f7fde;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hbffea8f2a6e1ecb4abed4dde41ae3582f8b0ebe03eb9d188ce6c7414;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hb8db16d9983e1961e6239463234e271cdf3afd082f32c93148f53bb;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1b72d86ea66545868ba1cb72a3747c66c546a3abb4d0d5bcdb82f0ba1;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1d555540c1f33b4c4d9eef7fc8b974f7965b2b4888d183d8791a3539e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h9a56b22718b46e2a62d6bf31ca665b80d83bdbada605d98295aad7e9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1ef9ae1f99130b1dd22604d050bd2e86f33a91dcbc08fd0a9e6928e7a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h15b392156d900c33fa92543af5ab8adf760f603a8f81f19b55b4f5da8;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'heca9f9359564cb3e07a8ea8ffd310795922bdcd54ca62e6bbe7de162;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h11f4b6e0bc278909daa752792d649def4b50234f159b2ad108d97c124;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h366c8ce386485a5841e1070b4a3f230f93701e6d592a05edf4a74d00;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hb4f65b6ebd430d9f4ab027a50adba61ab6c3b2e45828dfcee700217f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hf65910cbd26850ecd598104de901252896071344d3b3bee7cf8ffabc;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1f1267ef0b8ff1ccd020bf27f5b13f85cf94d38465a552169a610002d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h12eae87f071c593941bff07b5c532878594111aa5f7cbc018fa7ae02c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h58b56d3717329fc872fd72aff0314cf022ab5ff327029c1120e6f201;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1b7f5798af322035bf5d6e8a1776a0f6ba378a2da96f4edc705c18e20;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1998011a69559fb65f7dad37366c38dd10a03cd4efc143d73277cfcbe;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h6267dbfd6372f01de0af909a456135b71d6090ffe1793729667b202c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h360dd520d1302127c04120bfe5db6d92a8eec15c92a6b96e4c796092;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h9e76de4efd35251ed58b5c270ece903e98fa1798a34fd121b79c9862;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1a513dbdbfe136e0b431fa23ef0a70cc9047004258e93e8cf1c368731;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hc020333eded52665bf8a6188cd0862b5bf3ca4ccb93d5a3012f3cc2d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h10fb9af41d7185b64789d4fecb8727593a8b684f0eba90daaf43e789a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1c5eca16478d416f68ed9c45d3e97bac672baaa6b143fefafd7d0266d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hce70fa0e7f7fd3c9bf4d5b41849e79f2923f1f0d942f3d0dce8403ac;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h4ea056f85b3c9c850a60677c22f01dd2a040c73fde18ecfe5cc8b46b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h8d6dee9c0c80fdf04c8dff4ea267c5955365e6afd86d8db01464ce0a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hc900e657697c29f58ed01cd2d0c9c0f9d89360ef8b681b8d167c4804;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1f68cb71c933a9a88356d2e531e0810c08c9d5105eb23215c7593cc77;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h2beb18e38eb59c6587393dd26855231408ca4470cf2a3aa7979fd14d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h29a9da130c9f620c8345193ad01d4fcebe85385d54bc74d1bb02b328;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hbb6f100ea5d33abfe47884f98c7239ae8017096957f30460fcdf5295;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h18db31886c34169bc50963491c2b6903cb753ad798dd2a9daa4374b6e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h3280dd732e67896bd14ad8678a27e9c112e70c2aa5e13a9dc15a44e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h114e03ce1edc6ad0ad975180ebf928287537a0399ce508a57472cd54d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h14f50b3881fd2b513c421cafd1f32e0299480f63ce95b92b2cdd5dc8f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h11b322ad12dcaf0ac2e1c14cdeca6eb682452954411e3f225beda3025;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h5507b7ac01df81921c67540023c5d9bc7eed9712cfa7e468088b759d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h10c84f3e8a487ab3361fc08813a76834826aabe25fb3dda2d7761ff30;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h125ac558898316bfe4404018506934239c791599f2f4645e1ce0d9b3c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1780e01d2b928091bd244933923e90f1c69a88fc3789892014a525ce9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h29864648c6f693c2f6d28aafc6fead28fabde36f4f83438502589d4e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1f630cc0d053b4f0775742a42d311564cd543703fe052e2393dde70cd;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hff84817717912e5c727b8cf4d26e1a3ac8b6429088191fded2baebc0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1539c0a576203dce00d3b3c7eb1a7a9352ae3335f360e0fb6e90c0f5c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1e7dd0d79662c9acbc75ddd3d76abb1047952a2bde588bed0e8a8bca3;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1baa393011d5d358489c0462b76c7567f34ba9732d3aef11370816bf7;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1f78466571eaccf6596ce1f54c44ef40c61070226e430f93fb020c001;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h10fb4bc0843a8978e0b9c86bf5df20982dbb6c61138f6c5c94f572946;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h18c3030f6f22bef9a308df4591ebb6e0c1d12bc20eea90641eb844f40;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1621d50bf03cfce0337e322defa544c44fdffefe0450d534249a86cb3;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h5009df5db00c104556ca2204c08711ad7033a6dac8e83c49d3516834;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'he4f1826ebb4d13112f22603df1dd3582c69d526017fc40688f827ddf;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h530f58d18d26e1d35f1d2499bb2acdc2f49b804f8b12d2f213c009e3;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hb716b8f456b954ee46f2053d5f41d25324b77284aa554666d4125ee1;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h182a1e15d87e6def139ac6a1bea0eba2b45c32209e9dd533fc9b526a0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'he746966241f6787834e3aa78167d402e7ac9df334c8aaaee9d230961;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1458dac85bcceb55688eb8cf44e1b10cf55831d3af9866630431349c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1486e4897b78732bb4aa7c20ef6cb0c2991748f96698677089bf12de9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'ha7562bcf56a606c3efa85a36164283581a12a4c80b40d45301e1b7e5;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h18f3654fce4ef4af3b1ac0cb444ddc191c06580ce962ec124d9e37dc9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1089874915e99f199c7b0bdb63dc111f7cc10b860cf165024a0261271;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1a45f920e96c4314aef8d9c2f2d94da44b1e3809ed2372c519c86ea67;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hb91ce7f6e3fbf6faf76124d865089aa73314aef85e210be115b39230;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1e30c4736fba3a3ef5cddb8e31f1930042909e7c259047cdeb9b6ebe5;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1f594e87e8edb50774acd04c2d284131c94b3d89ad600f7ed4a0eecee;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h60843ca3a6ab05ba99f58d7b78a3a5cda28e05501e046633374bdf12;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h10b39e42f7b0e5684814a3c8d5a18e62dae70c4b8dbf95b87b58bb124;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h3fa8224586ef443f3d89338719834e90c67398306d388091278b2818;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h175e0f7a03865b5423166fb9c69283a0c03375d1553fec7ba36ad96ba;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1ef9510b82de520e4f9a7bee30926b700624b2574569b703d625a2345;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h9e8e386b4bb10a422e5ef0f4a3146165d0302a7d75d86de1e4a816fd;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h104947accdc0b40b9a0e1a7b8510297864ab74af7733436f839583621;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hed2e446a3530933487b2f05649ccbdbf9d46ad3fa72b6c3b1343c8c8;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1388416baf1ac76329803b3abbfd11cb99fa9bab9ff277a9e11b2bc7;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h119aa87d3b443ddda05a778145e97cc4209268f1ff2ac014f354be694;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hcb9a9dcad7ef735454ca10c71580a7c3e684d9d2b0b74682ff7e983;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h135492e84be555036d0c5440099dbc17c669f6e4eb14d06a6bb45cd16;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h24257d0f32a6906187599a8cd4492f06836232f372f93415bd1ba4a7;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1d6013ee66d9a4f9dc49b73d9adcba8a21e7b86912b88d1faccc6f461;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h4585592a00765391a07097a6f4389952b69588dde4672f28d96921ae;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1bc6b65fcf74338b64a8ce05c64b55cb1d0ef1490fe9c344140572d44;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1600f2f5f00118012dd61b11f3ed300d28a696374c17b2e1ddbd7f784;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h82c3f3b1d99b150062a1d1cebab8da8766d9068b88281b67d7c02995;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hd9e1cc4c4a66850f2b63394633578077e0733d9526383092b5f43bab;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h16794b885ec4cbe52fe60684aaae2a69ea986061ea2daa5030155de15;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h11b2812876b23ef68e6dcee179b0f2af2e769303b36650ab7648f30b2;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1866d4fa18d4cdb3d7c9d989a8eff2e3cda63b292f709f47595758971;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h7b54a1572ab12253667f5190306ddbdd67cb7bab5d777ce296de3295;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h80cd9665c2b8e001bdf04f84be3d0ed8b3b6cad8161fa58e99388790;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h10d6bb1aacb7916f0d4169d1324075977a21bb4739b71bac9f5b5e25a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h15bfb09030b8e7c2463e0d5bc6e0d2f0cdb56ef5a16f660e9ee4e7d8f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h5561ab4a5725ea74c74a70fca035e44bba7e738d88df4672e7bf2d81;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hfd5a34eabdfa438e27aae3146f0baeecee67ea883952d16fffa8ce66;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h25a06e7b6dbd6271c0ea7166522cb4199e6cc9cbea2af1b7e5b8dc4e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h44e2e38a8b89e54b5c399bd60d0aee8bbd95dde3beab9a6d04592594;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'ha758ed2c3d967312a8f5326879ebe81dbdb12912fbf930bd2adb10b9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hb989e8049cf70dfe3d02ef65966b4db6c48a5061cd2d3b26e911d700;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1ce403aa7966f87a1784bdc10cce40bc75433ffa67eabd3c170e4f8ba;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1a142210f1294d1cb6778f45fb88e3f90dcdb622a45ba1c88b4b51455;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1d737e44e16da3da396c6a7358793c9c2017855936288f379e18bc444;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hb614bba6abb17f9992c617d7ac6ea158413b5ff72b14c30328f2cd14;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hb49058634d276b9b2fe4d66db4279aefcb2e2760ac5752c45a247a0b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1639891326c83660ed10bb7a19bea13efca5e1a4bab6a9bbe19540fa;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1693c745e19a1edc99788c830cf49078c52c132803f7f3b0d040906f8;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hb45a2d69faec394512e5f019f74dc954b6dda39707f402226557d87e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'he0566e7a1f07e5313aeb1c4e60636b17d58ea09223e134195022d572;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1ec1466470a234978aaf53b723f0f9e45f60bb38078ce96f737ddc2ed;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h18946816660c62d547b0e088344f742602007c27ad4e6da2872658ab2;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h13ebe25b8c61fddc6dcf0c289ed93b797b9728266fa9d53cb93e7e34c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hb00282fdde1e5fd70a909a384556cf2f2b11cdece95a5be00cd06ca2;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h14653bd3274dce6cb56b0aae0a946694f554a4c3995a5a40cdd86b1f3;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h8e2b0b372befea68008318122832a78156798e18ea79e7f1df6696d9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1edfeea48c660266a63463414dae0dbc1b906200934395988d234aa94;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hf69ee27257674d96bc7fa0cb8cfbeec2aa2ff65c4fb5fa7d5c25173c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1ab6f458d00cf53a92540fac75602eb10004f1bdabf4ecce617d35e0d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hd3e4b6ea9cd4d8712ce535e2230fbd6232e88a86cb519682dbd7a09a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h55ff71656cbd0ea6ef8bd3f5031460d45c5de702b4bdbd22d462b01a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h446f10b4e3015f3b658be71387068334813a9c807a26c4433f7499b5;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h79f449629ed609a5b3be34ef51031633ab7f6b1c79e3a08e94aae6e0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h26d0c97d13f0021c5c3372f3bf92acf1a42b21dad92fb4a9d5d09c84;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hfe477bdb2ccb9343a365c29cecfb9b25eca2cdfb2e34083cdac82630;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h3610204331aef847a4bab2ac5a57ddd3c9eec22cc67abacedb722658;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h895dbc48b6015a9d815cad80cb21b2f9a1b10bcea230ac4fc5754aeb;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h10990528f4ddc204efec7c96000b8833235e8acd46ca276a2c8ec6e2d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hb36b254f3e9f3c9343333754e89df2578fb6af5bda7709932e44cf3;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h19fa3e23235b81f28a27d3dc32bdac38cc2ac83947bb785dc92dbbabc;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h3d4e0a76de41d81bd27492f9168e52aab99a8fd5d0c2452d42cabdf;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hb46c82ade73ec777d56e5a8e589b48336070ab1a66dbe049bf18e2cb;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h86317dac3e8032010a8cc342d39c2c16c81f59b9ad2153d2a28b076a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h14f162ebbebc6f815230804ce4978bcf85c063489349250e7bd68783c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1dcb34f3eb9969adead9b35ea92eba4313c68b0cf1b923a9825215159;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1c4feb0fa2b496aca997303ad22d88a55891dd50b7bf50628b923e602;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h120699c14d7012a839101373ec4716a96c31320f009fa5976963b2de6;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h8769445bfea14b7b5d2238bf29b7ba08ada712392bba5053922f71e5;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h13f9e1de1e951470b6a349db5b78f3a76aac503cb6185ab19a997bce1;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1056a2b49434cdb7a7ba078d603c0d954d269b821e74732e65d84dd0a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h3c103275cb54dcfaafb21fcea6b02f291be23676dcacc2418c86bdcd;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1aa096e0093e79002746f20d8ee56c2bb215e8e26271ff2c808710539;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hae3c0bfabd07db8e00e93fea011ca3ddec614eedefac108f4bcc5149;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h19e2a19048fe6227049a9c4642c833bb3d85abc8b82d75ad885ca8113;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h3545cc9f88e88274ff8eaec59592ea00f841f4ebdf03da3e75264ed7;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h2ebf2b29f35b5f70511d0b095e50a4b5312d7c8f957a6fc62e52b005;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h2e0e14acd39a0f6315369510db6e1750aa3777ede7f445608eae399d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h115d58da89c3273529584be213e90e08c6a6712a9e33e407d15fcebbe;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h105dedb2052ec7c7ed7f64dfb3286d400e4947866285c317a7cac2537;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h32cea4e5f1c9b9d985d3bf9c3471eacbbe5a9919ccd5d299188c0734;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h7300b9f02355c6f6a0adb45c34b3c591e7d8d034fd99dbdbe5d5211d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hab628cf7255f6f2b2304acfc1eab78e4b175237d70ac586374f2699a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h2d8ad702a08582b286a8409bbec7cd8b2b613433e662e33b97837628;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h91c7e446dbd8d54e0f46d67c9b65aa51c12c495a4cd6b513c206cc4c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hae8de96c57d0bf694dcc39e28739be498317b3be07cdef9be1565d5b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1399a27061592137d9adc5b818515f65dd3566b008c920f708482230;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1b4dcc25af92a924f1d9ac7ed44ceb0848b96c1debe485f5ae54b5f32;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1fe247d80bf06ab320fd6b99f60af5a99ede554413e86ba22013c8c3b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h871095d59f5bf0c9f5e5c310f68d766ff00b96ed6358ffa27e0c0645;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h117f936c8c3244bc9b3a0d2f7e57734728f8cefa58f9078f321d08a81;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'ha6edba51670d34742bad7407dd2b050627f72e8c25740b64897eccd8;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h6f05554efacf8b7d1994bcc8bd5a9442c02a9fb76dc84a4d2f4e83f2;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'ha929ee32d7145622674980ca013fed187131c17c84b4650b783871f5;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hd1e5f030473dc494db0c2023a8f3b8b26e3eac0963980436ad4735f6;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h24cb6bc353689bd15ca4f2f65ec9eec9f5755415814db6f89a5ae86b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1299a5566cc82f18b7ffbf95d32f657147c4e9092b2f598680eaf17ca;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h9d0dfc709b35f5dc276566ab0fad64033c6f6cdc272e05fb108ca468;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h85e03f557262e0055fdb73afac4ccdc03184e07e89241d6b3fd5dd3b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h124e62ca474c5d215a8f5e3bae9f8f852c9c83b001fe27fccd3b272d3;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1e9139246e021b8176f1ce6b5b668d4dda2efa50365c1e40759ae9bdb;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1442313c8887a6e72e37d13ef55093e4b78db10fdf17fc8ca3e30abcf;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'he036fe83731891e01c744ec01be5804dd765b263f6ee6253d0fb459a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h15eaa127c41c2505748105495d3f85c2c94c221f4d4b0aa3336f8229c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h81a7adf7c8278dc194eaea82a32955a0fe536e64a90d5d0b66e98e41;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h8bc7d4c16615539ba3f9801afb368330fa4f3a16e632828c7d70e0fc;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h9b9261eb80ee7879b90ce3620bff05e8f1f8ec904c6931e5291fd473;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h4dbbf75dbfbc768ddc12d55fe02af4506e7fa90e09eca4c683c46925;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h79d408c4b08afcac39c80fb7c08af3c24e5d55ce61691c780d3ddd02;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h15b1e2f29e0742b43701c7719d5b7e094266dc6446c35c84517074655;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1cd66668fccc054399950215a6f6643f76526bbad56f14b03d72744fb;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1609f1af607af3d0b5833b5a1ec4fb93b2c1397df83da3f7c5dc0a884;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h14b15d4c5aec9a173ba0652947e1fffe77f29197984633390d6215323;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hc0ef555a5a2205dab106568b3014d785a34298f1a5da42ae13ac3692;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1e0a35f1e63f0d200c25cfdaa89f65f3263d8b021c368b2a72aab237a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h5b47a31e4dea97694d5660588d4e46103d944d92eba02360225b8d62;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1f8442ba2de231f3de5b018284c4643ef6c963c55514197714c3e09ed;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h12d6416a6915df85d9fedc4b0a05128bea0adc723c25ec6edb32b1cea;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h20640359a48a5d3278dd096ddf2515e19457bb990b1c913eb0eb0455;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h168997c92ad473b3835761385256668e362cbb2417fd824416f140f4b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1c6d84d0c096b86614905cfd56f2764eaa9ab3cccdea9a86c2ad17568;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h198897e58a98a17c30ade6689f42fcf854993b0d04c24004e4f6e3404;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1bdd8091582ce0b60fad37ea4a6d8c94a7ff189e468836a61daf37e23;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h52d03e769aa8d04368e968f1ce8a545d6dcd92d0dbe7c470545bca7e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'ha787d185e3b72c8ddb1b92cc9a1a0597001a3df7a53ed75f42d05a69;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h66ab5824b233492eabbb48a9ecf6420645a7ddd41c9272683ef89261;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'ha07731ee99c0028e11dd2cde466698a7524ed161a7c5ee7a28a55130;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1bd71673ff9de5461472e513a4957d5e056bf52d7e06b85a6f1b18e03;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h16fd5bffaca6e450c09c034d23f230d8b19858650b300555be6dd0b0f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h2378344974ed7f321b15238372cf78368efb6a014ce7ba15b33aa71f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h924e8c1bb2e13f2dad4821c214af99d3144818f4f8d8fe5dd0a1d437;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h94d584e33b655b1867c7861eae99355ea0f0a5ef4d83dcb2bed8fce2;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h29b1daf23d85a64497b992d0f635712812de30dbffb220a87accbfb;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h173688946fc62b97df66db8aceb8f73c37701d5a3e0e20c346b48dac7;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h18db5296ac258ccf7abea93c79a49599e88b058f58fefe7f9572ecf6d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hbc3f120dc4ed4b07bdefb71b78429c3d8a8850f2c45425f2d20052e9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hbc8f0f01acbca4262235a60a46a8c1ac5201e66b2b80329ff46e222e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'ha7aeda6f85b95bd2be41a617be32768831d58d8dfa7d4b33d0899da9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h139c37a5bc0aa0a36f549b6ac83902ee5bfbb2c0032607723639577b3;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h198bf7640b506ecc9f5c638b9cc095d494e8760eef82d9e5623d92d8c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h123a55a629c3dc7c9213c3f9adce1b5fca24bf8630c61186860136fb8;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h10df1d4841e8c68496d152c644a43720840b425217fe57dbd4264c0b6;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h10f9ba1acbaccc9be170a7318f7ca2d883a238ddedc12c80ac755a59e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h177eb9c30e10bbd9c0e5434bff1cb5b1aed373c78d48cd96295239456;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h18b750a99b20b0c0ef6eae67c922c324b06635c05a38959677fb84dda;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'he7dbe5205499932b214969495f91f644d5d8f6fcf1e4f8d346a0c13b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1a91dc44d765007a603f9a87c67125d3ab3b0d607d3fe8421e2857eb3;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1f3dc3f0eebdbcc62b9e843eb2ef890a87530adce8d8f29c687f991da;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1b170939897d4c5c7a0205f1a81fce77ba0644329f0a738faafc444a0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h8a8eb16a099076634c1645307dca044aea7a15dcfb05313c9ef090d9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hb3f034d32a4ff4037e866105000a27dea251c119508511d8b1360c2c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hd48c1c12ec7255bdb01a087188daf08cfa0c6c8400cf82f14dc232d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1e06184cf0533f8443c7ba1a6d4b67ef2c2d6044da16ffb30028d7a59;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h14de902a2f342b555b56ab7937633750cbab024e879d5159b5d9853cb;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h26b5dc3456d53303676def8eabfc0f65b7174299744f0c7111646056;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1c2670295656ac908602ed50fd85c28d027eab1713cb9168ed28d954f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hafb8bf1f2f0cc0c989bc054ddfc0af9d2f93bed8bb643adea10b0f80;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h6f9af8991ba00405043904d05cd1966988b48316526dc4fbf6f1f279;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h280213727904cf5bb277dd6a67e72eaa46a6178a7398da754cc7c815;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h43f9c9248d7e2900c2f8cb85c7682d5f70b23810bfb14df7bfac1994;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h2d1e2b606de7165f9f870df968178d45225500aac5366ba162c4d62b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h40f55f518b1562a18bd2ecb312beac032f3f845c9b18df4394e4d10;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h19398799c1ae59d981cf739105a293a9fab086bdf4610c9ca9a6b19f6;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h15d0c7ae86e9d0dd0a1299b584cddc4bc5f65eecf2caa2888daa61f6;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h687031a0bbec4a32848523252eb81ec5c5bf7e9a148359ef110eb6fe;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h97c5a797445a3a6c5821cc1d0b948ae6314096c9b3c5ac6e6901063c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h165ceccfa54a7ea52f6901da6db341dbc26feebaf25a09fe66369a788;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1800691a7ed72f513d462debbecc85aa1545276efe1fe2c0eddbef0ab;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hfe6efac8358eb1fc8c7ec8effbb022e562e50c8f3b22233ec3c1ae20;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1f39b7e09ab340ed8e3a5f635f9576edfca0b3ef3f86bc6ddae923fb7;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'ha8e4f97446516c6c1adc309f85235b9c617b2c078457010f598bfdb2;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1a01d7e228c18471c867dcef1fba0fd260f65566f9983e1d05fdaa229;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h117b4d10a275380b1c74486dd3955f207203cdd7e1d5d11755e376d34;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hd2c2d83c8fbd8e41fa76d1c82775fc61a3ae1f263896c04c5ffaf064;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1151863ae642edf2a6dcd3d2bb633c65bf293ceecb0b41a0356924eef;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h12cf0c6b277748737557382f708a0a1841aa72d901b4af2362e3870cc;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hc63af9edaf286fbcd25595c6b1d2b60d443cf99420b2d8b6b5327d5;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1400b8375782084323607180208929bbbaa5c599be6711d352eb3973b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h194a62e20dc52823b96f715fe0bc154f5d7b18a27d4e7c616fc9b98a5;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1f071edfe1876f6414aff1d7e738efb7b1b01f5c84d94f63dbe78cb21;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h85f369839f02522c4f8cca18426489522c6c7009999eff87802e7e1a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h12516a8e437549cc10709483bbfe07802ed5effe5f78867cad08703ec;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h15f7eddfe7d0b7ca55184d6c7996465399cb12c80a7ea08921fc05255;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h5fb9d4c2bf598b46d75bf21fb8cff685fc745c8b949a3faf8827d718;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hb10127364f139b67c63e70d81b2dd492477f4f70d3b549f860a3f5f8;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h18d9cfa4d960c11801bcc397eeabcf6de5717774aca280b941a62fc1a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1cfa4ad0e6dbfaa75aea33bef4732c5060b4f6b07416e92cb372768e9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1438ad677645265c52c80a02e9959be2bdd90afdef2d7ae14888c51f9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h55f872966f9b8054b2407deac28e0a9d46cc540768fbdbaf7c84b022;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h191f0e7d2ef17dcc19fa6ccc34ce33ce54b928249324ca2cd6a9f7241;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hef23d8edc78fe93688e70acbac100dc767606043d0912e26d05c31b8;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h15475cb1856c11a54d5b6d5b72c4fb288599c2bdc7a62d4faf15ca046;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h18f48bf5fe06afaad9191b90caff9466c099cea3497258cce0428fd8f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h18db057deedead90e56cb8304f6e84f6316c1e7f2b97267cff5a227e9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h52cf56ff1fdae519db29854efacd1d70e001f7c6f66172db5f8fbe4d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1d34524051ffafd9dcead1594751c4c0cfea09d706539a41ea212b738;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hfa8c3724f04c0fc499eea93b2586a65c9f19f237dc9c2af1bc0aea26;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hf50c908028f7f7151db3d39d82ee5da924d825e78b16ef9acfe27319;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1028684edc6cb8b12826322270dd9d441d7e3a5b3c9cf114661925efa;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h17281238204e5cfac9dbbac1b164de1a9015b5a128c0aefcd2ea2890a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h2fa6c57c8dc1c1b06f2caac351f3d860cc79e151d99c6075e3beecd0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h3871f001f0d47021c8e51d131f816aaa7b1bdae707d59cd53ab8a4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h13f0ab42fac77026e11b52735dd197718abfdba7ef78597c826b7c1be;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hdc9dc05438335bc4366cbc88db869e230f212e8845281c8db8b29332;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h7ab206b709e804f9a3191e63579423bb42a02596011c7fc5e3ebb523;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h530f667c49ecdb579ffa3b19c77b0d69fe76b90dbaee4ac63b2fec8c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h14acfb29ae7626db30824ff1a4f01d6c4d7481e0856ef3fcb16e0d042;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1b8f25f60e892c08052e34a9e1c5bdbca6b795759ac6919fbc212b3f7;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h17b6bdf427ae87177cbd9aedd2cf8fbc92e8a61a232736028b90ba0aa;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h2645de40782bcf6177b4c806c50e61302ec547fe9b60b3726cb60958;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'haf8bca8de1a12ac7e80b8944ce9c63ec9d570e1b78da7a9c9703f39;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h192ea235efad953571936e6c6ae98df8b7fa33d6dffa74dfb7ad4148;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h179c7e2786062e8da98fbd511841115f4ba2d0de7cc84a094d0abce1e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h7a1bd42ad5028adeda34018dadcc8bc5769993821f35fce6ee8f950b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h8c6691526e2ef585a62379dcd2ad458e1843a743b5c2e839c1368b71;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h402fa9b859eac46c453fbc3c6f189b836df7f86b19f2cdc9260ce11b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hd97eca16dc6a370a3b010bc048da641f86a9653c62c242286d1e779e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h15edf6f90bdc7ebb0a62fb6f83508c13dab0a1a647cf1e763f76ac1f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hdc1a000706a704bec95cb2e36afb089085b67d56e80e59594b4ebf4e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hefd5e32c41ba44ee34d7d23f8991076f08453767e9d1df045ca4423e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1b2e984ccef853b11419c0229a96a35e92723a5c8b680e5da910ed6e3;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h744c5598ae83cdfe53e2e735c42de7702675e13715833f5b86380e00;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h53c6b5524d8cd828bb898f983e487cf6ce48bc30fecab082d532bb88;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h150dca8da04ac2278f864533dd81c13e3b0a3e933c7081c8ca60adbb2;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h643965ff3020e8d18cd040d64614651d53aef6edaae11f969c15e6d0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1a37ea08a004adfc7cd2ac656ec3796856bce73a6b13860b7653cf9e9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1c56e73a97797103bc70e56e5cd98f1643f52a3903650e53e8141b5da;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h13c3c5fc823c7dd38b1806460aaab089b32ccc4d34285bad0577ebe18;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1da7120b58797cb42b3d148e48ddd393f85d0a94668b23377c2dff830;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h16f6a9c5329d9b073efe9d02900370c2b0648e06113145c846a762a51;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1be2a18b58eca7868e52eee09fe4de158646d387224e8866ae29f5fab;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hdc876ac0fe2e8859a3b93ae7a2c05d1f8e583ef1175cc7da693d251d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h17613838131adc71edf765f2a66a705e6f4a2bc079e67d21fc314b70f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h191e3cdb9e45b5e71ba426af48765d777f65593b32b74519b076db618;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1e7ecc12940394edae951fc2e493d8f07c1a241472697f10b81a699d6;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h192416cc1b81372cec303096491775ca135e7643a867d613007e7e958;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h526d5c2ed639dc2d8559a2fd5c27400a28ff2453cc1ba2433760790d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1bccff02fcd137390d18ecc3ab68b7da454c354cb6b70076b0ec8967;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hd5f266d4a2016a57f2eeb8765328aab3b07b6c2043f3d7b0a6702107;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'he294126155fbd0620b1ba13c18dfaba0427771f776a22f3a6bfbca54;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hf5202ed2d19e898030157dd54abba32404af783d514502e7908163b6;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h12e9e734adc59fd2e16e84dc1721c0fbabd4caba3cc50cdc401deaf47;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h86d2029e3ce6a8999f62fdec1821f7a1a7bde0fb0a5aa39641100c34;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1a656bdd155ed5c356c5fd8d9e98ff4e27cc193afeff8999beaa86973;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h82dfca7c403e2a35f119eea9c216592290a129282d3a359bc5bf1599;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hbd69fc9b3ef3cea4f3450605f9e628d32858b28f167de660e39ed315;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hf3a6365b2f49f5020d12b7c8e225f29d5c909ff842169b23e2c778b6;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h6137e5e08c9811bbeeeb5d79c535a1a3012c9a5a23fd4e961a4b3fe5;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h14ae0d54955030e8e5ffdaa6dd62cbe0131a01ccbb155873a88b3671e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h11c1bb1dda8f89d6599609bc7ac273f433fac60252efb142ee71b8c05;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h14a521730ff9d191b64fcbb7fe4b668884aecbdf166f754dddd4eaef0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1e64ed22de1211d292ee2d21c50fcf0bd4d82be0caf56ab3269544205;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h379460bd923521e3d76c4b55e6199b6453986e8c0bb5afd89cf497ff;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hbedf4fdc95fddf383684ee72167b17b44fc6543fec5c3a3d7d518186;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hd0e03d9e7319fc91d5b00cfc66677f349b040b78a8a40be854bf16b1;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h443d3be167ad47fa94103fee01a028f91e5ffa61fa5b092869d2116f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h103a5778fa4d2fb3d49d0d2d0daa08f0ec1d3c4e087a5dfa9e3003033;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h11d8ad74a8155ef2d300d337ae9fe2fb2fc9d4b3eef310b6eaad870ea;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1fc8434e172da5992bb99e5b2462f5af57ad37ab2e27e18fc414f1a07;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h163bc8b5696d7593507259127b3563dc65df3f6b8ae7a7d8806a0e67d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h62f4c5fbddea3ab5e6ac7aefecade7b6fcba43326acadb202fdcbdc2;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h81b10b01f4ffea0553cbc5d45eb63317cae27e28cef9a2a923dcefef;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h14b14b40d4ff4984db1a45848a643c97e714d2fc88b86f8bcbee45f7c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h14bc3c10f00bed4d08928c70345886c14bb7118d59e31a178fbe668f3;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1dad4ea137b6366fa846962af9678920fc580b504b4fe279e78accaa;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h11be41bd7120046242ad05655df58b2dc6df0ceae3c47c92fe0b25e01;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h5f5010de6e49c6b5fa68c8d3086244fd26aa4b1067a81ad083c3b77d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hec5d650d3c1d68d52a59c7d5b8b3226fe8aa54789711a8eada36024e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1c47e7cc978a2c9798e5aa87731c0068615d1e20ce1292849306f27ed;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h16353c2b63b8fe44a5fa4f0338ccab1ccf64cc3c14b20136147dc687f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h15dbdf91bc5ac98294d475b4b7b8fba6641674bbbbdc2faa703ae94b6;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1d4001233e7e0004dc89ec914e634da6daa4f05770e6382bd6b134976;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h7d539ab867049710481ad95f7b9cf8f4621b52f5821da1dd2de86165;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hcb224601e603eb118a96f66eaaee34af01628954ec452a9e293b8f3f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h168f42b961deee1d1cc477d7eeceac5877aa830056c7dd2b9ff8f605d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h9d096651399e088cd28b110a3d1b2f43c27ff83fd9c63f91be7af3ea;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h11ccd2257bd665cf34b44cb50124843881c85fc390f1ca9e095c51045;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1a4bd731391b2c5fa5a60f6c68effe54ceab60aecdd672be77d3c0b90;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1bf19c361cc2ea4301d62177613c39a4ed1d1aa3020f8fdc08b1689dc;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1ae3ea4809fb8b6b43d2b6338a518adf968f25eb2ec9319f2957c7b38;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h617bd162c2b0cf0080ddd4e384e42263bf4bfe195a3c369edf2a543f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hda11a93685deb5f2066e5056a3c1cf0df039f37adf284e141c5792b0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hc2c454cc22afa60644cc26435764caf24f0c34aa717a334105281833;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h10637541b59a8aae9c7d5ac9314085d6a2d0b2e3667893024be34e4b6;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h21acc1116915a5c3545da0158eb5dc4a5c1498fc21093d428e7d9321;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h82dc260dea439feac8df4cd15d65a2056b08042f4cf892e111c2abe4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'he6d6f8253148fec7402d402728c337492a8d0870f7b5178159b141fa;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h2014bffd9e1bfaaaf37694d26ef1325fd1a83f399d6b748738f34d35;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hf63a7d686c71b8a47b80a415a3151b6d20b6f2e284cbbb8544be7da4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hd54453397c65c806deb1b658ee4dfeec572a7d102a2a263c745627f4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h900d38251057f2faea7dbad82c4fca46f6bbcf5e75495341f74552ce;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h444de318525c0083bb67afdfe6d05a92ae76a7d08e55b0af361c8a25;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h63f7d93b1ea3ab7883c276fa7c75887d4fb4d48a4613ae44f1744ed8;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h185bbb18dcd17661ae36ec3b2e3a8aff685824ba3fbb953c326b235d4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h11324e855b64ed108b991c794900cf9f28ffe880f5cf1939dafa6124f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1d36c27fa580beb09789f324023e7c81150978e66c805aa961c3f6d3a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h9b2c505d8b9672456147a39d7467a6132a7f1bbe2be4b0978d455aa7;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'had3d95cfaa068eeaf78b8e4af2f5fb08b86a2005d728ea4da3f8acd8;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h16831b43fca570a89c25adea1863f5abf42cfa767033ea5a5f04d3b4a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h11a7eb09d9de8895e926d85bf0bc3609389815c3847ab4162fa936d81;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hc70e3ab988ebeb621f4931f90e057f77eb8e1765a8160a3c54caa41;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h12e77d85a4e2742f1b612f5a45428af45ec7b2609c4e6b3198ff256bb;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h86560a33ca4ef5b29789a2764876caaeb690ecd0483fb399dbd162e0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1442d5a27c82b65f3ea34411c3c1145472764644089f3b1dbeefb3918;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h13ad64c658eddce8c02dfe4327f374fc25c40db3eb8ef7d7e49996d03;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h7e9009211629ce08ece1ffe3ba6857820b8d677d296bb92a454ec570;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h191dc4c773d3322980a0fb2b52ee801f2a6d7bca2e943e5ff3ae299be;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h39d2c2716f81265c7221ca33d7b2472e0e7ad13a6f9d539059870e23;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1bd1ae7d45d1329fbb654d3835db1ba417c6c57cdcc302970a5328f89;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h16c2b27987167d2ef0c7c20cc31cd71a1910ee87dfe10949fe7fa2eab;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h8043c3152ccc64c166cfa979ef3683dc81b3014fbf554481324afef6;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h179c9f870649a9e313e7c4d1085c665c34b4f02db14f63a8c533795cc;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1f2ce0f1b08e9bc11182040345a15bf73dfe0541e2ca741d84054e965;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1542e8d60ad448519c39180885f62d7c3dd4688c537da17dccbb8279f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h684454e61184b6685869dd6e3aa17d6109bd8b78e561381b245496b1;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h2e9147f7de45e830c2ba3369da6069be57281e368ffb9d46b6ad63a2;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h10e173f7d7e0c02475fe1e3086ce40d39a47a0020cb751bb6ed520b21;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h43c454a728fbcc23278789336c7a73d0e797495087e22a13af15606c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h58157d4f6beb8cb3041c2e0a690bb27e1247e691075b6e9ab72bae4d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h332ea23ad6241b3c2b2a77331fe1c70fad42739153d83f9fa464e996;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h7e7f17c32c2c071c84c9b8a7a19072be207aa4a52c54c039ee34928c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h155e10e91eba1f60117857fb3a29bcca39c5fe650a0ad40dd99587d2;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h16e70ef5f9ab3729a6d04a1b7d1b3c27f90f0d94867fef155a3951d9a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hd6491b6f4e42762075bc58fc1ef2b7b33bf9874d0fe90da654859da1;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h5aedbaf079cfb46d0c8687a320d5444925ece45f7ad986d23f218234;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h503e0e22ab15f71f99de655f347287af8fde554d6cd5cd8807ce8b21;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h120389711548cd974b58cf8741b93bbc88562709cda0cd3c1a5b4ee02;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'ha85b63d1f09c823af076718ad8aab83546f0866885c1ef33b22d735;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h5326a1d30ba1fba108d2ce53ac72c59b9664f0276dce24edde1bac68;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h11a54b5961201c5353a455f57697f64599fd0b83015ca57261c0d10d0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h11104b5cb48471a247c4685fa8c91416a5209cae4f1fadbd3c0a64f17;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h114058851b1d0f9ffc6e407bfba07eb0b46560ef7748846d22b839408;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1dad376bf5bab3a699b5a3c942cf33a93ae7da7ea8e025806a15fea2;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1ebbae64a69d997d613640ff9964543dddff40ebf518f94e3e32a300;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hf6366be0e3c76f128e81b55bcf1d277ba60aa9f83312c1299fd589e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hdab04448f1ff5d08d6c50156a5336637caf7ec7fa24494e6e7f34993;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'ha45947d1efffc3066573b2613bda31ef94f536c3b1a8491b35512c30;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h6ba014df3e26da4cffcfe59df8730960b79c7ecd63182c277df203c;
        #1
        $finish();
    end
endmodule
