module shift_register(
        input wire clk,
        input wire src0_,
        input wire src1_,
        input wire src2_,
        input wire src3_,
        input wire src4_,
        input wire src5_,
        input wire src6_,
        input wire src7_,
        input wire src8_,
        input wire src9_,
        input wire src10_,
        input wire src11_,
        input wire src12_,
        input wire src13_,
        input wire src14_,
        input wire src15_,
        input wire src16_,
        input wire src17_,
        input wire src18_,
        input wire src19_,
        input wire src20_,
        input wire src21_,
        input wire src22_,
        input wire src23_,
        input wire src24_,
        input wire src25_,
        input wire src26_,
        input wire src27_,
        input wire src28_,
        input wire src29_,
        input wire src30_,
        input wire src31_,
        output wire [0:0] dst0,
        output wire [0:0] dst1,
        output wire [0:0] dst2,
        output wire [0:0] dst3,
        output wire [0:0] dst4,
        output wire [0:0] dst5,
        output wire [0:0] dst6,
        output wire [0:0] dst7,
        output wire [0:0] dst8,
        output wire [0:0] dst9,
        output wire [0:0] dst10,
        output wire [0:0] dst11,
        output wire [0:0] dst12,
        output wire [0:0] dst13,
        output wire [0:0] dst14,
        output wire [0:0] dst15,
        output wire [0:0] dst16,
        output wire [0:0] dst17,
        output wire [0:0] dst18,
        output wire [0:0] dst19,
        output wire [0:0] dst20,
        output wire [0:0] dst21,
        output wire [0:0] dst22,
        output wire [0:0] dst23,
        output wire [0:0] dst24,
        output wire [0:0] dst25,
        output wire [0:0] dst26,
        output wire [0:0] dst27,
        output wire [0:0] dst28,
        output wire [0:0] dst29,
        output wire [0:0] dst30,
        output wire [0:0] dst31,
        output wire [0:0] dst32,
        output wire [0:0] dst33,
        output wire [0:0] dst34,
        output wire [0:0] dst35,
        output wire [0:0] dst36,
        output wire [0:0] dst37,
        output wire [0:0] dst38,
        output wire [0:0] dst39);
    reg [161:0] src0;
    reg [161:0] src1;
    reg [161:0] src2;
    reg [161:0] src3;
    reg [161:0] src4;
    reg [161:0] src5;
    reg [161:0] src6;
    reg [161:0] src7;
    reg [161:0] src8;
    reg [161:0] src9;
    reg [161:0] src10;
    reg [161:0] src11;
    reg [161:0] src12;
    reg [161:0] src13;
    reg [161:0] src14;
    reg [161:0] src15;
    reg [161:0] src16;
    reg [161:0] src17;
    reg [161:0] src18;
    reg [161:0] src19;
    reg [161:0] src20;
    reg [161:0] src21;
    reg [161:0] src22;
    reg [161:0] src23;
    reg [161:0] src24;
    reg [161:0] src25;
    reg [161:0] src26;
    reg [161:0] src27;
    reg [161:0] src28;
    reg [161:0] src29;
    reg [161:0] src30;
    reg [161:0] src31;
    compressor2_1_162_32 compressor2_1_162_32(
            .src0(src0),
            .src1(src1),
            .src2(src2),
            .src3(src3),
            .src4(src4),
            .src5(src5),
            .src6(src6),
            .src7(src7),
            .src8(src8),
            .src9(src9),
            .src10(src10),
            .src11(src11),
            .src12(src12),
            .src13(src13),
            .src14(src14),
            .src15(src15),
            .src16(src16),
            .src17(src17),
            .src18(src18),
            .src19(src19),
            .src20(src20),
            .src21(src21),
            .src22(src22),
            .src23(src23),
            .src24(src24),
            .src25(src25),
            .src26(src26),
            .src27(src27),
            .src28(src28),
            .src29(src29),
            .src30(src30),
            .src31(src31),
            .dst0(dst0),
            .dst1(dst1),
            .dst2(dst2),
            .dst3(dst3),
            .dst4(dst4),
            .dst5(dst5),
            .dst6(dst6),
            .dst7(dst7),
            .dst8(dst8),
            .dst9(dst9),
            .dst10(dst10),
            .dst11(dst11),
            .dst12(dst12),
            .dst13(dst13),
            .dst14(dst14),
            .dst15(dst15),
            .dst16(dst16),
            .dst17(dst17),
            .dst18(dst18),
            .dst19(dst19),
            .dst20(dst20),
            .dst21(dst21),
            .dst22(dst22),
            .dst23(dst23),
            .dst24(dst24),
            .dst25(dst25),
            .dst26(dst26),
            .dst27(dst27),
            .dst28(dst28),
            .dst29(dst29),
            .dst30(dst30),
            .dst31(dst31),
            .dst32(dst32),
            .dst33(dst33),
            .dst34(dst34),
            .dst35(dst35),
            .dst36(dst36),
            .dst37(dst37),
            .dst38(dst38),
            .dst39(dst39));
    initial begin
        src0 <= 162'h0;
        src1 <= 162'h0;
        src2 <= 162'h0;
        src3 <= 162'h0;
        src4 <= 162'h0;
        src5 <= 162'h0;
        src6 <= 162'h0;
        src7 <= 162'h0;
        src8 <= 162'h0;
        src9 <= 162'h0;
        src10 <= 162'h0;
        src11 <= 162'h0;
        src12 <= 162'h0;
        src13 <= 162'h0;
        src14 <= 162'h0;
        src15 <= 162'h0;
        src16 <= 162'h0;
        src17 <= 162'h0;
        src18 <= 162'h0;
        src19 <= 162'h0;
        src20 <= 162'h0;
        src21 <= 162'h0;
        src22 <= 162'h0;
        src23 <= 162'h0;
        src24 <= 162'h0;
        src25 <= 162'h0;
        src26 <= 162'h0;
        src27 <= 162'h0;
        src28 <= 162'h0;
        src29 <= 162'h0;
        src30 <= 162'h0;
        src31 <= 162'h0;
    end
    always @(posedge clk) begin
        src0 <= {src0, src0_};
        src1 <= {src1, src1_};
        src2 <= {src2, src2_};
        src3 <= {src3, src3_};
        src4 <= {src4, src4_};
        src5 <= {src5, src5_};
        src6 <= {src6, src6_};
        src7 <= {src7, src7_};
        src8 <= {src8, src8_};
        src9 <= {src9, src9_};
        src10 <= {src10, src10_};
        src11 <= {src11, src11_};
        src12 <= {src12, src12_};
        src13 <= {src13, src13_};
        src14 <= {src14, src14_};
        src15 <= {src15, src15_};
        src16 <= {src16, src16_};
        src17 <= {src17, src17_};
        src18 <= {src18, src18_};
        src19 <= {src19, src19_};
        src20 <= {src20, src20_};
        src21 <= {src21, src21_};
        src22 <= {src22, src22_};
        src23 <= {src23, src23_};
        src24 <= {src24, src24_};
        src25 <= {src25, src25_};
        src26 <= {src26, src26_};
        src27 <= {src27, src27_};
        src28 <= {src28, src28_};
        src29 <= {src29, src29_};
        src30 <= {src30, src30_};
        src31 <= {src31, src31_};
    end
endmodule
module compressor2_1_162_32(
    input [161:0]src0,
    input [161:0]src1,
    input [161:0]src2,
    input [161:0]src3,
    input [161:0]src4,
    input [161:0]src5,
    input [161:0]src6,
    input [161:0]src7,
    input [161:0]src8,
    input [161:0]src9,
    input [161:0]src10,
    input [161:0]src11,
    input [161:0]src12,
    input [161:0]src13,
    input [161:0]src14,
    input [161:0]src15,
    input [161:0]src16,
    input [161:0]src17,
    input [161:0]src18,
    input [161:0]src19,
    input [161:0]src20,
    input [161:0]src21,
    input [161:0]src22,
    input [161:0]src23,
    input [161:0]src24,
    input [161:0]src25,
    input [161:0]src26,
    input [161:0]src27,
    input [161:0]src28,
    input [161:0]src29,
    input [161:0]src30,
    input [161:0]src31,
    output dst0,
    output dst1,
    output dst2,
    output dst3,
    output dst4,
    output dst5,
    output dst6,
    output dst7,
    output dst8,
    output dst9,
    output dst10,
    output dst11,
    output dst12,
    output dst13,
    output dst14,
    output dst15,
    output dst16,
    output dst17,
    output dst18,
    output dst19,
    output dst20,
    output dst21,
    output dst22,
    output dst23,
    output dst24,
    output dst25,
    output dst26,
    output dst27,
    output dst28,
    output dst29,
    output dst30,
    output dst31,
    output dst32,
    output dst33,
    output dst34,
    output dst35,
    output dst36,
    output dst37,
    output dst38,
    output dst39);

    wire [1:0] comp_out0;
    wire [1:0] comp_out1;
    wire [1:0] comp_out2;
    wire [1:0] comp_out3;
    wire [1:0] comp_out4;
    wire [1:0] comp_out5;
    wire [1:0] comp_out6;
    wire [1:0] comp_out7;
    wire [1:0] comp_out8;
    wire [1:0] comp_out9;
    wire [1:0] comp_out10;
    wire [1:0] comp_out11;
    wire [1:0] comp_out12;
    wire [1:0] comp_out13;
    wire [1:0] comp_out14;
    wire [1:0] comp_out15;
    wire [1:0] comp_out16;
    wire [1:0] comp_out17;
    wire [1:0] comp_out18;
    wire [1:0] comp_out19;
    wire [1:0] comp_out20;
    wire [1:0] comp_out21;
    wire [1:0] comp_out22;
    wire [1:0] comp_out23;
    wire [1:0] comp_out24;
    wire [1:0] comp_out25;
    wire [1:0] comp_out26;
    wire [1:0] comp_out27;
    wire [1:0] comp_out28;
    wire [1:0] comp_out29;
    wire [1:0] comp_out30;
    wire [1:0] comp_out31;
    wire [1:0] comp_out32;
    wire [1:0] comp_out33;
    wire [1:0] comp_out34;
    wire [1:0] comp_out35;
    wire [1:0] comp_out36;
    wire [1:0] comp_out37;
    wire [1:0] comp_out38;
    compressor compressor_inst(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .src31(src31),
        .dst0(comp_out0),
        .dst1(comp_out1),
        .dst2(comp_out2),
        .dst3(comp_out3),
        .dst4(comp_out4),
        .dst5(comp_out5),
        .dst6(comp_out6),
        .dst7(comp_out7),
        .dst8(comp_out8),
        .dst9(comp_out9),
        .dst10(comp_out10),
        .dst11(comp_out11),
        .dst12(comp_out12),
        .dst13(comp_out13),
        .dst14(comp_out14),
        .dst15(comp_out15),
        .dst16(comp_out16),
        .dst17(comp_out17),
        .dst18(comp_out18),
        .dst19(comp_out19),
        .dst20(comp_out20),
        .dst21(comp_out21),
        .dst22(comp_out22),
        .dst23(comp_out23),
        .dst24(comp_out24),
        .dst25(comp_out25),
        .dst26(comp_out26),
        .dst27(comp_out27),
        .dst28(comp_out28),
        .dst29(comp_out29),
        .dst30(comp_out30),
        .dst31(comp_out31),
        .dst32(comp_out32),
        .dst33(comp_out33),
        .dst34(comp_out34),
        .dst35(comp_out35),
        .dst36(comp_out36),
        .dst37(comp_out37),
        .dst38(comp_out38)
    );
    rowadder2_1_39 rowadder2_1inst(
        .src0({comp_out38[0], comp_out37[0], comp_out36[0], comp_out35[0], comp_out34[0], comp_out33[0], comp_out32[0], comp_out31[0], comp_out30[0], comp_out29[0], comp_out28[0], comp_out27[0], comp_out26[0], comp_out25[0], comp_out24[0], comp_out23[0], comp_out22[0], comp_out21[0], comp_out20[0], comp_out19[0], comp_out18[0], comp_out17[0], comp_out16[0], comp_out15[0], comp_out14[0], comp_out13[0], comp_out12[0], comp_out11[0], comp_out10[0], comp_out9[0], comp_out8[0], comp_out7[0], comp_out6[0], comp_out5[0], comp_out4[0], comp_out3[0], comp_out2[0], comp_out1[0], comp_out0[0]}),
        .src1({comp_out38[1], comp_out37[1], comp_out36[1], comp_out35[1], comp_out34[1], comp_out33[1], comp_out32[1], comp_out31[1], comp_out30[1], comp_out29[1], comp_out28[1], comp_out27[1], comp_out26[1], comp_out25[1], comp_out24[1], comp_out23[1], comp_out22[1], comp_out21[1], comp_out20[1], comp_out19[1], comp_out18[1], comp_out17[1], comp_out16[1], comp_out15[1], comp_out14[1], comp_out13[1], comp_out12[1], comp_out11[1], comp_out10[1], comp_out9[1], comp_out8[1], comp_out7[1], comp_out6[1], comp_out5[1], comp_out4[1], comp_out3[1], comp_out2[1], comp_out1[1], comp_out0[1]}),
        .dst0({dst39, dst38, dst37, dst36, dst35, dst34, dst33, dst32, dst31, dst30, dst29, dst28, dst27, dst26, dst25, dst24, dst23, dst22, dst21, dst20, dst19, dst18, dst17, dst16, dst15, dst14, dst13, dst12, dst11, dst10, dst9, dst8, dst7, dst6, dst5, dst4, dst3, dst2, dst1, dst0})
    );
endmodule
module compressor (
      input wire [161:0] src0,
      input wire [161:0] src1,
      input wire [161:0] src2,
      input wire [161:0] src3,
      input wire [161:0] src4,
      input wire [161:0] src5,
      input wire [161:0] src6,
      input wire [161:0] src7,
      input wire [161:0] src8,
      input wire [161:0] src9,
      input wire [161:0] src10,
      input wire [161:0] src11,
      input wire [161:0] src12,
      input wire [161:0] src13,
      input wire [161:0] src14,
      input wire [161:0] src15,
      input wire [161:0] src16,
      input wire [161:0] src17,
      input wire [161:0] src18,
      input wire [161:0] src19,
      input wire [161:0] src20,
      input wire [161:0] src21,
      input wire [161:0] src22,
      input wire [161:0] src23,
      input wire [161:0] src24,
      input wire [161:0] src25,
      input wire [161:0] src26,
      input wire [161:0] src27,
      input wire [161:0] src28,
      input wire [161:0] src29,
      input wire [161:0] src30,
      input wire [161:0] src31,
      output wire [1:0] dst0,
      output wire [1:0] dst1,
      output wire [1:0] dst2,
      output wire [1:0] dst3,
      output wire [1:0] dst4,
      output wire [1:0] dst5,
      output wire [1:0] dst6,
      output wire [1:0] dst7,
      output wire [1:0] dst8,
      output wire [1:0] dst9,
      output wire [1:0] dst10,
      output wire [1:0] dst11,
      output wire [1:0] dst12,
      output wire [1:0] dst13,
      output wire [1:0] dst14,
      output wire [1:0] dst15,
      output wire [1:0] dst16,
      output wire [1:0] dst17,
      output wire [1:0] dst18,
      output wire [1:0] dst19,
      output wire [1:0] dst20,
      output wire [1:0] dst21,
      output wire [1:0] dst22,
      output wire [1:0] dst23,
      output wire [1:0] dst24,
      output wire [1:0] dst25,
      output wire [1:0] dst26,
      output wire [1:0] dst27,
      output wire [1:0] dst28,
      output wire [1:0] dst29,
      output wire [1:0] dst30,
      output wire [1:0] dst31,
      output wire [1:0] dst32,
      output wire [1:0] dst33,
      output wire [1:0] dst34,
      output wire [1:0] dst35,
      output wire [1:0] dst36,
      output wire [1:0] dst37,
      output wire [1:0] dst38);

   wire [161:0] stage0_0;
   wire [161:0] stage0_1;
   wire [161:0] stage0_2;
   wire [161:0] stage0_3;
   wire [161:0] stage0_4;
   wire [161:0] stage0_5;
   wire [161:0] stage0_6;
   wire [161:0] stage0_7;
   wire [161:0] stage0_8;
   wire [161:0] stage0_9;
   wire [161:0] stage0_10;
   wire [161:0] stage0_11;
   wire [161:0] stage0_12;
   wire [161:0] stage0_13;
   wire [161:0] stage0_14;
   wire [161:0] stage0_15;
   wire [161:0] stage0_16;
   wire [161:0] stage0_17;
   wire [161:0] stage0_18;
   wire [161:0] stage0_19;
   wire [161:0] stage0_20;
   wire [161:0] stage0_21;
   wire [161:0] stage0_22;
   wire [161:0] stage0_23;
   wire [161:0] stage0_24;
   wire [161:0] stage0_25;
   wire [161:0] stage0_26;
   wire [161:0] stage0_27;
   wire [161:0] stage0_28;
   wire [161:0] stage0_29;
   wire [161:0] stage0_30;
   wire [161:0] stage0_31;
   wire [49:0] stage1_0;
   wire [55:0] stage1_1;
   wire [55:0] stage1_2;
   wire [75:0] stage1_3;
   wire [94:0] stage1_4;
   wire [53:0] stage1_5;
   wire [105:0] stage1_6;
   wire [65:0] stage1_7;
   wire [53:0] stage1_8;
   wire [76:0] stage1_9;
   wire [92:0] stage1_10;
   wire [66:0] stage1_11;
   wire [55:0] stage1_12;
   wire [85:0] stage1_13;
   wire [68:0] stage1_14;
   wire [59:0] stage1_15;
   wire [106:0] stage1_16;
   wire [63:0] stage1_17;
   wire [81:0] stage1_18;
   wire [66:0] stage1_19;
   wire [60:0] stage1_20;
   wire [79:0] stage1_21;
   wire [81:0] stage1_22;
   wire [90:0] stage1_23;
   wire [66:0] stage1_24;
   wire [77:0] stage1_25;
   wire [54:0] stage1_26;
   wire [66:0] stage1_27;
   wire [77:0] stage1_28;
   wire [74:0] stage1_29;
   wire [62:0] stage1_30;
   wire [97:0] stage1_31;
   wire [44:0] stage1_32;
   wire [18:0] stage1_33;
   wire [10:0] stage2_0;
   wire [16:0] stage2_1;
   wire [16:0] stage2_2;
   wire [34:0] stage2_3;
   wire [40:0] stage2_4;
   wire [27:0] stage2_5;
   wire [30:0] stage2_6;
   wire [33:0] stage2_7;
   wire [32:0] stage2_8;
   wire [31:0] stage2_9;
   wire [45:0] stage2_10;
   wire [38:0] stage2_11;
   wire [23:0] stage2_12;
   wire [44:0] stage2_13;
   wire [36:0] stage2_14;
   wire [33:0] stage2_15;
   wire [43:0] stage2_16;
   wire [36:0] stage2_17;
   wire [28:0] stage2_18;
   wire [27:0] stage2_19;
   wire [37:0] stage2_20;
   wire [27:0] stage2_21;
   wire [33:0] stage2_22;
   wire [43:0] stage2_23;
   wire [34:0] stage2_24;
   wire [30:0] stage2_25;
   wire [30:0] stage2_26;
   wire [32:0] stage2_27;
   wire [29:0] stage2_28;
   wire [32:0] stage2_29;
   wire [36:0] stage2_30;
   wire [35:0] stage2_31;
   wire [40:0] stage2_32;
   wire [23:0] stage2_33;
   wire [6:0] stage2_34;
   wire [1:0] stage2_35;
   wire [6:0] stage3_0;
   wire [9:0] stage3_1;
   wire [9:0] stage3_2;
   wire [22:0] stage3_3;
   wire [8:0] stage3_4;
   wire [11:0] stage3_5;
   wire [16:0] stage3_6;
   wire [18:0] stage3_7;
   wire [17:0] stage3_8;
   wire [18:0] stage3_9;
   wire [14:0] stage3_10;
   wire [14:0] stage3_11;
   wire [14:0] stage3_12;
   wire [17:0] stage3_13;
   wire [16:0] stage3_14;
   wire [15:0] stage3_15;
   wire [12:0] stage3_16;
   wire [16:0] stage3_17;
   wire [16:0] stage3_18;
   wire [11:0] stage3_19;
   wire [17:0] stage3_20;
   wire [14:0] stage3_21;
   wire [22:0] stage3_22;
   wire [12:0] stage3_23;
   wire [16:0] stage3_24;
   wire [16:0] stage3_25;
   wire [11:0] stage3_26;
   wire [12:0] stage3_27;
   wire [22:0] stage3_28;
   wire [10:0] stage3_29;
   wire [13:0] stage3_30;
   wire [16:0] stage3_31;
   wire [15:0] stage3_32;
   wire [16:0] stage3_33;
   wire [15:0] stage3_34;
   wire [4:0] stage3_35;
   wire [1:0] stage4_0;
   wire [5:0] stage4_1;
   wire [5:0] stage4_2;
   wire [10:0] stage4_3;
   wire [5:0] stage4_4;
   wire [3:0] stage4_5;
   wire [5:0] stage4_6;
   wire [7:0] stage4_7;
   wire [6:0] stage4_8;
   wire [7:0] stage4_9;
   wire [7:0] stage4_10;
   wire [9:0] stage4_11;
   wire [8:0] stage4_12;
   wire [4:0] stage4_13;
   wire [5:0] stage4_14;
   wire [9:0] stage4_15;
   wire [6:0] stage4_16;
   wire [12:0] stage4_17;
   wire [8:0] stage4_18;
   wire [11:0] stage4_19;
   wire [5:0] stage4_20;
   wire [5:0] stage4_21;
   wire [8:0] stage4_22;
   wire [6:0] stage4_23;
   wire [7:0] stage4_24;
   wire [8:0] stage4_25;
   wire [8:0] stage4_26;
   wire [4:0] stage4_27;
   wire [8:0] stage4_28;
   wire [5:0] stage4_29;
   wire [5:0] stage4_30;
   wire [5:0] stage4_31;
   wire [10:0] stage4_32;
   wire [7:0] stage4_33;
   wire [8:0] stage4_34;
   wire [3:0] stage4_35;
   wire [2:0] stage4_36;
   wire [1:0] stage4_37;
   wire [1:0] stage5_0;
   wire [3:0] stage5_1;
   wire [4:0] stage5_2;
   wire [3:0] stage5_3;
   wire [1:0] stage5_4;
   wire [4:0] stage5_5;
   wire [1:0] stage5_6;
   wire [6:0] stage5_7;
   wire [2:0] stage5_8;
   wire [2:0] stage5_9;
   wire [3:0] stage5_10;
   wire [5:0] stage5_11;
   wire [2:0] stage5_12;
   wire [2:0] stage5_13;
   wire [5:0] stage5_14;
   wire [5:0] stage5_15;
   wire [1:0] stage5_16;
   wire [5:0] stage5_17;
   wire [4:0] stage5_18;
   wire [2:0] stage5_19;
   wire [3:0] stage5_20;
   wire [4:0] stage5_21;
   wire [1:0] stage5_22;
   wire [3:0] stage5_23;
   wire [5:0] stage5_24;
   wire [1:0] stage5_25;
   wire [3:0] stage5_26;
   wire [3:0] stage5_27;
   wire [3:0] stage5_28;
   wire [5:0] stage5_29;
   wire [2:0] stage5_30;
   wire [1:0] stage5_31;
   wire [2:0] stage5_32;
   wire [4:0] stage5_33;
   wire [3:0] stage5_34;
   wire [5:0] stage5_35;
   wire [3:0] stage5_36;
   wire [0:0] stage5_37;
   wire [0:0] stage5_38;
   wire [1:0] stage6_0;
   wire [1:0] stage6_1;
   wire [1:0] stage6_2;
   wire [1:0] stage6_3;
   wire [1:0] stage6_4;
   wire [1:0] stage6_5;
   wire [1:0] stage6_6;
   wire [1:0] stage6_7;
   wire [1:0] stage6_8;
   wire [1:0] stage6_9;
   wire [1:0] stage6_10;
   wire [1:0] stage6_11;
   wire [1:0] stage6_12;
   wire [1:0] stage6_13;
   wire [1:0] stage6_14;
   wire [1:0] stage6_15;
   wire [1:0] stage6_16;
   wire [1:0] stage6_17;
   wire [1:0] stage6_18;
   wire [1:0] stage6_19;
   wire [1:0] stage6_20;
   wire [1:0] stage6_21;
   wire [1:0] stage6_22;
   wire [1:0] stage6_23;
   wire [1:0] stage6_24;
   wire [1:0] stage6_25;
   wire [1:0] stage6_26;
   wire [1:0] stage6_27;
   wire [1:0] stage6_28;
   wire [1:0] stage6_29;
   wire [1:0] stage6_30;
   wire [1:0] stage6_31;
   wire [1:0] stage6_32;
   wire [1:0] stage6_33;
   wire [1:0] stage6_34;
   wire [1:0] stage6_35;
   wire [1:0] stage6_36;
   wire [1:0] stage6_37;
   wire [1:0] stage6_38;

   assign stage0_0 = src0;
   assign stage0_1 = src1;
   assign stage0_2 = src2;
   assign stage0_3 = src3;
   assign stage0_4 = src4;
   assign stage0_5 = src5;
   assign stage0_6 = src6;
   assign stage0_7 = src7;
   assign stage0_8 = src8;
   assign stage0_9 = src9;
   assign stage0_10 = src10;
   assign stage0_11 = src11;
   assign stage0_12 = src12;
   assign stage0_13 = src13;
   assign stage0_14 = src14;
   assign stage0_15 = src15;
   assign stage0_16 = src16;
   assign stage0_17 = src17;
   assign stage0_18 = src18;
   assign stage0_19 = src19;
   assign stage0_20 = src20;
   assign stage0_21 = src21;
   assign stage0_22 = src22;
   assign stage0_23 = src23;
   assign stage0_24 = src24;
   assign stage0_25 = src25;
   assign stage0_26 = src26;
   assign stage0_27 = src27;
   assign stage0_28 = src28;
   assign stage0_29 = src29;
   assign stage0_30 = src30;
   assign stage0_31 = src31;
   assign dst0 = stage6_0;
   assign dst1 = stage6_1;
   assign dst2 = stage6_2;
   assign dst3 = stage6_3;
   assign dst4 = stage6_4;
   assign dst5 = stage6_5;
   assign dst6 = stage6_6;
   assign dst7 = stage6_7;
   assign dst8 = stage6_8;
   assign dst9 = stage6_9;
   assign dst10 = stage6_10;
   assign dst11 = stage6_11;
   assign dst12 = stage6_12;
   assign dst13 = stage6_13;
   assign dst14 = stage6_14;
   assign dst15 = stage6_15;
   assign dst16 = stage6_16;
   assign dst17 = stage6_17;
   assign dst18 = stage6_18;
   assign dst19 = stage6_19;
   assign dst20 = stage6_20;
   assign dst21 = stage6_21;
   assign dst22 = stage6_22;
   assign dst23 = stage6_23;
   assign dst24 = stage6_24;
   assign dst25 = stage6_25;
   assign dst26 = stage6_26;
   assign dst27 = stage6_27;
   assign dst28 = stage6_28;
   assign dst29 = stage6_29;
   assign dst30 = stage6_30;
   assign dst31 = stage6_31;
   assign dst32 = stage6_32;
   assign dst33 = stage6_33;
   assign dst34 = stage6_34;
   assign dst35 = stage6_35;
   assign dst36 = stage6_36;
   assign dst37 = stage6_37;
   assign dst38 = stage6_38;

   gpc2135_5 gpc0 (
      {stage0_0[0], stage0_0[1], stage0_0[2], stage0_0[3], stage0_0[4]},
      {stage0_1[0], stage0_1[1], stage0_1[2]},
      {stage0_2[0]},
      {stage0_3[0], stage0_3[1]},
      {stage1_4[0],stage1_3[0],stage1_2[0],stage1_1[0],stage1_0[0]}
   );
   gpc2135_5 gpc1 (
      {stage0_0[5], stage0_0[6], stage0_0[7], stage0_0[8], stage0_0[9]},
      {stage0_1[3], stage0_1[4], stage0_1[5]},
      {stage0_2[1]},
      {stage0_3[2], stage0_3[3]},
      {stage1_4[1],stage1_3[1],stage1_2[1],stage1_1[1],stage1_0[1]}
   );
   gpc2135_5 gpc2 (
      {stage0_0[10], stage0_0[11], stage0_0[12], stage0_0[13], stage0_0[14]},
      {stage0_1[6], stage0_1[7], stage0_1[8]},
      {stage0_2[2]},
      {stage0_3[4], stage0_3[5]},
      {stage1_4[2],stage1_3[2],stage1_2[2],stage1_1[2],stage1_0[2]}
   );
   gpc2135_5 gpc3 (
      {stage0_0[15], stage0_0[16], stage0_0[17], stage0_0[18], stage0_0[19]},
      {stage0_1[9], stage0_1[10], stage0_1[11]},
      {stage0_2[3]},
      {stage0_3[6], stage0_3[7]},
      {stage1_4[3],stage1_3[3],stage1_2[3],stage1_1[3],stage1_0[3]}
   );
   gpc2135_5 gpc4 (
      {stage0_0[20], stage0_0[21], stage0_0[22], stage0_0[23], stage0_0[24]},
      {stage0_1[12], stage0_1[13], stage0_1[14]},
      {stage0_2[4]},
      {stage0_3[8], stage0_3[9]},
      {stage1_4[4],stage1_3[4],stage1_2[4],stage1_1[4],stage1_0[4]}
   );
   gpc2135_5 gpc5 (
      {stage0_0[25], stage0_0[26], stage0_0[27], stage0_0[28], stage0_0[29]},
      {stage0_1[15], stage0_1[16], stage0_1[17]},
      {stage0_2[5]},
      {stage0_3[10], stage0_3[11]},
      {stage1_4[5],stage1_3[5],stage1_2[5],stage1_1[5],stage1_0[5]}
   );
   gpc2135_5 gpc6 (
      {stage0_0[30], stage0_0[31], stage0_0[32], stage0_0[33], stage0_0[34]},
      {stage0_1[18], stage0_1[19], stage0_1[20]},
      {stage0_2[6]},
      {stage0_3[12], stage0_3[13]},
      {stage1_4[6],stage1_3[6],stage1_2[6],stage1_1[6],stage1_0[6]}
   );
   gpc2135_5 gpc7 (
      {stage0_0[35], stage0_0[36], stage0_0[37], stage0_0[38], stage0_0[39]},
      {stage0_1[21], stage0_1[22], stage0_1[23]},
      {stage0_2[7]},
      {stage0_3[14], stage0_3[15]},
      {stage1_4[7],stage1_3[7],stage1_2[7],stage1_1[7],stage1_0[7]}
   );
   gpc2135_5 gpc8 (
      {stage0_0[40], stage0_0[41], stage0_0[42], stage0_0[43], stage0_0[44]},
      {stage0_1[24], stage0_1[25], stage0_1[26]},
      {stage0_2[8]},
      {stage0_3[16], stage0_3[17]},
      {stage1_4[8],stage1_3[8],stage1_2[8],stage1_1[8],stage1_0[8]}
   );
   gpc2135_5 gpc9 (
      {stage0_0[45], stage0_0[46], stage0_0[47], stage0_0[48], stage0_0[49]},
      {stage0_1[27], stage0_1[28], stage0_1[29]},
      {stage0_2[9]},
      {stage0_3[18], stage0_3[19]},
      {stage1_4[9],stage1_3[9],stage1_2[9],stage1_1[9],stage1_0[9]}
   );
   gpc2135_5 gpc10 (
      {stage0_0[50], stage0_0[51], stage0_0[52], stage0_0[53], stage0_0[54]},
      {stage0_1[30], stage0_1[31], stage0_1[32]},
      {stage0_2[10]},
      {stage0_3[20], stage0_3[21]},
      {stage1_4[10],stage1_3[10],stage1_2[10],stage1_1[10],stage1_0[10]}
   );
   gpc2135_5 gpc11 (
      {stage0_0[55], stage0_0[56], stage0_0[57], stage0_0[58], stage0_0[59]},
      {stage0_1[33], stage0_1[34], stage0_1[35]},
      {stage0_2[11]},
      {stage0_3[22], stage0_3[23]},
      {stage1_4[11],stage1_3[11],stage1_2[11],stage1_1[11],stage1_0[11]}
   );
   gpc1163_5 gpc12 (
      {stage0_0[60], stage0_0[61], stage0_0[62]},
      {stage0_1[36], stage0_1[37], stage0_1[38], stage0_1[39], stage0_1[40], stage0_1[41]},
      {stage0_2[12]},
      {stage0_3[24]},
      {stage1_4[12],stage1_3[12],stage1_2[12],stage1_1[12],stage1_0[12]}
   );
   gpc1163_5 gpc13 (
      {stage0_0[63], stage0_0[64], stage0_0[65]},
      {stage0_1[42], stage0_1[43], stage0_1[44], stage0_1[45], stage0_1[46], stage0_1[47]},
      {stage0_2[13]},
      {stage0_3[25]},
      {stage1_4[13],stage1_3[13],stage1_2[13],stage1_1[13],stage1_0[13]}
   );
   gpc1163_5 gpc14 (
      {stage0_0[66], stage0_0[67], stage0_0[68]},
      {stage0_1[48], stage0_1[49], stage0_1[50], stage0_1[51], stage0_1[52], stage0_1[53]},
      {stage0_2[14]},
      {stage0_3[26]},
      {stage1_4[14],stage1_3[14],stage1_2[14],stage1_1[14],stage1_0[14]}
   );
   gpc1163_5 gpc15 (
      {stage0_0[69], stage0_0[70], stage0_0[71]},
      {stage0_1[54], stage0_1[55], stage0_1[56], stage0_1[57], stage0_1[58], stage0_1[59]},
      {stage0_2[15]},
      {stage0_3[27]},
      {stage1_4[15],stage1_3[15],stage1_2[15],stage1_1[15],stage1_0[15]}
   );
   gpc1163_5 gpc16 (
      {stage0_0[72], stage0_0[73], stage0_0[74]},
      {stage0_1[60], stage0_1[61], stage0_1[62], stage0_1[63], stage0_1[64], stage0_1[65]},
      {stage0_2[16]},
      {stage0_3[28]},
      {stage1_4[16],stage1_3[16],stage1_2[16],stage1_1[16],stage1_0[16]}
   );
   gpc1163_5 gpc17 (
      {stage0_0[75], stage0_0[76], stage0_0[77]},
      {stage0_1[66], stage0_1[67], stage0_1[68], stage0_1[69], stage0_1[70], stage0_1[71]},
      {stage0_2[17]},
      {stage0_3[29]},
      {stage1_4[17],stage1_3[17],stage1_2[17],stage1_1[17],stage1_0[17]}
   );
   gpc1163_5 gpc18 (
      {stage0_0[78], stage0_0[79], stage0_0[80]},
      {stage0_1[72], stage0_1[73], stage0_1[74], stage0_1[75], stage0_1[76], stage0_1[77]},
      {stage0_2[18]},
      {stage0_3[30]},
      {stage1_4[18],stage1_3[18],stage1_2[18],stage1_1[18],stage1_0[18]}
   );
   gpc1163_5 gpc19 (
      {stage0_0[81], stage0_0[82], stage0_0[83]},
      {stage0_1[78], stage0_1[79], stage0_1[80], stage0_1[81], stage0_1[82], stage0_1[83]},
      {stage0_2[19]},
      {stage0_3[31]},
      {stage1_4[19],stage1_3[19],stage1_2[19],stage1_1[19],stage1_0[19]}
   );
   gpc1163_5 gpc20 (
      {stage0_0[84], stage0_0[85], stage0_0[86]},
      {stage0_1[84], stage0_1[85], stage0_1[86], stage0_1[87], stage0_1[88], stage0_1[89]},
      {stage0_2[20]},
      {stage0_3[32]},
      {stage1_4[20],stage1_3[20],stage1_2[20],stage1_1[20],stage1_0[20]}
   );
   gpc1163_5 gpc21 (
      {stage0_0[87], stage0_0[88], stage0_0[89]},
      {stage0_1[90], stage0_1[91], stage0_1[92], stage0_1[93], stage0_1[94], stage0_1[95]},
      {stage0_2[21]},
      {stage0_3[33]},
      {stage1_4[21],stage1_3[21],stage1_2[21],stage1_1[21],stage1_0[21]}
   );
   gpc1163_5 gpc22 (
      {stage0_0[90], stage0_0[91], stage0_0[92]},
      {stage0_1[96], stage0_1[97], stage0_1[98], stage0_1[99], stage0_1[100], stage0_1[101]},
      {stage0_2[22]},
      {stage0_3[34]},
      {stage1_4[22],stage1_3[22],stage1_2[22],stage1_1[22],stage1_0[22]}
   );
   gpc1163_5 gpc23 (
      {stage0_0[93], stage0_0[94], stage0_0[95]},
      {stage0_1[102], stage0_1[103], stage0_1[104], stage0_1[105], stage0_1[106], stage0_1[107]},
      {stage0_2[23]},
      {stage0_3[35]},
      {stage1_4[23],stage1_3[23],stage1_2[23],stage1_1[23],stage1_0[23]}
   );
   gpc606_5 gpc24 (
      {stage0_0[96], stage0_0[97], stage0_0[98], stage0_0[99], stage0_0[100], stage0_0[101]},
      {stage0_2[24], stage0_2[25], stage0_2[26], stage0_2[27], stage0_2[28], stage0_2[29]},
      {stage1_4[24],stage1_3[24],stage1_2[24],stage1_1[24],stage1_0[24]}
   );
   gpc606_5 gpc25 (
      {stage0_0[102], stage0_0[103], stage0_0[104], stage0_0[105], stage0_0[106], stage0_0[107]},
      {stage0_2[30], stage0_2[31], stage0_2[32], stage0_2[33], stage0_2[34], stage0_2[35]},
      {stage1_4[25],stage1_3[25],stage1_2[25],stage1_1[25],stage1_0[25]}
   );
   gpc606_5 gpc26 (
      {stage0_0[108], stage0_0[109], stage0_0[110], stage0_0[111], stage0_0[112], stage0_0[113]},
      {stage0_2[36], stage0_2[37], stage0_2[38], stage0_2[39], stage0_2[40], stage0_2[41]},
      {stage1_4[26],stage1_3[26],stage1_2[26],stage1_1[26],stage1_0[26]}
   );
   gpc606_5 gpc27 (
      {stage0_0[114], stage0_0[115], stage0_0[116], stage0_0[117], stage0_0[118], stage0_0[119]},
      {stage0_2[42], stage0_2[43], stage0_2[44], stage0_2[45], stage0_2[46], stage0_2[47]},
      {stage1_4[27],stage1_3[27],stage1_2[27],stage1_1[27],stage1_0[27]}
   );
   gpc606_5 gpc28 (
      {stage0_0[120], stage0_0[121], stage0_0[122], stage0_0[123], stage0_0[124], stage0_0[125]},
      {stage0_2[48], stage0_2[49], stage0_2[50], stage0_2[51], stage0_2[52], stage0_2[53]},
      {stage1_4[28],stage1_3[28],stage1_2[28],stage1_1[28],stage1_0[28]}
   );
   gpc606_5 gpc29 (
      {stage0_0[126], stage0_0[127], stage0_0[128], stage0_0[129], stage0_0[130], stage0_0[131]},
      {stage0_2[54], stage0_2[55], stage0_2[56], stage0_2[57], stage0_2[58], stage0_2[59]},
      {stage1_4[29],stage1_3[29],stage1_2[29],stage1_1[29],stage1_0[29]}
   );
   gpc606_5 gpc30 (
      {stage0_0[132], stage0_0[133], stage0_0[134], stage0_0[135], stage0_0[136], stage0_0[137]},
      {stage0_2[60], stage0_2[61], stage0_2[62], stage0_2[63], stage0_2[64], stage0_2[65]},
      {stage1_4[30],stage1_3[30],stage1_2[30],stage1_1[30],stage1_0[30]}
   );
   gpc606_5 gpc31 (
      {stage0_0[138], stage0_0[139], stage0_0[140], stage0_0[141], stage0_0[142], stage0_0[143]},
      {stage0_2[66], stage0_2[67], stage0_2[68], stage0_2[69], stage0_2[70], stage0_2[71]},
      {stage1_4[31],stage1_3[31],stage1_2[31],stage1_1[31],stage1_0[31]}
   );
   gpc606_5 gpc32 (
      {stage0_1[108], stage0_1[109], stage0_1[110], stage0_1[111], stage0_1[112], stage0_1[113]},
      {stage0_3[36], stage0_3[37], stage0_3[38], stage0_3[39], stage0_3[40], stage0_3[41]},
      {stage1_5[0],stage1_4[32],stage1_3[32],stage1_2[32],stage1_1[32]}
   );
   gpc606_5 gpc33 (
      {stage0_1[114], stage0_1[115], stage0_1[116], stage0_1[117], stage0_1[118], stage0_1[119]},
      {stage0_3[42], stage0_3[43], stage0_3[44], stage0_3[45], stage0_3[46], stage0_3[47]},
      {stage1_5[1],stage1_4[33],stage1_3[33],stage1_2[33],stage1_1[33]}
   );
   gpc606_5 gpc34 (
      {stage0_1[120], stage0_1[121], stage0_1[122], stage0_1[123], stage0_1[124], stage0_1[125]},
      {stage0_3[48], stage0_3[49], stage0_3[50], stage0_3[51], stage0_3[52], stage0_3[53]},
      {stage1_5[2],stage1_4[34],stage1_3[34],stage1_2[34],stage1_1[34]}
   );
   gpc606_5 gpc35 (
      {stage0_1[126], stage0_1[127], stage0_1[128], stage0_1[129], stage0_1[130], stage0_1[131]},
      {stage0_3[54], stage0_3[55], stage0_3[56], stage0_3[57], stage0_3[58], stage0_3[59]},
      {stage1_5[3],stage1_4[35],stage1_3[35],stage1_2[35],stage1_1[35]}
   );
   gpc606_5 gpc36 (
      {stage0_1[132], stage0_1[133], stage0_1[134], stage0_1[135], stage0_1[136], stage0_1[137]},
      {stage0_3[60], stage0_3[61], stage0_3[62], stage0_3[63], stage0_3[64], stage0_3[65]},
      {stage1_5[4],stage1_4[36],stage1_3[36],stage1_2[36],stage1_1[36]}
   );
   gpc606_5 gpc37 (
      {stage0_1[138], stage0_1[139], stage0_1[140], stage0_1[141], stage0_1[142], stage0_1[143]},
      {stage0_3[66], stage0_3[67], stage0_3[68], stage0_3[69], stage0_3[70], stage0_3[71]},
      {stage1_5[5],stage1_4[37],stage1_3[37],stage1_2[37],stage1_1[37]}
   );
   gpc615_5 gpc38 (
      {stage0_2[72], stage0_2[73], stage0_2[74], stage0_2[75], stage0_2[76]},
      {stage0_3[72]},
      {stage0_4[0], stage0_4[1], stage0_4[2], stage0_4[3], stage0_4[4], stage0_4[5]},
      {stage1_6[0],stage1_5[6],stage1_4[38],stage1_3[38],stage1_2[38]}
   );
   gpc615_5 gpc39 (
      {stage0_2[77], stage0_2[78], stage0_2[79], stage0_2[80], stage0_2[81]},
      {stage0_3[73]},
      {stage0_4[6], stage0_4[7], stage0_4[8], stage0_4[9], stage0_4[10], stage0_4[11]},
      {stage1_6[1],stage1_5[7],stage1_4[39],stage1_3[39],stage1_2[39]}
   );
   gpc615_5 gpc40 (
      {stage0_2[82], stage0_2[83], stage0_2[84], stage0_2[85], stage0_2[86]},
      {stage0_3[74]},
      {stage0_4[12], stage0_4[13], stage0_4[14], stage0_4[15], stage0_4[16], stage0_4[17]},
      {stage1_6[2],stage1_5[8],stage1_4[40],stage1_3[40],stage1_2[40]}
   );
   gpc615_5 gpc41 (
      {stage0_2[87], stage0_2[88], stage0_2[89], stage0_2[90], stage0_2[91]},
      {stage0_3[75]},
      {stage0_4[18], stage0_4[19], stage0_4[20], stage0_4[21], stage0_4[22], stage0_4[23]},
      {stage1_6[3],stage1_5[9],stage1_4[41],stage1_3[41],stage1_2[41]}
   );
   gpc615_5 gpc42 (
      {stage0_2[92], stage0_2[93], stage0_2[94], stage0_2[95], stage0_2[96]},
      {stage0_3[76]},
      {stage0_4[24], stage0_4[25], stage0_4[26], stage0_4[27], stage0_4[28], stage0_4[29]},
      {stage1_6[4],stage1_5[10],stage1_4[42],stage1_3[42],stage1_2[42]}
   );
   gpc615_5 gpc43 (
      {stage0_2[97], stage0_2[98], stage0_2[99], stage0_2[100], stage0_2[101]},
      {stage0_3[77]},
      {stage0_4[30], stage0_4[31], stage0_4[32], stage0_4[33], stage0_4[34], stage0_4[35]},
      {stage1_6[5],stage1_5[11],stage1_4[43],stage1_3[43],stage1_2[43]}
   );
   gpc615_5 gpc44 (
      {stage0_2[102], stage0_2[103], stage0_2[104], stage0_2[105], stage0_2[106]},
      {stage0_3[78]},
      {stage0_4[36], stage0_4[37], stage0_4[38], stage0_4[39], stage0_4[40], stage0_4[41]},
      {stage1_6[6],stage1_5[12],stage1_4[44],stage1_3[44],stage1_2[44]}
   );
   gpc615_5 gpc45 (
      {stage0_2[107], stage0_2[108], stage0_2[109], stage0_2[110], stage0_2[111]},
      {stage0_3[79]},
      {stage0_4[42], stage0_4[43], stage0_4[44], stage0_4[45], stage0_4[46], stage0_4[47]},
      {stage1_6[7],stage1_5[13],stage1_4[45],stage1_3[45],stage1_2[45]}
   );
   gpc615_5 gpc46 (
      {stage0_2[112], stage0_2[113], stage0_2[114], stage0_2[115], stage0_2[116]},
      {stage0_3[80]},
      {stage0_4[48], stage0_4[49], stage0_4[50], stage0_4[51], stage0_4[52], stage0_4[53]},
      {stage1_6[8],stage1_5[14],stage1_4[46],stage1_3[46],stage1_2[46]}
   );
   gpc615_5 gpc47 (
      {stage0_2[117], stage0_2[118], stage0_2[119], stage0_2[120], stage0_2[121]},
      {stage0_3[81]},
      {stage0_4[54], stage0_4[55], stage0_4[56], stage0_4[57], stage0_4[58], stage0_4[59]},
      {stage1_6[9],stage1_5[15],stage1_4[47],stage1_3[47],stage1_2[47]}
   );
   gpc615_5 gpc48 (
      {stage0_2[122], stage0_2[123], stage0_2[124], stage0_2[125], stage0_2[126]},
      {stage0_3[82]},
      {stage0_4[60], stage0_4[61], stage0_4[62], stage0_4[63], stage0_4[64], stage0_4[65]},
      {stage1_6[10],stage1_5[16],stage1_4[48],stage1_3[48],stage1_2[48]}
   );
   gpc615_5 gpc49 (
      {stage0_2[127], stage0_2[128], stage0_2[129], stage0_2[130], stage0_2[131]},
      {stage0_3[83]},
      {stage0_4[66], stage0_4[67], stage0_4[68], stage0_4[69], stage0_4[70], stage0_4[71]},
      {stage1_6[11],stage1_5[17],stage1_4[49],stage1_3[49],stage1_2[49]}
   );
   gpc615_5 gpc50 (
      {stage0_2[132], stage0_2[133], stage0_2[134], stage0_2[135], stage0_2[136]},
      {stage0_3[84]},
      {stage0_4[72], stage0_4[73], stage0_4[74], stage0_4[75], stage0_4[76], stage0_4[77]},
      {stage1_6[12],stage1_5[18],stage1_4[50],stage1_3[50],stage1_2[50]}
   );
   gpc615_5 gpc51 (
      {stage0_2[137], stage0_2[138], stage0_2[139], stage0_2[140], stage0_2[141]},
      {stage0_3[85]},
      {stage0_4[78], stage0_4[79], stage0_4[80], stage0_4[81], stage0_4[82], stage0_4[83]},
      {stage1_6[13],stage1_5[19],stage1_4[51],stage1_3[51],stage1_2[51]}
   );
   gpc615_5 gpc52 (
      {stage0_2[142], stage0_2[143], stage0_2[144], stage0_2[145], stage0_2[146]},
      {stage0_3[86]},
      {stage0_4[84], stage0_4[85], stage0_4[86], stage0_4[87], stage0_4[88], stage0_4[89]},
      {stage1_6[14],stage1_5[20],stage1_4[52],stage1_3[52],stage1_2[52]}
   );
   gpc615_5 gpc53 (
      {stage0_2[147], stage0_2[148], stage0_2[149], stage0_2[150], stage0_2[151]},
      {stage0_3[87]},
      {stage0_4[90], stage0_4[91], stage0_4[92], stage0_4[93], stage0_4[94], stage0_4[95]},
      {stage1_6[15],stage1_5[21],stage1_4[53],stage1_3[53],stage1_2[53]}
   );
   gpc615_5 gpc54 (
      {stage0_2[152], stage0_2[153], stage0_2[154], stage0_2[155], stage0_2[156]},
      {stage0_3[88]},
      {stage0_4[96], stage0_4[97], stage0_4[98], stage0_4[99], stage0_4[100], stage0_4[101]},
      {stage1_6[16],stage1_5[22],stage1_4[54],stage1_3[54],stage1_2[54]}
   );
   gpc615_5 gpc55 (
      {stage0_2[157], stage0_2[158], stage0_2[159], stage0_2[160], stage0_2[161]},
      {stage0_3[89]},
      {stage0_4[102], stage0_4[103], stage0_4[104], stage0_4[105], stage0_4[106], stage0_4[107]},
      {stage1_6[17],stage1_5[23],stage1_4[55],stage1_3[55],stage1_2[55]}
   );
   gpc615_5 gpc56 (
      {stage0_3[90], stage0_3[91], stage0_3[92], stage0_3[93], stage0_3[94]},
      {stage0_4[108]},
      {stage0_5[0], stage0_5[1], stage0_5[2], stage0_5[3], stage0_5[4], stage0_5[5]},
      {stage1_7[0],stage1_6[18],stage1_5[24],stage1_4[56],stage1_3[56]}
   );
   gpc615_5 gpc57 (
      {stage0_3[95], stage0_3[96], stage0_3[97], stage0_3[98], stage0_3[99]},
      {stage0_4[109]},
      {stage0_5[6], stage0_5[7], stage0_5[8], stage0_5[9], stage0_5[10], stage0_5[11]},
      {stage1_7[1],stage1_6[19],stage1_5[25],stage1_4[57],stage1_3[57]}
   );
   gpc615_5 gpc58 (
      {stage0_3[100], stage0_3[101], stage0_3[102], stage0_3[103], stage0_3[104]},
      {stage0_4[110]},
      {stage0_5[12], stage0_5[13], stage0_5[14], stage0_5[15], stage0_5[16], stage0_5[17]},
      {stage1_7[2],stage1_6[20],stage1_5[26],stage1_4[58],stage1_3[58]}
   );
   gpc615_5 gpc59 (
      {stage0_3[105], stage0_3[106], stage0_3[107], stage0_3[108], stage0_3[109]},
      {stage0_4[111]},
      {stage0_5[18], stage0_5[19], stage0_5[20], stage0_5[21], stage0_5[22], stage0_5[23]},
      {stage1_7[3],stage1_6[21],stage1_5[27],stage1_4[59],stage1_3[59]}
   );
   gpc615_5 gpc60 (
      {stage0_3[110], stage0_3[111], stage0_3[112], stage0_3[113], stage0_3[114]},
      {stage0_4[112]},
      {stage0_5[24], stage0_5[25], stage0_5[26], stage0_5[27], stage0_5[28], stage0_5[29]},
      {stage1_7[4],stage1_6[22],stage1_5[28],stage1_4[60],stage1_3[60]}
   );
   gpc615_5 gpc61 (
      {stage0_3[115], stage0_3[116], stage0_3[117], stage0_3[118], stage0_3[119]},
      {stage0_4[113]},
      {stage0_5[30], stage0_5[31], stage0_5[32], stage0_5[33], stage0_5[34], stage0_5[35]},
      {stage1_7[5],stage1_6[23],stage1_5[29],stage1_4[61],stage1_3[61]}
   );
   gpc615_5 gpc62 (
      {stage0_3[120], stage0_3[121], stage0_3[122], stage0_3[123], stage0_3[124]},
      {stage0_4[114]},
      {stage0_5[36], stage0_5[37], stage0_5[38], stage0_5[39], stage0_5[40], stage0_5[41]},
      {stage1_7[6],stage1_6[24],stage1_5[30],stage1_4[62],stage1_3[62]}
   );
   gpc615_5 gpc63 (
      {stage0_3[125], stage0_3[126], stage0_3[127], stage0_3[128], stage0_3[129]},
      {stage0_4[115]},
      {stage0_5[42], stage0_5[43], stage0_5[44], stage0_5[45], stage0_5[46], stage0_5[47]},
      {stage1_7[7],stage1_6[25],stage1_5[31],stage1_4[63],stage1_3[63]}
   );
   gpc615_5 gpc64 (
      {stage0_3[130], stage0_3[131], stage0_3[132], stage0_3[133], stage0_3[134]},
      {stage0_4[116]},
      {stage0_5[48], stage0_5[49], stage0_5[50], stage0_5[51], stage0_5[52], stage0_5[53]},
      {stage1_7[8],stage1_6[26],stage1_5[32],stage1_4[64],stage1_3[64]}
   );
   gpc615_5 gpc65 (
      {stage0_3[135], stage0_3[136], stage0_3[137], stage0_3[138], stage0_3[139]},
      {stage0_4[117]},
      {stage0_5[54], stage0_5[55], stage0_5[56], stage0_5[57], stage0_5[58], stage0_5[59]},
      {stage1_7[9],stage1_6[27],stage1_5[33],stage1_4[65],stage1_3[65]}
   );
   gpc615_5 gpc66 (
      {stage0_3[140], stage0_3[141], stage0_3[142], stage0_3[143], stage0_3[144]},
      {stage0_4[118]},
      {stage0_5[60], stage0_5[61], stage0_5[62], stage0_5[63], stage0_5[64], stage0_5[65]},
      {stage1_7[10],stage1_6[28],stage1_5[34],stage1_4[66],stage1_3[66]}
   );
   gpc615_5 gpc67 (
      {stage0_3[145], stage0_3[146], stage0_3[147], stage0_3[148], stage0_3[149]},
      {stage0_4[119]},
      {stage0_5[66], stage0_5[67], stage0_5[68], stage0_5[69], stage0_5[70], stage0_5[71]},
      {stage1_7[11],stage1_6[29],stage1_5[35],stage1_4[67],stage1_3[67]}
   );
   gpc615_5 gpc68 (
      {stage0_3[150], stage0_3[151], stage0_3[152], stage0_3[153], stage0_3[154]},
      {stage0_4[120]},
      {stage0_5[72], stage0_5[73], stage0_5[74], stage0_5[75], stage0_5[76], stage0_5[77]},
      {stage1_7[12],stage1_6[30],stage1_5[36],stage1_4[68],stage1_3[68]}
   );
   gpc606_5 gpc69 (
      {stage0_4[121], stage0_4[122], stage0_4[123], stage0_4[124], stage0_4[125], stage0_4[126]},
      {stage0_6[0], stage0_6[1], stage0_6[2], stage0_6[3], stage0_6[4], stage0_6[5]},
      {stage1_8[0],stage1_7[13],stage1_6[31],stage1_5[37],stage1_4[69]}
   );
   gpc606_5 gpc70 (
      {stage0_4[127], stage0_4[128], stage0_4[129], stage0_4[130], stage0_4[131], stage0_4[132]},
      {stage0_6[6], stage0_6[7], stage0_6[8], stage0_6[9], stage0_6[10], stage0_6[11]},
      {stage1_8[1],stage1_7[14],stage1_6[32],stage1_5[38],stage1_4[70]}
   );
   gpc606_5 gpc71 (
      {stage0_4[133], stage0_4[134], stage0_4[135], stage0_4[136], stage0_4[137], stage0_4[138]},
      {stage0_6[12], stage0_6[13], stage0_6[14], stage0_6[15], stage0_6[16], stage0_6[17]},
      {stage1_8[2],stage1_7[15],stage1_6[33],stage1_5[39],stage1_4[71]}
   );
   gpc606_5 gpc72 (
      {stage0_5[78], stage0_5[79], stage0_5[80], stage0_5[81], stage0_5[82], stage0_5[83]},
      {stage0_7[0], stage0_7[1], stage0_7[2], stage0_7[3], stage0_7[4], stage0_7[5]},
      {stage1_9[0],stage1_8[3],stage1_7[16],stage1_6[34],stage1_5[40]}
   );
   gpc606_5 gpc73 (
      {stage0_5[84], stage0_5[85], stage0_5[86], stage0_5[87], stage0_5[88], stage0_5[89]},
      {stage0_7[6], stage0_7[7], stage0_7[8], stage0_7[9], stage0_7[10], stage0_7[11]},
      {stage1_9[1],stage1_8[4],stage1_7[17],stage1_6[35],stage1_5[41]}
   );
   gpc606_5 gpc74 (
      {stage0_5[90], stage0_5[91], stage0_5[92], stage0_5[93], stage0_5[94], stage0_5[95]},
      {stage0_7[12], stage0_7[13], stage0_7[14], stage0_7[15], stage0_7[16], stage0_7[17]},
      {stage1_9[2],stage1_8[5],stage1_7[18],stage1_6[36],stage1_5[42]}
   );
   gpc606_5 gpc75 (
      {stage0_5[96], stage0_5[97], stage0_5[98], stage0_5[99], stage0_5[100], stage0_5[101]},
      {stage0_7[18], stage0_7[19], stage0_7[20], stage0_7[21], stage0_7[22], stage0_7[23]},
      {stage1_9[3],stage1_8[6],stage1_7[19],stage1_6[37],stage1_5[43]}
   );
   gpc606_5 gpc76 (
      {stage0_5[102], stage0_5[103], stage0_5[104], stage0_5[105], stage0_5[106], stage0_5[107]},
      {stage0_7[24], stage0_7[25], stage0_7[26], stage0_7[27], stage0_7[28], stage0_7[29]},
      {stage1_9[4],stage1_8[7],stage1_7[20],stage1_6[38],stage1_5[44]}
   );
   gpc606_5 gpc77 (
      {stage0_5[108], stage0_5[109], stage0_5[110], stage0_5[111], stage0_5[112], stage0_5[113]},
      {stage0_7[30], stage0_7[31], stage0_7[32], stage0_7[33], stage0_7[34], stage0_7[35]},
      {stage1_9[5],stage1_8[8],stage1_7[21],stage1_6[39],stage1_5[45]}
   );
   gpc606_5 gpc78 (
      {stage0_5[114], stage0_5[115], stage0_5[116], stage0_5[117], stage0_5[118], stage0_5[119]},
      {stage0_7[36], stage0_7[37], stage0_7[38], stage0_7[39], stage0_7[40], stage0_7[41]},
      {stage1_9[6],stage1_8[9],stage1_7[22],stage1_6[40],stage1_5[46]}
   );
   gpc606_5 gpc79 (
      {stage0_5[120], stage0_5[121], stage0_5[122], stage0_5[123], stage0_5[124], stage0_5[125]},
      {stage0_7[42], stage0_7[43], stage0_7[44], stage0_7[45], stage0_7[46], stage0_7[47]},
      {stage1_9[7],stage1_8[10],stage1_7[23],stage1_6[41],stage1_5[47]}
   );
   gpc606_5 gpc80 (
      {stage0_5[126], stage0_5[127], stage0_5[128], stage0_5[129], stage0_5[130], stage0_5[131]},
      {stage0_7[48], stage0_7[49], stage0_7[50], stage0_7[51], stage0_7[52], stage0_7[53]},
      {stage1_9[8],stage1_8[11],stage1_7[24],stage1_6[42],stage1_5[48]}
   );
   gpc606_5 gpc81 (
      {stage0_5[132], stage0_5[133], stage0_5[134], stage0_5[135], stage0_5[136], stage0_5[137]},
      {stage0_7[54], stage0_7[55], stage0_7[56], stage0_7[57], stage0_7[58], stage0_7[59]},
      {stage1_9[9],stage1_8[12],stage1_7[25],stage1_6[43],stage1_5[49]}
   );
   gpc606_5 gpc82 (
      {stage0_5[138], stage0_5[139], stage0_5[140], stage0_5[141], stage0_5[142], stage0_5[143]},
      {stage0_7[60], stage0_7[61], stage0_7[62], stage0_7[63], stage0_7[64], stage0_7[65]},
      {stage1_9[10],stage1_8[13],stage1_7[26],stage1_6[44],stage1_5[50]}
   );
   gpc606_5 gpc83 (
      {stage0_5[144], stage0_5[145], stage0_5[146], stage0_5[147], stage0_5[148], stage0_5[149]},
      {stage0_7[66], stage0_7[67], stage0_7[68], stage0_7[69], stage0_7[70], stage0_7[71]},
      {stage1_9[11],stage1_8[14],stage1_7[27],stage1_6[45],stage1_5[51]}
   );
   gpc606_5 gpc84 (
      {stage0_5[150], stage0_5[151], stage0_5[152], stage0_5[153], stage0_5[154], stage0_5[155]},
      {stage0_7[72], stage0_7[73], stage0_7[74], stage0_7[75], stage0_7[76], stage0_7[77]},
      {stage1_9[12],stage1_8[15],stage1_7[28],stage1_6[46],stage1_5[52]}
   );
   gpc606_5 gpc85 (
      {stage0_5[156], stage0_5[157], stage0_5[158], stage0_5[159], stage0_5[160], stage0_5[161]},
      {stage0_7[78], stage0_7[79], stage0_7[80], stage0_7[81], stage0_7[82], stage0_7[83]},
      {stage1_9[13],stage1_8[16],stage1_7[29],stage1_6[47],stage1_5[53]}
   );
   gpc606_5 gpc86 (
      {stage0_6[18], stage0_6[19], stage0_6[20], stage0_6[21], stage0_6[22], stage0_6[23]},
      {stage0_8[0], stage0_8[1], stage0_8[2], stage0_8[3], stage0_8[4], stage0_8[5]},
      {stage1_10[0],stage1_9[14],stage1_8[17],stage1_7[30],stage1_6[48]}
   );
   gpc606_5 gpc87 (
      {stage0_6[24], stage0_6[25], stage0_6[26], stage0_6[27], stage0_6[28], stage0_6[29]},
      {stage0_8[6], stage0_8[7], stage0_8[8], stage0_8[9], stage0_8[10], stage0_8[11]},
      {stage1_10[1],stage1_9[15],stage1_8[18],stage1_7[31],stage1_6[49]}
   );
   gpc606_5 gpc88 (
      {stage0_6[30], stage0_6[31], stage0_6[32], stage0_6[33], stage0_6[34], stage0_6[35]},
      {stage0_8[12], stage0_8[13], stage0_8[14], stage0_8[15], stage0_8[16], stage0_8[17]},
      {stage1_10[2],stage1_9[16],stage1_8[19],stage1_7[32],stage1_6[50]}
   );
   gpc606_5 gpc89 (
      {stage0_6[36], stage0_6[37], stage0_6[38], stage0_6[39], stage0_6[40], stage0_6[41]},
      {stage0_8[18], stage0_8[19], stage0_8[20], stage0_8[21], stage0_8[22], stage0_8[23]},
      {stage1_10[3],stage1_9[17],stage1_8[20],stage1_7[33],stage1_6[51]}
   );
   gpc606_5 gpc90 (
      {stage0_6[42], stage0_6[43], stage0_6[44], stage0_6[45], stage0_6[46], stage0_6[47]},
      {stage0_8[24], stage0_8[25], stage0_8[26], stage0_8[27], stage0_8[28], stage0_8[29]},
      {stage1_10[4],stage1_9[18],stage1_8[21],stage1_7[34],stage1_6[52]}
   );
   gpc606_5 gpc91 (
      {stage0_6[48], stage0_6[49], stage0_6[50], stage0_6[51], stage0_6[52], stage0_6[53]},
      {stage0_8[30], stage0_8[31], stage0_8[32], stage0_8[33], stage0_8[34], stage0_8[35]},
      {stage1_10[5],stage1_9[19],stage1_8[22],stage1_7[35],stage1_6[53]}
   );
   gpc615_5 gpc92 (
      {stage0_6[54], stage0_6[55], stage0_6[56], stage0_6[57], stage0_6[58]},
      {stage0_7[84]},
      {stage0_8[36], stage0_8[37], stage0_8[38], stage0_8[39], stage0_8[40], stage0_8[41]},
      {stage1_10[6],stage1_9[20],stage1_8[23],stage1_7[36],stage1_6[54]}
   );
   gpc615_5 gpc93 (
      {stage0_6[59], stage0_6[60], stage0_6[61], stage0_6[62], stage0_6[63]},
      {stage0_7[85]},
      {stage0_8[42], stage0_8[43], stage0_8[44], stage0_8[45], stage0_8[46], stage0_8[47]},
      {stage1_10[7],stage1_9[21],stage1_8[24],stage1_7[37],stage1_6[55]}
   );
   gpc615_5 gpc94 (
      {stage0_6[64], stage0_6[65], stage0_6[66], stage0_6[67], stage0_6[68]},
      {stage0_7[86]},
      {stage0_8[48], stage0_8[49], stage0_8[50], stage0_8[51], stage0_8[52], stage0_8[53]},
      {stage1_10[8],stage1_9[22],stage1_8[25],stage1_7[38],stage1_6[56]}
   );
   gpc615_5 gpc95 (
      {stage0_6[69], stage0_6[70], stage0_6[71], stage0_6[72], stage0_6[73]},
      {stage0_7[87]},
      {stage0_8[54], stage0_8[55], stage0_8[56], stage0_8[57], stage0_8[58], stage0_8[59]},
      {stage1_10[9],stage1_9[23],stage1_8[26],stage1_7[39],stage1_6[57]}
   );
   gpc615_5 gpc96 (
      {stage0_6[74], stage0_6[75], stage0_6[76], stage0_6[77], stage0_6[78]},
      {stage0_7[88]},
      {stage0_8[60], stage0_8[61], stage0_8[62], stage0_8[63], stage0_8[64], stage0_8[65]},
      {stage1_10[10],stage1_9[24],stage1_8[27],stage1_7[40],stage1_6[58]}
   );
   gpc615_5 gpc97 (
      {stage0_6[79], stage0_6[80], stage0_6[81], stage0_6[82], stage0_6[83]},
      {stage0_7[89]},
      {stage0_8[66], stage0_8[67], stage0_8[68], stage0_8[69], stage0_8[70], stage0_8[71]},
      {stage1_10[11],stage1_9[25],stage1_8[28],stage1_7[41],stage1_6[59]}
   );
   gpc615_5 gpc98 (
      {stage0_6[84], stage0_6[85], stage0_6[86], stage0_6[87], stage0_6[88]},
      {stage0_7[90]},
      {stage0_8[72], stage0_8[73], stage0_8[74], stage0_8[75], stage0_8[76], stage0_8[77]},
      {stage1_10[12],stage1_9[26],stage1_8[29],stage1_7[42],stage1_6[60]}
   );
   gpc615_5 gpc99 (
      {stage0_6[89], stage0_6[90], stage0_6[91], stage0_6[92], stage0_6[93]},
      {stage0_7[91]},
      {stage0_8[78], stage0_8[79], stage0_8[80], stage0_8[81], stage0_8[82], stage0_8[83]},
      {stage1_10[13],stage1_9[27],stage1_8[30],stage1_7[43],stage1_6[61]}
   );
   gpc615_5 gpc100 (
      {stage0_6[94], stage0_6[95], stage0_6[96], stage0_6[97], stage0_6[98]},
      {stage0_7[92]},
      {stage0_8[84], stage0_8[85], stage0_8[86], stage0_8[87], stage0_8[88], stage0_8[89]},
      {stage1_10[14],stage1_9[28],stage1_8[31],stage1_7[44],stage1_6[62]}
   );
   gpc615_5 gpc101 (
      {stage0_6[99], stage0_6[100], stage0_6[101], stage0_6[102], stage0_6[103]},
      {stage0_7[93]},
      {stage0_8[90], stage0_8[91], stage0_8[92], stage0_8[93], stage0_8[94], stage0_8[95]},
      {stage1_10[15],stage1_9[29],stage1_8[32],stage1_7[45],stage1_6[63]}
   );
   gpc615_5 gpc102 (
      {stage0_6[104], stage0_6[105], stage0_6[106], stage0_6[107], stage0_6[108]},
      {stage0_7[94]},
      {stage0_8[96], stage0_8[97], stage0_8[98], stage0_8[99], stage0_8[100], stage0_8[101]},
      {stage1_10[16],stage1_9[30],stage1_8[33],stage1_7[46],stage1_6[64]}
   );
   gpc615_5 gpc103 (
      {stage0_6[109], stage0_6[110], stage0_6[111], stage0_6[112], stage0_6[113]},
      {stage0_7[95]},
      {stage0_8[102], stage0_8[103], stage0_8[104], stage0_8[105], stage0_8[106], stage0_8[107]},
      {stage1_10[17],stage1_9[31],stage1_8[34],stage1_7[47],stage1_6[65]}
   );
   gpc615_5 gpc104 (
      {stage0_6[114], stage0_6[115], stage0_6[116], stage0_6[117], stage0_6[118]},
      {stage0_7[96]},
      {stage0_8[108], stage0_8[109], stage0_8[110], stage0_8[111], stage0_8[112], stage0_8[113]},
      {stage1_10[18],stage1_9[32],stage1_8[35],stage1_7[48],stage1_6[66]}
   );
   gpc615_5 gpc105 (
      {stage0_6[119], stage0_6[120], stage0_6[121], stage0_6[122], stage0_6[123]},
      {stage0_7[97]},
      {stage0_8[114], stage0_8[115], stage0_8[116], stage0_8[117], stage0_8[118], stage0_8[119]},
      {stage1_10[19],stage1_9[33],stage1_8[36],stage1_7[49],stage1_6[67]}
   );
   gpc615_5 gpc106 (
      {stage0_7[98], stage0_7[99], stage0_7[100], stage0_7[101], stage0_7[102]},
      {stage0_8[120]},
      {stage0_9[0], stage0_9[1], stage0_9[2], stage0_9[3], stage0_9[4], stage0_9[5]},
      {stage1_11[0],stage1_10[20],stage1_9[34],stage1_8[37],stage1_7[50]}
   );
   gpc615_5 gpc107 (
      {stage0_7[103], stage0_7[104], stage0_7[105], stage0_7[106], stage0_7[107]},
      {stage0_8[121]},
      {stage0_9[6], stage0_9[7], stage0_9[8], stage0_9[9], stage0_9[10], stage0_9[11]},
      {stage1_11[1],stage1_10[21],stage1_9[35],stage1_8[38],stage1_7[51]}
   );
   gpc615_5 gpc108 (
      {stage0_7[108], stage0_7[109], stage0_7[110], stage0_7[111], stage0_7[112]},
      {stage0_8[122]},
      {stage0_9[12], stage0_9[13], stage0_9[14], stage0_9[15], stage0_9[16], stage0_9[17]},
      {stage1_11[2],stage1_10[22],stage1_9[36],stage1_8[39],stage1_7[52]}
   );
   gpc615_5 gpc109 (
      {stage0_7[113], stage0_7[114], stage0_7[115], stage0_7[116], stage0_7[117]},
      {stage0_8[123]},
      {stage0_9[18], stage0_9[19], stage0_9[20], stage0_9[21], stage0_9[22], stage0_9[23]},
      {stage1_11[3],stage1_10[23],stage1_9[37],stage1_8[40],stage1_7[53]}
   );
   gpc615_5 gpc110 (
      {stage0_7[118], stage0_7[119], stage0_7[120], stage0_7[121], stage0_7[122]},
      {stage0_8[124]},
      {stage0_9[24], stage0_9[25], stage0_9[26], stage0_9[27], stage0_9[28], stage0_9[29]},
      {stage1_11[4],stage1_10[24],stage1_9[38],stage1_8[41],stage1_7[54]}
   );
   gpc615_5 gpc111 (
      {stage0_7[123], stage0_7[124], stage0_7[125], stage0_7[126], stage0_7[127]},
      {stage0_8[125]},
      {stage0_9[30], stage0_9[31], stage0_9[32], stage0_9[33], stage0_9[34], stage0_9[35]},
      {stage1_11[5],stage1_10[25],stage1_9[39],stage1_8[42],stage1_7[55]}
   );
   gpc615_5 gpc112 (
      {stage0_7[128], stage0_7[129], stage0_7[130], stage0_7[131], stage0_7[132]},
      {stage0_8[126]},
      {stage0_9[36], stage0_9[37], stage0_9[38], stage0_9[39], stage0_9[40], stage0_9[41]},
      {stage1_11[6],stage1_10[26],stage1_9[40],stage1_8[43],stage1_7[56]}
   );
   gpc615_5 gpc113 (
      {stage0_7[133], stage0_7[134], stage0_7[135], stage0_7[136], stage0_7[137]},
      {stage0_8[127]},
      {stage0_9[42], stage0_9[43], stage0_9[44], stage0_9[45], stage0_9[46], stage0_9[47]},
      {stage1_11[7],stage1_10[27],stage1_9[41],stage1_8[44],stage1_7[57]}
   );
   gpc615_5 gpc114 (
      {stage0_7[138], stage0_7[139], stage0_7[140], stage0_7[141], stage0_7[142]},
      {stage0_8[128]},
      {stage0_9[48], stage0_9[49], stage0_9[50], stage0_9[51], stage0_9[52], stage0_9[53]},
      {stage1_11[8],stage1_10[28],stage1_9[42],stage1_8[45],stage1_7[58]}
   );
   gpc615_5 gpc115 (
      {stage0_7[143], stage0_7[144], stage0_7[145], stage0_7[146], stage0_7[147]},
      {stage0_8[129]},
      {stage0_9[54], stage0_9[55], stage0_9[56], stage0_9[57], stage0_9[58], stage0_9[59]},
      {stage1_11[9],stage1_10[29],stage1_9[43],stage1_8[46],stage1_7[59]}
   );
   gpc615_5 gpc116 (
      {stage0_7[148], stage0_7[149], stage0_7[150], stage0_7[151], stage0_7[152]},
      {stage0_8[130]},
      {stage0_9[60], stage0_9[61], stage0_9[62], stage0_9[63], stage0_9[64], stage0_9[65]},
      {stage1_11[10],stage1_10[30],stage1_9[44],stage1_8[47],stage1_7[60]}
   );
   gpc615_5 gpc117 (
      {stage0_7[153], stage0_7[154], stage0_7[155], stage0_7[156], stage0_7[157]},
      {stage0_8[131]},
      {stage0_9[66], stage0_9[67], stage0_9[68], stage0_9[69], stage0_9[70], stage0_9[71]},
      {stage1_11[11],stage1_10[31],stage1_9[45],stage1_8[48],stage1_7[61]}
   );
   gpc606_5 gpc118 (
      {stage0_8[132], stage0_8[133], stage0_8[134], stage0_8[135], stage0_8[136], stage0_8[137]},
      {stage0_10[0], stage0_10[1], stage0_10[2], stage0_10[3], stage0_10[4], stage0_10[5]},
      {stage1_12[0],stage1_11[12],stage1_10[32],stage1_9[46],stage1_8[49]}
   );
   gpc606_5 gpc119 (
      {stage0_8[138], stage0_8[139], stage0_8[140], stage0_8[141], stage0_8[142], stage0_8[143]},
      {stage0_10[6], stage0_10[7], stage0_10[8], stage0_10[9], stage0_10[10], stage0_10[11]},
      {stage1_12[1],stage1_11[13],stage1_10[33],stage1_9[47],stage1_8[50]}
   );
   gpc606_5 gpc120 (
      {stage0_8[144], stage0_8[145], stage0_8[146], stage0_8[147], stage0_8[148], stage0_8[149]},
      {stage0_10[12], stage0_10[13], stage0_10[14], stage0_10[15], stage0_10[16], stage0_10[17]},
      {stage1_12[2],stage1_11[14],stage1_10[34],stage1_9[48],stage1_8[51]}
   );
   gpc606_5 gpc121 (
      {stage0_8[150], stage0_8[151], stage0_8[152], stage0_8[153], stage0_8[154], stage0_8[155]},
      {stage0_10[18], stage0_10[19], stage0_10[20], stage0_10[21], stage0_10[22], stage0_10[23]},
      {stage1_12[3],stage1_11[15],stage1_10[35],stage1_9[49],stage1_8[52]}
   );
   gpc606_5 gpc122 (
      {stage0_8[156], stage0_8[157], stage0_8[158], stage0_8[159], stage0_8[160], stage0_8[161]},
      {stage0_10[24], stage0_10[25], stage0_10[26], stage0_10[27], stage0_10[28], stage0_10[29]},
      {stage1_12[4],stage1_11[16],stage1_10[36],stage1_9[50],stage1_8[53]}
   );
   gpc615_5 gpc123 (
      {stage0_9[72], stage0_9[73], stage0_9[74], stage0_9[75], stage0_9[76]},
      {stage0_10[30]},
      {stage0_11[0], stage0_11[1], stage0_11[2], stage0_11[3], stage0_11[4], stage0_11[5]},
      {stage1_13[0],stage1_12[5],stage1_11[17],stage1_10[37],stage1_9[51]}
   );
   gpc615_5 gpc124 (
      {stage0_9[77], stage0_9[78], stage0_9[79], stage0_9[80], stage0_9[81]},
      {stage0_10[31]},
      {stage0_11[6], stage0_11[7], stage0_11[8], stage0_11[9], stage0_11[10], stage0_11[11]},
      {stage1_13[1],stage1_12[6],stage1_11[18],stage1_10[38],stage1_9[52]}
   );
   gpc615_5 gpc125 (
      {stage0_9[82], stage0_9[83], stage0_9[84], stage0_9[85], stage0_9[86]},
      {stage0_10[32]},
      {stage0_11[12], stage0_11[13], stage0_11[14], stage0_11[15], stage0_11[16], stage0_11[17]},
      {stage1_13[2],stage1_12[7],stage1_11[19],stage1_10[39],stage1_9[53]}
   );
   gpc615_5 gpc126 (
      {stage0_9[87], stage0_9[88], stage0_9[89], stage0_9[90], stage0_9[91]},
      {stage0_10[33]},
      {stage0_11[18], stage0_11[19], stage0_11[20], stage0_11[21], stage0_11[22], stage0_11[23]},
      {stage1_13[3],stage1_12[8],stage1_11[20],stage1_10[40],stage1_9[54]}
   );
   gpc615_5 gpc127 (
      {stage0_9[92], stage0_9[93], stage0_9[94], stage0_9[95], stage0_9[96]},
      {stage0_10[34]},
      {stage0_11[24], stage0_11[25], stage0_11[26], stage0_11[27], stage0_11[28], stage0_11[29]},
      {stage1_13[4],stage1_12[9],stage1_11[21],stage1_10[41],stage1_9[55]}
   );
   gpc615_5 gpc128 (
      {stage0_9[97], stage0_9[98], stage0_9[99], stage0_9[100], stage0_9[101]},
      {stage0_10[35]},
      {stage0_11[30], stage0_11[31], stage0_11[32], stage0_11[33], stage0_11[34], stage0_11[35]},
      {stage1_13[5],stage1_12[10],stage1_11[22],stage1_10[42],stage1_9[56]}
   );
   gpc615_5 gpc129 (
      {stage0_9[102], stage0_9[103], stage0_9[104], stage0_9[105], stage0_9[106]},
      {stage0_10[36]},
      {stage0_11[36], stage0_11[37], stage0_11[38], stage0_11[39], stage0_11[40], stage0_11[41]},
      {stage1_13[6],stage1_12[11],stage1_11[23],stage1_10[43],stage1_9[57]}
   );
   gpc615_5 gpc130 (
      {stage0_9[107], stage0_9[108], stage0_9[109], stage0_9[110], stage0_9[111]},
      {stage0_10[37]},
      {stage0_11[42], stage0_11[43], stage0_11[44], stage0_11[45], stage0_11[46], stage0_11[47]},
      {stage1_13[7],stage1_12[12],stage1_11[24],stage1_10[44],stage1_9[58]}
   );
   gpc615_5 gpc131 (
      {stage0_9[112], stage0_9[113], stage0_9[114], stage0_9[115], stage0_9[116]},
      {stage0_10[38]},
      {stage0_11[48], stage0_11[49], stage0_11[50], stage0_11[51], stage0_11[52], stage0_11[53]},
      {stage1_13[8],stage1_12[13],stage1_11[25],stage1_10[45],stage1_9[59]}
   );
   gpc615_5 gpc132 (
      {stage0_9[117], stage0_9[118], stage0_9[119], stage0_9[120], stage0_9[121]},
      {stage0_10[39]},
      {stage0_11[54], stage0_11[55], stage0_11[56], stage0_11[57], stage0_11[58], stage0_11[59]},
      {stage1_13[9],stage1_12[14],stage1_11[26],stage1_10[46],stage1_9[60]}
   );
   gpc615_5 gpc133 (
      {stage0_9[122], stage0_9[123], stage0_9[124], stage0_9[125], stage0_9[126]},
      {stage0_10[40]},
      {stage0_11[60], stage0_11[61], stage0_11[62], stage0_11[63], stage0_11[64], stage0_11[65]},
      {stage1_13[10],stage1_12[15],stage1_11[27],stage1_10[47],stage1_9[61]}
   );
   gpc615_5 gpc134 (
      {stage0_9[127], stage0_9[128], stage0_9[129], stage0_9[130], stage0_9[131]},
      {stage0_10[41]},
      {stage0_11[66], stage0_11[67], stage0_11[68], stage0_11[69], stage0_11[70], stage0_11[71]},
      {stage1_13[11],stage1_12[16],stage1_11[28],stage1_10[48],stage1_9[62]}
   );
   gpc615_5 gpc135 (
      {stage0_9[132], stage0_9[133], stage0_9[134], stage0_9[135], stage0_9[136]},
      {stage0_10[42]},
      {stage0_11[72], stage0_11[73], stage0_11[74], stage0_11[75], stage0_11[76], stage0_11[77]},
      {stage1_13[12],stage1_12[17],stage1_11[29],stage1_10[49],stage1_9[63]}
   );
   gpc615_5 gpc136 (
      {stage0_9[137], stage0_9[138], stage0_9[139], stage0_9[140], stage0_9[141]},
      {stage0_10[43]},
      {stage0_11[78], stage0_11[79], stage0_11[80], stage0_11[81], stage0_11[82], stage0_11[83]},
      {stage1_13[13],stage1_12[18],stage1_11[30],stage1_10[50],stage1_9[64]}
   );
   gpc615_5 gpc137 (
      {stage0_9[142], stage0_9[143], stage0_9[144], stage0_9[145], stage0_9[146]},
      {stage0_10[44]},
      {stage0_11[84], stage0_11[85], stage0_11[86], stage0_11[87], stage0_11[88], stage0_11[89]},
      {stage1_13[14],stage1_12[19],stage1_11[31],stage1_10[51],stage1_9[65]}
   );
   gpc615_5 gpc138 (
      {stage0_9[147], stage0_9[148], stage0_9[149], stage0_9[150], stage0_9[151]},
      {stage0_10[45]},
      {stage0_11[90], stage0_11[91], stage0_11[92], stage0_11[93], stage0_11[94], stage0_11[95]},
      {stage1_13[15],stage1_12[20],stage1_11[32],stage1_10[52],stage1_9[66]}
   );
   gpc615_5 gpc139 (
      {stage0_10[46], stage0_10[47], stage0_10[48], stage0_10[49], stage0_10[50]},
      {stage0_11[96]},
      {stage0_12[0], stage0_12[1], stage0_12[2], stage0_12[3], stage0_12[4], stage0_12[5]},
      {stage1_14[0],stage1_13[16],stage1_12[21],stage1_11[33],stage1_10[53]}
   );
   gpc615_5 gpc140 (
      {stage0_10[51], stage0_10[52], stage0_10[53], stage0_10[54], stage0_10[55]},
      {stage0_11[97]},
      {stage0_12[6], stage0_12[7], stage0_12[8], stage0_12[9], stage0_12[10], stage0_12[11]},
      {stage1_14[1],stage1_13[17],stage1_12[22],stage1_11[34],stage1_10[54]}
   );
   gpc615_5 gpc141 (
      {stage0_10[56], stage0_10[57], stage0_10[58], stage0_10[59], stage0_10[60]},
      {stage0_11[98]},
      {stage0_12[12], stage0_12[13], stage0_12[14], stage0_12[15], stage0_12[16], stage0_12[17]},
      {stage1_14[2],stage1_13[18],stage1_12[23],stage1_11[35],stage1_10[55]}
   );
   gpc615_5 gpc142 (
      {stage0_10[61], stage0_10[62], stage0_10[63], stage0_10[64], stage0_10[65]},
      {stage0_11[99]},
      {stage0_12[18], stage0_12[19], stage0_12[20], stage0_12[21], stage0_12[22], stage0_12[23]},
      {stage1_14[3],stage1_13[19],stage1_12[24],stage1_11[36],stage1_10[56]}
   );
   gpc615_5 gpc143 (
      {stage0_10[66], stage0_10[67], stage0_10[68], stage0_10[69], stage0_10[70]},
      {stage0_11[100]},
      {stage0_12[24], stage0_12[25], stage0_12[26], stage0_12[27], stage0_12[28], stage0_12[29]},
      {stage1_14[4],stage1_13[20],stage1_12[25],stage1_11[37],stage1_10[57]}
   );
   gpc615_5 gpc144 (
      {stage0_10[71], stage0_10[72], stage0_10[73], stage0_10[74], stage0_10[75]},
      {stage0_11[101]},
      {stage0_12[30], stage0_12[31], stage0_12[32], stage0_12[33], stage0_12[34], stage0_12[35]},
      {stage1_14[5],stage1_13[21],stage1_12[26],stage1_11[38],stage1_10[58]}
   );
   gpc615_5 gpc145 (
      {stage0_10[76], stage0_10[77], stage0_10[78], stage0_10[79], stage0_10[80]},
      {stage0_11[102]},
      {stage0_12[36], stage0_12[37], stage0_12[38], stage0_12[39], stage0_12[40], stage0_12[41]},
      {stage1_14[6],stage1_13[22],stage1_12[27],stage1_11[39],stage1_10[59]}
   );
   gpc615_5 gpc146 (
      {stage0_10[81], stage0_10[82], stage0_10[83], stage0_10[84], stage0_10[85]},
      {stage0_11[103]},
      {stage0_12[42], stage0_12[43], stage0_12[44], stage0_12[45], stage0_12[46], stage0_12[47]},
      {stage1_14[7],stage1_13[23],stage1_12[28],stage1_11[40],stage1_10[60]}
   );
   gpc615_5 gpc147 (
      {stage0_10[86], stage0_10[87], stage0_10[88], stage0_10[89], stage0_10[90]},
      {stage0_11[104]},
      {stage0_12[48], stage0_12[49], stage0_12[50], stage0_12[51], stage0_12[52], stage0_12[53]},
      {stage1_14[8],stage1_13[24],stage1_12[29],stage1_11[41],stage1_10[61]}
   );
   gpc615_5 gpc148 (
      {stage0_10[91], stage0_10[92], stage0_10[93], stage0_10[94], stage0_10[95]},
      {stage0_11[105]},
      {stage0_12[54], stage0_12[55], stage0_12[56], stage0_12[57], stage0_12[58], stage0_12[59]},
      {stage1_14[9],stage1_13[25],stage1_12[30],stage1_11[42],stage1_10[62]}
   );
   gpc615_5 gpc149 (
      {stage0_10[96], stage0_10[97], stage0_10[98], stage0_10[99], stage0_10[100]},
      {stage0_11[106]},
      {stage0_12[60], stage0_12[61], stage0_12[62], stage0_12[63], stage0_12[64], stage0_12[65]},
      {stage1_14[10],stage1_13[26],stage1_12[31],stage1_11[43],stage1_10[63]}
   );
   gpc615_5 gpc150 (
      {stage0_10[101], stage0_10[102], stage0_10[103], stage0_10[104], stage0_10[105]},
      {stage0_11[107]},
      {stage0_12[66], stage0_12[67], stage0_12[68], stage0_12[69], stage0_12[70], stage0_12[71]},
      {stage1_14[11],stage1_13[27],stage1_12[32],stage1_11[44],stage1_10[64]}
   );
   gpc615_5 gpc151 (
      {stage0_10[106], stage0_10[107], stage0_10[108], stage0_10[109], stage0_10[110]},
      {stage0_11[108]},
      {stage0_12[72], stage0_12[73], stage0_12[74], stage0_12[75], stage0_12[76], stage0_12[77]},
      {stage1_14[12],stage1_13[28],stage1_12[33],stage1_11[45],stage1_10[65]}
   );
   gpc615_5 gpc152 (
      {stage0_10[111], stage0_10[112], stage0_10[113], stage0_10[114], stage0_10[115]},
      {stage0_11[109]},
      {stage0_12[78], stage0_12[79], stage0_12[80], stage0_12[81], stage0_12[82], stage0_12[83]},
      {stage1_14[13],stage1_13[29],stage1_12[34],stage1_11[46],stage1_10[66]}
   );
   gpc615_5 gpc153 (
      {stage0_10[116], stage0_10[117], stage0_10[118], stage0_10[119], stage0_10[120]},
      {stage0_11[110]},
      {stage0_12[84], stage0_12[85], stage0_12[86], stage0_12[87], stage0_12[88], stage0_12[89]},
      {stage1_14[14],stage1_13[30],stage1_12[35],stage1_11[47],stage1_10[67]}
   );
   gpc615_5 gpc154 (
      {stage0_10[121], stage0_10[122], stage0_10[123], stage0_10[124], stage0_10[125]},
      {stage0_11[111]},
      {stage0_12[90], stage0_12[91], stage0_12[92], stage0_12[93], stage0_12[94], stage0_12[95]},
      {stage1_14[15],stage1_13[31],stage1_12[36],stage1_11[48],stage1_10[68]}
   );
   gpc615_5 gpc155 (
      {stage0_10[126], stage0_10[127], stage0_10[128], stage0_10[129], stage0_10[130]},
      {stage0_11[112]},
      {stage0_12[96], stage0_12[97], stage0_12[98], stage0_12[99], stage0_12[100], stage0_12[101]},
      {stage1_14[16],stage1_13[32],stage1_12[37],stage1_11[49],stage1_10[69]}
   );
   gpc615_5 gpc156 (
      {stage0_10[131], stage0_10[132], stage0_10[133], stage0_10[134], stage0_10[135]},
      {stage0_11[113]},
      {stage0_12[102], stage0_12[103], stage0_12[104], stage0_12[105], stage0_12[106], stage0_12[107]},
      {stage1_14[17],stage1_13[33],stage1_12[38],stage1_11[50],stage1_10[70]}
   );
   gpc615_5 gpc157 (
      {stage0_10[136], stage0_10[137], stage0_10[138], stage0_10[139], stage0_10[140]},
      {stage0_11[114]},
      {stage0_12[108], stage0_12[109], stage0_12[110], stage0_12[111], stage0_12[112], stage0_12[113]},
      {stage1_14[18],stage1_13[34],stage1_12[39],stage1_11[51],stage1_10[71]}
   );
   gpc615_5 gpc158 (
      {stage0_11[115], stage0_11[116], stage0_11[117], stage0_11[118], stage0_11[119]},
      {stage0_12[114]},
      {stage0_13[0], stage0_13[1], stage0_13[2], stage0_13[3], stage0_13[4], stage0_13[5]},
      {stage1_15[0],stage1_14[19],stage1_13[35],stage1_12[40],stage1_11[52]}
   );
   gpc615_5 gpc159 (
      {stage0_11[120], stage0_11[121], stage0_11[122], stage0_11[123], stage0_11[124]},
      {stage0_12[115]},
      {stage0_13[6], stage0_13[7], stage0_13[8], stage0_13[9], stage0_13[10], stage0_13[11]},
      {stage1_15[1],stage1_14[20],stage1_13[36],stage1_12[41],stage1_11[53]}
   );
   gpc615_5 gpc160 (
      {stage0_11[125], stage0_11[126], stage0_11[127], stage0_11[128], stage0_11[129]},
      {stage0_12[116]},
      {stage0_13[12], stage0_13[13], stage0_13[14], stage0_13[15], stage0_13[16], stage0_13[17]},
      {stage1_15[2],stage1_14[21],stage1_13[37],stage1_12[42],stage1_11[54]}
   );
   gpc615_5 gpc161 (
      {stage0_11[130], stage0_11[131], stage0_11[132], stage0_11[133], stage0_11[134]},
      {stage0_12[117]},
      {stage0_13[18], stage0_13[19], stage0_13[20], stage0_13[21], stage0_13[22], stage0_13[23]},
      {stage1_15[3],stage1_14[22],stage1_13[38],stage1_12[43],stage1_11[55]}
   );
   gpc615_5 gpc162 (
      {stage0_11[135], stage0_11[136], stage0_11[137], stage0_11[138], stage0_11[139]},
      {stage0_12[118]},
      {stage0_13[24], stage0_13[25], stage0_13[26], stage0_13[27], stage0_13[28], stage0_13[29]},
      {stage1_15[4],stage1_14[23],stage1_13[39],stage1_12[44],stage1_11[56]}
   );
   gpc615_5 gpc163 (
      {stage0_11[140], stage0_11[141], stage0_11[142], stage0_11[143], stage0_11[144]},
      {stage0_12[119]},
      {stage0_13[30], stage0_13[31], stage0_13[32], stage0_13[33], stage0_13[34], stage0_13[35]},
      {stage1_15[5],stage1_14[24],stage1_13[40],stage1_12[45],stage1_11[57]}
   );
   gpc615_5 gpc164 (
      {stage0_11[145], stage0_11[146], stage0_11[147], stage0_11[148], stage0_11[149]},
      {stage0_12[120]},
      {stage0_13[36], stage0_13[37], stage0_13[38], stage0_13[39], stage0_13[40], stage0_13[41]},
      {stage1_15[6],stage1_14[25],stage1_13[41],stage1_12[46],stage1_11[58]}
   );
   gpc615_5 gpc165 (
      {stage0_11[150], stage0_11[151], stage0_11[152], stage0_11[153], stage0_11[154]},
      {stage0_12[121]},
      {stage0_13[42], stage0_13[43], stage0_13[44], stage0_13[45], stage0_13[46], stage0_13[47]},
      {stage1_15[7],stage1_14[26],stage1_13[42],stage1_12[47],stage1_11[59]}
   );
   gpc615_5 gpc166 (
      {stage0_12[122], stage0_12[123], stage0_12[124], stage0_12[125], stage0_12[126]},
      {stage0_13[48]},
      {stage0_14[0], stage0_14[1], stage0_14[2], stage0_14[3], stage0_14[4], stage0_14[5]},
      {stage1_16[0],stage1_15[8],stage1_14[27],stage1_13[43],stage1_12[48]}
   );
   gpc615_5 gpc167 (
      {stage0_12[127], stage0_12[128], stage0_12[129], stage0_12[130], stage0_12[131]},
      {stage0_13[49]},
      {stage0_14[6], stage0_14[7], stage0_14[8], stage0_14[9], stage0_14[10], stage0_14[11]},
      {stage1_16[1],stage1_15[9],stage1_14[28],stage1_13[44],stage1_12[49]}
   );
   gpc615_5 gpc168 (
      {stage0_12[132], stage0_12[133], stage0_12[134], stage0_12[135], stage0_12[136]},
      {stage0_13[50]},
      {stage0_14[12], stage0_14[13], stage0_14[14], stage0_14[15], stage0_14[16], stage0_14[17]},
      {stage1_16[2],stage1_15[10],stage1_14[29],stage1_13[45],stage1_12[50]}
   );
   gpc615_5 gpc169 (
      {stage0_12[137], stage0_12[138], stage0_12[139], stage0_12[140], stage0_12[141]},
      {stage0_13[51]},
      {stage0_14[18], stage0_14[19], stage0_14[20], stage0_14[21], stage0_14[22], stage0_14[23]},
      {stage1_16[3],stage1_15[11],stage1_14[30],stage1_13[46],stage1_12[51]}
   );
   gpc615_5 gpc170 (
      {stage0_12[142], stage0_12[143], stage0_12[144], stage0_12[145], stage0_12[146]},
      {stage0_13[52]},
      {stage0_14[24], stage0_14[25], stage0_14[26], stage0_14[27], stage0_14[28], stage0_14[29]},
      {stage1_16[4],stage1_15[12],stage1_14[31],stage1_13[47],stage1_12[52]}
   );
   gpc615_5 gpc171 (
      {stage0_12[147], stage0_12[148], stage0_12[149], stage0_12[150], stage0_12[151]},
      {stage0_13[53]},
      {stage0_14[30], stage0_14[31], stage0_14[32], stage0_14[33], stage0_14[34], stage0_14[35]},
      {stage1_16[5],stage1_15[13],stage1_14[32],stage1_13[48],stage1_12[53]}
   );
   gpc615_5 gpc172 (
      {stage0_12[152], stage0_12[153], stage0_12[154], stage0_12[155], stage0_12[156]},
      {stage0_13[54]},
      {stage0_14[36], stage0_14[37], stage0_14[38], stage0_14[39], stage0_14[40], stage0_14[41]},
      {stage1_16[6],stage1_15[14],stage1_14[33],stage1_13[49],stage1_12[54]}
   );
   gpc615_5 gpc173 (
      {stage0_12[157], stage0_12[158], stage0_12[159], stage0_12[160], stage0_12[161]},
      {stage0_13[55]},
      {stage0_14[42], stage0_14[43], stage0_14[44], stage0_14[45], stage0_14[46], stage0_14[47]},
      {stage1_16[7],stage1_15[15],stage1_14[34],stage1_13[50],stage1_12[55]}
   );
   gpc606_5 gpc174 (
      {stage0_13[56], stage0_13[57], stage0_13[58], stage0_13[59], stage0_13[60], stage0_13[61]},
      {stage0_15[0], stage0_15[1], stage0_15[2], stage0_15[3], stage0_15[4], stage0_15[5]},
      {stage1_17[0],stage1_16[8],stage1_15[16],stage1_14[35],stage1_13[51]}
   );
   gpc606_5 gpc175 (
      {stage0_13[62], stage0_13[63], stage0_13[64], stage0_13[65], stage0_13[66], stage0_13[67]},
      {stage0_15[6], stage0_15[7], stage0_15[8], stage0_15[9], stage0_15[10], stage0_15[11]},
      {stage1_17[1],stage1_16[9],stage1_15[17],stage1_14[36],stage1_13[52]}
   );
   gpc606_5 gpc176 (
      {stage0_13[68], stage0_13[69], stage0_13[70], stage0_13[71], stage0_13[72], stage0_13[73]},
      {stage0_15[12], stage0_15[13], stage0_15[14], stage0_15[15], stage0_15[16], stage0_15[17]},
      {stage1_17[2],stage1_16[10],stage1_15[18],stage1_14[37],stage1_13[53]}
   );
   gpc615_5 gpc177 (
      {stage0_13[74], stage0_13[75], stage0_13[76], stage0_13[77], stage0_13[78]},
      {stage0_14[48]},
      {stage0_15[18], stage0_15[19], stage0_15[20], stage0_15[21], stage0_15[22], stage0_15[23]},
      {stage1_17[3],stage1_16[11],stage1_15[19],stage1_14[38],stage1_13[54]}
   );
   gpc615_5 gpc178 (
      {stage0_13[79], stage0_13[80], stage0_13[81], stage0_13[82], stage0_13[83]},
      {stage0_14[49]},
      {stage0_15[24], stage0_15[25], stage0_15[26], stage0_15[27], stage0_15[28], stage0_15[29]},
      {stage1_17[4],stage1_16[12],stage1_15[20],stage1_14[39],stage1_13[55]}
   );
   gpc615_5 gpc179 (
      {stage0_13[84], stage0_13[85], stage0_13[86], stage0_13[87], stage0_13[88]},
      {stage0_14[50]},
      {stage0_15[30], stage0_15[31], stage0_15[32], stage0_15[33], stage0_15[34], stage0_15[35]},
      {stage1_17[5],stage1_16[13],stage1_15[21],stage1_14[40],stage1_13[56]}
   );
   gpc615_5 gpc180 (
      {stage0_13[89], stage0_13[90], stage0_13[91], stage0_13[92], stage0_13[93]},
      {stage0_14[51]},
      {stage0_15[36], stage0_15[37], stage0_15[38], stage0_15[39], stage0_15[40], stage0_15[41]},
      {stage1_17[6],stage1_16[14],stage1_15[22],stage1_14[41],stage1_13[57]}
   );
   gpc615_5 gpc181 (
      {stage0_13[94], stage0_13[95], stage0_13[96], stage0_13[97], stage0_13[98]},
      {stage0_14[52]},
      {stage0_15[42], stage0_15[43], stage0_15[44], stage0_15[45], stage0_15[46], stage0_15[47]},
      {stage1_17[7],stage1_16[15],stage1_15[23],stage1_14[42],stage1_13[58]}
   );
   gpc615_5 gpc182 (
      {stage0_13[99], stage0_13[100], stage0_13[101], stage0_13[102], stage0_13[103]},
      {stage0_14[53]},
      {stage0_15[48], stage0_15[49], stage0_15[50], stage0_15[51], stage0_15[52], stage0_15[53]},
      {stage1_17[8],stage1_16[16],stage1_15[24],stage1_14[43],stage1_13[59]}
   );
   gpc615_5 gpc183 (
      {stage0_13[104], stage0_13[105], stage0_13[106], stage0_13[107], stage0_13[108]},
      {stage0_14[54]},
      {stage0_15[54], stage0_15[55], stage0_15[56], stage0_15[57], stage0_15[58], stage0_15[59]},
      {stage1_17[9],stage1_16[17],stage1_15[25],stage1_14[44],stage1_13[60]}
   );
   gpc615_5 gpc184 (
      {stage0_13[109], stage0_13[110], stage0_13[111], stage0_13[112], stage0_13[113]},
      {stage0_14[55]},
      {stage0_15[60], stage0_15[61], stage0_15[62], stage0_15[63], stage0_15[64], stage0_15[65]},
      {stage1_17[10],stage1_16[18],stage1_15[26],stage1_14[45],stage1_13[61]}
   );
   gpc615_5 gpc185 (
      {stage0_13[114], stage0_13[115], stage0_13[116], stage0_13[117], stage0_13[118]},
      {stage0_14[56]},
      {stage0_15[66], stage0_15[67], stage0_15[68], stage0_15[69], stage0_15[70], stage0_15[71]},
      {stage1_17[11],stage1_16[19],stage1_15[27],stage1_14[46],stage1_13[62]}
   );
   gpc615_5 gpc186 (
      {stage0_13[119], stage0_13[120], stage0_13[121], stage0_13[122], stage0_13[123]},
      {stage0_14[57]},
      {stage0_15[72], stage0_15[73], stage0_15[74], stage0_15[75], stage0_15[76], stage0_15[77]},
      {stage1_17[12],stage1_16[20],stage1_15[28],stage1_14[47],stage1_13[63]}
   );
   gpc615_5 gpc187 (
      {stage0_13[124], stage0_13[125], stage0_13[126], stage0_13[127], stage0_13[128]},
      {stage0_14[58]},
      {stage0_15[78], stage0_15[79], stage0_15[80], stage0_15[81], stage0_15[82], stage0_15[83]},
      {stage1_17[13],stage1_16[21],stage1_15[29],stage1_14[48],stage1_13[64]}
   );
   gpc615_5 gpc188 (
      {stage0_13[129], stage0_13[130], stage0_13[131], stage0_13[132], stage0_13[133]},
      {stage0_14[59]},
      {stage0_15[84], stage0_15[85], stage0_15[86], stage0_15[87], stage0_15[88], stage0_15[89]},
      {stage1_17[14],stage1_16[22],stage1_15[30],stage1_14[49],stage1_13[65]}
   );
   gpc615_5 gpc189 (
      {stage0_13[134], stage0_13[135], stage0_13[136], stage0_13[137], stage0_13[138]},
      {stage0_14[60]},
      {stage0_15[90], stage0_15[91], stage0_15[92], stage0_15[93], stage0_15[94], stage0_15[95]},
      {stage1_17[15],stage1_16[23],stage1_15[31],stage1_14[50],stage1_13[66]}
   );
   gpc615_5 gpc190 (
      {stage0_13[139], stage0_13[140], stage0_13[141], stage0_13[142], stage0_13[143]},
      {stage0_14[61]},
      {stage0_15[96], stage0_15[97], stage0_15[98], stage0_15[99], stage0_15[100], stage0_15[101]},
      {stage1_17[16],stage1_16[24],stage1_15[32],stage1_14[51],stage1_13[67]}
   );
   gpc117_4 gpc191 (
      {stage0_14[62], stage0_14[63], stage0_14[64], stage0_14[65], stage0_14[66], stage0_14[67], stage0_14[68]},
      {stage0_15[102]},
      {stage0_16[0]},
      {stage1_17[17],stage1_16[25],stage1_15[33],stage1_14[52]}
   );
   gpc117_4 gpc192 (
      {stage0_14[69], stage0_14[70], stage0_14[71], stage0_14[72], stage0_14[73], stage0_14[74], stage0_14[75]},
      {stage0_15[103]},
      {stage0_16[1]},
      {stage1_17[18],stage1_16[26],stage1_15[34],stage1_14[53]}
   );
   gpc117_4 gpc193 (
      {stage0_14[76], stage0_14[77], stage0_14[78], stage0_14[79], stage0_14[80], stage0_14[81], stage0_14[82]},
      {stage0_15[104]},
      {stage0_16[2]},
      {stage1_17[19],stage1_16[27],stage1_15[35],stage1_14[54]}
   );
   gpc117_4 gpc194 (
      {stage0_14[83], stage0_14[84], stage0_14[85], stage0_14[86], stage0_14[87], stage0_14[88], stage0_14[89]},
      {stage0_15[105]},
      {stage0_16[3]},
      {stage1_17[20],stage1_16[28],stage1_15[36],stage1_14[55]}
   );
   gpc606_5 gpc195 (
      {stage0_14[90], stage0_14[91], stage0_14[92], stage0_14[93], stage0_14[94], stage0_14[95]},
      {stage0_16[4], stage0_16[5], stage0_16[6], stage0_16[7], stage0_16[8], stage0_16[9]},
      {stage1_18[0],stage1_17[21],stage1_16[29],stage1_15[37],stage1_14[56]}
   );
   gpc606_5 gpc196 (
      {stage0_14[96], stage0_14[97], stage0_14[98], stage0_14[99], stage0_14[100], stage0_14[101]},
      {stage0_16[10], stage0_16[11], stage0_16[12], stage0_16[13], stage0_16[14], stage0_16[15]},
      {stage1_18[1],stage1_17[22],stage1_16[30],stage1_15[38],stage1_14[57]}
   );
   gpc606_5 gpc197 (
      {stage0_14[102], stage0_14[103], stage0_14[104], stage0_14[105], stage0_14[106], stage0_14[107]},
      {stage0_16[16], stage0_16[17], stage0_16[18], stage0_16[19], stage0_16[20], stage0_16[21]},
      {stage1_18[2],stage1_17[23],stage1_16[31],stage1_15[39],stage1_14[58]}
   );
   gpc606_5 gpc198 (
      {stage0_14[108], stage0_14[109], stage0_14[110], stage0_14[111], stage0_14[112], stage0_14[113]},
      {stage0_16[22], stage0_16[23], stage0_16[24], stage0_16[25], stage0_16[26], stage0_16[27]},
      {stage1_18[3],stage1_17[24],stage1_16[32],stage1_15[40],stage1_14[59]}
   );
   gpc606_5 gpc199 (
      {stage0_14[114], stage0_14[115], stage0_14[116], stage0_14[117], stage0_14[118], stage0_14[119]},
      {stage0_16[28], stage0_16[29], stage0_16[30], stage0_16[31], stage0_16[32], stage0_16[33]},
      {stage1_18[4],stage1_17[25],stage1_16[33],stage1_15[41],stage1_14[60]}
   );
   gpc606_5 gpc200 (
      {stage0_14[120], stage0_14[121], stage0_14[122], stage0_14[123], stage0_14[124], stage0_14[125]},
      {stage0_16[34], stage0_16[35], stage0_16[36], stage0_16[37], stage0_16[38], stage0_16[39]},
      {stage1_18[5],stage1_17[26],stage1_16[34],stage1_15[42],stage1_14[61]}
   );
   gpc606_5 gpc201 (
      {stage0_14[126], stage0_14[127], stage0_14[128], stage0_14[129], stage0_14[130], stage0_14[131]},
      {stage0_16[40], stage0_16[41], stage0_16[42], stage0_16[43], stage0_16[44], stage0_16[45]},
      {stage1_18[6],stage1_17[27],stage1_16[35],stage1_15[43],stage1_14[62]}
   );
   gpc606_5 gpc202 (
      {stage0_14[132], stage0_14[133], stage0_14[134], stage0_14[135], stage0_14[136], stage0_14[137]},
      {stage0_16[46], stage0_16[47], stage0_16[48], stage0_16[49], stage0_16[50], stage0_16[51]},
      {stage1_18[7],stage1_17[28],stage1_16[36],stage1_15[44],stage1_14[63]}
   );
   gpc606_5 gpc203 (
      {stage0_14[138], stage0_14[139], stage0_14[140], stage0_14[141], stage0_14[142], stage0_14[143]},
      {stage0_16[52], stage0_16[53], stage0_16[54], stage0_16[55], stage0_16[56], stage0_16[57]},
      {stage1_18[8],stage1_17[29],stage1_16[37],stage1_15[45],stage1_14[64]}
   );
   gpc606_5 gpc204 (
      {stage0_14[144], stage0_14[145], stage0_14[146], stage0_14[147], stage0_14[148], stage0_14[149]},
      {stage0_16[58], stage0_16[59], stage0_16[60], stage0_16[61], stage0_16[62], stage0_16[63]},
      {stage1_18[9],stage1_17[30],stage1_16[38],stage1_15[46],stage1_14[65]}
   );
   gpc606_5 gpc205 (
      {stage0_14[150], stage0_14[151], stage0_14[152], stage0_14[153], stage0_14[154], stage0_14[155]},
      {stage0_16[64], stage0_16[65], stage0_16[66], stage0_16[67], stage0_16[68], stage0_16[69]},
      {stage1_18[10],stage1_17[31],stage1_16[39],stage1_15[47],stage1_14[66]}
   );
   gpc615_5 gpc206 (
      {stage0_14[156], stage0_14[157], stage0_14[158], stage0_14[159], stage0_14[160]},
      {stage0_15[106]},
      {stage0_16[70], stage0_16[71], stage0_16[72], stage0_16[73], stage0_16[74], stage0_16[75]},
      {stage1_18[11],stage1_17[32],stage1_16[40],stage1_15[48],stage1_14[67]}
   );
   gpc615_5 gpc207 (
      {stage0_15[107], stage0_15[108], stage0_15[109], stage0_15[110], stage0_15[111]},
      {stage0_16[76]},
      {stage0_17[0], stage0_17[1], stage0_17[2], stage0_17[3], stage0_17[4], stage0_17[5]},
      {stage1_19[0],stage1_18[12],stage1_17[33],stage1_16[41],stage1_15[49]}
   );
   gpc615_5 gpc208 (
      {stage0_15[112], stage0_15[113], stage0_15[114], stage0_15[115], stage0_15[116]},
      {stage0_16[77]},
      {stage0_17[6], stage0_17[7], stage0_17[8], stage0_17[9], stage0_17[10], stage0_17[11]},
      {stage1_19[1],stage1_18[13],stage1_17[34],stage1_16[42],stage1_15[50]}
   );
   gpc615_5 gpc209 (
      {stage0_15[117], stage0_15[118], stage0_15[119], stage0_15[120], stage0_15[121]},
      {stage0_16[78]},
      {stage0_17[12], stage0_17[13], stage0_17[14], stage0_17[15], stage0_17[16], stage0_17[17]},
      {stage1_19[2],stage1_18[14],stage1_17[35],stage1_16[43],stage1_15[51]}
   );
   gpc615_5 gpc210 (
      {stage0_15[122], stage0_15[123], stage0_15[124], stage0_15[125], stage0_15[126]},
      {stage0_16[79]},
      {stage0_17[18], stage0_17[19], stage0_17[20], stage0_17[21], stage0_17[22], stage0_17[23]},
      {stage1_19[3],stage1_18[15],stage1_17[36],stage1_16[44],stage1_15[52]}
   );
   gpc615_5 gpc211 (
      {stage0_15[127], stage0_15[128], stage0_15[129], stage0_15[130], stage0_15[131]},
      {stage0_16[80]},
      {stage0_17[24], stage0_17[25], stage0_17[26], stage0_17[27], stage0_17[28], stage0_17[29]},
      {stage1_19[4],stage1_18[16],stage1_17[37],stage1_16[45],stage1_15[53]}
   );
   gpc615_5 gpc212 (
      {stage0_15[132], stage0_15[133], stage0_15[134], stage0_15[135], stage0_15[136]},
      {stage0_16[81]},
      {stage0_17[30], stage0_17[31], stage0_17[32], stage0_17[33], stage0_17[34], stage0_17[35]},
      {stage1_19[5],stage1_18[17],stage1_17[38],stage1_16[46],stage1_15[54]}
   );
   gpc615_5 gpc213 (
      {stage0_15[137], stage0_15[138], stage0_15[139], stage0_15[140], stage0_15[141]},
      {stage0_16[82]},
      {stage0_17[36], stage0_17[37], stage0_17[38], stage0_17[39], stage0_17[40], stage0_17[41]},
      {stage1_19[6],stage1_18[18],stage1_17[39],stage1_16[47],stage1_15[55]}
   );
   gpc615_5 gpc214 (
      {stage0_15[142], stage0_15[143], stage0_15[144], stage0_15[145], stage0_15[146]},
      {stage0_16[83]},
      {stage0_17[42], stage0_17[43], stage0_17[44], stage0_17[45], stage0_17[46], stage0_17[47]},
      {stage1_19[7],stage1_18[19],stage1_17[40],stage1_16[48],stage1_15[56]}
   );
   gpc615_5 gpc215 (
      {stage0_15[147], stage0_15[148], stage0_15[149], stage0_15[150], stage0_15[151]},
      {stage0_16[84]},
      {stage0_17[48], stage0_17[49], stage0_17[50], stage0_17[51], stage0_17[52], stage0_17[53]},
      {stage1_19[8],stage1_18[20],stage1_17[41],stage1_16[49],stage1_15[57]}
   );
   gpc615_5 gpc216 (
      {stage0_15[152], stage0_15[153], stage0_15[154], stage0_15[155], stage0_15[156]},
      {stage0_16[85]},
      {stage0_17[54], stage0_17[55], stage0_17[56], stage0_17[57], stage0_17[58], stage0_17[59]},
      {stage1_19[9],stage1_18[21],stage1_17[42],stage1_16[50],stage1_15[58]}
   );
   gpc615_5 gpc217 (
      {stage0_15[157], stage0_15[158], stage0_15[159], stage0_15[160], stage0_15[161]},
      {stage0_16[86]},
      {stage0_17[60], stage0_17[61], stage0_17[62], stage0_17[63], stage0_17[64], stage0_17[65]},
      {stage1_19[10],stage1_18[22],stage1_17[43],stage1_16[51],stage1_15[59]}
   );
   gpc606_5 gpc218 (
      {stage0_16[87], stage0_16[88], stage0_16[89], stage0_16[90], stage0_16[91], stage0_16[92]},
      {stage0_18[0], stage0_18[1], stage0_18[2], stage0_18[3], stage0_18[4], stage0_18[5]},
      {stage1_20[0],stage1_19[11],stage1_18[23],stage1_17[44],stage1_16[52]}
   );
   gpc606_5 gpc219 (
      {stage0_16[93], stage0_16[94], stage0_16[95], stage0_16[96], stage0_16[97], stage0_16[98]},
      {stage0_18[6], stage0_18[7], stage0_18[8], stage0_18[9], stage0_18[10], stage0_18[11]},
      {stage1_20[1],stage1_19[12],stage1_18[24],stage1_17[45],stage1_16[53]}
   );
   gpc606_5 gpc220 (
      {stage0_16[99], stage0_16[100], stage0_16[101], stage0_16[102], stage0_16[103], stage0_16[104]},
      {stage0_18[12], stage0_18[13], stage0_18[14], stage0_18[15], stage0_18[16], stage0_18[17]},
      {stage1_20[2],stage1_19[13],stage1_18[25],stage1_17[46],stage1_16[54]}
   );
   gpc606_5 gpc221 (
      {stage0_16[105], stage0_16[106], stage0_16[107], stage0_16[108], stage0_16[109], stage0_16[110]},
      {stage0_18[18], stage0_18[19], stage0_18[20], stage0_18[21], stage0_18[22], stage0_18[23]},
      {stage1_20[3],stage1_19[14],stage1_18[26],stage1_17[47],stage1_16[55]}
   );
   gpc606_5 gpc222 (
      {stage0_17[66], stage0_17[67], stage0_17[68], stage0_17[69], stage0_17[70], stage0_17[71]},
      {stage0_19[0], stage0_19[1], stage0_19[2], stage0_19[3], stage0_19[4], stage0_19[5]},
      {stage1_21[0],stage1_20[4],stage1_19[15],stage1_18[27],stage1_17[48]}
   );
   gpc606_5 gpc223 (
      {stage0_17[72], stage0_17[73], stage0_17[74], stage0_17[75], stage0_17[76], stage0_17[77]},
      {stage0_19[6], stage0_19[7], stage0_19[8], stage0_19[9], stage0_19[10], stage0_19[11]},
      {stage1_21[1],stage1_20[5],stage1_19[16],stage1_18[28],stage1_17[49]}
   );
   gpc606_5 gpc224 (
      {stage0_17[78], stage0_17[79], stage0_17[80], stage0_17[81], stage0_17[82], stage0_17[83]},
      {stage0_19[12], stage0_19[13], stage0_19[14], stage0_19[15], stage0_19[16], stage0_19[17]},
      {stage1_21[2],stage1_20[6],stage1_19[17],stage1_18[29],stage1_17[50]}
   );
   gpc606_5 gpc225 (
      {stage0_17[84], stage0_17[85], stage0_17[86], stage0_17[87], stage0_17[88], stage0_17[89]},
      {stage0_19[18], stage0_19[19], stage0_19[20], stage0_19[21], stage0_19[22], stage0_19[23]},
      {stage1_21[3],stage1_20[7],stage1_19[18],stage1_18[30],stage1_17[51]}
   );
   gpc606_5 gpc226 (
      {stage0_17[90], stage0_17[91], stage0_17[92], stage0_17[93], stage0_17[94], stage0_17[95]},
      {stage0_19[24], stage0_19[25], stage0_19[26], stage0_19[27], stage0_19[28], stage0_19[29]},
      {stage1_21[4],stage1_20[8],stage1_19[19],stage1_18[31],stage1_17[52]}
   );
   gpc606_5 gpc227 (
      {stage0_17[96], stage0_17[97], stage0_17[98], stage0_17[99], stage0_17[100], stage0_17[101]},
      {stage0_19[30], stage0_19[31], stage0_19[32], stage0_19[33], stage0_19[34], stage0_19[35]},
      {stage1_21[5],stage1_20[9],stage1_19[20],stage1_18[32],stage1_17[53]}
   );
   gpc606_5 gpc228 (
      {stage0_17[102], stage0_17[103], stage0_17[104], stage0_17[105], stage0_17[106], stage0_17[107]},
      {stage0_19[36], stage0_19[37], stage0_19[38], stage0_19[39], stage0_19[40], stage0_19[41]},
      {stage1_21[6],stage1_20[10],stage1_19[21],stage1_18[33],stage1_17[54]}
   );
   gpc606_5 gpc229 (
      {stage0_17[108], stage0_17[109], stage0_17[110], stage0_17[111], stage0_17[112], stage0_17[113]},
      {stage0_19[42], stage0_19[43], stage0_19[44], stage0_19[45], stage0_19[46], stage0_19[47]},
      {stage1_21[7],stage1_20[11],stage1_19[22],stage1_18[34],stage1_17[55]}
   );
   gpc606_5 gpc230 (
      {stage0_17[114], stage0_17[115], stage0_17[116], stage0_17[117], stage0_17[118], stage0_17[119]},
      {stage0_19[48], stage0_19[49], stage0_19[50], stage0_19[51], stage0_19[52], stage0_19[53]},
      {stage1_21[8],stage1_20[12],stage1_19[23],stage1_18[35],stage1_17[56]}
   );
   gpc606_5 gpc231 (
      {stage0_17[120], stage0_17[121], stage0_17[122], stage0_17[123], stage0_17[124], stage0_17[125]},
      {stage0_19[54], stage0_19[55], stage0_19[56], stage0_19[57], stage0_19[58], stage0_19[59]},
      {stage1_21[9],stage1_20[13],stage1_19[24],stage1_18[36],stage1_17[57]}
   );
   gpc606_5 gpc232 (
      {stage0_17[126], stage0_17[127], stage0_17[128], stage0_17[129], stage0_17[130], stage0_17[131]},
      {stage0_19[60], stage0_19[61], stage0_19[62], stage0_19[63], stage0_19[64], stage0_19[65]},
      {stage1_21[10],stage1_20[14],stage1_19[25],stage1_18[37],stage1_17[58]}
   );
   gpc606_5 gpc233 (
      {stage0_17[132], stage0_17[133], stage0_17[134], stage0_17[135], stage0_17[136], stage0_17[137]},
      {stage0_19[66], stage0_19[67], stage0_19[68], stage0_19[69], stage0_19[70], stage0_19[71]},
      {stage1_21[11],stage1_20[15],stage1_19[26],stage1_18[38],stage1_17[59]}
   );
   gpc606_5 gpc234 (
      {stage0_17[138], stage0_17[139], stage0_17[140], stage0_17[141], stage0_17[142], stage0_17[143]},
      {stage0_19[72], stage0_19[73], stage0_19[74], stage0_19[75], stage0_19[76], stage0_19[77]},
      {stage1_21[12],stage1_20[16],stage1_19[27],stage1_18[39],stage1_17[60]}
   );
   gpc606_5 gpc235 (
      {stage0_17[144], stage0_17[145], stage0_17[146], stage0_17[147], stage0_17[148], stage0_17[149]},
      {stage0_19[78], stage0_19[79], stage0_19[80], stage0_19[81], stage0_19[82], stage0_19[83]},
      {stage1_21[13],stage1_20[17],stage1_19[28],stage1_18[40],stage1_17[61]}
   );
   gpc606_5 gpc236 (
      {stage0_17[150], stage0_17[151], stage0_17[152], stage0_17[153], stage0_17[154], stage0_17[155]},
      {stage0_19[84], stage0_19[85], stage0_19[86], stage0_19[87], stage0_19[88], stage0_19[89]},
      {stage1_21[14],stage1_20[18],stage1_19[29],stage1_18[41],stage1_17[62]}
   );
   gpc606_5 gpc237 (
      {stage0_17[156], stage0_17[157], stage0_17[158], stage0_17[159], stage0_17[160], stage0_17[161]},
      {stage0_19[90], stage0_19[91], stage0_19[92], stage0_19[93], stage0_19[94], stage0_19[95]},
      {stage1_21[15],stage1_20[19],stage1_19[30],stage1_18[42],stage1_17[63]}
   );
   gpc117_4 gpc238 (
      {stage0_18[24], stage0_18[25], stage0_18[26], stage0_18[27], stage0_18[28], stage0_18[29], stage0_18[30]},
      {stage0_19[96]},
      {stage0_20[0]},
      {stage1_21[16],stage1_20[20],stage1_19[31],stage1_18[43]}
   );
   gpc117_4 gpc239 (
      {stage0_18[31], stage0_18[32], stage0_18[33], stage0_18[34], stage0_18[35], stage0_18[36], stage0_18[37]},
      {stage0_19[97]},
      {stage0_20[1]},
      {stage1_21[17],stage1_20[21],stage1_19[32],stage1_18[44]}
   );
   gpc117_4 gpc240 (
      {stage0_18[38], stage0_18[39], stage0_18[40], stage0_18[41], stage0_18[42], stage0_18[43], stage0_18[44]},
      {stage0_19[98]},
      {stage0_20[2]},
      {stage1_21[18],stage1_20[22],stage1_19[33],stage1_18[45]}
   );
   gpc117_4 gpc241 (
      {stage0_18[45], stage0_18[46], stage0_18[47], stage0_18[48], stage0_18[49], stage0_18[50], stage0_18[51]},
      {stage0_19[99]},
      {stage0_20[3]},
      {stage1_21[19],stage1_20[23],stage1_19[34],stage1_18[46]}
   );
   gpc606_5 gpc242 (
      {stage0_18[52], stage0_18[53], stage0_18[54], stage0_18[55], stage0_18[56], stage0_18[57]},
      {stage0_20[4], stage0_20[5], stage0_20[6], stage0_20[7], stage0_20[8], stage0_20[9]},
      {stage1_22[0],stage1_21[20],stage1_20[24],stage1_19[35],stage1_18[47]}
   );
   gpc606_5 gpc243 (
      {stage0_18[58], stage0_18[59], stage0_18[60], stage0_18[61], stage0_18[62], stage0_18[63]},
      {stage0_20[10], stage0_20[11], stage0_20[12], stage0_20[13], stage0_20[14], stage0_20[15]},
      {stage1_22[1],stage1_21[21],stage1_20[25],stage1_19[36],stage1_18[48]}
   );
   gpc606_5 gpc244 (
      {stage0_18[64], stage0_18[65], stage0_18[66], stage0_18[67], stage0_18[68], stage0_18[69]},
      {stage0_20[16], stage0_20[17], stage0_20[18], stage0_20[19], stage0_20[20], stage0_20[21]},
      {stage1_22[2],stage1_21[22],stage1_20[26],stage1_19[37],stage1_18[49]}
   );
   gpc606_5 gpc245 (
      {stage0_18[70], stage0_18[71], stage0_18[72], stage0_18[73], stage0_18[74], stage0_18[75]},
      {stage0_20[22], stage0_20[23], stage0_20[24], stage0_20[25], stage0_20[26], stage0_20[27]},
      {stage1_22[3],stage1_21[23],stage1_20[27],stage1_19[38],stage1_18[50]}
   );
   gpc606_5 gpc246 (
      {stage0_18[76], stage0_18[77], stage0_18[78], stage0_18[79], stage0_18[80], stage0_18[81]},
      {stage0_20[28], stage0_20[29], stage0_20[30], stage0_20[31], stage0_20[32], stage0_20[33]},
      {stage1_22[4],stage1_21[24],stage1_20[28],stage1_19[39],stage1_18[51]}
   );
   gpc606_5 gpc247 (
      {stage0_18[82], stage0_18[83], stage0_18[84], stage0_18[85], stage0_18[86], stage0_18[87]},
      {stage0_20[34], stage0_20[35], stage0_20[36], stage0_20[37], stage0_20[38], stage0_20[39]},
      {stage1_22[5],stage1_21[25],stage1_20[29],stage1_19[40],stage1_18[52]}
   );
   gpc606_5 gpc248 (
      {stage0_18[88], stage0_18[89], stage0_18[90], stage0_18[91], stage0_18[92], stage0_18[93]},
      {stage0_20[40], stage0_20[41], stage0_20[42], stage0_20[43], stage0_20[44], stage0_20[45]},
      {stage1_22[6],stage1_21[26],stage1_20[30],stage1_19[41],stage1_18[53]}
   );
   gpc606_5 gpc249 (
      {stage0_18[94], stage0_18[95], stage0_18[96], stage0_18[97], stage0_18[98], stage0_18[99]},
      {stage0_20[46], stage0_20[47], stage0_20[48], stage0_20[49], stage0_20[50], stage0_20[51]},
      {stage1_22[7],stage1_21[27],stage1_20[31],stage1_19[42],stage1_18[54]}
   );
   gpc606_5 gpc250 (
      {stage0_18[100], stage0_18[101], stage0_18[102], stage0_18[103], stage0_18[104], stage0_18[105]},
      {stage0_20[52], stage0_20[53], stage0_20[54], stage0_20[55], stage0_20[56], stage0_20[57]},
      {stage1_22[8],stage1_21[28],stage1_20[32],stage1_19[43],stage1_18[55]}
   );
   gpc606_5 gpc251 (
      {stage0_18[106], stage0_18[107], stage0_18[108], stage0_18[109], stage0_18[110], stage0_18[111]},
      {stage0_20[58], stage0_20[59], stage0_20[60], stage0_20[61], stage0_20[62], stage0_20[63]},
      {stage1_22[9],stage1_21[29],stage1_20[33],stage1_19[44],stage1_18[56]}
   );
   gpc606_5 gpc252 (
      {stage0_18[112], stage0_18[113], stage0_18[114], stage0_18[115], stage0_18[116], stage0_18[117]},
      {stage0_20[64], stage0_20[65], stage0_20[66], stage0_20[67], stage0_20[68], stage0_20[69]},
      {stage1_22[10],stage1_21[30],stage1_20[34],stage1_19[45],stage1_18[57]}
   );
   gpc606_5 gpc253 (
      {stage0_18[118], stage0_18[119], stage0_18[120], stage0_18[121], stage0_18[122], stage0_18[123]},
      {stage0_20[70], stage0_20[71], stage0_20[72], stage0_20[73], stage0_20[74], stage0_20[75]},
      {stage1_22[11],stage1_21[31],stage1_20[35],stage1_19[46],stage1_18[58]}
   );
   gpc606_5 gpc254 (
      {stage0_18[124], stage0_18[125], stage0_18[126], stage0_18[127], stage0_18[128], stage0_18[129]},
      {stage0_20[76], stage0_20[77], stage0_20[78], stage0_20[79], stage0_20[80], stage0_20[81]},
      {stage1_22[12],stage1_21[32],stage1_20[36],stage1_19[47],stage1_18[59]}
   );
   gpc606_5 gpc255 (
      {stage0_18[130], stage0_18[131], stage0_18[132], stage0_18[133], stage0_18[134], stage0_18[135]},
      {stage0_20[82], stage0_20[83], stage0_20[84], stage0_20[85], stage0_20[86], stage0_20[87]},
      {stage1_22[13],stage1_21[33],stage1_20[37],stage1_19[48],stage1_18[60]}
   );
   gpc606_5 gpc256 (
      {stage0_18[136], stage0_18[137], stage0_18[138], stage0_18[139], stage0_18[140], stage0_18[141]},
      {stage0_20[88], stage0_20[89], stage0_20[90], stage0_20[91], stage0_20[92], stage0_20[93]},
      {stage1_22[14],stage1_21[34],stage1_20[38],stage1_19[49],stage1_18[61]}
   );
   gpc606_5 gpc257 (
      {stage0_19[100], stage0_19[101], stage0_19[102], stage0_19[103], stage0_19[104], stage0_19[105]},
      {stage0_21[0], stage0_21[1], stage0_21[2], stage0_21[3], stage0_21[4], stage0_21[5]},
      {stage1_23[0],stage1_22[15],stage1_21[35],stage1_20[39],stage1_19[50]}
   );
   gpc606_5 gpc258 (
      {stage0_19[106], stage0_19[107], stage0_19[108], stage0_19[109], stage0_19[110], stage0_19[111]},
      {stage0_21[6], stage0_21[7], stage0_21[8], stage0_21[9], stage0_21[10], stage0_21[11]},
      {stage1_23[1],stage1_22[16],stage1_21[36],stage1_20[40],stage1_19[51]}
   );
   gpc606_5 gpc259 (
      {stage0_19[112], stage0_19[113], stage0_19[114], stage0_19[115], stage0_19[116], stage0_19[117]},
      {stage0_21[12], stage0_21[13], stage0_21[14], stage0_21[15], stage0_21[16], stage0_21[17]},
      {stage1_23[2],stage1_22[17],stage1_21[37],stage1_20[41],stage1_19[52]}
   );
   gpc606_5 gpc260 (
      {stage0_19[118], stage0_19[119], stage0_19[120], stage0_19[121], stage0_19[122], stage0_19[123]},
      {stage0_21[18], stage0_21[19], stage0_21[20], stage0_21[21], stage0_21[22], stage0_21[23]},
      {stage1_23[3],stage1_22[18],stage1_21[38],stage1_20[42],stage1_19[53]}
   );
   gpc606_5 gpc261 (
      {stage0_19[124], stage0_19[125], stage0_19[126], stage0_19[127], stage0_19[128], stage0_19[129]},
      {stage0_21[24], stage0_21[25], stage0_21[26], stage0_21[27], stage0_21[28], stage0_21[29]},
      {stage1_23[4],stage1_22[19],stage1_21[39],stage1_20[43],stage1_19[54]}
   );
   gpc606_5 gpc262 (
      {stage0_19[130], stage0_19[131], stage0_19[132], stage0_19[133], stage0_19[134], stage0_19[135]},
      {stage0_21[30], stage0_21[31], stage0_21[32], stage0_21[33], stage0_21[34], stage0_21[35]},
      {stage1_23[5],stage1_22[20],stage1_21[40],stage1_20[44],stage1_19[55]}
   );
   gpc606_5 gpc263 (
      {stage0_19[136], stage0_19[137], stage0_19[138], stage0_19[139], stage0_19[140], stage0_19[141]},
      {stage0_21[36], stage0_21[37], stage0_21[38], stage0_21[39], stage0_21[40], stage0_21[41]},
      {stage1_23[6],stage1_22[21],stage1_21[41],stage1_20[45],stage1_19[56]}
   );
   gpc606_5 gpc264 (
      {stage0_19[142], stage0_19[143], stage0_19[144], stage0_19[145], stage0_19[146], stage0_19[147]},
      {stage0_21[42], stage0_21[43], stage0_21[44], stage0_21[45], stage0_21[46], stage0_21[47]},
      {stage1_23[7],stage1_22[22],stage1_21[42],stage1_20[46],stage1_19[57]}
   );
   gpc606_5 gpc265 (
      {stage0_19[148], stage0_19[149], stage0_19[150], stage0_19[151], stage0_19[152], stage0_19[153]},
      {stage0_21[48], stage0_21[49], stage0_21[50], stage0_21[51], stage0_21[52], stage0_21[53]},
      {stage1_23[8],stage1_22[23],stage1_21[43],stage1_20[47],stage1_19[58]}
   );
   gpc606_5 gpc266 (
      {stage0_20[94], stage0_20[95], stage0_20[96], stage0_20[97], stage0_20[98], stage0_20[99]},
      {stage0_22[0], stage0_22[1], stage0_22[2], stage0_22[3], stage0_22[4], stage0_22[5]},
      {stage1_24[0],stage1_23[9],stage1_22[24],stage1_21[44],stage1_20[48]}
   );
   gpc606_5 gpc267 (
      {stage0_20[100], stage0_20[101], stage0_20[102], stage0_20[103], stage0_20[104], stage0_20[105]},
      {stage0_22[6], stage0_22[7], stage0_22[8], stage0_22[9], stage0_22[10], stage0_22[11]},
      {stage1_24[1],stage1_23[10],stage1_22[25],stage1_21[45],stage1_20[49]}
   );
   gpc606_5 gpc268 (
      {stage0_20[106], stage0_20[107], stage0_20[108], stage0_20[109], stage0_20[110], stage0_20[111]},
      {stage0_22[12], stage0_22[13], stage0_22[14], stage0_22[15], stage0_22[16], stage0_22[17]},
      {stage1_24[2],stage1_23[11],stage1_22[26],stage1_21[46],stage1_20[50]}
   );
   gpc615_5 gpc269 (
      {stage0_20[112], stage0_20[113], stage0_20[114], stage0_20[115], stage0_20[116]},
      {stage0_21[54]},
      {stage0_22[18], stage0_22[19], stage0_22[20], stage0_22[21], stage0_22[22], stage0_22[23]},
      {stage1_24[3],stage1_23[12],stage1_22[27],stage1_21[47],stage1_20[51]}
   );
   gpc615_5 gpc270 (
      {stage0_20[117], stage0_20[118], stage0_20[119], stage0_20[120], stage0_20[121]},
      {stage0_21[55]},
      {stage0_22[24], stage0_22[25], stage0_22[26], stage0_22[27], stage0_22[28], stage0_22[29]},
      {stage1_24[4],stage1_23[13],stage1_22[28],stage1_21[48],stage1_20[52]}
   );
   gpc615_5 gpc271 (
      {stage0_20[122], stage0_20[123], stage0_20[124], stage0_20[125], stage0_20[126]},
      {stage0_21[56]},
      {stage0_22[30], stage0_22[31], stage0_22[32], stage0_22[33], stage0_22[34], stage0_22[35]},
      {stage1_24[5],stage1_23[14],stage1_22[29],stage1_21[49],stage1_20[53]}
   );
   gpc615_5 gpc272 (
      {stage0_20[127], stage0_20[128], stage0_20[129], stage0_20[130], stage0_20[131]},
      {stage0_21[57]},
      {stage0_22[36], stage0_22[37], stage0_22[38], stage0_22[39], stage0_22[40], stage0_22[41]},
      {stage1_24[6],stage1_23[15],stage1_22[30],stage1_21[50],stage1_20[54]}
   );
   gpc615_5 gpc273 (
      {stage0_20[132], stage0_20[133], stage0_20[134], stage0_20[135], stage0_20[136]},
      {stage0_21[58]},
      {stage0_22[42], stage0_22[43], stage0_22[44], stage0_22[45], stage0_22[46], stage0_22[47]},
      {stage1_24[7],stage1_23[16],stage1_22[31],stage1_21[51],stage1_20[55]}
   );
   gpc615_5 gpc274 (
      {stage0_20[137], stage0_20[138], stage0_20[139], stage0_20[140], stage0_20[141]},
      {stage0_21[59]},
      {stage0_22[48], stage0_22[49], stage0_22[50], stage0_22[51], stage0_22[52], stage0_22[53]},
      {stage1_24[8],stage1_23[17],stage1_22[32],stage1_21[52],stage1_20[56]}
   );
   gpc615_5 gpc275 (
      {stage0_20[142], stage0_20[143], stage0_20[144], stage0_20[145], stage0_20[146]},
      {stage0_21[60]},
      {stage0_22[54], stage0_22[55], stage0_22[56], stage0_22[57], stage0_22[58], stage0_22[59]},
      {stage1_24[9],stage1_23[18],stage1_22[33],stage1_21[53],stage1_20[57]}
   );
   gpc615_5 gpc276 (
      {stage0_20[147], stage0_20[148], stage0_20[149], stage0_20[150], stage0_20[151]},
      {stage0_21[61]},
      {stage0_22[60], stage0_22[61], stage0_22[62], stage0_22[63], stage0_22[64], stage0_22[65]},
      {stage1_24[10],stage1_23[19],stage1_22[34],stage1_21[54],stage1_20[58]}
   );
   gpc615_5 gpc277 (
      {stage0_20[152], stage0_20[153], stage0_20[154], stage0_20[155], stage0_20[156]},
      {stage0_21[62]},
      {stage0_22[66], stage0_22[67], stage0_22[68], stage0_22[69], stage0_22[70], stage0_22[71]},
      {stage1_24[11],stage1_23[20],stage1_22[35],stage1_21[55],stage1_20[59]}
   );
   gpc615_5 gpc278 (
      {stage0_20[157], stage0_20[158], stage0_20[159], stage0_20[160], stage0_20[161]},
      {stage0_21[63]},
      {stage0_22[72], stage0_22[73], stage0_22[74], stage0_22[75], stage0_22[76], stage0_22[77]},
      {stage1_24[12],stage1_23[21],stage1_22[36],stage1_21[56],stage1_20[60]}
   );
   gpc1163_5 gpc279 (
      {stage0_21[64], stage0_21[65], stage0_21[66]},
      {stage0_22[78], stage0_22[79], stage0_22[80], stage0_22[81], stage0_22[82], stage0_22[83]},
      {stage0_23[0]},
      {stage0_24[0]},
      {stage1_25[0],stage1_24[13],stage1_23[22],stage1_22[37],stage1_21[57]}
   );
   gpc1163_5 gpc280 (
      {stage0_21[67], stage0_21[68], stage0_21[69]},
      {stage0_22[84], stage0_22[85], stage0_22[86], stage0_22[87], stage0_22[88], stage0_22[89]},
      {stage0_23[1]},
      {stage0_24[1]},
      {stage1_25[1],stage1_24[14],stage1_23[23],stage1_22[38],stage1_21[58]}
   );
   gpc1163_5 gpc281 (
      {stage0_21[70], stage0_21[71], stage0_21[72]},
      {stage0_22[90], stage0_22[91], stage0_22[92], stage0_22[93], stage0_22[94], stage0_22[95]},
      {stage0_23[2]},
      {stage0_24[2]},
      {stage1_25[2],stage1_24[15],stage1_23[24],stage1_22[39],stage1_21[59]}
   );
   gpc1163_5 gpc282 (
      {stage0_21[73], stage0_21[74], stage0_21[75]},
      {stage0_22[96], stage0_22[97], stage0_22[98], stage0_22[99], stage0_22[100], stage0_22[101]},
      {stage0_23[3]},
      {stage0_24[3]},
      {stage1_25[3],stage1_24[16],stage1_23[25],stage1_22[40],stage1_21[60]}
   );
   gpc1163_5 gpc283 (
      {stage0_21[76], stage0_21[77], stage0_21[78]},
      {stage0_22[102], stage0_22[103], stage0_22[104], stage0_22[105], stage0_22[106], stage0_22[107]},
      {stage0_23[4]},
      {stage0_24[4]},
      {stage1_25[4],stage1_24[17],stage1_23[26],stage1_22[41],stage1_21[61]}
   );
   gpc1163_5 gpc284 (
      {stage0_21[79], stage0_21[80], stage0_21[81]},
      {stage0_22[108], stage0_22[109], stage0_22[110], stage0_22[111], stage0_22[112], stage0_22[113]},
      {stage0_23[5]},
      {stage0_24[5]},
      {stage1_25[5],stage1_24[18],stage1_23[27],stage1_22[42],stage1_21[62]}
   );
   gpc1163_5 gpc285 (
      {stage0_21[82], stage0_21[83], stage0_21[84]},
      {stage0_22[114], stage0_22[115], stage0_22[116], stage0_22[117], stage0_22[118], stage0_22[119]},
      {stage0_23[6]},
      {stage0_24[6]},
      {stage1_25[6],stage1_24[19],stage1_23[28],stage1_22[43],stage1_21[63]}
   );
   gpc1163_5 gpc286 (
      {stage0_21[85], stage0_21[86], stage0_21[87]},
      {stage0_22[120], stage0_22[121], stage0_22[122], stage0_22[123], stage0_22[124], stage0_22[125]},
      {stage0_23[7]},
      {stage0_24[7]},
      {stage1_25[7],stage1_24[20],stage1_23[29],stage1_22[44],stage1_21[64]}
   );
   gpc1163_5 gpc287 (
      {stage0_21[88], stage0_21[89], stage0_21[90]},
      {stage0_22[126], stage0_22[127], stage0_22[128], stage0_22[129], stage0_22[130], stage0_22[131]},
      {stage0_23[8]},
      {stage0_24[8]},
      {stage1_25[8],stage1_24[21],stage1_23[30],stage1_22[45],stage1_21[65]}
   );
   gpc1163_5 gpc288 (
      {stage0_21[91], stage0_21[92], stage0_21[93]},
      {stage0_22[132], stage0_22[133], stage0_22[134], stage0_22[135], stage0_22[136], stage0_22[137]},
      {stage0_23[9]},
      {stage0_24[9]},
      {stage1_25[9],stage1_24[22],stage1_23[31],stage1_22[46],stage1_21[66]}
   );
   gpc606_5 gpc289 (
      {stage0_21[94], stage0_21[95], stage0_21[96], stage0_21[97], stage0_21[98], stage0_21[99]},
      {stage0_23[10], stage0_23[11], stage0_23[12], stage0_23[13], stage0_23[14], stage0_23[15]},
      {stage1_25[10],stage1_24[23],stage1_23[32],stage1_22[47],stage1_21[67]}
   );
   gpc606_5 gpc290 (
      {stage0_21[100], stage0_21[101], stage0_21[102], stage0_21[103], stage0_21[104], stage0_21[105]},
      {stage0_23[16], stage0_23[17], stage0_23[18], stage0_23[19], stage0_23[20], stage0_23[21]},
      {stage1_25[11],stage1_24[24],stage1_23[33],stage1_22[48],stage1_21[68]}
   );
   gpc606_5 gpc291 (
      {stage0_21[106], stage0_21[107], stage0_21[108], stage0_21[109], stage0_21[110], stage0_21[111]},
      {stage0_23[22], stage0_23[23], stage0_23[24], stage0_23[25], stage0_23[26], stage0_23[27]},
      {stage1_25[12],stage1_24[25],stage1_23[34],stage1_22[49],stage1_21[69]}
   );
   gpc606_5 gpc292 (
      {stage0_21[112], stage0_21[113], stage0_21[114], stage0_21[115], stage0_21[116], stage0_21[117]},
      {stage0_23[28], stage0_23[29], stage0_23[30], stage0_23[31], stage0_23[32], stage0_23[33]},
      {stage1_25[13],stage1_24[26],stage1_23[35],stage1_22[50],stage1_21[70]}
   );
   gpc606_5 gpc293 (
      {stage0_21[118], stage0_21[119], stage0_21[120], stage0_21[121], stage0_21[122], stage0_21[123]},
      {stage0_23[34], stage0_23[35], stage0_23[36], stage0_23[37], stage0_23[38], stage0_23[39]},
      {stage1_25[14],stage1_24[27],stage1_23[36],stage1_22[51],stage1_21[71]}
   );
   gpc606_5 gpc294 (
      {stage0_21[124], stage0_21[125], stage0_21[126], stage0_21[127], stage0_21[128], stage0_21[129]},
      {stage0_23[40], stage0_23[41], stage0_23[42], stage0_23[43], stage0_23[44], stage0_23[45]},
      {stage1_25[15],stage1_24[28],stage1_23[37],stage1_22[52],stage1_21[72]}
   );
   gpc606_5 gpc295 (
      {stage0_21[130], stage0_21[131], stage0_21[132], stage0_21[133], stage0_21[134], stage0_21[135]},
      {stage0_23[46], stage0_23[47], stage0_23[48], stage0_23[49], stage0_23[50], stage0_23[51]},
      {stage1_25[16],stage1_24[29],stage1_23[38],stage1_22[53],stage1_21[73]}
   );
   gpc606_5 gpc296 (
      {stage0_21[136], stage0_21[137], stage0_21[138], stage0_21[139], stage0_21[140], stage0_21[141]},
      {stage0_23[52], stage0_23[53], stage0_23[54], stage0_23[55], stage0_23[56], stage0_23[57]},
      {stage1_25[17],stage1_24[30],stage1_23[39],stage1_22[54],stage1_21[74]}
   );
   gpc606_5 gpc297 (
      {stage0_21[142], stage0_21[143], stage0_21[144], stage0_21[145], stage0_21[146], stage0_21[147]},
      {stage0_23[58], stage0_23[59], stage0_23[60], stage0_23[61], stage0_23[62], stage0_23[63]},
      {stage1_25[18],stage1_24[31],stage1_23[40],stage1_22[55],stage1_21[75]}
   );
   gpc606_5 gpc298 (
      {stage0_21[148], stage0_21[149], stage0_21[150], stage0_21[151], stage0_21[152], stage0_21[153]},
      {stage0_23[64], stage0_23[65], stage0_23[66], stage0_23[67], stage0_23[68], stage0_23[69]},
      {stage1_25[19],stage1_24[32],stage1_23[41],stage1_22[56],stage1_21[76]}
   );
   gpc606_5 gpc299 (
      {stage0_21[154], stage0_21[155], stage0_21[156], stage0_21[157], stage0_21[158], stage0_21[159]},
      {stage0_23[70], stage0_23[71], stage0_23[72], stage0_23[73], stage0_23[74], stage0_23[75]},
      {stage1_25[20],stage1_24[33],stage1_23[42],stage1_22[57],stage1_21[77]}
   );
   gpc606_5 gpc300 (
      {stage0_23[76], stage0_23[77], stage0_23[78], stage0_23[79], stage0_23[80], stage0_23[81]},
      {stage0_25[0], stage0_25[1], stage0_25[2], stage0_25[3], stage0_25[4], stage0_25[5]},
      {stage1_27[0],stage1_26[0],stage1_25[21],stage1_24[34],stage1_23[43]}
   );
   gpc606_5 gpc301 (
      {stage0_23[82], stage0_23[83], stage0_23[84], stage0_23[85], stage0_23[86], stage0_23[87]},
      {stage0_25[6], stage0_25[7], stage0_25[8], stage0_25[9], stage0_25[10], stage0_25[11]},
      {stage1_27[1],stage1_26[1],stage1_25[22],stage1_24[35],stage1_23[44]}
   );
   gpc606_5 gpc302 (
      {stage0_23[88], stage0_23[89], stage0_23[90], stage0_23[91], stage0_23[92], stage0_23[93]},
      {stage0_25[12], stage0_25[13], stage0_25[14], stage0_25[15], stage0_25[16], stage0_25[17]},
      {stage1_27[2],stage1_26[2],stage1_25[23],stage1_24[36],stage1_23[45]}
   );
   gpc606_5 gpc303 (
      {stage0_23[94], stage0_23[95], stage0_23[96], stage0_23[97], stage0_23[98], stage0_23[99]},
      {stage0_25[18], stage0_25[19], stage0_25[20], stage0_25[21], stage0_25[22], stage0_25[23]},
      {stage1_27[3],stage1_26[3],stage1_25[24],stage1_24[37],stage1_23[46]}
   );
   gpc606_5 gpc304 (
      {stage0_23[100], stage0_23[101], stage0_23[102], stage0_23[103], stage0_23[104], stage0_23[105]},
      {stage0_25[24], stage0_25[25], stage0_25[26], stage0_25[27], stage0_25[28], stage0_25[29]},
      {stage1_27[4],stage1_26[4],stage1_25[25],stage1_24[38],stage1_23[47]}
   );
   gpc606_5 gpc305 (
      {stage0_23[106], stage0_23[107], stage0_23[108], stage0_23[109], stage0_23[110], stage0_23[111]},
      {stage0_25[30], stage0_25[31], stage0_25[32], stage0_25[33], stage0_25[34], stage0_25[35]},
      {stage1_27[5],stage1_26[5],stage1_25[26],stage1_24[39],stage1_23[48]}
   );
   gpc615_5 gpc306 (
      {stage0_23[112], stage0_23[113], stage0_23[114], stage0_23[115], stage0_23[116]},
      {stage0_24[10]},
      {stage0_25[36], stage0_25[37], stage0_25[38], stage0_25[39], stage0_25[40], stage0_25[41]},
      {stage1_27[6],stage1_26[6],stage1_25[27],stage1_24[40],stage1_23[49]}
   );
   gpc615_5 gpc307 (
      {stage0_23[117], stage0_23[118], stage0_23[119], stage0_23[120], stage0_23[121]},
      {stage0_24[11]},
      {stage0_25[42], stage0_25[43], stage0_25[44], stage0_25[45], stage0_25[46], stage0_25[47]},
      {stage1_27[7],stage1_26[7],stage1_25[28],stage1_24[41],stage1_23[50]}
   );
   gpc606_5 gpc308 (
      {stage0_24[12], stage0_24[13], stage0_24[14], stage0_24[15], stage0_24[16], stage0_24[17]},
      {stage0_26[0], stage0_26[1], stage0_26[2], stage0_26[3], stage0_26[4], stage0_26[5]},
      {stage1_28[0],stage1_27[8],stage1_26[8],stage1_25[29],stage1_24[42]}
   );
   gpc606_5 gpc309 (
      {stage0_24[18], stage0_24[19], stage0_24[20], stage0_24[21], stage0_24[22], stage0_24[23]},
      {stage0_26[6], stage0_26[7], stage0_26[8], stage0_26[9], stage0_26[10], stage0_26[11]},
      {stage1_28[1],stage1_27[9],stage1_26[9],stage1_25[30],stage1_24[43]}
   );
   gpc606_5 gpc310 (
      {stage0_24[24], stage0_24[25], stage0_24[26], stage0_24[27], stage0_24[28], stage0_24[29]},
      {stage0_26[12], stage0_26[13], stage0_26[14], stage0_26[15], stage0_26[16], stage0_26[17]},
      {stage1_28[2],stage1_27[10],stage1_26[10],stage1_25[31],stage1_24[44]}
   );
   gpc606_5 gpc311 (
      {stage0_24[30], stage0_24[31], stage0_24[32], stage0_24[33], stage0_24[34], stage0_24[35]},
      {stage0_26[18], stage0_26[19], stage0_26[20], stage0_26[21], stage0_26[22], stage0_26[23]},
      {stage1_28[3],stage1_27[11],stage1_26[11],stage1_25[32],stage1_24[45]}
   );
   gpc606_5 gpc312 (
      {stage0_24[36], stage0_24[37], stage0_24[38], stage0_24[39], stage0_24[40], stage0_24[41]},
      {stage0_26[24], stage0_26[25], stage0_26[26], stage0_26[27], stage0_26[28], stage0_26[29]},
      {stage1_28[4],stage1_27[12],stage1_26[12],stage1_25[33],stage1_24[46]}
   );
   gpc606_5 gpc313 (
      {stage0_24[42], stage0_24[43], stage0_24[44], stage0_24[45], stage0_24[46], stage0_24[47]},
      {stage0_26[30], stage0_26[31], stage0_26[32], stage0_26[33], stage0_26[34], stage0_26[35]},
      {stage1_28[5],stage1_27[13],stage1_26[13],stage1_25[34],stage1_24[47]}
   );
   gpc606_5 gpc314 (
      {stage0_24[48], stage0_24[49], stage0_24[50], stage0_24[51], stage0_24[52], stage0_24[53]},
      {stage0_26[36], stage0_26[37], stage0_26[38], stage0_26[39], stage0_26[40], stage0_26[41]},
      {stage1_28[6],stage1_27[14],stage1_26[14],stage1_25[35],stage1_24[48]}
   );
   gpc606_5 gpc315 (
      {stage0_24[54], stage0_24[55], stage0_24[56], stage0_24[57], stage0_24[58], stage0_24[59]},
      {stage0_26[42], stage0_26[43], stage0_26[44], stage0_26[45], stage0_26[46], stage0_26[47]},
      {stage1_28[7],stage1_27[15],stage1_26[15],stage1_25[36],stage1_24[49]}
   );
   gpc606_5 gpc316 (
      {stage0_24[60], stage0_24[61], stage0_24[62], stage0_24[63], stage0_24[64], stage0_24[65]},
      {stage0_26[48], stage0_26[49], stage0_26[50], stage0_26[51], stage0_26[52], stage0_26[53]},
      {stage1_28[8],stage1_27[16],stage1_26[16],stage1_25[37],stage1_24[50]}
   );
   gpc606_5 gpc317 (
      {stage0_24[66], stage0_24[67], stage0_24[68], stage0_24[69], stage0_24[70], stage0_24[71]},
      {stage0_26[54], stage0_26[55], stage0_26[56], stage0_26[57], stage0_26[58], stage0_26[59]},
      {stage1_28[9],stage1_27[17],stage1_26[17],stage1_25[38],stage1_24[51]}
   );
   gpc606_5 gpc318 (
      {stage0_24[72], stage0_24[73], stage0_24[74], stage0_24[75], stage0_24[76], stage0_24[77]},
      {stage0_26[60], stage0_26[61], stage0_26[62], stage0_26[63], stage0_26[64], stage0_26[65]},
      {stage1_28[10],stage1_27[18],stage1_26[18],stage1_25[39],stage1_24[52]}
   );
   gpc606_5 gpc319 (
      {stage0_24[78], stage0_24[79], stage0_24[80], stage0_24[81], stage0_24[82], stage0_24[83]},
      {stage0_26[66], stage0_26[67], stage0_26[68], stage0_26[69], stage0_26[70], stage0_26[71]},
      {stage1_28[11],stage1_27[19],stage1_26[19],stage1_25[40],stage1_24[53]}
   );
   gpc606_5 gpc320 (
      {stage0_24[84], stage0_24[85], stage0_24[86], stage0_24[87], stage0_24[88], stage0_24[89]},
      {stage0_26[72], stage0_26[73], stage0_26[74], stage0_26[75], stage0_26[76], stage0_26[77]},
      {stage1_28[12],stage1_27[20],stage1_26[20],stage1_25[41],stage1_24[54]}
   );
   gpc606_5 gpc321 (
      {stage0_24[90], stage0_24[91], stage0_24[92], stage0_24[93], stage0_24[94], stage0_24[95]},
      {stage0_26[78], stage0_26[79], stage0_26[80], stage0_26[81], stage0_26[82], stage0_26[83]},
      {stage1_28[13],stage1_27[21],stage1_26[21],stage1_25[42],stage1_24[55]}
   );
   gpc606_5 gpc322 (
      {stage0_24[96], stage0_24[97], stage0_24[98], stage0_24[99], stage0_24[100], stage0_24[101]},
      {stage0_26[84], stage0_26[85], stage0_26[86], stage0_26[87], stage0_26[88], stage0_26[89]},
      {stage1_28[14],stage1_27[22],stage1_26[22],stage1_25[43],stage1_24[56]}
   );
   gpc606_5 gpc323 (
      {stage0_24[102], stage0_24[103], stage0_24[104], stage0_24[105], stage0_24[106], stage0_24[107]},
      {stage0_26[90], stage0_26[91], stage0_26[92], stage0_26[93], stage0_26[94], stage0_26[95]},
      {stage1_28[15],stage1_27[23],stage1_26[23],stage1_25[44],stage1_24[57]}
   );
   gpc606_5 gpc324 (
      {stage0_24[108], stage0_24[109], stage0_24[110], stage0_24[111], stage0_24[112], stage0_24[113]},
      {stage0_26[96], stage0_26[97], stage0_26[98], stage0_26[99], stage0_26[100], stage0_26[101]},
      {stage1_28[16],stage1_27[24],stage1_26[24],stage1_25[45],stage1_24[58]}
   );
   gpc606_5 gpc325 (
      {stage0_24[114], stage0_24[115], stage0_24[116], stage0_24[117], stage0_24[118], stage0_24[119]},
      {stage0_26[102], stage0_26[103], stage0_26[104], stage0_26[105], stage0_26[106], stage0_26[107]},
      {stage1_28[17],stage1_27[25],stage1_26[25],stage1_25[46],stage1_24[59]}
   );
   gpc606_5 gpc326 (
      {stage0_24[120], stage0_24[121], stage0_24[122], stage0_24[123], stage0_24[124], stage0_24[125]},
      {stage0_26[108], stage0_26[109], stage0_26[110], stage0_26[111], stage0_26[112], stage0_26[113]},
      {stage1_28[18],stage1_27[26],stage1_26[26],stage1_25[47],stage1_24[60]}
   );
   gpc606_5 gpc327 (
      {stage0_24[126], stage0_24[127], stage0_24[128], stage0_24[129], stage0_24[130], stage0_24[131]},
      {stage0_26[114], stage0_26[115], stage0_26[116], stage0_26[117], stage0_26[118], stage0_26[119]},
      {stage1_28[19],stage1_27[27],stage1_26[27],stage1_25[48],stage1_24[61]}
   );
   gpc606_5 gpc328 (
      {stage0_24[132], stage0_24[133], stage0_24[134], stage0_24[135], stage0_24[136], stage0_24[137]},
      {stage0_26[120], stage0_26[121], stage0_26[122], stage0_26[123], stage0_26[124], stage0_26[125]},
      {stage1_28[20],stage1_27[28],stage1_26[28],stage1_25[49],stage1_24[62]}
   );
   gpc606_5 gpc329 (
      {stage0_24[138], stage0_24[139], stage0_24[140], stage0_24[141], stage0_24[142], stage0_24[143]},
      {stage0_26[126], stage0_26[127], stage0_26[128], stage0_26[129], stage0_26[130], stage0_26[131]},
      {stage1_28[21],stage1_27[29],stage1_26[29],stage1_25[50],stage1_24[63]}
   );
   gpc606_5 gpc330 (
      {stage0_24[144], stage0_24[145], stage0_24[146], stage0_24[147], stage0_24[148], stage0_24[149]},
      {stage0_26[132], stage0_26[133], stage0_26[134], stage0_26[135], stage0_26[136], stage0_26[137]},
      {stage1_28[22],stage1_27[30],stage1_26[30],stage1_25[51],stage1_24[64]}
   );
   gpc606_5 gpc331 (
      {stage0_24[150], stage0_24[151], stage0_24[152], stage0_24[153], stage0_24[154], stage0_24[155]},
      {stage0_26[138], stage0_26[139], stage0_26[140], stage0_26[141], stage0_26[142], stage0_26[143]},
      {stage1_28[23],stage1_27[31],stage1_26[31],stage1_25[52],stage1_24[65]}
   );
   gpc606_5 gpc332 (
      {stage0_24[156], stage0_24[157], stage0_24[158], stage0_24[159], stage0_24[160], stage0_24[161]},
      {stage0_26[144], stage0_26[145], stage0_26[146], stage0_26[147], stage0_26[148], stage0_26[149]},
      {stage1_28[24],stage1_27[32],stage1_26[32],stage1_25[53],stage1_24[66]}
   );
   gpc606_5 gpc333 (
      {stage0_25[48], stage0_25[49], stage0_25[50], stage0_25[51], stage0_25[52], stage0_25[53]},
      {stage0_27[0], stage0_27[1], stage0_27[2], stage0_27[3], stage0_27[4], stage0_27[5]},
      {stage1_29[0],stage1_28[25],stage1_27[33],stage1_26[33],stage1_25[54]}
   );
   gpc606_5 gpc334 (
      {stage0_25[54], stage0_25[55], stage0_25[56], stage0_25[57], stage0_25[58], stage0_25[59]},
      {stage0_27[6], stage0_27[7], stage0_27[8], stage0_27[9], stage0_27[10], stage0_27[11]},
      {stage1_29[1],stage1_28[26],stage1_27[34],stage1_26[34],stage1_25[55]}
   );
   gpc606_5 gpc335 (
      {stage0_25[60], stage0_25[61], stage0_25[62], stage0_25[63], stage0_25[64], stage0_25[65]},
      {stage0_27[12], stage0_27[13], stage0_27[14], stage0_27[15], stage0_27[16], stage0_27[17]},
      {stage1_29[2],stage1_28[27],stage1_27[35],stage1_26[35],stage1_25[56]}
   );
   gpc606_5 gpc336 (
      {stage0_25[66], stage0_25[67], stage0_25[68], stage0_25[69], stage0_25[70], stage0_25[71]},
      {stage0_27[18], stage0_27[19], stage0_27[20], stage0_27[21], stage0_27[22], stage0_27[23]},
      {stage1_29[3],stage1_28[28],stage1_27[36],stage1_26[36],stage1_25[57]}
   );
   gpc606_5 gpc337 (
      {stage0_25[72], stage0_25[73], stage0_25[74], stage0_25[75], stage0_25[76], stage0_25[77]},
      {stage0_27[24], stage0_27[25], stage0_27[26], stage0_27[27], stage0_27[28], stage0_27[29]},
      {stage1_29[4],stage1_28[29],stage1_27[37],stage1_26[37],stage1_25[58]}
   );
   gpc606_5 gpc338 (
      {stage0_25[78], stage0_25[79], stage0_25[80], stage0_25[81], stage0_25[82], stage0_25[83]},
      {stage0_27[30], stage0_27[31], stage0_27[32], stage0_27[33], stage0_27[34], stage0_27[35]},
      {stage1_29[5],stage1_28[30],stage1_27[38],stage1_26[38],stage1_25[59]}
   );
   gpc606_5 gpc339 (
      {stage0_25[84], stage0_25[85], stage0_25[86], stage0_25[87], stage0_25[88], stage0_25[89]},
      {stage0_27[36], stage0_27[37], stage0_27[38], stage0_27[39], stage0_27[40], stage0_27[41]},
      {stage1_29[6],stage1_28[31],stage1_27[39],stage1_26[39],stage1_25[60]}
   );
   gpc606_5 gpc340 (
      {stage0_25[90], stage0_25[91], stage0_25[92], stage0_25[93], stage0_25[94], stage0_25[95]},
      {stage0_27[42], stage0_27[43], stage0_27[44], stage0_27[45], stage0_27[46], stage0_27[47]},
      {stage1_29[7],stage1_28[32],stage1_27[40],stage1_26[40],stage1_25[61]}
   );
   gpc606_5 gpc341 (
      {stage0_25[96], stage0_25[97], stage0_25[98], stage0_25[99], stage0_25[100], stage0_25[101]},
      {stage0_27[48], stage0_27[49], stage0_27[50], stage0_27[51], stage0_27[52], stage0_27[53]},
      {stage1_29[8],stage1_28[33],stage1_27[41],stage1_26[41],stage1_25[62]}
   );
   gpc606_5 gpc342 (
      {stage0_25[102], stage0_25[103], stage0_25[104], stage0_25[105], stage0_25[106], stage0_25[107]},
      {stage0_27[54], stage0_27[55], stage0_27[56], stage0_27[57], stage0_27[58], stage0_27[59]},
      {stage1_29[9],stage1_28[34],stage1_27[42],stage1_26[42],stage1_25[63]}
   );
   gpc615_5 gpc343 (
      {stage0_25[108], stage0_25[109], stage0_25[110], stage0_25[111], stage0_25[112]},
      {stage0_26[150]},
      {stage0_27[60], stage0_27[61], stage0_27[62], stage0_27[63], stage0_27[64], stage0_27[65]},
      {stage1_29[10],stage1_28[35],stage1_27[43],stage1_26[43],stage1_25[64]}
   );
   gpc615_5 gpc344 (
      {stage0_25[113], stage0_25[114], stage0_25[115], stage0_25[116], stage0_25[117]},
      {stage0_26[151]},
      {stage0_27[66], stage0_27[67], stage0_27[68], stage0_27[69], stage0_27[70], stage0_27[71]},
      {stage1_29[11],stage1_28[36],stage1_27[44],stage1_26[44],stage1_25[65]}
   );
   gpc615_5 gpc345 (
      {stage0_25[118], stage0_25[119], stage0_25[120], stage0_25[121], stage0_25[122]},
      {stage0_26[152]},
      {stage0_27[72], stage0_27[73], stage0_27[74], stage0_27[75], stage0_27[76], stage0_27[77]},
      {stage1_29[12],stage1_28[37],stage1_27[45],stage1_26[45],stage1_25[66]}
   );
   gpc615_5 gpc346 (
      {stage0_25[123], stage0_25[124], stage0_25[125], stage0_25[126], stage0_25[127]},
      {stage0_26[153]},
      {stage0_27[78], stage0_27[79], stage0_27[80], stage0_27[81], stage0_27[82], stage0_27[83]},
      {stage1_29[13],stage1_28[38],stage1_27[46],stage1_26[46],stage1_25[67]}
   );
   gpc615_5 gpc347 (
      {stage0_25[128], stage0_25[129], stage0_25[130], stage0_25[131], stage0_25[132]},
      {stage0_26[154]},
      {stage0_27[84], stage0_27[85], stage0_27[86], stage0_27[87], stage0_27[88], stage0_27[89]},
      {stage1_29[14],stage1_28[39],stage1_27[47],stage1_26[47],stage1_25[68]}
   );
   gpc615_5 gpc348 (
      {stage0_25[133], stage0_25[134], stage0_25[135], stage0_25[136], stage0_25[137]},
      {stage0_26[155]},
      {stage0_27[90], stage0_27[91], stage0_27[92], stage0_27[93], stage0_27[94], stage0_27[95]},
      {stage1_29[15],stage1_28[40],stage1_27[48],stage1_26[48],stage1_25[69]}
   );
   gpc615_5 gpc349 (
      {stage0_25[138], stage0_25[139], stage0_25[140], stage0_25[141], stage0_25[142]},
      {stage0_26[156]},
      {stage0_27[96], stage0_27[97], stage0_27[98], stage0_27[99], stage0_27[100], stage0_27[101]},
      {stage1_29[16],stage1_28[41],stage1_27[49],stage1_26[49],stage1_25[70]}
   );
   gpc615_5 gpc350 (
      {stage0_25[143], stage0_25[144], stage0_25[145], stage0_25[146], stage0_25[147]},
      {stage0_26[157]},
      {stage0_27[102], stage0_27[103], stage0_27[104], stage0_27[105], stage0_27[106], stage0_27[107]},
      {stage1_29[17],stage1_28[42],stage1_27[50],stage1_26[50],stage1_25[71]}
   );
   gpc615_5 gpc351 (
      {stage0_25[148], stage0_25[149], stage0_25[150], stage0_25[151], stage0_25[152]},
      {stage0_26[158]},
      {stage0_27[108], stage0_27[109], stage0_27[110], stage0_27[111], stage0_27[112], stage0_27[113]},
      {stage1_29[18],stage1_28[43],stage1_27[51],stage1_26[51],stage1_25[72]}
   );
   gpc615_5 gpc352 (
      {stage0_25[153], stage0_25[154], stage0_25[155], stage0_25[156], stage0_25[157]},
      {stage0_26[159]},
      {stage0_27[114], stage0_27[115], stage0_27[116], stage0_27[117], stage0_27[118], stage0_27[119]},
      {stage1_29[19],stage1_28[44],stage1_27[52],stage1_26[52],stage1_25[73]}
   );
   gpc615_5 gpc353 (
      {stage0_27[120], stage0_27[121], stage0_27[122], stage0_27[123], stage0_27[124]},
      {stage0_28[0]},
      {stage0_29[0], stage0_29[1], stage0_29[2], stage0_29[3], stage0_29[4], stage0_29[5]},
      {stage1_31[0],stage1_30[0],stage1_29[20],stage1_28[45],stage1_27[53]}
   );
   gpc615_5 gpc354 (
      {stage0_27[125], stage0_27[126], stage0_27[127], stage0_27[128], stage0_27[129]},
      {stage0_28[1]},
      {stage0_29[6], stage0_29[7], stage0_29[8], stage0_29[9], stage0_29[10], stage0_29[11]},
      {stage1_31[1],stage1_30[1],stage1_29[21],stage1_28[46],stage1_27[54]}
   );
   gpc615_5 gpc355 (
      {stage0_27[130], stage0_27[131], stage0_27[132], stage0_27[133], stage0_27[134]},
      {stage0_28[2]},
      {stage0_29[12], stage0_29[13], stage0_29[14], stage0_29[15], stage0_29[16], stage0_29[17]},
      {stage1_31[2],stage1_30[2],stage1_29[22],stage1_28[47],stage1_27[55]}
   );
   gpc615_5 gpc356 (
      {stage0_27[135], stage0_27[136], stage0_27[137], stage0_27[138], stage0_27[139]},
      {stage0_28[3]},
      {stage0_29[18], stage0_29[19], stage0_29[20], stage0_29[21], stage0_29[22], stage0_29[23]},
      {stage1_31[3],stage1_30[3],stage1_29[23],stage1_28[48],stage1_27[56]}
   );
   gpc615_5 gpc357 (
      {stage0_27[140], stage0_27[141], stage0_27[142], stage0_27[143], stage0_27[144]},
      {stage0_28[4]},
      {stage0_29[24], stage0_29[25], stage0_29[26], stage0_29[27], stage0_29[28], stage0_29[29]},
      {stage1_31[4],stage1_30[4],stage1_29[24],stage1_28[49],stage1_27[57]}
   );
   gpc615_5 gpc358 (
      {stage0_27[145], stage0_27[146], stage0_27[147], stage0_27[148], stage0_27[149]},
      {stage0_28[5]},
      {stage0_29[30], stage0_29[31], stage0_29[32], stage0_29[33], stage0_29[34], stage0_29[35]},
      {stage1_31[5],stage1_30[5],stage1_29[25],stage1_28[50],stage1_27[58]}
   );
   gpc615_5 gpc359 (
      {stage0_27[150], stage0_27[151], stage0_27[152], stage0_27[153], stage0_27[154]},
      {stage0_28[6]},
      {stage0_29[36], stage0_29[37], stage0_29[38], stage0_29[39], stage0_29[40], stage0_29[41]},
      {stage1_31[6],stage1_30[6],stage1_29[26],stage1_28[51],stage1_27[59]}
   );
   gpc2135_5 gpc360 (
      {stage0_28[7], stage0_28[8], stage0_28[9], stage0_28[10], stage0_28[11]},
      {stage0_29[42], stage0_29[43], stage0_29[44]},
      {stage0_30[0]},
      {stage0_31[0], stage0_31[1]},
      {stage1_32[0],stage1_31[7],stage1_30[7],stage1_29[27],stage1_28[52]}
   );
   gpc606_5 gpc361 (
      {stage0_28[12], stage0_28[13], stage0_28[14], stage0_28[15], stage0_28[16], stage0_28[17]},
      {stage0_30[1], stage0_30[2], stage0_30[3], stage0_30[4], stage0_30[5], stage0_30[6]},
      {stage1_32[1],stage1_31[8],stage1_30[8],stage1_29[28],stage1_28[53]}
   );
   gpc606_5 gpc362 (
      {stage0_28[18], stage0_28[19], stage0_28[20], stage0_28[21], stage0_28[22], stage0_28[23]},
      {stage0_30[7], stage0_30[8], stage0_30[9], stage0_30[10], stage0_30[11], stage0_30[12]},
      {stage1_32[2],stage1_31[9],stage1_30[9],stage1_29[29],stage1_28[54]}
   );
   gpc606_5 gpc363 (
      {stage0_28[24], stage0_28[25], stage0_28[26], stage0_28[27], stage0_28[28], stage0_28[29]},
      {stage0_30[13], stage0_30[14], stage0_30[15], stage0_30[16], stage0_30[17], stage0_30[18]},
      {stage1_32[3],stage1_31[10],stage1_30[10],stage1_29[30],stage1_28[55]}
   );
   gpc606_5 gpc364 (
      {stage0_28[30], stage0_28[31], stage0_28[32], stage0_28[33], stage0_28[34], stage0_28[35]},
      {stage0_30[19], stage0_30[20], stage0_30[21], stage0_30[22], stage0_30[23], stage0_30[24]},
      {stage1_32[4],stage1_31[11],stage1_30[11],stage1_29[31],stage1_28[56]}
   );
   gpc606_5 gpc365 (
      {stage0_28[36], stage0_28[37], stage0_28[38], stage0_28[39], stage0_28[40], stage0_28[41]},
      {stage0_30[25], stage0_30[26], stage0_30[27], stage0_30[28], stage0_30[29], stage0_30[30]},
      {stage1_32[5],stage1_31[12],stage1_30[12],stage1_29[32],stage1_28[57]}
   );
   gpc606_5 gpc366 (
      {stage0_28[42], stage0_28[43], stage0_28[44], stage0_28[45], stage0_28[46], stage0_28[47]},
      {stage0_30[31], stage0_30[32], stage0_30[33], stage0_30[34], stage0_30[35], stage0_30[36]},
      {stage1_32[6],stage1_31[13],stage1_30[13],stage1_29[33],stage1_28[58]}
   );
   gpc606_5 gpc367 (
      {stage0_28[48], stage0_28[49], stage0_28[50], stage0_28[51], stage0_28[52], stage0_28[53]},
      {stage0_30[37], stage0_30[38], stage0_30[39], stage0_30[40], stage0_30[41], stage0_30[42]},
      {stage1_32[7],stage1_31[14],stage1_30[14],stage1_29[34],stage1_28[59]}
   );
   gpc606_5 gpc368 (
      {stage0_28[54], stage0_28[55], stage0_28[56], stage0_28[57], stage0_28[58], stage0_28[59]},
      {stage0_30[43], stage0_30[44], stage0_30[45], stage0_30[46], stage0_30[47], stage0_30[48]},
      {stage1_32[8],stage1_31[15],stage1_30[15],stage1_29[35],stage1_28[60]}
   );
   gpc606_5 gpc369 (
      {stage0_28[60], stage0_28[61], stage0_28[62], stage0_28[63], stage0_28[64], stage0_28[65]},
      {stage0_30[49], stage0_30[50], stage0_30[51], stage0_30[52], stage0_30[53], stage0_30[54]},
      {stage1_32[9],stage1_31[16],stage1_30[16],stage1_29[36],stage1_28[61]}
   );
   gpc606_5 gpc370 (
      {stage0_28[66], stage0_28[67], stage0_28[68], stage0_28[69], stage0_28[70], stage0_28[71]},
      {stage0_30[55], stage0_30[56], stage0_30[57], stage0_30[58], stage0_30[59], stage0_30[60]},
      {stage1_32[10],stage1_31[17],stage1_30[17],stage1_29[37],stage1_28[62]}
   );
   gpc606_5 gpc371 (
      {stage0_28[72], stage0_28[73], stage0_28[74], stage0_28[75], stage0_28[76], stage0_28[77]},
      {stage0_30[61], stage0_30[62], stage0_30[63], stage0_30[64], stage0_30[65], stage0_30[66]},
      {stage1_32[11],stage1_31[18],stage1_30[18],stage1_29[38],stage1_28[63]}
   );
   gpc606_5 gpc372 (
      {stage0_28[78], stage0_28[79], stage0_28[80], stage0_28[81], stage0_28[82], stage0_28[83]},
      {stage0_30[67], stage0_30[68], stage0_30[69], stage0_30[70], stage0_30[71], stage0_30[72]},
      {stage1_32[12],stage1_31[19],stage1_30[19],stage1_29[39],stage1_28[64]}
   );
   gpc606_5 gpc373 (
      {stage0_28[84], stage0_28[85], stage0_28[86], stage0_28[87], stage0_28[88], stage0_28[89]},
      {stage0_30[73], stage0_30[74], stage0_30[75], stage0_30[76], stage0_30[77], stage0_30[78]},
      {stage1_32[13],stage1_31[20],stage1_30[20],stage1_29[40],stage1_28[65]}
   );
   gpc606_5 gpc374 (
      {stage0_28[90], stage0_28[91], stage0_28[92], stage0_28[93], stage0_28[94], stage0_28[95]},
      {stage0_30[79], stage0_30[80], stage0_30[81], stage0_30[82], stage0_30[83], stage0_30[84]},
      {stage1_32[14],stage1_31[21],stage1_30[21],stage1_29[41],stage1_28[66]}
   );
   gpc606_5 gpc375 (
      {stage0_28[96], stage0_28[97], stage0_28[98], stage0_28[99], stage0_28[100], stage0_28[101]},
      {stage0_30[85], stage0_30[86], stage0_30[87], stage0_30[88], stage0_30[89], stage0_30[90]},
      {stage1_32[15],stage1_31[22],stage1_30[22],stage1_29[42],stage1_28[67]}
   );
   gpc606_5 gpc376 (
      {stage0_28[102], stage0_28[103], stage0_28[104], stage0_28[105], stage0_28[106], stage0_28[107]},
      {stage0_30[91], stage0_30[92], stage0_30[93], stage0_30[94], stage0_30[95], stage0_30[96]},
      {stage1_32[16],stage1_31[23],stage1_30[23],stage1_29[43],stage1_28[68]}
   );
   gpc606_5 gpc377 (
      {stage0_28[108], stage0_28[109], stage0_28[110], stage0_28[111], stage0_28[112], stage0_28[113]},
      {stage0_30[97], stage0_30[98], stage0_30[99], stage0_30[100], stage0_30[101], stage0_30[102]},
      {stage1_32[17],stage1_31[24],stage1_30[24],stage1_29[44],stage1_28[69]}
   );
   gpc606_5 gpc378 (
      {stage0_28[114], stage0_28[115], stage0_28[116], stage0_28[117], stage0_28[118], stage0_28[119]},
      {stage0_30[103], stage0_30[104], stage0_30[105], stage0_30[106], stage0_30[107], stage0_30[108]},
      {stage1_32[18],stage1_31[25],stage1_30[25],stage1_29[45],stage1_28[70]}
   );
   gpc606_5 gpc379 (
      {stage0_28[120], stage0_28[121], stage0_28[122], stage0_28[123], stage0_28[124], stage0_28[125]},
      {stage0_30[109], stage0_30[110], stage0_30[111], stage0_30[112], stage0_30[113], stage0_30[114]},
      {stage1_32[19],stage1_31[26],stage1_30[26],stage1_29[46],stage1_28[71]}
   );
   gpc606_5 gpc380 (
      {stage0_28[126], stage0_28[127], stage0_28[128], stage0_28[129], stage0_28[130], stage0_28[131]},
      {stage0_30[115], stage0_30[116], stage0_30[117], stage0_30[118], stage0_30[119], stage0_30[120]},
      {stage1_32[20],stage1_31[27],stage1_30[27],stage1_29[47],stage1_28[72]}
   );
   gpc606_5 gpc381 (
      {stage0_28[132], stage0_28[133], stage0_28[134], stage0_28[135], stage0_28[136], stage0_28[137]},
      {stage0_30[121], stage0_30[122], stage0_30[123], stage0_30[124], stage0_30[125], stage0_30[126]},
      {stage1_32[21],stage1_31[28],stage1_30[28],stage1_29[48],stage1_28[73]}
   );
   gpc606_5 gpc382 (
      {stage0_28[138], stage0_28[139], stage0_28[140], stage0_28[141], stage0_28[142], stage0_28[143]},
      {stage0_30[127], stage0_30[128], stage0_30[129], stage0_30[130], stage0_30[131], stage0_30[132]},
      {stage1_32[22],stage1_31[29],stage1_30[29],stage1_29[49],stage1_28[74]}
   );
   gpc606_5 gpc383 (
      {stage0_28[144], stage0_28[145], stage0_28[146], stage0_28[147], stage0_28[148], stage0_28[149]},
      {stage0_30[133], stage0_30[134], stage0_30[135], stage0_30[136], stage0_30[137], stage0_30[138]},
      {stage1_32[23],stage1_31[30],stage1_30[30],stage1_29[50],stage1_28[75]}
   );
   gpc606_5 gpc384 (
      {stage0_28[150], stage0_28[151], stage0_28[152], stage0_28[153], stage0_28[154], stage0_28[155]},
      {stage0_30[139], stage0_30[140], stage0_30[141], stage0_30[142], stage0_30[143], stage0_30[144]},
      {stage1_32[24],stage1_31[31],stage1_30[31],stage1_29[51],stage1_28[76]}
   );
   gpc606_5 gpc385 (
      {stage0_28[156], stage0_28[157], stage0_28[158], stage0_28[159], stage0_28[160], stage0_28[161]},
      {stage0_30[145], stage0_30[146], stage0_30[147], stage0_30[148], stage0_30[149], stage0_30[150]},
      {stage1_32[25],stage1_31[32],stage1_30[32],stage1_29[52],stage1_28[77]}
   );
   gpc606_5 gpc386 (
      {stage0_29[45], stage0_29[46], stage0_29[47], stage0_29[48], stage0_29[49], stage0_29[50]},
      {stage0_31[2], stage0_31[3], stage0_31[4], stage0_31[5], stage0_31[6], stage0_31[7]},
      {stage1_33[0],stage1_32[26],stage1_31[33],stage1_30[33],stage1_29[53]}
   );
   gpc606_5 gpc387 (
      {stage0_29[51], stage0_29[52], stage0_29[53], stage0_29[54], stage0_29[55], stage0_29[56]},
      {stage0_31[8], stage0_31[9], stage0_31[10], stage0_31[11], stage0_31[12], stage0_31[13]},
      {stage1_33[1],stage1_32[27],stage1_31[34],stage1_30[34],stage1_29[54]}
   );
   gpc606_5 gpc388 (
      {stage0_29[57], stage0_29[58], stage0_29[59], stage0_29[60], stage0_29[61], stage0_29[62]},
      {stage0_31[14], stage0_31[15], stage0_31[16], stage0_31[17], stage0_31[18], stage0_31[19]},
      {stage1_33[2],stage1_32[28],stage1_31[35],stage1_30[35],stage1_29[55]}
   );
   gpc606_5 gpc389 (
      {stage0_29[63], stage0_29[64], stage0_29[65], stage0_29[66], stage0_29[67], stage0_29[68]},
      {stage0_31[20], stage0_31[21], stage0_31[22], stage0_31[23], stage0_31[24], stage0_31[25]},
      {stage1_33[3],stage1_32[29],stage1_31[36],stage1_30[36],stage1_29[56]}
   );
   gpc606_5 gpc390 (
      {stage0_29[69], stage0_29[70], stage0_29[71], stage0_29[72], stage0_29[73], stage0_29[74]},
      {stage0_31[26], stage0_31[27], stage0_31[28], stage0_31[29], stage0_31[30], stage0_31[31]},
      {stage1_33[4],stage1_32[30],stage1_31[37],stage1_30[37],stage1_29[57]}
   );
   gpc606_5 gpc391 (
      {stage0_29[75], stage0_29[76], stage0_29[77], stage0_29[78], stage0_29[79], stage0_29[80]},
      {stage0_31[32], stage0_31[33], stage0_31[34], stage0_31[35], stage0_31[36], stage0_31[37]},
      {stage1_33[5],stage1_32[31],stage1_31[38],stage1_30[38],stage1_29[58]}
   );
   gpc606_5 gpc392 (
      {stage0_29[81], stage0_29[82], stage0_29[83], stage0_29[84], stage0_29[85], stage0_29[86]},
      {stage0_31[38], stage0_31[39], stage0_31[40], stage0_31[41], stage0_31[42], stage0_31[43]},
      {stage1_33[6],stage1_32[32],stage1_31[39],stage1_30[39],stage1_29[59]}
   );
   gpc606_5 gpc393 (
      {stage0_29[87], stage0_29[88], stage0_29[89], stage0_29[90], stage0_29[91], stage0_29[92]},
      {stage0_31[44], stage0_31[45], stage0_31[46], stage0_31[47], stage0_31[48], stage0_31[49]},
      {stage1_33[7],stage1_32[33],stage1_31[40],stage1_30[40],stage1_29[60]}
   );
   gpc606_5 gpc394 (
      {stage0_29[93], stage0_29[94], stage0_29[95], stage0_29[96], stage0_29[97], stage0_29[98]},
      {stage0_31[50], stage0_31[51], stage0_31[52], stage0_31[53], stage0_31[54], stage0_31[55]},
      {stage1_33[8],stage1_32[34],stage1_31[41],stage1_30[41],stage1_29[61]}
   );
   gpc606_5 gpc395 (
      {stage0_29[99], stage0_29[100], stage0_29[101], stage0_29[102], stage0_29[103], stage0_29[104]},
      {stage0_31[56], stage0_31[57], stage0_31[58], stage0_31[59], stage0_31[60], stage0_31[61]},
      {stage1_33[9],stage1_32[35],stage1_31[42],stage1_30[42],stage1_29[62]}
   );
   gpc606_5 gpc396 (
      {stage0_29[105], stage0_29[106], stage0_29[107], stage0_29[108], stage0_29[109], stage0_29[110]},
      {stage0_31[62], stage0_31[63], stage0_31[64], stage0_31[65], stage0_31[66], stage0_31[67]},
      {stage1_33[10],stage1_32[36],stage1_31[43],stage1_30[43],stage1_29[63]}
   );
   gpc606_5 gpc397 (
      {stage0_29[111], stage0_29[112], stage0_29[113], stage0_29[114], stage0_29[115], stage0_29[116]},
      {stage0_31[68], stage0_31[69], stage0_31[70], stage0_31[71], stage0_31[72], stage0_31[73]},
      {stage1_33[11],stage1_32[37],stage1_31[44],stage1_30[44],stage1_29[64]}
   );
   gpc606_5 gpc398 (
      {stage0_29[117], stage0_29[118], stage0_29[119], stage0_29[120], stage0_29[121], stage0_29[122]},
      {stage0_31[74], stage0_31[75], stage0_31[76], stage0_31[77], stage0_31[78], stage0_31[79]},
      {stage1_33[12],stage1_32[38],stage1_31[45],stage1_30[45],stage1_29[65]}
   );
   gpc606_5 gpc399 (
      {stage0_29[123], stage0_29[124], stage0_29[125], stage0_29[126], stage0_29[127], stage0_29[128]},
      {stage0_31[80], stage0_31[81], stage0_31[82], stage0_31[83], stage0_31[84], stage0_31[85]},
      {stage1_33[13],stage1_32[39],stage1_31[46],stage1_30[46],stage1_29[66]}
   );
   gpc606_5 gpc400 (
      {stage0_29[129], stage0_29[130], stage0_29[131], stage0_29[132], stage0_29[133], stage0_29[134]},
      {stage0_31[86], stage0_31[87], stage0_31[88], stage0_31[89], stage0_31[90], stage0_31[91]},
      {stage1_33[14],stage1_32[40],stage1_31[47],stage1_30[47],stage1_29[67]}
   );
   gpc606_5 gpc401 (
      {stage0_29[135], stage0_29[136], stage0_29[137], stage0_29[138], stage0_29[139], stage0_29[140]},
      {stage0_31[92], stage0_31[93], stage0_31[94], stage0_31[95], stage0_31[96], stage0_31[97]},
      {stage1_33[15],stage1_32[41],stage1_31[48],stage1_30[48],stage1_29[68]}
   );
   gpc606_5 gpc402 (
      {stage0_29[141], stage0_29[142], stage0_29[143], stage0_29[144], stage0_29[145], stage0_29[146]},
      {stage0_31[98], stage0_31[99], stage0_31[100], stage0_31[101], stage0_31[102], stage0_31[103]},
      {stage1_33[16],stage1_32[42],stage1_31[49],stage1_30[49],stage1_29[69]}
   );
   gpc606_5 gpc403 (
      {stage0_29[147], stage0_29[148], stage0_29[149], stage0_29[150], stage0_29[151], stage0_29[152]},
      {stage0_31[104], stage0_31[105], stage0_31[106], stage0_31[107], stage0_31[108], stage0_31[109]},
      {stage1_33[17],stage1_32[43],stage1_31[50],stage1_30[50],stage1_29[70]}
   );
   gpc606_5 gpc404 (
      {stage0_29[153], stage0_29[154], stage0_29[155], stage0_29[156], stage0_29[157], stage0_29[158]},
      {stage0_31[110], stage0_31[111], stage0_31[112], stage0_31[113], stage0_31[114], stage0_31[115]},
      {stage1_33[18],stage1_32[44],stage1_31[51],stage1_30[51],stage1_29[71]}
   );
   gpc1_1 gpc405 (
      {stage0_0[144]},
      {stage1_0[32]}
   );
   gpc1_1 gpc406 (
      {stage0_0[145]},
      {stage1_0[33]}
   );
   gpc1_1 gpc407 (
      {stage0_0[146]},
      {stage1_0[34]}
   );
   gpc1_1 gpc408 (
      {stage0_0[147]},
      {stage1_0[35]}
   );
   gpc1_1 gpc409 (
      {stage0_0[148]},
      {stage1_0[36]}
   );
   gpc1_1 gpc410 (
      {stage0_0[149]},
      {stage1_0[37]}
   );
   gpc1_1 gpc411 (
      {stage0_0[150]},
      {stage1_0[38]}
   );
   gpc1_1 gpc412 (
      {stage0_0[151]},
      {stage1_0[39]}
   );
   gpc1_1 gpc413 (
      {stage0_0[152]},
      {stage1_0[40]}
   );
   gpc1_1 gpc414 (
      {stage0_0[153]},
      {stage1_0[41]}
   );
   gpc1_1 gpc415 (
      {stage0_0[154]},
      {stage1_0[42]}
   );
   gpc1_1 gpc416 (
      {stage0_0[155]},
      {stage1_0[43]}
   );
   gpc1_1 gpc417 (
      {stage0_0[156]},
      {stage1_0[44]}
   );
   gpc1_1 gpc418 (
      {stage0_0[157]},
      {stage1_0[45]}
   );
   gpc1_1 gpc419 (
      {stage0_0[158]},
      {stage1_0[46]}
   );
   gpc1_1 gpc420 (
      {stage0_0[159]},
      {stage1_0[47]}
   );
   gpc1_1 gpc421 (
      {stage0_0[160]},
      {stage1_0[48]}
   );
   gpc1_1 gpc422 (
      {stage0_0[161]},
      {stage1_0[49]}
   );
   gpc1_1 gpc423 (
      {stage0_1[144]},
      {stage1_1[38]}
   );
   gpc1_1 gpc424 (
      {stage0_1[145]},
      {stage1_1[39]}
   );
   gpc1_1 gpc425 (
      {stage0_1[146]},
      {stage1_1[40]}
   );
   gpc1_1 gpc426 (
      {stage0_1[147]},
      {stage1_1[41]}
   );
   gpc1_1 gpc427 (
      {stage0_1[148]},
      {stage1_1[42]}
   );
   gpc1_1 gpc428 (
      {stage0_1[149]},
      {stage1_1[43]}
   );
   gpc1_1 gpc429 (
      {stage0_1[150]},
      {stage1_1[44]}
   );
   gpc1_1 gpc430 (
      {stage0_1[151]},
      {stage1_1[45]}
   );
   gpc1_1 gpc431 (
      {stage0_1[152]},
      {stage1_1[46]}
   );
   gpc1_1 gpc432 (
      {stage0_1[153]},
      {stage1_1[47]}
   );
   gpc1_1 gpc433 (
      {stage0_1[154]},
      {stage1_1[48]}
   );
   gpc1_1 gpc434 (
      {stage0_1[155]},
      {stage1_1[49]}
   );
   gpc1_1 gpc435 (
      {stage0_1[156]},
      {stage1_1[50]}
   );
   gpc1_1 gpc436 (
      {stage0_1[157]},
      {stage1_1[51]}
   );
   gpc1_1 gpc437 (
      {stage0_1[158]},
      {stage1_1[52]}
   );
   gpc1_1 gpc438 (
      {stage0_1[159]},
      {stage1_1[53]}
   );
   gpc1_1 gpc439 (
      {stage0_1[160]},
      {stage1_1[54]}
   );
   gpc1_1 gpc440 (
      {stage0_1[161]},
      {stage1_1[55]}
   );
   gpc1_1 gpc441 (
      {stage0_3[155]},
      {stage1_3[69]}
   );
   gpc1_1 gpc442 (
      {stage0_3[156]},
      {stage1_3[70]}
   );
   gpc1_1 gpc443 (
      {stage0_3[157]},
      {stage1_3[71]}
   );
   gpc1_1 gpc444 (
      {stage0_3[158]},
      {stage1_3[72]}
   );
   gpc1_1 gpc445 (
      {stage0_3[159]},
      {stage1_3[73]}
   );
   gpc1_1 gpc446 (
      {stage0_3[160]},
      {stage1_3[74]}
   );
   gpc1_1 gpc447 (
      {stage0_3[161]},
      {stage1_3[75]}
   );
   gpc1_1 gpc448 (
      {stage0_4[139]},
      {stage1_4[72]}
   );
   gpc1_1 gpc449 (
      {stage0_4[140]},
      {stage1_4[73]}
   );
   gpc1_1 gpc450 (
      {stage0_4[141]},
      {stage1_4[74]}
   );
   gpc1_1 gpc451 (
      {stage0_4[142]},
      {stage1_4[75]}
   );
   gpc1_1 gpc452 (
      {stage0_4[143]},
      {stage1_4[76]}
   );
   gpc1_1 gpc453 (
      {stage0_4[144]},
      {stage1_4[77]}
   );
   gpc1_1 gpc454 (
      {stage0_4[145]},
      {stage1_4[78]}
   );
   gpc1_1 gpc455 (
      {stage0_4[146]},
      {stage1_4[79]}
   );
   gpc1_1 gpc456 (
      {stage0_4[147]},
      {stage1_4[80]}
   );
   gpc1_1 gpc457 (
      {stage0_4[148]},
      {stage1_4[81]}
   );
   gpc1_1 gpc458 (
      {stage0_4[149]},
      {stage1_4[82]}
   );
   gpc1_1 gpc459 (
      {stage0_4[150]},
      {stage1_4[83]}
   );
   gpc1_1 gpc460 (
      {stage0_4[151]},
      {stage1_4[84]}
   );
   gpc1_1 gpc461 (
      {stage0_4[152]},
      {stage1_4[85]}
   );
   gpc1_1 gpc462 (
      {stage0_4[153]},
      {stage1_4[86]}
   );
   gpc1_1 gpc463 (
      {stage0_4[154]},
      {stage1_4[87]}
   );
   gpc1_1 gpc464 (
      {stage0_4[155]},
      {stage1_4[88]}
   );
   gpc1_1 gpc465 (
      {stage0_4[156]},
      {stage1_4[89]}
   );
   gpc1_1 gpc466 (
      {stage0_4[157]},
      {stage1_4[90]}
   );
   gpc1_1 gpc467 (
      {stage0_4[158]},
      {stage1_4[91]}
   );
   gpc1_1 gpc468 (
      {stage0_4[159]},
      {stage1_4[92]}
   );
   gpc1_1 gpc469 (
      {stage0_4[160]},
      {stage1_4[93]}
   );
   gpc1_1 gpc470 (
      {stage0_4[161]},
      {stage1_4[94]}
   );
   gpc1_1 gpc471 (
      {stage0_6[124]},
      {stage1_6[68]}
   );
   gpc1_1 gpc472 (
      {stage0_6[125]},
      {stage1_6[69]}
   );
   gpc1_1 gpc473 (
      {stage0_6[126]},
      {stage1_6[70]}
   );
   gpc1_1 gpc474 (
      {stage0_6[127]},
      {stage1_6[71]}
   );
   gpc1_1 gpc475 (
      {stage0_6[128]},
      {stage1_6[72]}
   );
   gpc1_1 gpc476 (
      {stage0_6[129]},
      {stage1_6[73]}
   );
   gpc1_1 gpc477 (
      {stage0_6[130]},
      {stage1_6[74]}
   );
   gpc1_1 gpc478 (
      {stage0_6[131]},
      {stage1_6[75]}
   );
   gpc1_1 gpc479 (
      {stage0_6[132]},
      {stage1_6[76]}
   );
   gpc1_1 gpc480 (
      {stage0_6[133]},
      {stage1_6[77]}
   );
   gpc1_1 gpc481 (
      {stage0_6[134]},
      {stage1_6[78]}
   );
   gpc1_1 gpc482 (
      {stage0_6[135]},
      {stage1_6[79]}
   );
   gpc1_1 gpc483 (
      {stage0_6[136]},
      {stage1_6[80]}
   );
   gpc1_1 gpc484 (
      {stage0_6[137]},
      {stage1_6[81]}
   );
   gpc1_1 gpc485 (
      {stage0_6[138]},
      {stage1_6[82]}
   );
   gpc1_1 gpc486 (
      {stage0_6[139]},
      {stage1_6[83]}
   );
   gpc1_1 gpc487 (
      {stage0_6[140]},
      {stage1_6[84]}
   );
   gpc1_1 gpc488 (
      {stage0_6[141]},
      {stage1_6[85]}
   );
   gpc1_1 gpc489 (
      {stage0_6[142]},
      {stage1_6[86]}
   );
   gpc1_1 gpc490 (
      {stage0_6[143]},
      {stage1_6[87]}
   );
   gpc1_1 gpc491 (
      {stage0_6[144]},
      {stage1_6[88]}
   );
   gpc1_1 gpc492 (
      {stage0_6[145]},
      {stage1_6[89]}
   );
   gpc1_1 gpc493 (
      {stage0_6[146]},
      {stage1_6[90]}
   );
   gpc1_1 gpc494 (
      {stage0_6[147]},
      {stage1_6[91]}
   );
   gpc1_1 gpc495 (
      {stage0_6[148]},
      {stage1_6[92]}
   );
   gpc1_1 gpc496 (
      {stage0_6[149]},
      {stage1_6[93]}
   );
   gpc1_1 gpc497 (
      {stage0_6[150]},
      {stage1_6[94]}
   );
   gpc1_1 gpc498 (
      {stage0_6[151]},
      {stage1_6[95]}
   );
   gpc1_1 gpc499 (
      {stage0_6[152]},
      {stage1_6[96]}
   );
   gpc1_1 gpc500 (
      {stage0_6[153]},
      {stage1_6[97]}
   );
   gpc1_1 gpc501 (
      {stage0_6[154]},
      {stage1_6[98]}
   );
   gpc1_1 gpc502 (
      {stage0_6[155]},
      {stage1_6[99]}
   );
   gpc1_1 gpc503 (
      {stage0_6[156]},
      {stage1_6[100]}
   );
   gpc1_1 gpc504 (
      {stage0_6[157]},
      {stage1_6[101]}
   );
   gpc1_1 gpc505 (
      {stage0_6[158]},
      {stage1_6[102]}
   );
   gpc1_1 gpc506 (
      {stage0_6[159]},
      {stage1_6[103]}
   );
   gpc1_1 gpc507 (
      {stage0_6[160]},
      {stage1_6[104]}
   );
   gpc1_1 gpc508 (
      {stage0_6[161]},
      {stage1_6[105]}
   );
   gpc1_1 gpc509 (
      {stage0_7[158]},
      {stage1_7[62]}
   );
   gpc1_1 gpc510 (
      {stage0_7[159]},
      {stage1_7[63]}
   );
   gpc1_1 gpc511 (
      {stage0_7[160]},
      {stage1_7[64]}
   );
   gpc1_1 gpc512 (
      {stage0_7[161]},
      {stage1_7[65]}
   );
   gpc1_1 gpc513 (
      {stage0_9[152]},
      {stage1_9[67]}
   );
   gpc1_1 gpc514 (
      {stage0_9[153]},
      {stage1_9[68]}
   );
   gpc1_1 gpc515 (
      {stage0_9[154]},
      {stage1_9[69]}
   );
   gpc1_1 gpc516 (
      {stage0_9[155]},
      {stage1_9[70]}
   );
   gpc1_1 gpc517 (
      {stage0_9[156]},
      {stage1_9[71]}
   );
   gpc1_1 gpc518 (
      {stage0_9[157]},
      {stage1_9[72]}
   );
   gpc1_1 gpc519 (
      {stage0_9[158]},
      {stage1_9[73]}
   );
   gpc1_1 gpc520 (
      {stage0_9[159]},
      {stage1_9[74]}
   );
   gpc1_1 gpc521 (
      {stage0_9[160]},
      {stage1_9[75]}
   );
   gpc1_1 gpc522 (
      {stage0_9[161]},
      {stage1_9[76]}
   );
   gpc1_1 gpc523 (
      {stage0_10[141]},
      {stage1_10[72]}
   );
   gpc1_1 gpc524 (
      {stage0_10[142]},
      {stage1_10[73]}
   );
   gpc1_1 gpc525 (
      {stage0_10[143]},
      {stage1_10[74]}
   );
   gpc1_1 gpc526 (
      {stage0_10[144]},
      {stage1_10[75]}
   );
   gpc1_1 gpc527 (
      {stage0_10[145]},
      {stage1_10[76]}
   );
   gpc1_1 gpc528 (
      {stage0_10[146]},
      {stage1_10[77]}
   );
   gpc1_1 gpc529 (
      {stage0_10[147]},
      {stage1_10[78]}
   );
   gpc1_1 gpc530 (
      {stage0_10[148]},
      {stage1_10[79]}
   );
   gpc1_1 gpc531 (
      {stage0_10[149]},
      {stage1_10[80]}
   );
   gpc1_1 gpc532 (
      {stage0_10[150]},
      {stage1_10[81]}
   );
   gpc1_1 gpc533 (
      {stage0_10[151]},
      {stage1_10[82]}
   );
   gpc1_1 gpc534 (
      {stage0_10[152]},
      {stage1_10[83]}
   );
   gpc1_1 gpc535 (
      {stage0_10[153]},
      {stage1_10[84]}
   );
   gpc1_1 gpc536 (
      {stage0_10[154]},
      {stage1_10[85]}
   );
   gpc1_1 gpc537 (
      {stage0_10[155]},
      {stage1_10[86]}
   );
   gpc1_1 gpc538 (
      {stage0_10[156]},
      {stage1_10[87]}
   );
   gpc1_1 gpc539 (
      {stage0_10[157]},
      {stage1_10[88]}
   );
   gpc1_1 gpc540 (
      {stage0_10[158]},
      {stage1_10[89]}
   );
   gpc1_1 gpc541 (
      {stage0_10[159]},
      {stage1_10[90]}
   );
   gpc1_1 gpc542 (
      {stage0_10[160]},
      {stage1_10[91]}
   );
   gpc1_1 gpc543 (
      {stage0_10[161]},
      {stage1_10[92]}
   );
   gpc1_1 gpc544 (
      {stage0_11[155]},
      {stage1_11[60]}
   );
   gpc1_1 gpc545 (
      {stage0_11[156]},
      {stage1_11[61]}
   );
   gpc1_1 gpc546 (
      {stage0_11[157]},
      {stage1_11[62]}
   );
   gpc1_1 gpc547 (
      {stage0_11[158]},
      {stage1_11[63]}
   );
   gpc1_1 gpc548 (
      {stage0_11[159]},
      {stage1_11[64]}
   );
   gpc1_1 gpc549 (
      {stage0_11[160]},
      {stage1_11[65]}
   );
   gpc1_1 gpc550 (
      {stage0_11[161]},
      {stage1_11[66]}
   );
   gpc1_1 gpc551 (
      {stage0_13[144]},
      {stage1_13[68]}
   );
   gpc1_1 gpc552 (
      {stage0_13[145]},
      {stage1_13[69]}
   );
   gpc1_1 gpc553 (
      {stage0_13[146]},
      {stage1_13[70]}
   );
   gpc1_1 gpc554 (
      {stage0_13[147]},
      {stage1_13[71]}
   );
   gpc1_1 gpc555 (
      {stage0_13[148]},
      {stage1_13[72]}
   );
   gpc1_1 gpc556 (
      {stage0_13[149]},
      {stage1_13[73]}
   );
   gpc1_1 gpc557 (
      {stage0_13[150]},
      {stage1_13[74]}
   );
   gpc1_1 gpc558 (
      {stage0_13[151]},
      {stage1_13[75]}
   );
   gpc1_1 gpc559 (
      {stage0_13[152]},
      {stage1_13[76]}
   );
   gpc1_1 gpc560 (
      {stage0_13[153]},
      {stage1_13[77]}
   );
   gpc1_1 gpc561 (
      {stage0_13[154]},
      {stage1_13[78]}
   );
   gpc1_1 gpc562 (
      {stage0_13[155]},
      {stage1_13[79]}
   );
   gpc1_1 gpc563 (
      {stage0_13[156]},
      {stage1_13[80]}
   );
   gpc1_1 gpc564 (
      {stage0_13[157]},
      {stage1_13[81]}
   );
   gpc1_1 gpc565 (
      {stage0_13[158]},
      {stage1_13[82]}
   );
   gpc1_1 gpc566 (
      {stage0_13[159]},
      {stage1_13[83]}
   );
   gpc1_1 gpc567 (
      {stage0_13[160]},
      {stage1_13[84]}
   );
   gpc1_1 gpc568 (
      {stage0_13[161]},
      {stage1_13[85]}
   );
   gpc1_1 gpc569 (
      {stage0_14[161]},
      {stage1_14[68]}
   );
   gpc1_1 gpc570 (
      {stage0_16[111]},
      {stage1_16[56]}
   );
   gpc1_1 gpc571 (
      {stage0_16[112]},
      {stage1_16[57]}
   );
   gpc1_1 gpc572 (
      {stage0_16[113]},
      {stage1_16[58]}
   );
   gpc1_1 gpc573 (
      {stage0_16[114]},
      {stage1_16[59]}
   );
   gpc1_1 gpc574 (
      {stage0_16[115]},
      {stage1_16[60]}
   );
   gpc1_1 gpc575 (
      {stage0_16[116]},
      {stage1_16[61]}
   );
   gpc1_1 gpc576 (
      {stage0_16[117]},
      {stage1_16[62]}
   );
   gpc1_1 gpc577 (
      {stage0_16[118]},
      {stage1_16[63]}
   );
   gpc1_1 gpc578 (
      {stage0_16[119]},
      {stage1_16[64]}
   );
   gpc1_1 gpc579 (
      {stage0_16[120]},
      {stage1_16[65]}
   );
   gpc1_1 gpc580 (
      {stage0_16[121]},
      {stage1_16[66]}
   );
   gpc1_1 gpc581 (
      {stage0_16[122]},
      {stage1_16[67]}
   );
   gpc1_1 gpc582 (
      {stage0_16[123]},
      {stage1_16[68]}
   );
   gpc1_1 gpc583 (
      {stage0_16[124]},
      {stage1_16[69]}
   );
   gpc1_1 gpc584 (
      {stage0_16[125]},
      {stage1_16[70]}
   );
   gpc1_1 gpc585 (
      {stage0_16[126]},
      {stage1_16[71]}
   );
   gpc1_1 gpc586 (
      {stage0_16[127]},
      {stage1_16[72]}
   );
   gpc1_1 gpc587 (
      {stage0_16[128]},
      {stage1_16[73]}
   );
   gpc1_1 gpc588 (
      {stage0_16[129]},
      {stage1_16[74]}
   );
   gpc1_1 gpc589 (
      {stage0_16[130]},
      {stage1_16[75]}
   );
   gpc1_1 gpc590 (
      {stage0_16[131]},
      {stage1_16[76]}
   );
   gpc1_1 gpc591 (
      {stage0_16[132]},
      {stage1_16[77]}
   );
   gpc1_1 gpc592 (
      {stage0_16[133]},
      {stage1_16[78]}
   );
   gpc1_1 gpc593 (
      {stage0_16[134]},
      {stage1_16[79]}
   );
   gpc1_1 gpc594 (
      {stage0_16[135]},
      {stage1_16[80]}
   );
   gpc1_1 gpc595 (
      {stage0_16[136]},
      {stage1_16[81]}
   );
   gpc1_1 gpc596 (
      {stage0_16[137]},
      {stage1_16[82]}
   );
   gpc1_1 gpc597 (
      {stage0_16[138]},
      {stage1_16[83]}
   );
   gpc1_1 gpc598 (
      {stage0_16[139]},
      {stage1_16[84]}
   );
   gpc1_1 gpc599 (
      {stage0_16[140]},
      {stage1_16[85]}
   );
   gpc1_1 gpc600 (
      {stage0_16[141]},
      {stage1_16[86]}
   );
   gpc1_1 gpc601 (
      {stage0_16[142]},
      {stage1_16[87]}
   );
   gpc1_1 gpc602 (
      {stage0_16[143]},
      {stage1_16[88]}
   );
   gpc1_1 gpc603 (
      {stage0_16[144]},
      {stage1_16[89]}
   );
   gpc1_1 gpc604 (
      {stage0_16[145]},
      {stage1_16[90]}
   );
   gpc1_1 gpc605 (
      {stage0_16[146]},
      {stage1_16[91]}
   );
   gpc1_1 gpc606 (
      {stage0_16[147]},
      {stage1_16[92]}
   );
   gpc1_1 gpc607 (
      {stage0_16[148]},
      {stage1_16[93]}
   );
   gpc1_1 gpc608 (
      {stage0_16[149]},
      {stage1_16[94]}
   );
   gpc1_1 gpc609 (
      {stage0_16[150]},
      {stage1_16[95]}
   );
   gpc1_1 gpc610 (
      {stage0_16[151]},
      {stage1_16[96]}
   );
   gpc1_1 gpc611 (
      {stage0_16[152]},
      {stage1_16[97]}
   );
   gpc1_1 gpc612 (
      {stage0_16[153]},
      {stage1_16[98]}
   );
   gpc1_1 gpc613 (
      {stage0_16[154]},
      {stage1_16[99]}
   );
   gpc1_1 gpc614 (
      {stage0_16[155]},
      {stage1_16[100]}
   );
   gpc1_1 gpc615 (
      {stage0_16[156]},
      {stage1_16[101]}
   );
   gpc1_1 gpc616 (
      {stage0_16[157]},
      {stage1_16[102]}
   );
   gpc1_1 gpc617 (
      {stage0_16[158]},
      {stage1_16[103]}
   );
   gpc1_1 gpc618 (
      {stage0_16[159]},
      {stage1_16[104]}
   );
   gpc1_1 gpc619 (
      {stage0_16[160]},
      {stage1_16[105]}
   );
   gpc1_1 gpc620 (
      {stage0_16[161]},
      {stage1_16[106]}
   );
   gpc1_1 gpc621 (
      {stage0_18[142]},
      {stage1_18[62]}
   );
   gpc1_1 gpc622 (
      {stage0_18[143]},
      {stage1_18[63]}
   );
   gpc1_1 gpc623 (
      {stage0_18[144]},
      {stage1_18[64]}
   );
   gpc1_1 gpc624 (
      {stage0_18[145]},
      {stage1_18[65]}
   );
   gpc1_1 gpc625 (
      {stage0_18[146]},
      {stage1_18[66]}
   );
   gpc1_1 gpc626 (
      {stage0_18[147]},
      {stage1_18[67]}
   );
   gpc1_1 gpc627 (
      {stage0_18[148]},
      {stage1_18[68]}
   );
   gpc1_1 gpc628 (
      {stage0_18[149]},
      {stage1_18[69]}
   );
   gpc1_1 gpc629 (
      {stage0_18[150]},
      {stage1_18[70]}
   );
   gpc1_1 gpc630 (
      {stage0_18[151]},
      {stage1_18[71]}
   );
   gpc1_1 gpc631 (
      {stage0_18[152]},
      {stage1_18[72]}
   );
   gpc1_1 gpc632 (
      {stage0_18[153]},
      {stage1_18[73]}
   );
   gpc1_1 gpc633 (
      {stage0_18[154]},
      {stage1_18[74]}
   );
   gpc1_1 gpc634 (
      {stage0_18[155]},
      {stage1_18[75]}
   );
   gpc1_1 gpc635 (
      {stage0_18[156]},
      {stage1_18[76]}
   );
   gpc1_1 gpc636 (
      {stage0_18[157]},
      {stage1_18[77]}
   );
   gpc1_1 gpc637 (
      {stage0_18[158]},
      {stage1_18[78]}
   );
   gpc1_1 gpc638 (
      {stage0_18[159]},
      {stage1_18[79]}
   );
   gpc1_1 gpc639 (
      {stage0_18[160]},
      {stage1_18[80]}
   );
   gpc1_1 gpc640 (
      {stage0_18[161]},
      {stage1_18[81]}
   );
   gpc1_1 gpc641 (
      {stage0_19[154]},
      {stage1_19[59]}
   );
   gpc1_1 gpc642 (
      {stage0_19[155]},
      {stage1_19[60]}
   );
   gpc1_1 gpc643 (
      {stage0_19[156]},
      {stage1_19[61]}
   );
   gpc1_1 gpc644 (
      {stage0_19[157]},
      {stage1_19[62]}
   );
   gpc1_1 gpc645 (
      {stage0_19[158]},
      {stage1_19[63]}
   );
   gpc1_1 gpc646 (
      {stage0_19[159]},
      {stage1_19[64]}
   );
   gpc1_1 gpc647 (
      {stage0_19[160]},
      {stage1_19[65]}
   );
   gpc1_1 gpc648 (
      {stage0_19[161]},
      {stage1_19[66]}
   );
   gpc1_1 gpc649 (
      {stage0_21[160]},
      {stage1_21[78]}
   );
   gpc1_1 gpc650 (
      {stage0_21[161]},
      {stage1_21[79]}
   );
   gpc1_1 gpc651 (
      {stage0_22[138]},
      {stage1_22[58]}
   );
   gpc1_1 gpc652 (
      {stage0_22[139]},
      {stage1_22[59]}
   );
   gpc1_1 gpc653 (
      {stage0_22[140]},
      {stage1_22[60]}
   );
   gpc1_1 gpc654 (
      {stage0_22[141]},
      {stage1_22[61]}
   );
   gpc1_1 gpc655 (
      {stage0_22[142]},
      {stage1_22[62]}
   );
   gpc1_1 gpc656 (
      {stage0_22[143]},
      {stage1_22[63]}
   );
   gpc1_1 gpc657 (
      {stage0_22[144]},
      {stage1_22[64]}
   );
   gpc1_1 gpc658 (
      {stage0_22[145]},
      {stage1_22[65]}
   );
   gpc1_1 gpc659 (
      {stage0_22[146]},
      {stage1_22[66]}
   );
   gpc1_1 gpc660 (
      {stage0_22[147]},
      {stage1_22[67]}
   );
   gpc1_1 gpc661 (
      {stage0_22[148]},
      {stage1_22[68]}
   );
   gpc1_1 gpc662 (
      {stage0_22[149]},
      {stage1_22[69]}
   );
   gpc1_1 gpc663 (
      {stage0_22[150]},
      {stage1_22[70]}
   );
   gpc1_1 gpc664 (
      {stage0_22[151]},
      {stage1_22[71]}
   );
   gpc1_1 gpc665 (
      {stage0_22[152]},
      {stage1_22[72]}
   );
   gpc1_1 gpc666 (
      {stage0_22[153]},
      {stage1_22[73]}
   );
   gpc1_1 gpc667 (
      {stage0_22[154]},
      {stage1_22[74]}
   );
   gpc1_1 gpc668 (
      {stage0_22[155]},
      {stage1_22[75]}
   );
   gpc1_1 gpc669 (
      {stage0_22[156]},
      {stage1_22[76]}
   );
   gpc1_1 gpc670 (
      {stage0_22[157]},
      {stage1_22[77]}
   );
   gpc1_1 gpc671 (
      {stage0_22[158]},
      {stage1_22[78]}
   );
   gpc1_1 gpc672 (
      {stage0_22[159]},
      {stage1_22[79]}
   );
   gpc1_1 gpc673 (
      {stage0_22[160]},
      {stage1_22[80]}
   );
   gpc1_1 gpc674 (
      {stage0_22[161]},
      {stage1_22[81]}
   );
   gpc1_1 gpc675 (
      {stage0_23[122]},
      {stage1_23[51]}
   );
   gpc1_1 gpc676 (
      {stage0_23[123]},
      {stage1_23[52]}
   );
   gpc1_1 gpc677 (
      {stage0_23[124]},
      {stage1_23[53]}
   );
   gpc1_1 gpc678 (
      {stage0_23[125]},
      {stage1_23[54]}
   );
   gpc1_1 gpc679 (
      {stage0_23[126]},
      {stage1_23[55]}
   );
   gpc1_1 gpc680 (
      {stage0_23[127]},
      {stage1_23[56]}
   );
   gpc1_1 gpc681 (
      {stage0_23[128]},
      {stage1_23[57]}
   );
   gpc1_1 gpc682 (
      {stage0_23[129]},
      {stage1_23[58]}
   );
   gpc1_1 gpc683 (
      {stage0_23[130]},
      {stage1_23[59]}
   );
   gpc1_1 gpc684 (
      {stage0_23[131]},
      {stage1_23[60]}
   );
   gpc1_1 gpc685 (
      {stage0_23[132]},
      {stage1_23[61]}
   );
   gpc1_1 gpc686 (
      {stage0_23[133]},
      {stage1_23[62]}
   );
   gpc1_1 gpc687 (
      {stage0_23[134]},
      {stage1_23[63]}
   );
   gpc1_1 gpc688 (
      {stage0_23[135]},
      {stage1_23[64]}
   );
   gpc1_1 gpc689 (
      {stage0_23[136]},
      {stage1_23[65]}
   );
   gpc1_1 gpc690 (
      {stage0_23[137]},
      {stage1_23[66]}
   );
   gpc1_1 gpc691 (
      {stage0_23[138]},
      {stage1_23[67]}
   );
   gpc1_1 gpc692 (
      {stage0_23[139]},
      {stage1_23[68]}
   );
   gpc1_1 gpc693 (
      {stage0_23[140]},
      {stage1_23[69]}
   );
   gpc1_1 gpc694 (
      {stage0_23[141]},
      {stage1_23[70]}
   );
   gpc1_1 gpc695 (
      {stage0_23[142]},
      {stage1_23[71]}
   );
   gpc1_1 gpc696 (
      {stage0_23[143]},
      {stage1_23[72]}
   );
   gpc1_1 gpc697 (
      {stage0_23[144]},
      {stage1_23[73]}
   );
   gpc1_1 gpc698 (
      {stage0_23[145]},
      {stage1_23[74]}
   );
   gpc1_1 gpc699 (
      {stage0_23[146]},
      {stage1_23[75]}
   );
   gpc1_1 gpc700 (
      {stage0_23[147]},
      {stage1_23[76]}
   );
   gpc1_1 gpc701 (
      {stage0_23[148]},
      {stage1_23[77]}
   );
   gpc1_1 gpc702 (
      {stage0_23[149]},
      {stage1_23[78]}
   );
   gpc1_1 gpc703 (
      {stage0_23[150]},
      {stage1_23[79]}
   );
   gpc1_1 gpc704 (
      {stage0_23[151]},
      {stage1_23[80]}
   );
   gpc1_1 gpc705 (
      {stage0_23[152]},
      {stage1_23[81]}
   );
   gpc1_1 gpc706 (
      {stage0_23[153]},
      {stage1_23[82]}
   );
   gpc1_1 gpc707 (
      {stage0_23[154]},
      {stage1_23[83]}
   );
   gpc1_1 gpc708 (
      {stage0_23[155]},
      {stage1_23[84]}
   );
   gpc1_1 gpc709 (
      {stage0_23[156]},
      {stage1_23[85]}
   );
   gpc1_1 gpc710 (
      {stage0_23[157]},
      {stage1_23[86]}
   );
   gpc1_1 gpc711 (
      {stage0_23[158]},
      {stage1_23[87]}
   );
   gpc1_1 gpc712 (
      {stage0_23[159]},
      {stage1_23[88]}
   );
   gpc1_1 gpc713 (
      {stage0_23[160]},
      {stage1_23[89]}
   );
   gpc1_1 gpc714 (
      {stage0_23[161]},
      {stage1_23[90]}
   );
   gpc1_1 gpc715 (
      {stage0_25[158]},
      {stage1_25[74]}
   );
   gpc1_1 gpc716 (
      {stage0_25[159]},
      {stage1_25[75]}
   );
   gpc1_1 gpc717 (
      {stage0_25[160]},
      {stage1_25[76]}
   );
   gpc1_1 gpc718 (
      {stage0_25[161]},
      {stage1_25[77]}
   );
   gpc1_1 gpc719 (
      {stage0_26[160]},
      {stage1_26[53]}
   );
   gpc1_1 gpc720 (
      {stage0_26[161]},
      {stage1_26[54]}
   );
   gpc1_1 gpc721 (
      {stage0_27[155]},
      {stage1_27[60]}
   );
   gpc1_1 gpc722 (
      {stage0_27[156]},
      {stage1_27[61]}
   );
   gpc1_1 gpc723 (
      {stage0_27[157]},
      {stage1_27[62]}
   );
   gpc1_1 gpc724 (
      {stage0_27[158]},
      {stage1_27[63]}
   );
   gpc1_1 gpc725 (
      {stage0_27[159]},
      {stage1_27[64]}
   );
   gpc1_1 gpc726 (
      {stage0_27[160]},
      {stage1_27[65]}
   );
   gpc1_1 gpc727 (
      {stage0_27[161]},
      {stage1_27[66]}
   );
   gpc1_1 gpc728 (
      {stage0_29[159]},
      {stage1_29[72]}
   );
   gpc1_1 gpc729 (
      {stage0_29[160]},
      {stage1_29[73]}
   );
   gpc1_1 gpc730 (
      {stage0_29[161]},
      {stage1_29[74]}
   );
   gpc1_1 gpc731 (
      {stage0_30[151]},
      {stage1_30[52]}
   );
   gpc1_1 gpc732 (
      {stage0_30[152]},
      {stage1_30[53]}
   );
   gpc1_1 gpc733 (
      {stage0_30[153]},
      {stage1_30[54]}
   );
   gpc1_1 gpc734 (
      {stage0_30[154]},
      {stage1_30[55]}
   );
   gpc1_1 gpc735 (
      {stage0_30[155]},
      {stage1_30[56]}
   );
   gpc1_1 gpc736 (
      {stage0_30[156]},
      {stage1_30[57]}
   );
   gpc1_1 gpc737 (
      {stage0_30[157]},
      {stage1_30[58]}
   );
   gpc1_1 gpc738 (
      {stage0_30[158]},
      {stage1_30[59]}
   );
   gpc1_1 gpc739 (
      {stage0_30[159]},
      {stage1_30[60]}
   );
   gpc1_1 gpc740 (
      {stage0_30[160]},
      {stage1_30[61]}
   );
   gpc1_1 gpc741 (
      {stage0_30[161]},
      {stage1_30[62]}
   );
   gpc1_1 gpc742 (
      {stage0_31[116]},
      {stage1_31[52]}
   );
   gpc1_1 gpc743 (
      {stage0_31[117]},
      {stage1_31[53]}
   );
   gpc1_1 gpc744 (
      {stage0_31[118]},
      {stage1_31[54]}
   );
   gpc1_1 gpc745 (
      {stage0_31[119]},
      {stage1_31[55]}
   );
   gpc1_1 gpc746 (
      {stage0_31[120]},
      {stage1_31[56]}
   );
   gpc1_1 gpc747 (
      {stage0_31[121]},
      {stage1_31[57]}
   );
   gpc1_1 gpc748 (
      {stage0_31[122]},
      {stage1_31[58]}
   );
   gpc1_1 gpc749 (
      {stage0_31[123]},
      {stage1_31[59]}
   );
   gpc1_1 gpc750 (
      {stage0_31[124]},
      {stage1_31[60]}
   );
   gpc1_1 gpc751 (
      {stage0_31[125]},
      {stage1_31[61]}
   );
   gpc1_1 gpc752 (
      {stage0_31[126]},
      {stage1_31[62]}
   );
   gpc1_1 gpc753 (
      {stage0_31[127]},
      {stage1_31[63]}
   );
   gpc1_1 gpc754 (
      {stage0_31[128]},
      {stage1_31[64]}
   );
   gpc1_1 gpc755 (
      {stage0_31[129]},
      {stage1_31[65]}
   );
   gpc1_1 gpc756 (
      {stage0_31[130]},
      {stage1_31[66]}
   );
   gpc1_1 gpc757 (
      {stage0_31[131]},
      {stage1_31[67]}
   );
   gpc1_1 gpc758 (
      {stage0_31[132]},
      {stage1_31[68]}
   );
   gpc1_1 gpc759 (
      {stage0_31[133]},
      {stage1_31[69]}
   );
   gpc1_1 gpc760 (
      {stage0_31[134]},
      {stage1_31[70]}
   );
   gpc1_1 gpc761 (
      {stage0_31[135]},
      {stage1_31[71]}
   );
   gpc1_1 gpc762 (
      {stage0_31[136]},
      {stage1_31[72]}
   );
   gpc1_1 gpc763 (
      {stage0_31[137]},
      {stage1_31[73]}
   );
   gpc1_1 gpc764 (
      {stage0_31[138]},
      {stage1_31[74]}
   );
   gpc1_1 gpc765 (
      {stage0_31[139]},
      {stage1_31[75]}
   );
   gpc1_1 gpc766 (
      {stage0_31[140]},
      {stage1_31[76]}
   );
   gpc1_1 gpc767 (
      {stage0_31[141]},
      {stage1_31[77]}
   );
   gpc1_1 gpc768 (
      {stage0_31[142]},
      {stage1_31[78]}
   );
   gpc1_1 gpc769 (
      {stage0_31[143]},
      {stage1_31[79]}
   );
   gpc1_1 gpc770 (
      {stage0_31[144]},
      {stage1_31[80]}
   );
   gpc1_1 gpc771 (
      {stage0_31[145]},
      {stage1_31[81]}
   );
   gpc1_1 gpc772 (
      {stage0_31[146]},
      {stage1_31[82]}
   );
   gpc1_1 gpc773 (
      {stage0_31[147]},
      {stage1_31[83]}
   );
   gpc1_1 gpc774 (
      {stage0_31[148]},
      {stage1_31[84]}
   );
   gpc1_1 gpc775 (
      {stage0_31[149]},
      {stage1_31[85]}
   );
   gpc1_1 gpc776 (
      {stage0_31[150]},
      {stage1_31[86]}
   );
   gpc1_1 gpc777 (
      {stage0_31[151]},
      {stage1_31[87]}
   );
   gpc1_1 gpc778 (
      {stage0_31[152]},
      {stage1_31[88]}
   );
   gpc1_1 gpc779 (
      {stage0_31[153]},
      {stage1_31[89]}
   );
   gpc1_1 gpc780 (
      {stage0_31[154]},
      {stage1_31[90]}
   );
   gpc1_1 gpc781 (
      {stage0_31[155]},
      {stage1_31[91]}
   );
   gpc1_1 gpc782 (
      {stage0_31[156]},
      {stage1_31[92]}
   );
   gpc1_1 gpc783 (
      {stage0_31[157]},
      {stage1_31[93]}
   );
   gpc1_1 gpc784 (
      {stage0_31[158]},
      {stage1_31[94]}
   );
   gpc1_1 gpc785 (
      {stage0_31[159]},
      {stage1_31[95]}
   );
   gpc1_1 gpc786 (
      {stage0_31[160]},
      {stage1_31[96]}
   );
   gpc1_1 gpc787 (
      {stage0_31[161]},
      {stage1_31[97]}
   );
   gpc1163_5 gpc788 (
      {stage1_0[0], stage1_0[1], stage1_0[2]},
      {stage1_1[0], stage1_1[1], stage1_1[2], stage1_1[3], stage1_1[4], stage1_1[5]},
      {stage1_2[0]},
      {stage1_3[0]},
      {stage2_4[0],stage2_3[0],stage2_2[0],stage2_1[0],stage2_0[0]}
   );
   gpc1163_5 gpc789 (
      {stage1_0[3], stage1_0[4], stage1_0[5]},
      {stage1_1[6], stage1_1[7], stage1_1[8], stage1_1[9], stage1_1[10], stage1_1[11]},
      {stage1_2[1]},
      {stage1_3[1]},
      {stage2_4[1],stage2_3[1],stage2_2[1],stage2_1[1],stage2_0[1]}
   );
   gpc1163_5 gpc790 (
      {stage1_0[6], stage1_0[7], stage1_0[8]},
      {stage1_1[12], stage1_1[13], stage1_1[14], stage1_1[15], stage1_1[16], stage1_1[17]},
      {stage1_2[2]},
      {stage1_3[2]},
      {stage2_4[2],stage2_3[2],stage2_2[2],stage2_1[2],stage2_0[2]}
   );
   gpc606_5 gpc791 (
      {stage1_0[9], stage1_0[10], stage1_0[11], stage1_0[12], stage1_0[13], stage1_0[14]},
      {stage1_2[3], stage1_2[4], stage1_2[5], stage1_2[6], stage1_2[7], stage1_2[8]},
      {stage2_4[3],stage2_3[3],stage2_2[3],stage2_1[3],stage2_0[3]}
   );
   gpc615_5 gpc792 (
      {stage1_0[15], stage1_0[16], stage1_0[17], stage1_0[18], stage1_0[19]},
      {stage1_1[18]},
      {stage1_2[9], stage1_2[10], stage1_2[11], stage1_2[12], stage1_2[13], stage1_2[14]},
      {stage2_4[4],stage2_3[4],stage2_2[4],stage2_1[4],stage2_0[4]}
   );
   gpc615_5 gpc793 (
      {stage1_0[20], stage1_0[21], stage1_0[22], stage1_0[23], stage1_0[24]},
      {stage1_1[19]},
      {stage1_2[15], stage1_2[16], stage1_2[17], stage1_2[18], stage1_2[19], stage1_2[20]},
      {stage2_4[5],stage2_3[5],stage2_2[5],stage2_1[5],stage2_0[5]}
   );
   gpc615_5 gpc794 (
      {stage1_0[25], stage1_0[26], stage1_0[27], stage1_0[28], stage1_0[29]},
      {stage1_1[20]},
      {stage1_2[21], stage1_2[22], stage1_2[23], stage1_2[24], stage1_2[25], stage1_2[26]},
      {stage2_4[6],stage2_3[6],stage2_2[6],stage2_1[6],stage2_0[6]}
   );
   gpc615_5 gpc795 (
      {stage1_0[30], stage1_0[31], stage1_0[32], stage1_0[33], stage1_0[34]},
      {stage1_1[21]},
      {stage1_2[27], stage1_2[28], stage1_2[29], stage1_2[30], stage1_2[31], stage1_2[32]},
      {stage2_4[7],stage2_3[7],stage2_2[7],stage2_1[7],stage2_0[7]}
   );
   gpc615_5 gpc796 (
      {stage1_0[35], stage1_0[36], stage1_0[37], stage1_0[38], stage1_0[39]},
      {stage1_1[22]},
      {stage1_2[33], stage1_2[34], stage1_2[35], stage1_2[36], stage1_2[37], stage1_2[38]},
      {stage2_4[8],stage2_3[8],stage2_2[8],stage2_1[8],stage2_0[8]}
   );
   gpc615_5 gpc797 (
      {stage1_0[40], stage1_0[41], stage1_0[42], stage1_0[43], stage1_0[44]},
      {stage1_1[23]},
      {stage1_2[39], stage1_2[40], stage1_2[41], stage1_2[42], stage1_2[43], stage1_2[44]},
      {stage2_4[9],stage2_3[9],stage2_2[9],stage2_1[9],stage2_0[9]}
   );
   gpc615_5 gpc798 (
      {stage1_0[45], stage1_0[46], stage1_0[47], stage1_0[48], stage1_0[49]},
      {stage1_1[24]},
      {stage1_2[45], stage1_2[46], stage1_2[47], stage1_2[48], stage1_2[49], stage1_2[50]},
      {stage2_4[10],stage2_3[10],stage2_2[10],stage2_1[10],stage2_0[10]}
   );
   gpc606_5 gpc799 (
      {stage1_1[25], stage1_1[26], stage1_1[27], stage1_1[28], stage1_1[29], stage1_1[30]},
      {stage1_3[3], stage1_3[4], stage1_3[5], stage1_3[6], stage1_3[7], stage1_3[8]},
      {stage2_5[0],stage2_4[11],stage2_3[11],stage2_2[11],stage2_1[11]}
   );
   gpc606_5 gpc800 (
      {stage1_1[31], stage1_1[32], stage1_1[33], stage1_1[34], stage1_1[35], stage1_1[36]},
      {stage1_3[9], stage1_3[10], stage1_3[11], stage1_3[12], stage1_3[13], stage1_3[14]},
      {stage2_5[1],stage2_4[12],stage2_3[12],stage2_2[12],stage2_1[12]}
   );
   gpc606_5 gpc801 (
      {stage1_1[37], stage1_1[38], stage1_1[39], stage1_1[40], stage1_1[41], stage1_1[42]},
      {stage1_3[15], stage1_3[16], stage1_3[17], stage1_3[18], stage1_3[19], stage1_3[20]},
      {stage2_5[2],stage2_4[13],stage2_3[13],stage2_2[13],stage2_1[13]}
   );
   gpc606_5 gpc802 (
      {stage1_1[43], stage1_1[44], stage1_1[45], stage1_1[46], stage1_1[47], stage1_1[48]},
      {stage1_3[21], stage1_3[22], stage1_3[23], stage1_3[24], stage1_3[25], stage1_3[26]},
      {stage2_5[3],stage2_4[14],stage2_3[14],stage2_2[14],stage2_1[14]}
   );
   gpc606_5 gpc803 (
      {stage1_1[49], stage1_1[50], stage1_1[51], stage1_1[52], stage1_1[53], stage1_1[54]},
      {stage1_3[27], stage1_3[28], stage1_3[29], stage1_3[30], stage1_3[31], stage1_3[32]},
      {stage2_5[4],stage2_4[15],stage2_3[15],stage2_2[15],stage2_1[15]}
   );
   gpc615_5 gpc804 (
      {stage1_2[51], stage1_2[52], stage1_2[53], stage1_2[54], stage1_2[55]},
      {stage1_3[33]},
      {stage1_4[0], stage1_4[1], stage1_4[2], stage1_4[3], stage1_4[4], stage1_4[5]},
      {stage2_6[0],stage2_5[5],stage2_4[16],stage2_3[16],stage2_2[16]}
   );
   gpc615_5 gpc805 (
      {stage1_3[34], stage1_3[35], stage1_3[36], stage1_3[37], stage1_3[38]},
      {stage1_4[6]},
      {stage1_5[0], stage1_5[1], stage1_5[2], stage1_5[3], stage1_5[4], stage1_5[5]},
      {stage2_7[0],stage2_6[1],stage2_5[6],stage2_4[17],stage2_3[17]}
   );
   gpc615_5 gpc806 (
      {stage1_3[39], stage1_3[40], stage1_3[41], stage1_3[42], stage1_3[43]},
      {stage1_4[7]},
      {stage1_5[6], stage1_5[7], stage1_5[8], stage1_5[9], stage1_5[10], stage1_5[11]},
      {stage2_7[1],stage2_6[2],stage2_5[7],stage2_4[18],stage2_3[18]}
   );
   gpc615_5 gpc807 (
      {stage1_3[44], stage1_3[45], stage1_3[46], stage1_3[47], stage1_3[48]},
      {stage1_4[8]},
      {stage1_5[12], stage1_5[13], stage1_5[14], stage1_5[15], stage1_5[16], stage1_5[17]},
      {stage2_7[2],stage2_6[3],stage2_5[8],stage2_4[19],stage2_3[19]}
   );
   gpc615_5 gpc808 (
      {stage1_3[49], stage1_3[50], stage1_3[51], stage1_3[52], stage1_3[53]},
      {stage1_4[9]},
      {stage1_5[18], stage1_5[19], stage1_5[20], stage1_5[21], stage1_5[22], stage1_5[23]},
      {stage2_7[3],stage2_6[4],stage2_5[9],stage2_4[20],stage2_3[20]}
   );
   gpc615_5 gpc809 (
      {stage1_3[54], stage1_3[55], stage1_3[56], stage1_3[57], stage1_3[58]},
      {stage1_4[10]},
      {stage1_5[24], stage1_5[25], stage1_5[26], stage1_5[27], stage1_5[28], stage1_5[29]},
      {stage2_7[4],stage2_6[5],stage2_5[10],stage2_4[21],stage2_3[21]}
   );
   gpc615_5 gpc810 (
      {stage1_3[59], stage1_3[60], stage1_3[61], stage1_3[62], stage1_3[63]},
      {stage1_4[11]},
      {stage1_5[30], stage1_5[31], stage1_5[32], stage1_5[33], stage1_5[34], stage1_5[35]},
      {stage2_7[5],stage2_6[6],stage2_5[11],stage2_4[22],stage2_3[22]}
   );
   gpc606_5 gpc811 (
      {stage1_4[12], stage1_4[13], stage1_4[14], stage1_4[15], stage1_4[16], stage1_4[17]},
      {stage1_6[0], stage1_6[1], stage1_6[2], stage1_6[3], stage1_6[4], stage1_6[5]},
      {stage2_8[0],stage2_7[6],stage2_6[7],stage2_5[12],stage2_4[23]}
   );
   gpc606_5 gpc812 (
      {stage1_4[18], stage1_4[19], stage1_4[20], stage1_4[21], stage1_4[22], stage1_4[23]},
      {stage1_6[6], stage1_6[7], stage1_6[8], stage1_6[9], stage1_6[10], stage1_6[11]},
      {stage2_8[1],stage2_7[7],stage2_6[8],stage2_5[13],stage2_4[24]}
   );
   gpc606_5 gpc813 (
      {stage1_4[24], stage1_4[25], stage1_4[26], stage1_4[27], stage1_4[28], stage1_4[29]},
      {stage1_6[12], stage1_6[13], stage1_6[14], stage1_6[15], stage1_6[16], stage1_6[17]},
      {stage2_8[2],stage2_7[8],stage2_6[9],stage2_5[14],stage2_4[25]}
   );
   gpc606_5 gpc814 (
      {stage1_4[30], stage1_4[31], stage1_4[32], stage1_4[33], stage1_4[34], stage1_4[35]},
      {stage1_6[18], stage1_6[19], stage1_6[20], stage1_6[21], stage1_6[22], stage1_6[23]},
      {stage2_8[3],stage2_7[9],stage2_6[10],stage2_5[15],stage2_4[26]}
   );
   gpc606_5 gpc815 (
      {stage1_4[36], stage1_4[37], stage1_4[38], stage1_4[39], stage1_4[40], stage1_4[41]},
      {stage1_6[24], stage1_6[25], stage1_6[26], stage1_6[27], stage1_6[28], stage1_6[29]},
      {stage2_8[4],stage2_7[10],stage2_6[11],stage2_5[16],stage2_4[27]}
   );
   gpc606_5 gpc816 (
      {stage1_4[42], stage1_4[43], stage1_4[44], stage1_4[45], stage1_4[46], stage1_4[47]},
      {stage1_6[30], stage1_6[31], stage1_6[32], stage1_6[33], stage1_6[34], stage1_6[35]},
      {stage2_8[5],stage2_7[11],stage2_6[12],stage2_5[17],stage2_4[28]}
   );
   gpc606_5 gpc817 (
      {stage1_4[48], stage1_4[49], stage1_4[50], stage1_4[51], stage1_4[52], stage1_4[53]},
      {stage1_6[36], stage1_6[37], stage1_6[38], stage1_6[39], stage1_6[40], stage1_6[41]},
      {stage2_8[6],stage2_7[12],stage2_6[13],stage2_5[18],stage2_4[29]}
   );
   gpc606_5 gpc818 (
      {stage1_4[54], stage1_4[55], stage1_4[56], stage1_4[57], stage1_4[58], stage1_4[59]},
      {stage1_6[42], stage1_6[43], stage1_6[44], stage1_6[45], stage1_6[46], stage1_6[47]},
      {stage2_8[7],stage2_7[13],stage2_6[14],stage2_5[19],stage2_4[30]}
   );
   gpc606_5 gpc819 (
      {stage1_4[60], stage1_4[61], stage1_4[62], stage1_4[63], stage1_4[64], stage1_4[65]},
      {stage1_6[48], stage1_6[49], stage1_6[50], stage1_6[51], stage1_6[52], stage1_6[53]},
      {stage2_8[8],stage2_7[14],stage2_6[15],stage2_5[20],stage2_4[31]}
   );
   gpc606_5 gpc820 (
      {stage1_4[66], stage1_4[67], stage1_4[68], stage1_4[69], stage1_4[70], stage1_4[71]},
      {stage1_6[54], stage1_6[55], stage1_6[56], stage1_6[57], stage1_6[58], stage1_6[59]},
      {stage2_8[9],stage2_7[15],stage2_6[16],stage2_5[21],stage2_4[32]}
   );
   gpc606_5 gpc821 (
      {stage1_4[72], stage1_4[73], stage1_4[74], stage1_4[75], stage1_4[76], stage1_4[77]},
      {stage1_6[60], stage1_6[61], stage1_6[62], stage1_6[63], stage1_6[64], stage1_6[65]},
      {stage2_8[10],stage2_7[16],stage2_6[17],stage2_5[22],stage2_4[33]}
   );
   gpc606_5 gpc822 (
      {stage1_4[78], stage1_4[79], stage1_4[80], stage1_4[81], stage1_4[82], stage1_4[83]},
      {stage1_6[66], stage1_6[67], stage1_6[68], stage1_6[69], stage1_6[70], stage1_6[71]},
      {stage2_8[11],stage2_7[17],stage2_6[18],stage2_5[23],stage2_4[34]}
   );
   gpc606_5 gpc823 (
      {stage1_4[84], stage1_4[85], stage1_4[86], stage1_4[87], stage1_4[88], stage1_4[89]},
      {stage1_6[72], stage1_6[73], stage1_6[74], stage1_6[75], stage1_6[76], stage1_6[77]},
      {stage2_8[12],stage2_7[18],stage2_6[19],stage2_5[24],stage2_4[35]}
   );
   gpc606_5 gpc824 (
      {stage1_5[36], stage1_5[37], stage1_5[38], stage1_5[39], stage1_5[40], stage1_5[41]},
      {stage1_7[0], stage1_7[1], stage1_7[2], stage1_7[3], stage1_7[4], stage1_7[5]},
      {stage2_9[0],stage2_8[13],stage2_7[19],stage2_6[20],stage2_5[25]}
   );
   gpc606_5 gpc825 (
      {stage1_5[42], stage1_5[43], stage1_5[44], stage1_5[45], stage1_5[46], stage1_5[47]},
      {stage1_7[6], stage1_7[7], stage1_7[8], stage1_7[9], stage1_7[10], stage1_7[11]},
      {stage2_9[1],stage2_8[14],stage2_7[20],stage2_6[21],stage2_5[26]}
   );
   gpc606_5 gpc826 (
      {stage1_5[48], stage1_5[49], stage1_5[50], stage1_5[51], stage1_5[52], stage1_5[53]},
      {stage1_7[12], stage1_7[13], stage1_7[14], stage1_7[15], stage1_7[16], stage1_7[17]},
      {stage2_9[2],stage2_8[15],stage2_7[21],stage2_6[22],stage2_5[27]}
   );
   gpc606_5 gpc827 (
      {stage1_6[78], stage1_6[79], stage1_6[80], stage1_6[81], stage1_6[82], stage1_6[83]},
      {stage1_8[0], stage1_8[1], stage1_8[2], stage1_8[3], stage1_8[4], stage1_8[5]},
      {stage2_10[0],stage2_9[3],stage2_8[16],stage2_7[22],stage2_6[23]}
   );
   gpc606_5 gpc828 (
      {stage1_6[84], stage1_6[85], stage1_6[86], stage1_6[87], stage1_6[88], stage1_6[89]},
      {stage1_8[6], stage1_8[7], stage1_8[8], stage1_8[9], stage1_8[10], stage1_8[11]},
      {stage2_10[1],stage2_9[4],stage2_8[17],stage2_7[23],stage2_6[24]}
   );
   gpc606_5 gpc829 (
      {stage1_6[90], stage1_6[91], stage1_6[92], stage1_6[93], stage1_6[94], stage1_6[95]},
      {stage1_8[12], stage1_8[13], stage1_8[14], stage1_8[15], stage1_8[16], stage1_8[17]},
      {stage2_10[2],stage2_9[5],stage2_8[18],stage2_7[24],stage2_6[25]}
   );
   gpc606_5 gpc830 (
      {stage1_6[96], stage1_6[97], stage1_6[98], stage1_6[99], stage1_6[100], stage1_6[101]},
      {stage1_8[18], stage1_8[19], stage1_8[20], stage1_8[21], stage1_8[22], stage1_8[23]},
      {stage2_10[3],stage2_9[6],stage2_8[19],stage2_7[25],stage2_6[26]}
   );
   gpc606_5 gpc831 (
      {stage1_7[18], stage1_7[19], stage1_7[20], stage1_7[21], stage1_7[22], stage1_7[23]},
      {stage1_9[0], stage1_9[1], stage1_9[2], stage1_9[3], stage1_9[4], stage1_9[5]},
      {stage2_11[0],stage2_10[4],stage2_9[7],stage2_8[20],stage2_7[26]}
   );
   gpc606_5 gpc832 (
      {stage1_7[24], stage1_7[25], stage1_7[26], stage1_7[27], stage1_7[28], stage1_7[29]},
      {stage1_9[6], stage1_9[7], stage1_9[8], stage1_9[9], stage1_9[10], stage1_9[11]},
      {stage2_11[1],stage2_10[5],stage2_9[8],stage2_8[21],stage2_7[27]}
   );
   gpc606_5 gpc833 (
      {stage1_7[30], stage1_7[31], stage1_7[32], stage1_7[33], stage1_7[34], stage1_7[35]},
      {stage1_9[12], stage1_9[13], stage1_9[14], stage1_9[15], stage1_9[16], stage1_9[17]},
      {stage2_11[2],stage2_10[6],stage2_9[9],stage2_8[22],stage2_7[28]}
   );
   gpc606_5 gpc834 (
      {stage1_7[36], stage1_7[37], stage1_7[38], stage1_7[39], stage1_7[40], stage1_7[41]},
      {stage1_9[18], stage1_9[19], stage1_9[20], stage1_9[21], stage1_9[22], stage1_9[23]},
      {stage2_11[3],stage2_10[7],stage2_9[10],stage2_8[23],stage2_7[29]}
   );
   gpc606_5 gpc835 (
      {stage1_7[42], stage1_7[43], stage1_7[44], stage1_7[45], stage1_7[46], stage1_7[47]},
      {stage1_9[24], stage1_9[25], stage1_9[26], stage1_9[27], stage1_9[28], stage1_9[29]},
      {stage2_11[4],stage2_10[8],stage2_9[11],stage2_8[24],stage2_7[30]}
   );
   gpc606_5 gpc836 (
      {stage1_7[48], stage1_7[49], stage1_7[50], stage1_7[51], stage1_7[52], stage1_7[53]},
      {stage1_9[30], stage1_9[31], stage1_9[32], stage1_9[33], stage1_9[34], stage1_9[35]},
      {stage2_11[5],stage2_10[9],stage2_9[12],stage2_8[25],stage2_7[31]}
   );
   gpc606_5 gpc837 (
      {stage1_7[54], stage1_7[55], stage1_7[56], stage1_7[57], stage1_7[58], stage1_7[59]},
      {stage1_9[36], stage1_9[37], stage1_9[38], stage1_9[39], stage1_9[40], stage1_9[41]},
      {stage2_11[6],stage2_10[10],stage2_9[13],stage2_8[26],stage2_7[32]}
   );
   gpc606_5 gpc838 (
      {stage1_7[60], stage1_7[61], stage1_7[62], stage1_7[63], stage1_7[64], stage1_7[65]},
      {stage1_9[42], stage1_9[43], stage1_9[44], stage1_9[45], stage1_9[46], stage1_9[47]},
      {stage2_11[7],stage2_10[11],stage2_9[14],stage2_8[27],stage2_7[33]}
   );
   gpc606_5 gpc839 (
      {stage1_8[24], stage1_8[25], stage1_8[26], stage1_8[27], stage1_8[28], stage1_8[29]},
      {stage1_10[0], stage1_10[1], stage1_10[2], stage1_10[3], stage1_10[4], stage1_10[5]},
      {stage2_12[0],stage2_11[8],stage2_10[12],stage2_9[15],stage2_8[28]}
   );
   gpc606_5 gpc840 (
      {stage1_8[30], stage1_8[31], stage1_8[32], stage1_8[33], stage1_8[34], stage1_8[35]},
      {stage1_10[6], stage1_10[7], stage1_10[8], stage1_10[9], stage1_10[10], stage1_10[11]},
      {stage2_12[1],stage2_11[9],stage2_10[13],stage2_9[16],stage2_8[29]}
   );
   gpc606_5 gpc841 (
      {stage1_8[36], stage1_8[37], stage1_8[38], stage1_8[39], stage1_8[40], stage1_8[41]},
      {stage1_10[12], stage1_10[13], stage1_10[14], stage1_10[15], stage1_10[16], stage1_10[17]},
      {stage2_12[2],stage2_11[10],stage2_10[14],stage2_9[17],stage2_8[30]}
   );
   gpc606_5 gpc842 (
      {stage1_8[42], stage1_8[43], stage1_8[44], stage1_8[45], stage1_8[46], stage1_8[47]},
      {stage1_10[18], stage1_10[19], stage1_10[20], stage1_10[21], stage1_10[22], stage1_10[23]},
      {stage2_12[3],stage2_11[11],stage2_10[15],stage2_9[18],stage2_8[31]}
   );
   gpc606_5 gpc843 (
      {stage1_8[48], stage1_8[49], stage1_8[50], stage1_8[51], stage1_8[52], stage1_8[53]},
      {stage1_10[24], stage1_10[25], stage1_10[26], stage1_10[27], stage1_10[28], stage1_10[29]},
      {stage2_12[4],stage2_11[12],stage2_10[16],stage2_9[19],stage2_8[32]}
   );
   gpc606_5 gpc844 (
      {stage1_9[48], stage1_9[49], stage1_9[50], stage1_9[51], stage1_9[52], stage1_9[53]},
      {stage1_11[0], stage1_11[1], stage1_11[2], stage1_11[3], stage1_11[4], stage1_11[5]},
      {stage2_13[0],stage2_12[5],stage2_11[13],stage2_10[17],stage2_9[20]}
   );
   gpc615_5 gpc845 (
      {stage1_9[54], stage1_9[55], stage1_9[56], stage1_9[57], stage1_9[58]},
      {stage1_10[30]},
      {stage1_11[6], stage1_11[7], stage1_11[8], stage1_11[9], stage1_11[10], stage1_11[11]},
      {stage2_13[1],stage2_12[6],stage2_11[14],stage2_10[18],stage2_9[21]}
   );
   gpc615_5 gpc846 (
      {stage1_9[59], stage1_9[60], stage1_9[61], stage1_9[62], stage1_9[63]},
      {stage1_10[31]},
      {stage1_11[12], stage1_11[13], stage1_11[14], stage1_11[15], stage1_11[16], stage1_11[17]},
      {stage2_13[2],stage2_12[7],stage2_11[15],stage2_10[19],stage2_9[22]}
   );
   gpc615_5 gpc847 (
      {stage1_9[64], stage1_9[65], stage1_9[66], stage1_9[67], stage1_9[68]},
      {stage1_10[32]},
      {stage1_11[18], stage1_11[19], stage1_11[20], stage1_11[21], stage1_11[22], stage1_11[23]},
      {stage2_13[3],stage2_12[8],stage2_11[16],stage2_10[20],stage2_9[23]}
   );
   gpc606_5 gpc848 (
      {stage1_10[33], stage1_10[34], stage1_10[35], stage1_10[36], stage1_10[37], stage1_10[38]},
      {stage1_12[0], stage1_12[1], stage1_12[2], stage1_12[3], stage1_12[4], stage1_12[5]},
      {stage2_14[0],stage2_13[4],stage2_12[9],stage2_11[17],stage2_10[21]}
   );
   gpc606_5 gpc849 (
      {stage1_10[39], stage1_10[40], stage1_10[41], stage1_10[42], stage1_10[43], stage1_10[44]},
      {stage1_12[6], stage1_12[7], stage1_12[8], stage1_12[9], stage1_12[10], stage1_12[11]},
      {stage2_14[1],stage2_13[5],stage2_12[10],stage2_11[18],stage2_10[22]}
   );
   gpc606_5 gpc850 (
      {stage1_10[45], stage1_10[46], stage1_10[47], stage1_10[48], stage1_10[49], stage1_10[50]},
      {stage1_12[12], stage1_12[13], stage1_12[14], stage1_12[15], stage1_12[16], stage1_12[17]},
      {stage2_14[2],stage2_13[6],stage2_12[11],stage2_11[19],stage2_10[23]}
   );
   gpc606_5 gpc851 (
      {stage1_10[51], stage1_10[52], stage1_10[53], stage1_10[54], stage1_10[55], stage1_10[56]},
      {stage1_12[18], stage1_12[19], stage1_12[20], stage1_12[21], stage1_12[22], stage1_12[23]},
      {stage2_14[3],stage2_13[7],stage2_12[12],stage2_11[20],stage2_10[24]}
   );
   gpc606_5 gpc852 (
      {stage1_10[57], stage1_10[58], stage1_10[59], stage1_10[60], stage1_10[61], stage1_10[62]},
      {stage1_12[24], stage1_12[25], stage1_12[26], stage1_12[27], stage1_12[28], stage1_12[29]},
      {stage2_14[4],stage2_13[8],stage2_12[13],stage2_11[21],stage2_10[25]}
   );
   gpc606_5 gpc853 (
      {stage1_10[63], stage1_10[64], stage1_10[65], stage1_10[66], stage1_10[67], stage1_10[68]},
      {stage1_12[30], stage1_12[31], stage1_12[32], stage1_12[33], stage1_12[34], stage1_12[35]},
      {stage2_14[5],stage2_13[9],stage2_12[14],stage2_11[22],stage2_10[26]}
   );
   gpc606_5 gpc854 (
      {stage1_10[69], stage1_10[70], stage1_10[71], stage1_10[72], stage1_10[73], stage1_10[74]},
      {stage1_12[36], stage1_12[37], stage1_12[38], stage1_12[39], stage1_12[40], stage1_12[41]},
      {stage2_14[6],stage2_13[10],stage2_12[15],stage2_11[23],stage2_10[27]}
   );
   gpc606_5 gpc855 (
      {stage1_11[24], stage1_11[25], stage1_11[26], stage1_11[27], stage1_11[28], stage1_11[29]},
      {stage1_13[0], stage1_13[1], stage1_13[2], stage1_13[3], stage1_13[4], stage1_13[5]},
      {stage2_15[0],stage2_14[7],stage2_13[11],stage2_12[16],stage2_11[24]}
   );
   gpc606_5 gpc856 (
      {stage1_11[30], stage1_11[31], stage1_11[32], stage1_11[33], stage1_11[34], stage1_11[35]},
      {stage1_13[6], stage1_13[7], stage1_13[8], stage1_13[9], stage1_13[10], stage1_13[11]},
      {stage2_15[1],stage2_14[8],stage2_13[12],stage2_12[17],stage2_11[25]}
   );
   gpc606_5 gpc857 (
      {stage1_11[36], stage1_11[37], stage1_11[38], stage1_11[39], stage1_11[40], stage1_11[41]},
      {stage1_13[12], stage1_13[13], stage1_13[14], stage1_13[15], stage1_13[16], stage1_13[17]},
      {stage2_15[2],stage2_14[9],stage2_13[13],stage2_12[18],stage2_11[26]}
   );
   gpc606_5 gpc858 (
      {stage1_11[42], stage1_11[43], stage1_11[44], stage1_11[45], stage1_11[46], stage1_11[47]},
      {stage1_13[18], stage1_13[19], stage1_13[20], stage1_13[21], stage1_13[22], stage1_13[23]},
      {stage2_15[3],stage2_14[10],stage2_13[14],stage2_12[19],stage2_11[27]}
   );
   gpc615_5 gpc859 (
      {stage1_11[48], stage1_11[49], stage1_11[50], stage1_11[51], stage1_11[52]},
      {stage1_12[42]},
      {stage1_13[24], stage1_13[25], stage1_13[26], stage1_13[27], stage1_13[28], stage1_13[29]},
      {stage2_15[4],stage2_14[11],stage2_13[15],stage2_12[20],stage2_11[28]}
   );
   gpc615_5 gpc860 (
      {stage1_11[53], stage1_11[54], stage1_11[55], stage1_11[56], stage1_11[57]},
      {stage1_12[43]},
      {stage1_13[30], stage1_13[31], stage1_13[32], stage1_13[33], stage1_13[34], stage1_13[35]},
      {stage2_15[5],stage2_14[12],stage2_13[16],stage2_12[21],stage2_11[29]}
   );
   gpc606_5 gpc861 (
      {stage1_12[44], stage1_12[45], stage1_12[46], stage1_12[47], stage1_12[48], stage1_12[49]},
      {stage1_14[0], stage1_14[1], stage1_14[2], stage1_14[3], stage1_14[4], stage1_14[5]},
      {stage2_16[0],stage2_15[6],stage2_14[13],stage2_13[17],stage2_12[22]}
   );
   gpc606_5 gpc862 (
      {stage1_12[50], stage1_12[51], stage1_12[52], stage1_12[53], stage1_12[54], stage1_12[55]},
      {stage1_14[6], stage1_14[7], stage1_14[8], stage1_14[9], stage1_14[10], stage1_14[11]},
      {stage2_16[1],stage2_15[7],stage2_14[14],stage2_13[18],stage2_12[23]}
   );
   gpc1415_5 gpc863 (
      {stage1_13[36], stage1_13[37], stage1_13[38], stage1_13[39], stage1_13[40]},
      {stage1_14[12]},
      {stage1_15[0], stage1_15[1], stage1_15[2], stage1_15[3]},
      {stage1_16[0]},
      {stage2_17[0],stage2_16[2],stage2_15[8],stage2_14[15],stage2_13[19]}
   );
   gpc615_5 gpc864 (
      {stage1_13[41], stage1_13[42], stage1_13[43], stage1_13[44], stage1_13[45]},
      {stage1_14[13]},
      {stage1_15[4], stage1_15[5], stage1_15[6], stage1_15[7], stage1_15[8], stage1_15[9]},
      {stage2_17[1],stage2_16[3],stage2_15[9],stage2_14[16],stage2_13[20]}
   );
   gpc615_5 gpc865 (
      {stage1_13[46], stage1_13[47], stage1_13[48], stage1_13[49], stage1_13[50]},
      {stage1_14[14]},
      {stage1_15[10], stage1_15[11], stage1_15[12], stage1_15[13], stage1_15[14], stage1_15[15]},
      {stage2_17[2],stage2_16[4],stage2_15[10],stage2_14[17],stage2_13[21]}
   );
   gpc615_5 gpc866 (
      {stage1_13[51], stage1_13[52], stage1_13[53], stage1_13[54], stage1_13[55]},
      {stage1_14[15]},
      {stage1_15[16], stage1_15[17], stage1_15[18], stage1_15[19], stage1_15[20], stage1_15[21]},
      {stage2_17[3],stage2_16[5],stage2_15[11],stage2_14[18],stage2_13[22]}
   );
   gpc615_5 gpc867 (
      {stage1_13[56], stage1_13[57], stage1_13[58], stage1_13[59], stage1_13[60]},
      {stage1_14[16]},
      {stage1_15[22], stage1_15[23], stage1_15[24], stage1_15[25], stage1_15[26], stage1_15[27]},
      {stage2_17[4],stage2_16[6],stage2_15[12],stage2_14[19],stage2_13[23]}
   );
   gpc615_5 gpc868 (
      {stage1_13[61], stage1_13[62], stage1_13[63], stage1_13[64], stage1_13[65]},
      {stage1_14[17]},
      {stage1_15[28], stage1_15[29], stage1_15[30], stage1_15[31], stage1_15[32], stage1_15[33]},
      {stage2_17[5],stage2_16[7],stage2_15[13],stage2_14[20],stage2_13[24]}
   );
   gpc606_5 gpc869 (
      {stage1_14[18], stage1_14[19], stage1_14[20], stage1_14[21], stage1_14[22], stage1_14[23]},
      {stage1_16[1], stage1_16[2], stage1_16[3], stage1_16[4], stage1_16[5], stage1_16[6]},
      {stage2_18[0],stage2_17[6],stage2_16[8],stage2_15[14],stage2_14[21]}
   );
   gpc606_5 gpc870 (
      {stage1_14[24], stage1_14[25], stage1_14[26], stage1_14[27], stage1_14[28], stage1_14[29]},
      {stage1_16[7], stage1_16[8], stage1_16[9], stage1_16[10], stage1_16[11], stage1_16[12]},
      {stage2_18[1],stage2_17[7],stage2_16[9],stage2_15[15],stage2_14[22]}
   );
   gpc606_5 gpc871 (
      {stage1_14[30], stage1_14[31], stage1_14[32], stage1_14[33], stage1_14[34], stage1_14[35]},
      {stage1_16[13], stage1_16[14], stage1_16[15], stage1_16[16], stage1_16[17], stage1_16[18]},
      {stage2_18[2],stage2_17[8],stage2_16[10],stage2_15[16],stage2_14[23]}
   );
   gpc606_5 gpc872 (
      {stage1_14[36], stage1_14[37], stage1_14[38], stage1_14[39], stage1_14[40], stage1_14[41]},
      {stage1_16[19], stage1_16[20], stage1_16[21], stage1_16[22], stage1_16[23], stage1_16[24]},
      {stage2_18[3],stage2_17[9],stage2_16[11],stage2_15[17],stage2_14[24]}
   );
   gpc606_5 gpc873 (
      {stage1_14[42], stage1_14[43], stage1_14[44], stage1_14[45], stage1_14[46], stage1_14[47]},
      {stage1_16[25], stage1_16[26], stage1_16[27], stage1_16[28], stage1_16[29], stage1_16[30]},
      {stage2_18[4],stage2_17[10],stage2_16[12],stage2_15[18],stage2_14[25]}
   );
   gpc606_5 gpc874 (
      {stage1_14[48], stage1_14[49], stage1_14[50], stage1_14[51], stage1_14[52], stage1_14[53]},
      {stage1_16[31], stage1_16[32], stage1_16[33], stage1_16[34], stage1_16[35], stage1_16[36]},
      {stage2_18[5],stage2_17[11],stage2_16[13],stage2_15[19],stage2_14[26]}
   );
   gpc606_5 gpc875 (
      {stage1_14[54], stage1_14[55], stage1_14[56], stage1_14[57], stage1_14[58], stage1_14[59]},
      {stage1_16[37], stage1_16[38], stage1_16[39], stage1_16[40], stage1_16[41], stage1_16[42]},
      {stage2_18[6],stage2_17[12],stage2_16[14],stage2_15[20],stage2_14[27]}
   );
   gpc1406_5 gpc876 (
      {stage1_15[34], stage1_15[35], stage1_15[36], stage1_15[37], stage1_15[38], stage1_15[39]},
      {stage1_17[0], stage1_17[1], stage1_17[2], stage1_17[3]},
      {stage1_18[0]},
      {stage2_19[0],stage2_18[7],stage2_17[13],stage2_16[15],stage2_15[21]}
   );
   gpc615_5 gpc877 (
      {stage1_15[40], stage1_15[41], stage1_15[42], stage1_15[43], stage1_15[44]},
      {stage1_16[43]},
      {stage1_17[4], stage1_17[5], stage1_17[6], stage1_17[7], stage1_17[8], stage1_17[9]},
      {stage2_19[1],stage2_18[8],stage2_17[14],stage2_16[16],stage2_15[22]}
   );
   gpc615_5 gpc878 (
      {stage1_15[45], stage1_15[46], stage1_15[47], stage1_15[48], stage1_15[49]},
      {stage1_16[44]},
      {stage1_17[10], stage1_17[11], stage1_17[12], stage1_17[13], stage1_17[14], stage1_17[15]},
      {stage2_19[2],stage2_18[9],stage2_17[15],stage2_16[17],stage2_15[23]}
   );
   gpc615_5 gpc879 (
      {stage1_16[45], stage1_16[46], stage1_16[47], stage1_16[48], stage1_16[49]},
      {stage1_17[16]},
      {stage1_18[1], stage1_18[2], stage1_18[3], stage1_18[4], stage1_18[5], stage1_18[6]},
      {stage2_20[0],stage2_19[3],stage2_18[10],stage2_17[16],stage2_16[18]}
   );
   gpc615_5 gpc880 (
      {stage1_16[50], stage1_16[51], stage1_16[52], stage1_16[53], stage1_16[54]},
      {stage1_17[17]},
      {stage1_18[7], stage1_18[8], stage1_18[9], stage1_18[10], stage1_18[11], stage1_18[12]},
      {stage2_20[1],stage2_19[4],stage2_18[11],stage2_17[17],stage2_16[19]}
   );
   gpc615_5 gpc881 (
      {stage1_16[55], stage1_16[56], stage1_16[57], stage1_16[58], stage1_16[59]},
      {stage1_17[18]},
      {stage1_18[13], stage1_18[14], stage1_18[15], stage1_18[16], stage1_18[17], stage1_18[18]},
      {stage2_20[2],stage2_19[5],stage2_18[12],stage2_17[18],stage2_16[20]}
   );
   gpc615_5 gpc882 (
      {stage1_16[60], stage1_16[61], stage1_16[62], stage1_16[63], stage1_16[64]},
      {stage1_17[19]},
      {stage1_18[19], stage1_18[20], stage1_18[21], stage1_18[22], stage1_18[23], stage1_18[24]},
      {stage2_20[3],stage2_19[6],stage2_18[13],stage2_17[19],stage2_16[21]}
   );
   gpc615_5 gpc883 (
      {stage1_16[65], stage1_16[66], stage1_16[67], stage1_16[68], stage1_16[69]},
      {stage1_17[20]},
      {stage1_18[25], stage1_18[26], stage1_18[27], stage1_18[28], stage1_18[29], stage1_18[30]},
      {stage2_20[4],stage2_19[7],stage2_18[14],stage2_17[20],stage2_16[22]}
   );
   gpc615_5 gpc884 (
      {stage1_16[70], stage1_16[71], stage1_16[72], stage1_16[73], stage1_16[74]},
      {stage1_17[21]},
      {stage1_18[31], stage1_18[32], stage1_18[33], stage1_18[34], stage1_18[35], stage1_18[36]},
      {stage2_20[5],stage2_19[8],stage2_18[15],stage2_17[21],stage2_16[23]}
   );
   gpc615_5 gpc885 (
      {stage1_16[75], stage1_16[76], stage1_16[77], stage1_16[78], stage1_16[79]},
      {stage1_17[22]},
      {stage1_18[37], stage1_18[38], stage1_18[39], stage1_18[40], stage1_18[41], stage1_18[42]},
      {stage2_20[6],stage2_19[9],stage2_18[16],stage2_17[22],stage2_16[24]}
   );
   gpc615_5 gpc886 (
      {stage1_16[80], stage1_16[81], stage1_16[82], stage1_16[83], stage1_16[84]},
      {stage1_17[23]},
      {stage1_18[43], stage1_18[44], stage1_18[45], stage1_18[46], stage1_18[47], stage1_18[48]},
      {stage2_20[7],stage2_19[10],stage2_18[17],stage2_17[23],stage2_16[25]}
   );
   gpc615_5 gpc887 (
      {stage1_16[85], stage1_16[86], stage1_16[87], stage1_16[88], stage1_16[89]},
      {stage1_17[24]},
      {stage1_18[49], stage1_18[50], stage1_18[51], stage1_18[52], stage1_18[53], stage1_18[54]},
      {stage2_20[8],stage2_19[11],stage2_18[18],stage2_17[24],stage2_16[26]}
   );
   gpc606_5 gpc888 (
      {stage1_17[25], stage1_17[26], stage1_17[27], stage1_17[28], stage1_17[29], stage1_17[30]},
      {stage1_19[0], stage1_19[1], stage1_19[2], stage1_19[3], stage1_19[4], stage1_19[5]},
      {stage2_21[0],stage2_20[9],stage2_19[12],stage2_18[19],stage2_17[25]}
   );
   gpc606_5 gpc889 (
      {stage1_17[31], stage1_17[32], stage1_17[33], stage1_17[34], stage1_17[35], stage1_17[36]},
      {stage1_19[6], stage1_19[7], stage1_19[8], stage1_19[9], stage1_19[10], stage1_19[11]},
      {stage2_21[1],stage2_20[10],stage2_19[13],stage2_18[20],stage2_17[26]}
   );
   gpc606_5 gpc890 (
      {stage1_17[37], stage1_17[38], stage1_17[39], stage1_17[40], stage1_17[41], stage1_17[42]},
      {stage1_19[12], stage1_19[13], stage1_19[14], stage1_19[15], stage1_19[16], stage1_19[17]},
      {stage2_21[2],stage2_20[11],stage2_19[14],stage2_18[21],stage2_17[27]}
   );
   gpc615_5 gpc891 (
      {stage1_17[43], stage1_17[44], stage1_17[45], stage1_17[46], stage1_17[47]},
      {stage1_18[55]},
      {stage1_19[18], stage1_19[19], stage1_19[20], stage1_19[21], stage1_19[22], stage1_19[23]},
      {stage2_21[3],stage2_20[12],stage2_19[15],stage2_18[22],stage2_17[28]}
   );
   gpc615_5 gpc892 (
      {stage1_17[48], stage1_17[49], stage1_17[50], stage1_17[51], stage1_17[52]},
      {stage1_18[56]},
      {stage1_19[24], stage1_19[25], stage1_19[26], stage1_19[27], stage1_19[28], stage1_19[29]},
      {stage2_21[4],stage2_20[13],stage2_19[16],stage2_18[23],stage2_17[29]}
   );
   gpc615_5 gpc893 (
      {stage1_17[53], stage1_17[54], stage1_17[55], stage1_17[56], stage1_17[57]},
      {stage1_18[57]},
      {stage1_19[30], stage1_19[31], stage1_19[32], stage1_19[33], stage1_19[34], stage1_19[35]},
      {stage2_21[5],stage2_20[14],stage2_19[17],stage2_18[24],stage2_17[30]}
   );
   gpc606_5 gpc894 (
      {stage1_18[58], stage1_18[59], stage1_18[60], stage1_18[61], stage1_18[62], stage1_18[63]},
      {stage1_20[0], stage1_20[1], stage1_20[2], stage1_20[3], stage1_20[4], stage1_20[5]},
      {stage2_22[0],stage2_21[6],stage2_20[15],stage2_19[18],stage2_18[25]}
   );
   gpc606_5 gpc895 (
      {stage1_18[64], stage1_18[65], stage1_18[66], stage1_18[67], stage1_18[68], stage1_18[69]},
      {stage1_20[6], stage1_20[7], stage1_20[8], stage1_20[9], stage1_20[10], stage1_20[11]},
      {stage2_22[1],stage2_21[7],stage2_20[16],stage2_19[19],stage2_18[26]}
   );
   gpc606_5 gpc896 (
      {stage1_18[70], stage1_18[71], stage1_18[72], stage1_18[73], stage1_18[74], stage1_18[75]},
      {stage1_20[12], stage1_20[13], stage1_20[14], stage1_20[15], stage1_20[16], stage1_20[17]},
      {stage2_22[2],stage2_21[8],stage2_20[17],stage2_19[20],stage2_18[27]}
   );
   gpc606_5 gpc897 (
      {stage1_18[76], stage1_18[77], stage1_18[78], stage1_18[79], stage1_18[80], stage1_18[81]},
      {stage1_20[18], stage1_20[19], stage1_20[20], stage1_20[21], stage1_20[22], stage1_20[23]},
      {stage2_22[3],stage2_21[9],stage2_20[18],stage2_19[21],stage2_18[28]}
   );
   gpc606_5 gpc898 (
      {stage1_19[36], stage1_19[37], stage1_19[38], stage1_19[39], stage1_19[40], stage1_19[41]},
      {stage1_21[0], stage1_21[1], stage1_21[2], stage1_21[3], stage1_21[4], stage1_21[5]},
      {stage2_23[0],stage2_22[4],stage2_21[10],stage2_20[19],stage2_19[22]}
   );
   gpc606_5 gpc899 (
      {stage1_19[42], stage1_19[43], stage1_19[44], stage1_19[45], stage1_19[46], stage1_19[47]},
      {stage1_21[6], stage1_21[7], stage1_21[8], stage1_21[9], stage1_21[10], stage1_21[11]},
      {stage2_23[1],stage2_22[5],stage2_21[11],stage2_20[20],stage2_19[23]}
   );
   gpc606_5 gpc900 (
      {stage1_19[48], stage1_19[49], stage1_19[50], stage1_19[51], stage1_19[52], stage1_19[53]},
      {stage1_21[12], stage1_21[13], stage1_21[14], stage1_21[15], stage1_21[16], stage1_21[17]},
      {stage2_23[2],stage2_22[6],stage2_21[12],stage2_20[21],stage2_19[24]}
   );
   gpc606_5 gpc901 (
      {stage1_19[54], stage1_19[55], stage1_19[56], stage1_19[57], stage1_19[58], stage1_19[59]},
      {stage1_21[18], stage1_21[19], stage1_21[20], stage1_21[21], stage1_21[22], stage1_21[23]},
      {stage2_23[3],stage2_22[7],stage2_21[13],stage2_20[22],stage2_19[25]}
   );
   gpc606_5 gpc902 (
      {stage1_19[60], stage1_19[61], stage1_19[62], stage1_19[63], stage1_19[64], stage1_19[65]},
      {stage1_21[24], stage1_21[25], stage1_21[26], stage1_21[27], stage1_21[28], stage1_21[29]},
      {stage2_23[4],stage2_22[8],stage2_21[14],stage2_20[23],stage2_19[26]}
   );
   gpc606_5 gpc903 (
      {stage1_20[24], stage1_20[25], stage1_20[26], stage1_20[27], stage1_20[28], stage1_20[29]},
      {stage1_22[0], stage1_22[1], stage1_22[2], stage1_22[3], stage1_22[4], stage1_22[5]},
      {stage2_24[0],stage2_23[5],stage2_22[9],stage2_21[15],stage2_20[24]}
   );
   gpc606_5 gpc904 (
      {stage1_20[30], stage1_20[31], stage1_20[32], stage1_20[33], stage1_20[34], stage1_20[35]},
      {stage1_22[6], stage1_22[7], stage1_22[8], stage1_22[9], stage1_22[10], stage1_22[11]},
      {stage2_24[1],stage2_23[6],stage2_22[10],stage2_21[16],stage2_20[25]}
   );
   gpc606_5 gpc905 (
      {stage1_20[36], stage1_20[37], stage1_20[38], stage1_20[39], stage1_20[40], stage1_20[41]},
      {stage1_22[12], stage1_22[13], stage1_22[14], stage1_22[15], stage1_22[16], stage1_22[17]},
      {stage2_24[2],stage2_23[7],stage2_22[11],stage2_21[17],stage2_20[26]}
   );
   gpc615_5 gpc906 (
      {stage1_20[42], stage1_20[43], stage1_20[44], stage1_20[45], stage1_20[46]},
      {stage1_21[30]},
      {stage1_22[18], stage1_22[19], stage1_22[20], stage1_22[21], stage1_22[22], stage1_22[23]},
      {stage2_24[3],stage2_23[8],stage2_22[12],stage2_21[18],stage2_20[27]}
   );
   gpc615_5 gpc907 (
      {stage1_20[47], stage1_20[48], stage1_20[49], stage1_20[50], stage1_20[51]},
      {stage1_21[31]},
      {stage1_22[24], stage1_22[25], stage1_22[26], stage1_22[27], stage1_22[28], stage1_22[29]},
      {stage2_24[4],stage2_23[9],stage2_22[13],stage2_21[19],stage2_20[28]}
   );
   gpc606_5 gpc908 (
      {stage1_21[32], stage1_21[33], stage1_21[34], stage1_21[35], stage1_21[36], stage1_21[37]},
      {stage1_23[0], stage1_23[1], stage1_23[2], stage1_23[3], stage1_23[4], stage1_23[5]},
      {stage2_25[0],stage2_24[5],stage2_23[10],stage2_22[14],stage2_21[20]}
   );
   gpc606_5 gpc909 (
      {stage1_21[38], stage1_21[39], stage1_21[40], stage1_21[41], stage1_21[42], stage1_21[43]},
      {stage1_23[6], stage1_23[7], stage1_23[8], stage1_23[9], stage1_23[10], stage1_23[11]},
      {stage2_25[1],stage2_24[6],stage2_23[11],stage2_22[15],stage2_21[21]}
   );
   gpc606_5 gpc910 (
      {stage1_21[44], stage1_21[45], stage1_21[46], stage1_21[47], stage1_21[48], stage1_21[49]},
      {stage1_23[12], stage1_23[13], stage1_23[14], stage1_23[15], stage1_23[16], stage1_23[17]},
      {stage2_25[2],stage2_24[7],stage2_23[12],stage2_22[16],stage2_21[22]}
   );
   gpc606_5 gpc911 (
      {stage1_21[50], stage1_21[51], stage1_21[52], stage1_21[53], stage1_21[54], stage1_21[55]},
      {stage1_23[18], stage1_23[19], stage1_23[20], stage1_23[21], stage1_23[22], stage1_23[23]},
      {stage2_25[3],stage2_24[8],stage2_23[13],stage2_22[17],stage2_21[23]}
   );
   gpc606_5 gpc912 (
      {stage1_21[56], stage1_21[57], stage1_21[58], stage1_21[59], stage1_21[60], stage1_21[61]},
      {stage1_23[24], stage1_23[25], stage1_23[26], stage1_23[27], stage1_23[28], stage1_23[29]},
      {stage2_25[4],stage2_24[9],stage2_23[14],stage2_22[18],stage2_21[24]}
   );
   gpc606_5 gpc913 (
      {stage1_21[62], stage1_21[63], stage1_21[64], stage1_21[65], stage1_21[66], stage1_21[67]},
      {stage1_23[30], stage1_23[31], stage1_23[32], stage1_23[33], stage1_23[34], stage1_23[35]},
      {stage2_25[5],stage2_24[10],stage2_23[15],stage2_22[19],stage2_21[25]}
   );
   gpc606_5 gpc914 (
      {stage1_21[68], stage1_21[69], stage1_21[70], stage1_21[71], stage1_21[72], stage1_21[73]},
      {stage1_23[36], stage1_23[37], stage1_23[38], stage1_23[39], stage1_23[40], stage1_23[41]},
      {stage2_25[6],stage2_24[11],stage2_23[16],stage2_22[20],stage2_21[26]}
   );
   gpc606_5 gpc915 (
      {stage1_21[74], stage1_21[75], stage1_21[76], stage1_21[77], stage1_21[78], stage1_21[79]},
      {stage1_23[42], stage1_23[43], stage1_23[44], stage1_23[45], stage1_23[46], stage1_23[47]},
      {stage2_25[7],stage2_24[12],stage2_23[17],stage2_22[21],stage2_21[27]}
   );
   gpc606_5 gpc916 (
      {stage1_22[30], stage1_22[31], stage1_22[32], stage1_22[33], stage1_22[34], stage1_22[35]},
      {stage1_24[0], stage1_24[1], stage1_24[2], stage1_24[3], stage1_24[4], stage1_24[5]},
      {stage2_26[0],stage2_25[8],stage2_24[13],stage2_23[18],stage2_22[22]}
   );
   gpc606_5 gpc917 (
      {stage1_22[36], stage1_22[37], stage1_22[38], stage1_22[39], stage1_22[40], stage1_22[41]},
      {stage1_24[6], stage1_24[7], stage1_24[8], stage1_24[9], stage1_24[10], stage1_24[11]},
      {stage2_26[1],stage2_25[9],stage2_24[14],stage2_23[19],stage2_22[23]}
   );
   gpc606_5 gpc918 (
      {stage1_22[42], stage1_22[43], stage1_22[44], stage1_22[45], stage1_22[46], stage1_22[47]},
      {stage1_24[12], stage1_24[13], stage1_24[14], stage1_24[15], stage1_24[16], stage1_24[17]},
      {stage2_26[2],stage2_25[10],stage2_24[15],stage2_23[20],stage2_22[24]}
   );
   gpc606_5 gpc919 (
      {stage1_22[48], stage1_22[49], stage1_22[50], stage1_22[51], stage1_22[52], stage1_22[53]},
      {stage1_24[18], stage1_24[19], stage1_24[20], stage1_24[21], stage1_24[22], stage1_24[23]},
      {stage2_26[3],stage2_25[11],stage2_24[16],stage2_23[21],stage2_22[25]}
   );
   gpc606_5 gpc920 (
      {stage1_22[54], stage1_22[55], stage1_22[56], stage1_22[57], stage1_22[58], stage1_22[59]},
      {stage1_24[24], stage1_24[25], stage1_24[26], stage1_24[27], stage1_24[28], stage1_24[29]},
      {stage2_26[4],stage2_25[12],stage2_24[17],stage2_23[22],stage2_22[26]}
   );
   gpc606_5 gpc921 (
      {stage1_22[60], stage1_22[61], stage1_22[62], stage1_22[63], stage1_22[64], stage1_22[65]},
      {stage1_24[30], stage1_24[31], stage1_24[32], stage1_24[33], stage1_24[34], stage1_24[35]},
      {stage2_26[5],stage2_25[13],stage2_24[18],stage2_23[23],stage2_22[27]}
   );
   gpc606_5 gpc922 (
      {stage1_22[66], stage1_22[67], stage1_22[68], stage1_22[69], stage1_22[70], stage1_22[71]},
      {stage1_24[36], stage1_24[37], stage1_24[38], stage1_24[39], stage1_24[40], stage1_24[41]},
      {stage2_26[6],stage2_25[14],stage2_24[19],stage2_23[24],stage2_22[28]}
   );
   gpc606_5 gpc923 (
      {stage1_22[72], stage1_22[73], stage1_22[74], stage1_22[75], stage1_22[76], stage1_22[77]},
      {stage1_24[42], stage1_24[43], stage1_24[44], stage1_24[45], stage1_24[46], stage1_24[47]},
      {stage2_26[7],stage2_25[15],stage2_24[20],stage2_23[25],stage2_22[29]}
   );
   gpc606_5 gpc924 (
      {stage1_23[48], stage1_23[49], stage1_23[50], stage1_23[51], stage1_23[52], stage1_23[53]},
      {stage1_25[0], stage1_25[1], stage1_25[2], stage1_25[3], stage1_25[4], stage1_25[5]},
      {stage2_27[0],stage2_26[8],stage2_25[16],stage2_24[21],stage2_23[26]}
   );
   gpc606_5 gpc925 (
      {stage1_23[54], stage1_23[55], stage1_23[56], stage1_23[57], stage1_23[58], stage1_23[59]},
      {stage1_25[6], stage1_25[7], stage1_25[8], stage1_25[9], stage1_25[10], stage1_25[11]},
      {stage2_27[1],stage2_26[9],stage2_25[17],stage2_24[22],stage2_23[27]}
   );
   gpc606_5 gpc926 (
      {stage1_23[60], stage1_23[61], stage1_23[62], stage1_23[63], stage1_23[64], stage1_23[65]},
      {stage1_25[12], stage1_25[13], stage1_25[14], stage1_25[15], stage1_25[16], stage1_25[17]},
      {stage2_27[2],stage2_26[10],stage2_25[18],stage2_24[23],stage2_23[28]}
   );
   gpc606_5 gpc927 (
      {stage1_23[66], stage1_23[67], stage1_23[68], stage1_23[69], stage1_23[70], stage1_23[71]},
      {stage1_25[18], stage1_25[19], stage1_25[20], stage1_25[21], stage1_25[22], stage1_25[23]},
      {stage2_27[3],stage2_26[11],stage2_25[19],stage2_24[24],stage2_23[29]}
   );
   gpc606_5 gpc928 (
      {stage1_23[72], stage1_23[73], stage1_23[74], stage1_23[75], stage1_23[76], stage1_23[77]},
      {stage1_25[24], stage1_25[25], stage1_25[26], stage1_25[27], stage1_25[28], stage1_25[29]},
      {stage2_27[4],stage2_26[12],stage2_25[20],stage2_24[25],stage2_23[30]}
   );
   gpc606_5 gpc929 (
      {stage1_24[48], stage1_24[49], stage1_24[50], stage1_24[51], stage1_24[52], stage1_24[53]},
      {stage1_26[0], stage1_26[1], stage1_26[2], stage1_26[3], stage1_26[4], stage1_26[5]},
      {stage2_28[0],stage2_27[5],stage2_26[13],stage2_25[21],stage2_24[26]}
   );
   gpc606_5 gpc930 (
      {stage1_24[54], stage1_24[55], stage1_24[56], stage1_24[57], stage1_24[58], stage1_24[59]},
      {stage1_26[6], stage1_26[7], stage1_26[8], stage1_26[9], stage1_26[10], stage1_26[11]},
      {stage2_28[1],stage2_27[6],stage2_26[14],stage2_25[22],stage2_24[27]}
   );
   gpc606_5 gpc931 (
      {stage1_25[30], stage1_25[31], stage1_25[32], stage1_25[33], stage1_25[34], stage1_25[35]},
      {stage1_27[0], stage1_27[1], stage1_27[2], stage1_27[3], stage1_27[4], stage1_27[5]},
      {stage2_29[0],stage2_28[2],stage2_27[7],stage2_26[15],stage2_25[23]}
   );
   gpc606_5 gpc932 (
      {stage1_25[36], stage1_25[37], stage1_25[38], stage1_25[39], stage1_25[40], stage1_25[41]},
      {stage1_27[6], stage1_27[7], stage1_27[8], stage1_27[9], stage1_27[10], stage1_27[11]},
      {stage2_29[1],stage2_28[3],stage2_27[8],stage2_26[16],stage2_25[24]}
   );
   gpc606_5 gpc933 (
      {stage1_25[42], stage1_25[43], stage1_25[44], stage1_25[45], stage1_25[46], stage1_25[47]},
      {stage1_27[12], stage1_27[13], stage1_27[14], stage1_27[15], stage1_27[16], stage1_27[17]},
      {stage2_29[2],stage2_28[4],stage2_27[9],stage2_26[17],stage2_25[25]}
   );
   gpc606_5 gpc934 (
      {stage1_25[48], stage1_25[49], stage1_25[50], stage1_25[51], stage1_25[52], stage1_25[53]},
      {stage1_27[18], stage1_27[19], stage1_27[20], stage1_27[21], stage1_27[22], stage1_27[23]},
      {stage2_29[3],stage2_28[5],stage2_27[10],stage2_26[18],stage2_25[26]}
   );
   gpc606_5 gpc935 (
      {stage1_25[54], stage1_25[55], stage1_25[56], stage1_25[57], stage1_25[58], stage1_25[59]},
      {stage1_27[24], stage1_27[25], stage1_27[26], stage1_27[27], stage1_27[28], stage1_27[29]},
      {stage2_29[4],stage2_28[6],stage2_27[11],stage2_26[19],stage2_25[27]}
   );
   gpc606_5 gpc936 (
      {stage1_25[60], stage1_25[61], stage1_25[62], stage1_25[63], stage1_25[64], stage1_25[65]},
      {stage1_27[30], stage1_27[31], stage1_27[32], stage1_27[33], stage1_27[34], stage1_27[35]},
      {stage2_29[5],stage2_28[7],stage2_27[12],stage2_26[20],stage2_25[28]}
   );
   gpc606_5 gpc937 (
      {stage1_25[66], stage1_25[67], stage1_25[68], stage1_25[69], stage1_25[70], stage1_25[71]},
      {stage1_27[36], stage1_27[37], stage1_27[38], stage1_27[39], stage1_27[40], stage1_27[41]},
      {stage2_29[6],stage2_28[8],stage2_27[13],stage2_26[21],stage2_25[29]}
   );
   gpc606_5 gpc938 (
      {stage1_25[72], stage1_25[73], stage1_25[74], stage1_25[75], stage1_25[76], stage1_25[77]},
      {stage1_27[42], stage1_27[43], stage1_27[44], stage1_27[45], stage1_27[46], stage1_27[47]},
      {stage2_29[7],stage2_28[9],stage2_27[14],stage2_26[22],stage2_25[30]}
   );
   gpc606_5 gpc939 (
      {stage1_26[12], stage1_26[13], stage1_26[14], stage1_26[15], stage1_26[16], stage1_26[17]},
      {stage1_28[0], stage1_28[1], stage1_28[2], stage1_28[3], stage1_28[4], stage1_28[5]},
      {stage2_30[0],stage2_29[8],stage2_28[10],stage2_27[15],stage2_26[23]}
   );
   gpc606_5 gpc940 (
      {stage1_26[18], stage1_26[19], stage1_26[20], stage1_26[21], stage1_26[22], stage1_26[23]},
      {stage1_28[6], stage1_28[7], stage1_28[8], stage1_28[9], stage1_28[10], stage1_28[11]},
      {stage2_30[1],stage2_29[9],stage2_28[11],stage2_27[16],stage2_26[24]}
   );
   gpc606_5 gpc941 (
      {stage1_26[24], stage1_26[25], stage1_26[26], stage1_26[27], stage1_26[28], stage1_26[29]},
      {stage1_28[12], stage1_28[13], stage1_28[14], stage1_28[15], stage1_28[16], stage1_28[17]},
      {stage2_30[2],stage2_29[10],stage2_28[12],stage2_27[17],stage2_26[25]}
   );
   gpc606_5 gpc942 (
      {stage1_26[30], stage1_26[31], stage1_26[32], stage1_26[33], stage1_26[34], stage1_26[35]},
      {stage1_28[18], stage1_28[19], stage1_28[20], stage1_28[21], stage1_28[22], stage1_28[23]},
      {stage2_30[3],stage2_29[11],stage2_28[13],stage2_27[18],stage2_26[26]}
   );
   gpc606_5 gpc943 (
      {stage1_26[36], stage1_26[37], stage1_26[38], stage1_26[39], stage1_26[40], stage1_26[41]},
      {stage1_28[24], stage1_28[25], stage1_28[26], stage1_28[27], stage1_28[28], stage1_28[29]},
      {stage2_30[4],stage2_29[12],stage2_28[14],stage2_27[19],stage2_26[27]}
   );
   gpc606_5 gpc944 (
      {stage1_26[42], stage1_26[43], stage1_26[44], stage1_26[45], stage1_26[46], stage1_26[47]},
      {stage1_28[30], stage1_28[31], stage1_28[32], stage1_28[33], stage1_28[34], stage1_28[35]},
      {stage2_30[5],stage2_29[13],stage2_28[15],stage2_27[20],stage2_26[28]}
   );
   gpc606_5 gpc945 (
      {stage1_26[48], stage1_26[49], stage1_26[50], stage1_26[51], stage1_26[52], stage1_26[53]},
      {stage1_28[36], stage1_28[37], stage1_28[38], stage1_28[39], stage1_28[40], stage1_28[41]},
      {stage2_30[6],stage2_29[14],stage2_28[16],stage2_27[21],stage2_26[29]}
   );
   gpc615_5 gpc946 (
      {stage1_27[48], stage1_27[49], stage1_27[50], stage1_27[51], stage1_27[52]},
      {stage1_28[42]},
      {stage1_29[0], stage1_29[1], stage1_29[2], stage1_29[3], stage1_29[4], stage1_29[5]},
      {stage2_31[0],stage2_30[7],stage2_29[15],stage2_28[17],stage2_27[22]}
   );
   gpc615_5 gpc947 (
      {stage1_27[53], stage1_27[54], stage1_27[55], stage1_27[56], stage1_27[57]},
      {stage1_28[43]},
      {stage1_29[6], stage1_29[7], stage1_29[8], stage1_29[9], stage1_29[10], stage1_29[11]},
      {stage2_31[1],stage2_30[8],stage2_29[16],stage2_28[18],stage2_27[23]}
   );
   gpc606_5 gpc948 (
      {stage1_28[44], stage1_28[45], stage1_28[46], stage1_28[47], stage1_28[48], stage1_28[49]},
      {stage1_30[0], stage1_30[1], stage1_30[2], stage1_30[3], stage1_30[4], stage1_30[5]},
      {stage2_32[0],stage2_31[2],stage2_30[9],stage2_29[17],stage2_28[19]}
   );
   gpc606_5 gpc949 (
      {stage1_28[50], stage1_28[51], stage1_28[52], stage1_28[53], stage1_28[54], stage1_28[55]},
      {stage1_30[6], stage1_30[7], stage1_30[8], stage1_30[9], stage1_30[10], stage1_30[11]},
      {stage2_32[1],stage2_31[3],stage2_30[10],stage2_29[18],stage2_28[20]}
   );
   gpc606_5 gpc950 (
      {stage1_28[56], stage1_28[57], stage1_28[58], stage1_28[59], stage1_28[60], stage1_28[61]},
      {stage1_30[12], stage1_30[13], stage1_30[14], stage1_30[15], stage1_30[16], stage1_30[17]},
      {stage2_32[2],stage2_31[4],stage2_30[11],stage2_29[19],stage2_28[21]}
   );
   gpc615_5 gpc951 (
      {stage1_28[62], stage1_28[63], stage1_28[64], stage1_28[65], stage1_28[66]},
      {stage1_29[12]},
      {stage1_30[18], stage1_30[19], stage1_30[20], stage1_30[21], stage1_30[22], stage1_30[23]},
      {stage2_32[3],stage2_31[5],stage2_30[12],stage2_29[20],stage2_28[22]}
   );
   gpc615_5 gpc952 (
      {stage1_28[67], stage1_28[68], stage1_28[69], stage1_28[70], stage1_28[71]},
      {stage1_29[13]},
      {stage1_30[24], stage1_30[25], stage1_30[26], stage1_30[27], stage1_30[28], stage1_30[29]},
      {stage2_32[4],stage2_31[6],stage2_30[13],stage2_29[21],stage2_28[23]}
   );
   gpc606_5 gpc953 (
      {stage1_29[14], stage1_29[15], stage1_29[16], stage1_29[17], stage1_29[18], stage1_29[19]},
      {stage1_31[0], stage1_31[1], stage1_31[2], stage1_31[3], stage1_31[4], stage1_31[5]},
      {stage2_33[0],stage2_32[5],stage2_31[7],stage2_30[14],stage2_29[22]}
   );
   gpc606_5 gpc954 (
      {stage1_29[20], stage1_29[21], stage1_29[22], stage1_29[23], stage1_29[24], stage1_29[25]},
      {stage1_31[6], stage1_31[7], stage1_31[8], stage1_31[9], stage1_31[10], stage1_31[11]},
      {stage2_33[1],stage2_32[6],stage2_31[8],stage2_30[15],stage2_29[23]}
   );
   gpc606_5 gpc955 (
      {stage1_29[26], stage1_29[27], stage1_29[28], stage1_29[29], stage1_29[30], stage1_29[31]},
      {stage1_31[12], stage1_31[13], stage1_31[14], stage1_31[15], stage1_31[16], stage1_31[17]},
      {stage2_33[2],stage2_32[7],stage2_31[9],stage2_30[16],stage2_29[24]}
   );
   gpc606_5 gpc956 (
      {stage1_29[32], stage1_29[33], stage1_29[34], stage1_29[35], stage1_29[36], stage1_29[37]},
      {stage1_31[18], stage1_31[19], stage1_31[20], stage1_31[21], stage1_31[22], stage1_31[23]},
      {stage2_33[3],stage2_32[8],stage2_31[10],stage2_30[17],stage2_29[25]}
   );
   gpc606_5 gpc957 (
      {stage1_29[38], stage1_29[39], stage1_29[40], stage1_29[41], stage1_29[42], stage1_29[43]},
      {stage1_31[24], stage1_31[25], stage1_31[26], stage1_31[27], stage1_31[28], stage1_31[29]},
      {stage2_33[4],stage2_32[9],stage2_31[11],stage2_30[18],stage2_29[26]}
   );
   gpc606_5 gpc958 (
      {stage1_29[44], stage1_29[45], stage1_29[46], stage1_29[47], stage1_29[48], stage1_29[49]},
      {stage1_31[30], stage1_31[31], stage1_31[32], stage1_31[33], stage1_31[34], stage1_31[35]},
      {stage2_33[5],stage2_32[10],stage2_31[12],stage2_30[19],stage2_29[27]}
   );
   gpc615_5 gpc959 (
      {stage1_29[50], stage1_29[51], stage1_29[52], stage1_29[53], stage1_29[54]},
      {stage1_30[30]},
      {stage1_31[36], stage1_31[37], stage1_31[38], stage1_31[39], stage1_31[40], stage1_31[41]},
      {stage2_33[6],stage2_32[11],stage2_31[13],stage2_30[20],stage2_29[28]}
   );
   gpc615_5 gpc960 (
      {stage1_29[55], stage1_29[56], stage1_29[57], stage1_29[58], stage1_29[59]},
      {stage1_30[31]},
      {stage1_31[42], stage1_31[43], stage1_31[44], stage1_31[45], stage1_31[46], stage1_31[47]},
      {stage2_33[7],stage2_32[12],stage2_31[14],stage2_30[21],stage2_29[29]}
   );
   gpc615_5 gpc961 (
      {stage1_29[60], stage1_29[61], stage1_29[62], stage1_29[63], stage1_29[64]},
      {stage1_30[32]},
      {stage1_31[48], stage1_31[49], stage1_31[50], stage1_31[51], stage1_31[52], stage1_31[53]},
      {stage2_33[8],stage2_32[13],stage2_31[15],stage2_30[22],stage2_29[30]}
   );
   gpc615_5 gpc962 (
      {stage1_29[65], stage1_29[66], stage1_29[67], stage1_29[68], stage1_29[69]},
      {stage1_30[33]},
      {stage1_31[54], stage1_31[55], stage1_31[56], stage1_31[57], stage1_31[58], stage1_31[59]},
      {stage2_33[9],stage2_32[14],stage2_31[16],stage2_30[23],stage2_29[31]}
   );
   gpc615_5 gpc963 (
      {stage1_29[70], stage1_29[71], stage1_29[72], stage1_29[73], stage1_29[74]},
      {stage1_30[34]},
      {stage1_31[60], stage1_31[61], stage1_31[62], stage1_31[63], stage1_31[64], stage1_31[65]},
      {stage2_33[10],stage2_32[15],stage2_31[17],stage2_30[24],stage2_29[32]}
   );
   gpc615_5 gpc964 (
      {stage1_30[35], stage1_30[36], stage1_30[37], stage1_30[38], stage1_30[39]},
      {stage1_31[66]},
      {stage1_32[0], stage1_32[1], stage1_32[2], stage1_32[3], stage1_32[4], stage1_32[5]},
      {stage2_34[0],stage2_33[11],stage2_32[16],stage2_31[18],stage2_30[25]}
   );
   gpc615_5 gpc965 (
      {stage1_30[40], stage1_30[41], stage1_30[42], stage1_30[43], stage1_30[44]},
      {stage1_31[67]},
      {stage1_32[6], stage1_32[7], stage1_32[8], stage1_32[9], stage1_32[10], stage1_32[11]},
      {stage2_34[1],stage2_33[12],stage2_32[17],stage2_31[19],stage2_30[26]}
   );
   gpc615_5 gpc966 (
      {stage1_30[45], stage1_30[46], stage1_30[47], stage1_30[48], stage1_30[49]},
      {stage1_31[68]},
      {stage1_32[12], stage1_32[13], stage1_32[14], stage1_32[15], stage1_32[16], stage1_32[17]},
      {stage2_34[2],stage2_33[13],stage2_32[18],stage2_31[20],stage2_30[27]}
   );
   gpc615_5 gpc967 (
      {stage1_30[50], stage1_30[51], stage1_30[52], stage1_30[53], stage1_30[54]},
      {stage1_31[69]},
      {stage1_32[18], stage1_32[19], stage1_32[20], stage1_32[21], stage1_32[22], stage1_32[23]},
      {stage2_34[3],stage2_33[14],stage2_32[19],stage2_31[21],stage2_30[28]}
   );
   gpc135_4 gpc968 (
      {stage1_31[70], stage1_31[71], stage1_31[72], stage1_31[73], stage1_31[74]},
      {stage1_32[24], stage1_32[25], stage1_32[26]},
      {stage1_33[0]},
      {stage2_34[4],stage2_33[15],stage2_32[20],stage2_31[22]}
   );
   gpc606_5 gpc969 (
      {stage1_31[75], stage1_31[76], stage1_31[77], stage1_31[78], stage1_31[79], stage1_31[80]},
      {stage1_33[1], stage1_33[2], stage1_33[3], stage1_33[4], stage1_33[5], stage1_33[6]},
      {stage2_35[0],stage2_34[5],stage2_33[16],stage2_32[21],stage2_31[23]}
   );
   gpc606_5 gpc970 (
      {stage1_31[81], stage1_31[82], stage1_31[83], stage1_31[84], stage1_31[85], stage1_31[86]},
      {stage1_33[7], stage1_33[8], stage1_33[9], stage1_33[10], stage1_33[11], stage1_33[12]},
      {stage2_35[1],stage2_34[6],stage2_33[17],stage2_32[22],stage2_31[24]}
   );
   gpc1_1 gpc971 (
      {stage1_1[55]},
      {stage2_1[16]}
   );
   gpc1_1 gpc972 (
      {stage1_3[64]},
      {stage2_3[23]}
   );
   gpc1_1 gpc973 (
      {stage1_3[65]},
      {stage2_3[24]}
   );
   gpc1_1 gpc974 (
      {stage1_3[66]},
      {stage2_3[25]}
   );
   gpc1_1 gpc975 (
      {stage1_3[67]},
      {stage2_3[26]}
   );
   gpc1_1 gpc976 (
      {stage1_3[68]},
      {stage2_3[27]}
   );
   gpc1_1 gpc977 (
      {stage1_3[69]},
      {stage2_3[28]}
   );
   gpc1_1 gpc978 (
      {stage1_3[70]},
      {stage2_3[29]}
   );
   gpc1_1 gpc979 (
      {stage1_3[71]},
      {stage2_3[30]}
   );
   gpc1_1 gpc980 (
      {stage1_3[72]},
      {stage2_3[31]}
   );
   gpc1_1 gpc981 (
      {stage1_3[73]},
      {stage2_3[32]}
   );
   gpc1_1 gpc982 (
      {stage1_3[74]},
      {stage2_3[33]}
   );
   gpc1_1 gpc983 (
      {stage1_3[75]},
      {stage2_3[34]}
   );
   gpc1_1 gpc984 (
      {stage1_4[90]},
      {stage2_4[36]}
   );
   gpc1_1 gpc985 (
      {stage1_4[91]},
      {stage2_4[37]}
   );
   gpc1_1 gpc986 (
      {stage1_4[92]},
      {stage2_4[38]}
   );
   gpc1_1 gpc987 (
      {stage1_4[93]},
      {stage2_4[39]}
   );
   gpc1_1 gpc988 (
      {stage1_4[94]},
      {stage2_4[40]}
   );
   gpc1_1 gpc989 (
      {stage1_6[102]},
      {stage2_6[27]}
   );
   gpc1_1 gpc990 (
      {stage1_6[103]},
      {stage2_6[28]}
   );
   gpc1_1 gpc991 (
      {stage1_6[104]},
      {stage2_6[29]}
   );
   gpc1_1 gpc992 (
      {stage1_6[105]},
      {stage2_6[30]}
   );
   gpc1_1 gpc993 (
      {stage1_9[69]},
      {stage2_9[24]}
   );
   gpc1_1 gpc994 (
      {stage1_9[70]},
      {stage2_9[25]}
   );
   gpc1_1 gpc995 (
      {stage1_9[71]},
      {stage2_9[26]}
   );
   gpc1_1 gpc996 (
      {stage1_9[72]},
      {stage2_9[27]}
   );
   gpc1_1 gpc997 (
      {stage1_9[73]},
      {stage2_9[28]}
   );
   gpc1_1 gpc998 (
      {stage1_9[74]},
      {stage2_9[29]}
   );
   gpc1_1 gpc999 (
      {stage1_9[75]},
      {stage2_9[30]}
   );
   gpc1_1 gpc1000 (
      {stage1_9[76]},
      {stage2_9[31]}
   );
   gpc1_1 gpc1001 (
      {stage1_10[75]},
      {stage2_10[28]}
   );
   gpc1_1 gpc1002 (
      {stage1_10[76]},
      {stage2_10[29]}
   );
   gpc1_1 gpc1003 (
      {stage1_10[77]},
      {stage2_10[30]}
   );
   gpc1_1 gpc1004 (
      {stage1_10[78]},
      {stage2_10[31]}
   );
   gpc1_1 gpc1005 (
      {stage1_10[79]},
      {stage2_10[32]}
   );
   gpc1_1 gpc1006 (
      {stage1_10[80]},
      {stage2_10[33]}
   );
   gpc1_1 gpc1007 (
      {stage1_10[81]},
      {stage2_10[34]}
   );
   gpc1_1 gpc1008 (
      {stage1_10[82]},
      {stage2_10[35]}
   );
   gpc1_1 gpc1009 (
      {stage1_10[83]},
      {stage2_10[36]}
   );
   gpc1_1 gpc1010 (
      {stage1_10[84]},
      {stage2_10[37]}
   );
   gpc1_1 gpc1011 (
      {stage1_10[85]},
      {stage2_10[38]}
   );
   gpc1_1 gpc1012 (
      {stage1_10[86]},
      {stage2_10[39]}
   );
   gpc1_1 gpc1013 (
      {stage1_10[87]},
      {stage2_10[40]}
   );
   gpc1_1 gpc1014 (
      {stage1_10[88]},
      {stage2_10[41]}
   );
   gpc1_1 gpc1015 (
      {stage1_10[89]},
      {stage2_10[42]}
   );
   gpc1_1 gpc1016 (
      {stage1_10[90]},
      {stage2_10[43]}
   );
   gpc1_1 gpc1017 (
      {stage1_10[91]},
      {stage2_10[44]}
   );
   gpc1_1 gpc1018 (
      {stage1_10[92]},
      {stage2_10[45]}
   );
   gpc1_1 gpc1019 (
      {stage1_11[58]},
      {stage2_11[30]}
   );
   gpc1_1 gpc1020 (
      {stage1_11[59]},
      {stage2_11[31]}
   );
   gpc1_1 gpc1021 (
      {stage1_11[60]},
      {stage2_11[32]}
   );
   gpc1_1 gpc1022 (
      {stage1_11[61]},
      {stage2_11[33]}
   );
   gpc1_1 gpc1023 (
      {stage1_11[62]},
      {stage2_11[34]}
   );
   gpc1_1 gpc1024 (
      {stage1_11[63]},
      {stage2_11[35]}
   );
   gpc1_1 gpc1025 (
      {stage1_11[64]},
      {stage2_11[36]}
   );
   gpc1_1 gpc1026 (
      {stage1_11[65]},
      {stage2_11[37]}
   );
   gpc1_1 gpc1027 (
      {stage1_11[66]},
      {stage2_11[38]}
   );
   gpc1_1 gpc1028 (
      {stage1_13[66]},
      {stage2_13[25]}
   );
   gpc1_1 gpc1029 (
      {stage1_13[67]},
      {stage2_13[26]}
   );
   gpc1_1 gpc1030 (
      {stage1_13[68]},
      {stage2_13[27]}
   );
   gpc1_1 gpc1031 (
      {stage1_13[69]},
      {stage2_13[28]}
   );
   gpc1_1 gpc1032 (
      {stage1_13[70]},
      {stage2_13[29]}
   );
   gpc1_1 gpc1033 (
      {stage1_13[71]},
      {stage2_13[30]}
   );
   gpc1_1 gpc1034 (
      {stage1_13[72]},
      {stage2_13[31]}
   );
   gpc1_1 gpc1035 (
      {stage1_13[73]},
      {stage2_13[32]}
   );
   gpc1_1 gpc1036 (
      {stage1_13[74]},
      {stage2_13[33]}
   );
   gpc1_1 gpc1037 (
      {stage1_13[75]},
      {stage2_13[34]}
   );
   gpc1_1 gpc1038 (
      {stage1_13[76]},
      {stage2_13[35]}
   );
   gpc1_1 gpc1039 (
      {stage1_13[77]},
      {stage2_13[36]}
   );
   gpc1_1 gpc1040 (
      {stage1_13[78]},
      {stage2_13[37]}
   );
   gpc1_1 gpc1041 (
      {stage1_13[79]},
      {stage2_13[38]}
   );
   gpc1_1 gpc1042 (
      {stage1_13[80]},
      {stage2_13[39]}
   );
   gpc1_1 gpc1043 (
      {stage1_13[81]},
      {stage2_13[40]}
   );
   gpc1_1 gpc1044 (
      {stage1_13[82]},
      {stage2_13[41]}
   );
   gpc1_1 gpc1045 (
      {stage1_13[83]},
      {stage2_13[42]}
   );
   gpc1_1 gpc1046 (
      {stage1_13[84]},
      {stage2_13[43]}
   );
   gpc1_1 gpc1047 (
      {stage1_13[85]},
      {stage2_13[44]}
   );
   gpc1_1 gpc1048 (
      {stage1_14[60]},
      {stage2_14[28]}
   );
   gpc1_1 gpc1049 (
      {stage1_14[61]},
      {stage2_14[29]}
   );
   gpc1_1 gpc1050 (
      {stage1_14[62]},
      {stage2_14[30]}
   );
   gpc1_1 gpc1051 (
      {stage1_14[63]},
      {stage2_14[31]}
   );
   gpc1_1 gpc1052 (
      {stage1_14[64]},
      {stage2_14[32]}
   );
   gpc1_1 gpc1053 (
      {stage1_14[65]},
      {stage2_14[33]}
   );
   gpc1_1 gpc1054 (
      {stage1_14[66]},
      {stage2_14[34]}
   );
   gpc1_1 gpc1055 (
      {stage1_14[67]},
      {stage2_14[35]}
   );
   gpc1_1 gpc1056 (
      {stage1_14[68]},
      {stage2_14[36]}
   );
   gpc1_1 gpc1057 (
      {stage1_15[50]},
      {stage2_15[24]}
   );
   gpc1_1 gpc1058 (
      {stage1_15[51]},
      {stage2_15[25]}
   );
   gpc1_1 gpc1059 (
      {stage1_15[52]},
      {stage2_15[26]}
   );
   gpc1_1 gpc1060 (
      {stage1_15[53]},
      {stage2_15[27]}
   );
   gpc1_1 gpc1061 (
      {stage1_15[54]},
      {stage2_15[28]}
   );
   gpc1_1 gpc1062 (
      {stage1_15[55]},
      {stage2_15[29]}
   );
   gpc1_1 gpc1063 (
      {stage1_15[56]},
      {stage2_15[30]}
   );
   gpc1_1 gpc1064 (
      {stage1_15[57]},
      {stage2_15[31]}
   );
   gpc1_1 gpc1065 (
      {stage1_15[58]},
      {stage2_15[32]}
   );
   gpc1_1 gpc1066 (
      {stage1_15[59]},
      {stage2_15[33]}
   );
   gpc1_1 gpc1067 (
      {stage1_16[90]},
      {stage2_16[27]}
   );
   gpc1_1 gpc1068 (
      {stage1_16[91]},
      {stage2_16[28]}
   );
   gpc1_1 gpc1069 (
      {stage1_16[92]},
      {stage2_16[29]}
   );
   gpc1_1 gpc1070 (
      {stage1_16[93]},
      {stage2_16[30]}
   );
   gpc1_1 gpc1071 (
      {stage1_16[94]},
      {stage2_16[31]}
   );
   gpc1_1 gpc1072 (
      {stage1_16[95]},
      {stage2_16[32]}
   );
   gpc1_1 gpc1073 (
      {stage1_16[96]},
      {stage2_16[33]}
   );
   gpc1_1 gpc1074 (
      {stage1_16[97]},
      {stage2_16[34]}
   );
   gpc1_1 gpc1075 (
      {stage1_16[98]},
      {stage2_16[35]}
   );
   gpc1_1 gpc1076 (
      {stage1_16[99]},
      {stage2_16[36]}
   );
   gpc1_1 gpc1077 (
      {stage1_16[100]},
      {stage2_16[37]}
   );
   gpc1_1 gpc1078 (
      {stage1_16[101]},
      {stage2_16[38]}
   );
   gpc1_1 gpc1079 (
      {stage1_16[102]},
      {stage2_16[39]}
   );
   gpc1_1 gpc1080 (
      {stage1_16[103]},
      {stage2_16[40]}
   );
   gpc1_1 gpc1081 (
      {stage1_16[104]},
      {stage2_16[41]}
   );
   gpc1_1 gpc1082 (
      {stage1_16[105]},
      {stage2_16[42]}
   );
   gpc1_1 gpc1083 (
      {stage1_16[106]},
      {stage2_16[43]}
   );
   gpc1_1 gpc1084 (
      {stage1_17[58]},
      {stage2_17[31]}
   );
   gpc1_1 gpc1085 (
      {stage1_17[59]},
      {stage2_17[32]}
   );
   gpc1_1 gpc1086 (
      {stage1_17[60]},
      {stage2_17[33]}
   );
   gpc1_1 gpc1087 (
      {stage1_17[61]},
      {stage2_17[34]}
   );
   gpc1_1 gpc1088 (
      {stage1_17[62]},
      {stage2_17[35]}
   );
   gpc1_1 gpc1089 (
      {stage1_17[63]},
      {stage2_17[36]}
   );
   gpc1_1 gpc1090 (
      {stage1_19[66]},
      {stage2_19[27]}
   );
   gpc1_1 gpc1091 (
      {stage1_20[52]},
      {stage2_20[29]}
   );
   gpc1_1 gpc1092 (
      {stage1_20[53]},
      {stage2_20[30]}
   );
   gpc1_1 gpc1093 (
      {stage1_20[54]},
      {stage2_20[31]}
   );
   gpc1_1 gpc1094 (
      {stage1_20[55]},
      {stage2_20[32]}
   );
   gpc1_1 gpc1095 (
      {stage1_20[56]},
      {stage2_20[33]}
   );
   gpc1_1 gpc1096 (
      {stage1_20[57]},
      {stage2_20[34]}
   );
   gpc1_1 gpc1097 (
      {stage1_20[58]},
      {stage2_20[35]}
   );
   gpc1_1 gpc1098 (
      {stage1_20[59]},
      {stage2_20[36]}
   );
   gpc1_1 gpc1099 (
      {stage1_20[60]},
      {stage2_20[37]}
   );
   gpc1_1 gpc1100 (
      {stage1_22[78]},
      {stage2_22[30]}
   );
   gpc1_1 gpc1101 (
      {stage1_22[79]},
      {stage2_22[31]}
   );
   gpc1_1 gpc1102 (
      {stage1_22[80]},
      {stage2_22[32]}
   );
   gpc1_1 gpc1103 (
      {stage1_22[81]},
      {stage2_22[33]}
   );
   gpc1_1 gpc1104 (
      {stage1_23[78]},
      {stage2_23[31]}
   );
   gpc1_1 gpc1105 (
      {stage1_23[79]},
      {stage2_23[32]}
   );
   gpc1_1 gpc1106 (
      {stage1_23[80]},
      {stage2_23[33]}
   );
   gpc1_1 gpc1107 (
      {stage1_23[81]},
      {stage2_23[34]}
   );
   gpc1_1 gpc1108 (
      {stage1_23[82]},
      {stage2_23[35]}
   );
   gpc1_1 gpc1109 (
      {stage1_23[83]},
      {stage2_23[36]}
   );
   gpc1_1 gpc1110 (
      {stage1_23[84]},
      {stage2_23[37]}
   );
   gpc1_1 gpc1111 (
      {stage1_23[85]},
      {stage2_23[38]}
   );
   gpc1_1 gpc1112 (
      {stage1_23[86]},
      {stage2_23[39]}
   );
   gpc1_1 gpc1113 (
      {stage1_23[87]},
      {stage2_23[40]}
   );
   gpc1_1 gpc1114 (
      {stage1_23[88]},
      {stage2_23[41]}
   );
   gpc1_1 gpc1115 (
      {stage1_23[89]},
      {stage2_23[42]}
   );
   gpc1_1 gpc1116 (
      {stage1_23[90]},
      {stage2_23[43]}
   );
   gpc1_1 gpc1117 (
      {stage1_24[60]},
      {stage2_24[28]}
   );
   gpc1_1 gpc1118 (
      {stage1_24[61]},
      {stage2_24[29]}
   );
   gpc1_1 gpc1119 (
      {stage1_24[62]},
      {stage2_24[30]}
   );
   gpc1_1 gpc1120 (
      {stage1_24[63]},
      {stage2_24[31]}
   );
   gpc1_1 gpc1121 (
      {stage1_24[64]},
      {stage2_24[32]}
   );
   gpc1_1 gpc1122 (
      {stage1_24[65]},
      {stage2_24[33]}
   );
   gpc1_1 gpc1123 (
      {stage1_24[66]},
      {stage2_24[34]}
   );
   gpc1_1 gpc1124 (
      {stage1_26[54]},
      {stage2_26[30]}
   );
   gpc1_1 gpc1125 (
      {stage1_27[58]},
      {stage2_27[24]}
   );
   gpc1_1 gpc1126 (
      {stage1_27[59]},
      {stage2_27[25]}
   );
   gpc1_1 gpc1127 (
      {stage1_27[60]},
      {stage2_27[26]}
   );
   gpc1_1 gpc1128 (
      {stage1_27[61]},
      {stage2_27[27]}
   );
   gpc1_1 gpc1129 (
      {stage1_27[62]},
      {stage2_27[28]}
   );
   gpc1_1 gpc1130 (
      {stage1_27[63]},
      {stage2_27[29]}
   );
   gpc1_1 gpc1131 (
      {stage1_27[64]},
      {stage2_27[30]}
   );
   gpc1_1 gpc1132 (
      {stage1_27[65]},
      {stage2_27[31]}
   );
   gpc1_1 gpc1133 (
      {stage1_27[66]},
      {stage2_27[32]}
   );
   gpc1_1 gpc1134 (
      {stage1_28[72]},
      {stage2_28[24]}
   );
   gpc1_1 gpc1135 (
      {stage1_28[73]},
      {stage2_28[25]}
   );
   gpc1_1 gpc1136 (
      {stage1_28[74]},
      {stage2_28[26]}
   );
   gpc1_1 gpc1137 (
      {stage1_28[75]},
      {stage2_28[27]}
   );
   gpc1_1 gpc1138 (
      {stage1_28[76]},
      {stage2_28[28]}
   );
   gpc1_1 gpc1139 (
      {stage1_28[77]},
      {stage2_28[29]}
   );
   gpc1_1 gpc1140 (
      {stage1_30[55]},
      {stage2_30[29]}
   );
   gpc1_1 gpc1141 (
      {stage1_30[56]},
      {stage2_30[30]}
   );
   gpc1_1 gpc1142 (
      {stage1_30[57]},
      {stage2_30[31]}
   );
   gpc1_1 gpc1143 (
      {stage1_30[58]},
      {stage2_30[32]}
   );
   gpc1_1 gpc1144 (
      {stage1_30[59]},
      {stage2_30[33]}
   );
   gpc1_1 gpc1145 (
      {stage1_30[60]},
      {stage2_30[34]}
   );
   gpc1_1 gpc1146 (
      {stage1_30[61]},
      {stage2_30[35]}
   );
   gpc1_1 gpc1147 (
      {stage1_30[62]},
      {stage2_30[36]}
   );
   gpc1_1 gpc1148 (
      {stage1_31[87]},
      {stage2_31[25]}
   );
   gpc1_1 gpc1149 (
      {stage1_31[88]},
      {stage2_31[26]}
   );
   gpc1_1 gpc1150 (
      {stage1_31[89]},
      {stage2_31[27]}
   );
   gpc1_1 gpc1151 (
      {stage1_31[90]},
      {stage2_31[28]}
   );
   gpc1_1 gpc1152 (
      {stage1_31[91]},
      {stage2_31[29]}
   );
   gpc1_1 gpc1153 (
      {stage1_31[92]},
      {stage2_31[30]}
   );
   gpc1_1 gpc1154 (
      {stage1_31[93]},
      {stage2_31[31]}
   );
   gpc1_1 gpc1155 (
      {stage1_31[94]},
      {stage2_31[32]}
   );
   gpc1_1 gpc1156 (
      {stage1_31[95]},
      {stage2_31[33]}
   );
   gpc1_1 gpc1157 (
      {stage1_31[96]},
      {stage2_31[34]}
   );
   gpc1_1 gpc1158 (
      {stage1_31[97]},
      {stage2_31[35]}
   );
   gpc1_1 gpc1159 (
      {stage1_32[27]},
      {stage2_32[23]}
   );
   gpc1_1 gpc1160 (
      {stage1_32[28]},
      {stage2_32[24]}
   );
   gpc1_1 gpc1161 (
      {stage1_32[29]},
      {stage2_32[25]}
   );
   gpc1_1 gpc1162 (
      {stage1_32[30]},
      {stage2_32[26]}
   );
   gpc1_1 gpc1163 (
      {stage1_32[31]},
      {stage2_32[27]}
   );
   gpc1_1 gpc1164 (
      {stage1_32[32]},
      {stage2_32[28]}
   );
   gpc1_1 gpc1165 (
      {stage1_32[33]},
      {stage2_32[29]}
   );
   gpc1_1 gpc1166 (
      {stage1_32[34]},
      {stage2_32[30]}
   );
   gpc1_1 gpc1167 (
      {stage1_32[35]},
      {stage2_32[31]}
   );
   gpc1_1 gpc1168 (
      {stage1_32[36]},
      {stage2_32[32]}
   );
   gpc1_1 gpc1169 (
      {stage1_32[37]},
      {stage2_32[33]}
   );
   gpc1_1 gpc1170 (
      {stage1_32[38]},
      {stage2_32[34]}
   );
   gpc1_1 gpc1171 (
      {stage1_32[39]},
      {stage2_32[35]}
   );
   gpc1_1 gpc1172 (
      {stage1_32[40]},
      {stage2_32[36]}
   );
   gpc1_1 gpc1173 (
      {stage1_32[41]},
      {stage2_32[37]}
   );
   gpc1_1 gpc1174 (
      {stage1_32[42]},
      {stage2_32[38]}
   );
   gpc1_1 gpc1175 (
      {stage1_32[43]},
      {stage2_32[39]}
   );
   gpc1_1 gpc1176 (
      {stage1_32[44]},
      {stage2_32[40]}
   );
   gpc1_1 gpc1177 (
      {stage1_33[13]},
      {stage2_33[18]}
   );
   gpc1_1 gpc1178 (
      {stage1_33[14]},
      {stage2_33[19]}
   );
   gpc1_1 gpc1179 (
      {stage1_33[15]},
      {stage2_33[20]}
   );
   gpc1_1 gpc1180 (
      {stage1_33[16]},
      {stage2_33[21]}
   );
   gpc1_1 gpc1181 (
      {stage1_33[17]},
      {stage2_33[22]}
   );
   gpc1_1 gpc1182 (
      {stage1_33[18]},
      {stage2_33[23]}
   );
   gpc135_4 gpc1183 (
      {stage2_0[0], stage2_0[1], stage2_0[2], stage2_0[3], stage2_0[4]},
      {stage2_1[0], stage2_1[1], stage2_1[2]},
      {stage2_2[0]},
      {stage3_3[0],stage3_2[0],stage3_1[0],stage3_0[0]}
   );
   gpc606_5 gpc1184 (
      {stage2_1[3], stage2_1[4], stage2_1[5], stage2_1[6], stage2_1[7], stage2_1[8]},
      {stage2_3[0], stage2_3[1], stage2_3[2], stage2_3[3], stage2_3[4], stage2_3[5]},
      {stage3_5[0],stage3_4[0],stage3_3[1],stage3_2[1],stage3_1[1]}
   );
   gpc615_5 gpc1185 (
      {stage2_2[1], stage2_2[2], stage2_2[3], stage2_2[4], stage2_2[5]},
      {stage2_3[6]},
      {stage2_4[0], stage2_4[1], stage2_4[2], stage2_4[3], stage2_4[4], stage2_4[5]},
      {stage3_6[0],stage3_5[1],stage3_4[1],stage3_3[2],stage3_2[2]}
   );
   gpc615_5 gpc1186 (
      {stage2_2[6], stage2_2[7], stage2_2[8], stage2_2[9], stage2_2[10]},
      {stage2_3[7]},
      {stage2_4[6], stage2_4[7], stage2_4[8], stage2_4[9], stage2_4[10], stage2_4[11]},
      {stage3_6[1],stage3_5[2],stage3_4[2],stage3_3[3],stage3_2[3]}
   );
   gpc1163_5 gpc1187 (
      {stage2_3[8], stage2_3[9], stage2_3[10]},
      {stage2_4[12], stage2_4[13], stage2_4[14], stage2_4[15], stage2_4[16], stage2_4[17]},
      {stage2_5[0]},
      {stage2_6[0]},
      {stage3_7[0],stage3_6[2],stage3_5[3],stage3_4[3],stage3_3[4]}
   );
   gpc1163_5 gpc1188 (
      {stage2_3[11], stage2_3[12], stage2_3[13]},
      {stage2_4[18], stage2_4[19], stage2_4[20], stage2_4[21], stage2_4[22], stage2_4[23]},
      {stage2_5[1]},
      {stage2_6[1]},
      {stage3_7[1],stage3_6[3],stage3_5[4],stage3_4[4],stage3_3[5]}
   );
   gpc1163_5 gpc1189 (
      {stage2_3[14], stage2_3[15], stage2_3[16]},
      {stage2_4[24], stage2_4[25], stage2_4[26], stage2_4[27], stage2_4[28], stage2_4[29]},
      {stage2_5[2]},
      {stage2_6[2]},
      {stage3_7[2],stage3_6[4],stage3_5[5],stage3_4[5],stage3_3[6]}
   );
   gpc623_5 gpc1190 (
      {stage2_3[17], stage2_3[18], stage2_3[19]},
      {stage2_4[30], stage2_4[31]},
      {stage2_5[3], stage2_5[4], stage2_5[5], stage2_5[6], stage2_5[7], stage2_5[8]},
      {stage3_7[3],stage3_6[5],stage3_5[6],stage3_4[6],stage3_3[7]}
   );
   gpc615_5 gpc1191 (
      {stage2_4[32], stage2_4[33], stage2_4[34], stage2_4[35], stage2_4[36]},
      {stage2_5[9]},
      {stage2_6[3], stage2_6[4], stage2_6[5], stage2_6[6], stage2_6[7], stage2_6[8]},
      {stage3_8[0],stage3_7[4],stage3_6[6],stage3_5[7],stage3_4[7]}
   );
   gpc615_5 gpc1192 (
      {stage2_4[37], stage2_4[38], stage2_4[39], stage2_4[40], 1'b0},
      {stage2_5[10]},
      {stage2_6[9], stage2_6[10], stage2_6[11], stage2_6[12], stage2_6[13], stage2_6[14]},
      {stage3_8[1],stage3_7[5],stage3_6[7],stage3_5[8],stage3_4[8]}
   );
   gpc606_5 gpc1193 (
      {stage2_5[11], stage2_5[12], stage2_5[13], stage2_5[14], stage2_5[15], stage2_5[16]},
      {stage2_7[0], stage2_7[1], stage2_7[2], stage2_7[3], stage2_7[4], stage2_7[5]},
      {stage3_9[0],stage3_8[2],stage3_7[6],stage3_6[8],stage3_5[9]}
   );
   gpc606_5 gpc1194 (
      {stage2_5[17], stage2_5[18], stage2_5[19], stage2_5[20], stage2_5[21], stage2_5[22]},
      {stage2_7[6], stage2_7[7], stage2_7[8], stage2_7[9], stage2_7[10], stage2_7[11]},
      {stage3_9[1],stage3_8[3],stage3_7[7],stage3_6[9],stage3_5[10]}
   );
   gpc606_5 gpc1195 (
      {stage2_5[23], stage2_5[24], stage2_5[25], stage2_5[26], stage2_5[27], 1'b0},
      {stage2_7[12], stage2_7[13], stage2_7[14], stage2_7[15], stage2_7[16], stage2_7[17]},
      {stage3_9[2],stage3_8[4],stage3_7[8],stage3_6[10],stage3_5[11]}
   );
   gpc606_5 gpc1196 (
      {stage2_6[15], stage2_6[16], stage2_6[17], stage2_6[18], stage2_6[19], stage2_6[20]},
      {stage2_8[0], stage2_8[1], stage2_8[2], stage2_8[3], stage2_8[4], stage2_8[5]},
      {stage3_10[0],stage3_9[3],stage3_8[5],stage3_7[9],stage3_6[11]}
   );
   gpc606_5 gpc1197 (
      {stage2_6[21], stage2_6[22], stage2_6[23], stage2_6[24], stage2_6[25], stage2_6[26]},
      {stage2_8[6], stage2_8[7], stage2_8[8], stage2_8[9], stage2_8[10], stage2_8[11]},
      {stage3_10[1],stage3_9[4],stage3_8[6],stage3_7[10],stage3_6[12]}
   );
   gpc615_5 gpc1198 (
      {stage2_7[18], stage2_7[19], stage2_7[20], stage2_7[21], stage2_7[22]},
      {stage2_8[12]},
      {stage2_9[0], stage2_9[1], stage2_9[2], stage2_9[3], stage2_9[4], stage2_9[5]},
      {stage3_11[0],stage3_10[2],stage3_9[5],stage3_8[7],stage3_7[11]}
   );
   gpc615_5 gpc1199 (
      {stage2_7[23], stage2_7[24], stage2_7[25], stage2_7[26], stage2_7[27]},
      {stage2_8[13]},
      {stage2_9[6], stage2_9[7], stage2_9[8], stage2_9[9], stage2_9[10], stage2_9[11]},
      {stage3_11[1],stage3_10[3],stage3_9[6],stage3_8[8],stage3_7[12]}
   );
   gpc606_5 gpc1200 (
      {stage2_8[14], stage2_8[15], stage2_8[16], stage2_8[17], stage2_8[18], stage2_8[19]},
      {stage2_10[0], stage2_10[1], stage2_10[2], stage2_10[3], stage2_10[4], stage2_10[5]},
      {stage3_12[0],stage3_11[2],stage3_10[4],stage3_9[7],stage3_8[9]}
   );
   gpc606_5 gpc1201 (
      {stage2_8[20], stage2_8[21], stage2_8[22], stage2_8[23], stage2_8[24], stage2_8[25]},
      {stage2_10[6], stage2_10[7], stage2_10[8], stage2_10[9], stage2_10[10], stage2_10[11]},
      {stage3_12[1],stage3_11[3],stage3_10[5],stage3_9[8],stage3_8[10]}
   );
   gpc1343_5 gpc1202 (
      {stage2_9[12], stage2_9[13], stage2_9[14]},
      {stage2_10[12], stage2_10[13], stage2_10[14], stage2_10[15]},
      {stage2_11[0], stage2_11[1], stage2_11[2]},
      {stage2_12[0]},
      {stage3_13[0],stage3_12[2],stage3_11[4],stage3_10[6],stage3_9[9]}
   );
   gpc1343_5 gpc1203 (
      {stage2_9[15], stage2_9[16], stage2_9[17]},
      {stage2_10[16], stage2_10[17], stage2_10[18], stage2_10[19]},
      {stage2_11[3], stage2_11[4], stage2_11[5]},
      {stage2_12[1]},
      {stage3_13[1],stage3_12[3],stage3_11[5],stage3_10[7],stage3_9[10]}
   );
   gpc1343_5 gpc1204 (
      {stage2_9[18], stage2_9[19], stage2_9[20]},
      {stage2_10[20], stage2_10[21], stage2_10[22], stage2_10[23]},
      {stage2_11[6], stage2_11[7], stage2_11[8]},
      {stage2_12[2]},
      {stage3_13[2],stage3_12[4],stage3_11[6],stage3_10[8],stage3_9[11]}
   );
   gpc1343_5 gpc1205 (
      {stage2_9[21], stage2_9[22], stage2_9[23]},
      {stage2_10[24], stage2_10[25], stage2_10[26], stage2_10[27]},
      {stage2_11[9], stage2_11[10], stage2_11[11]},
      {stage2_12[3]},
      {stage3_13[3],stage3_12[5],stage3_11[7],stage3_10[9],stage3_9[12]}
   );
   gpc1343_5 gpc1206 (
      {stage2_9[24], stage2_9[25], stage2_9[26]},
      {stage2_10[28], stage2_10[29], stage2_10[30], stage2_10[31]},
      {stage2_11[12], stage2_11[13], stage2_11[14]},
      {stage2_12[4]},
      {stage3_13[4],stage3_12[6],stage3_11[8],stage3_10[10],stage3_9[13]}
   );
   gpc606_5 gpc1207 (
      {stage2_10[32], stage2_10[33], stage2_10[34], stage2_10[35], stage2_10[36], stage2_10[37]},
      {stage2_12[5], stage2_12[6], stage2_12[7], stage2_12[8], stage2_12[9], stage2_12[10]},
      {stage3_14[0],stage3_13[5],stage3_12[7],stage3_11[9],stage3_10[11]}
   );
   gpc606_5 gpc1208 (
      {stage2_10[38], stage2_10[39], stage2_10[40], stage2_10[41], stage2_10[42], stage2_10[43]},
      {stage2_12[11], stage2_12[12], stage2_12[13], stage2_12[14], stage2_12[15], stage2_12[16]},
      {stage3_14[1],stage3_13[6],stage3_12[8],stage3_11[10],stage3_10[12]}
   );
   gpc606_5 gpc1209 (
      {stage2_11[15], stage2_11[16], stage2_11[17], stage2_11[18], stage2_11[19], stage2_11[20]},
      {stage2_13[0], stage2_13[1], stage2_13[2], stage2_13[3], stage2_13[4], stage2_13[5]},
      {stage3_15[0],stage3_14[2],stage3_13[7],stage3_12[9],stage3_11[11]}
   );
   gpc606_5 gpc1210 (
      {stage2_11[21], stage2_11[22], stage2_11[23], stage2_11[24], stage2_11[25], stage2_11[26]},
      {stage2_13[6], stage2_13[7], stage2_13[8], stage2_13[9], stage2_13[10], stage2_13[11]},
      {stage3_15[1],stage3_14[3],stage3_13[8],stage3_12[10],stage3_11[12]}
   );
   gpc606_5 gpc1211 (
      {stage2_11[27], stage2_11[28], stage2_11[29], stage2_11[30], stage2_11[31], stage2_11[32]},
      {stage2_13[12], stage2_13[13], stage2_13[14], stage2_13[15], stage2_13[16], stage2_13[17]},
      {stage3_15[2],stage3_14[4],stage3_13[9],stage3_12[11],stage3_11[13]}
   );
   gpc606_5 gpc1212 (
      {stage2_11[33], stage2_11[34], stage2_11[35], stage2_11[36], stage2_11[37], stage2_11[38]},
      {stage2_13[18], stage2_13[19], stage2_13[20], stage2_13[21], stage2_13[22], stage2_13[23]},
      {stage3_15[3],stage3_14[5],stage3_13[10],stage3_12[12],stage3_11[14]}
   );
   gpc606_5 gpc1213 (
      {stage2_12[17], stage2_12[18], stage2_12[19], stage2_12[20], stage2_12[21], stage2_12[22]},
      {stage2_14[0], stage2_14[1], stage2_14[2], stage2_14[3], stage2_14[4], stage2_14[5]},
      {stage3_16[0],stage3_15[4],stage3_14[6],stage3_13[11],stage3_12[13]}
   );
   gpc606_5 gpc1214 (
      {stage2_13[24], stage2_13[25], stage2_13[26], stage2_13[27], stage2_13[28], stage2_13[29]},
      {stage2_15[0], stage2_15[1], stage2_15[2], stage2_15[3], stage2_15[4], stage2_15[5]},
      {stage3_17[0],stage3_16[1],stage3_15[5],stage3_14[7],stage3_13[12]}
   );
   gpc606_5 gpc1215 (
      {stage2_13[30], stage2_13[31], stage2_13[32], stage2_13[33], stage2_13[34], stage2_13[35]},
      {stage2_15[6], stage2_15[7], stage2_15[8], stage2_15[9], stage2_15[10], stage2_15[11]},
      {stage3_17[1],stage3_16[2],stage3_15[6],stage3_14[8],stage3_13[13]}
   );
   gpc606_5 gpc1216 (
      {stage2_13[36], stage2_13[37], stage2_13[38], stage2_13[39], stage2_13[40], stage2_13[41]},
      {stage2_15[12], stage2_15[13], stage2_15[14], stage2_15[15], stage2_15[16], stage2_15[17]},
      {stage3_17[2],stage3_16[3],stage3_15[7],stage3_14[9],stage3_13[14]}
   );
   gpc615_5 gpc1217 (
      {stage2_14[6], stage2_14[7], stage2_14[8], stage2_14[9], stage2_14[10]},
      {stage2_15[18]},
      {stage2_16[0], stage2_16[1], stage2_16[2], stage2_16[3], stage2_16[4], stage2_16[5]},
      {stage3_18[0],stage3_17[3],stage3_16[4],stage3_15[8],stage3_14[10]}
   );
   gpc615_5 gpc1218 (
      {stage2_14[11], stage2_14[12], stage2_14[13], stage2_14[14], stage2_14[15]},
      {stage2_15[19]},
      {stage2_16[6], stage2_16[7], stage2_16[8], stage2_16[9], stage2_16[10], stage2_16[11]},
      {stage3_18[1],stage3_17[4],stage3_16[5],stage3_15[9],stage3_14[11]}
   );
   gpc615_5 gpc1219 (
      {stage2_14[16], stage2_14[17], stage2_14[18], stage2_14[19], stage2_14[20]},
      {stage2_15[20]},
      {stage2_16[12], stage2_16[13], stage2_16[14], stage2_16[15], stage2_16[16], stage2_16[17]},
      {stage3_18[2],stage3_17[5],stage3_16[6],stage3_15[10],stage3_14[12]}
   );
   gpc615_5 gpc1220 (
      {stage2_14[21], stage2_14[22], stage2_14[23], stage2_14[24], stage2_14[25]},
      {stage2_15[21]},
      {stage2_16[18], stage2_16[19], stage2_16[20], stage2_16[21], stage2_16[22], stage2_16[23]},
      {stage3_18[3],stage3_17[6],stage3_16[7],stage3_15[11],stage3_14[13]}
   );
   gpc615_5 gpc1221 (
      {stage2_14[26], stage2_14[27], stage2_14[28], stage2_14[29], stage2_14[30]},
      {stage2_15[22]},
      {stage2_16[24], stage2_16[25], stage2_16[26], stage2_16[27], stage2_16[28], stage2_16[29]},
      {stage3_18[4],stage3_17[7],stage3_16[8],stage3_15[12],stage3_14[14]}
   );
   gpc615_5 gpc1222 (
      {stage2_14[31], stage2_14[32], stage2_14[33], stage2_14[34], stage2_14[35]},
      {stage2_15[23]},
      {stage2_16[30], stage2_16[31], stage2_16[32], stage2_16[33], stage2_16[34], stage2_16[35]},
      {stage3_18[5],stage3_17[8],stage3_16[9],stage3_15[13],stage3_14[15]}
   );
   gpc615_5 gpc1223 (
      {stage2_15[24], stage2_15[25], stage2_15[26], stage2_15[27], stage2_15[28]},
      {stage2_16[36]},
      {stage2_17[0], stage2_17[1], stage2_17[2], stage2_17[3], stage2_17[4], stage2_17[5]},
      {stage3_19[0],stage3_18[6],stage3_17[9],stage3_16[10],stage3_15[14]}
   );
   gpc615_5 gpc1224 (
      {stage2_15[29], stage2_15[30], stage2_15[31], stage2_15[32], stage2_15[33]},
      {stage2_16[37]},
      {stage2_17[6], stage2_17[7], stage2_17[8], stage2_17[9], stage2_17[10], stage2_17[11]},
      {stage3_19[1],stage3_18[7],stage3_17[10],stage3_16[11],stage3_15[15]}
   );
   gpc606_5 gpc1225 (
      {stage2_16[38], stage2_16[39], stage2_16[40], stage2_16[41], stage2_16[42], stage2_16[43]},
      {stage2_18[0], stage2_18[1], stage2_18[2], stage2_18[3], stage2_18[4], stage2_18[5]},
      {stage3_20[0],stage3_19[2],stage3_18[8],stage3_17[11],stage3_16[12]}
   );
   gpc606_5 gpc1226 (
      {stage2_17[12], stage2_17[13], stage2_17[14], stage2_17[15], stage2_17[16], stage2_17[17]},
      {stage2_19[0], stage2_19[1], stage2_19[2], stage2_19[3], stage2_19[4], stage2_19[5]},
      {stage3_21[0],stage3_20[1],stage3_19[3],stage3_18[9],stage3_17[12]}
   );
   gpc606_5 gpc1227 (
      {stage2_17[18], stage2_17[19], stage2_17[20], stage2_17[21], stage2_17[22], stage2_17[23]},
      {stage2_19[6], stage2_19[7], stage2_19[8], stage2_19[9], stage2_19[10], stage2_19[11]},
      {stage3_21[1],stage3_20[2],stage3_19[4],stage3_18[10],stage3_17[13]}
   );
   gpc606_5 gpc1228 (
      {stage2_17[24], stage2_17[25], stage2_17[26], stage2_17[27], stage2_17[28], stage2_17[29]},
      {stage2_19[12], stage2_19[13], stage2_19[14], stage2_19[15], stage2_19[16], stage2_19[17]},
      {stage3_21[2],stage3_20[3],stage3_19[5],stage3_18[11],stage3_17[14]}
   );
   gpc606_5 gpc1229 (
      {stage2_17[30], stage2_17[31], stage2_17[32], stage2_17[33], stage2_17[34], stage2_17[35]},
      {stage2_19[18], stage2_19[19], stage2_19[20], stage2_19[21], stage2_19[22], stage2_19[23]},
      {stage3_21[3],stage3_20[4],stage3_19[6],stage3_18[12],stage3_17[15]}
   );
   gpc606_5 gpc1230 (
      {stage2_18[6], stage2_18[7], stage2_18[8], stage2_18[9], stage2_18[10], stage2_18[11]},
      {stage2_20[0], stage2_20[1], stage2_20[2], stage2_20[3], stage2_20[4], stage2_20[5]},
      {stage3_22[0],stage3_21[4],stage3_20[5],stage3_19[7],stage3_18[13]}
   );
   gpc606_5 gpc1231 (
      {stage2_18[12], stage2_18[13], stage2_18[14], stage2_18[15], stage2_18[16], stage2_18[17]},
      {stage2_20[6], stage2_20[7], stage2_20[8], stage2_20[9], stage2_20[10], stage2_20[11]},
      {stage3_22[1],stage3_21[5],stage3_20[6],stage3_19[8],stage3_18[14]}
   );
   gpc606_5 gpc1232 (
      {stage2_18[18], stage2_18[19], stage2_18[20], stage2_18[21], stage2_18[22], stage2_18[23]},
      {stage2_20[12], stage2_20[13], stage2_20[14], stage2_20[15], stage2_20[16], stage2_20[17]},
      {stage3_22[2],stage3_21[6],stage3_20[7],stage3_19[9],stage3_18[15]}
   );
   gpc615_5 gpc1233 (
      {stage2_18[24], stage2_18[25], stage2_18[26], stage2_18[27], stage2_18[28]},
      {stage2_19[24]},
      {stage2_20[18], stage2_20[19], stage2_20[20], stage2_20[21], stage2_20[22], stage2_20[23]},
      {stage3_22[3],stage3_21[7],stage3_20[8],stage3_19[10],stage3_18[16]}
   );
   gpc615_5 gpc1234 (
      {stage2_19[25], stage2_19[26], stage2_19[27], 1'b0, 1'b0},
      {stage2_20[24]},
      {stage2_21[0], stage2_21[1], stage2_21[2], stage2_21[3], stage2_21[4], stage2_21[5]},
      {stage3_23[0],stage3_22[4],stage3_21[8],stage3_20[9],stage3_19[11]}
   );
   gpc606_5 gpc1235 (
      {stage2_20[25], stage2_20[26], stage2_20[27], stage2_20[28], stage2_20[29], stage2_20[30]},
      {stage2_22[0], stage2_22[1], stage2_22[2], stage2_22[3], stage2_22[4], stage2_22[5]},
      {stage3_24[0],stage3_23[1],stage3_22[5],stage3_21[9],stage3_20[10]}
   );
   gpc615_5 gpc1236 (
      {stage2_21[6], stage2_21[7], stage2_21[8], stage2_21[9], stage2_21[10]},
      {stage2_22[6]},
      {stage2_23[0], stage2_23[1], stage2_23[2], stage2_23[3], stage2_23[4], stage2_23[5]},
      {stage3_25[0],stage3_24[1],stage3_23[2],stage3_22[6],stage3_21[10]}
   );
   gpc615_5 gpc1237 (
      {stage2_21[11], stage2_21[12], stage2_21[13], stage2_21[14], stage2_21[15]},
      {stage2_22[7]},
      {stage2_23[6], stage2_23[7], stage2_23[8], stage2_23[9], stage2_23[10], stage2_23[11]},
      {stage3_25[1],stage3_24[2],stage3_23[3],stage3_22[7],stage3_21[11]}
   );
   gpc615_5 gpc1238 (
      {stage2_21[16], stage2_21[17], stage2_21[18], stage2_21[19], stage2_21[20]},
      {stage2_22[8]},
      {stage2_23[12], stage2_23[13], stage2_23[14], stage2_23[15], stage2_23[16], stage2_23[17]},
      {stage3_25[2],stage3_24[3],stage3_23[4],stage3_22[8],stage3_21[12]}
   );
   gpc615_5 gpc1239 (
      {stage2_21[21], stage2_21[22], stage2_21[23], stage2_21[24], stage2_21[25]},
      {stage2_22[9]},
      {stage2_23[18], stage2_23[19], stage2_23[20], stage2_23[21], stage2_23[22], stage2_23[23]},
      {stage3_25[3],stage3_24[4],stage3_23[5],stage3_22[9],stage3_21[13]}
   );
   gpc615_5 gpc1240 (
      {stage2_21[26], stage2_21[27], 1'b0, 1'b0, 1'b0},
      {stage2_22[10]},
      {stage2_23[24], stage2_23[25], stage2_23[26], stage2_23[27], stage2_23[28], stage2_23[29]},
      {stage3_25[4],stage3_24[5],stage3_23[6],stage3_22[10],stage3_21[14]}
   );
   gpc207_4 gpc1241 (
      {stage2_22[11], stage2_22[12], stage2_22[13], stage2_22[14], stage2_22[15], stage2_22[16], stage2_22[17]},
      {stage2_24[0], stage2_24[1]},
      {stage3_25[5],stage3_24[6],stage3_23[7],stage3_22[11]}
   );
   gpc606_5 gpc1242 (
      {stage2_22[18], stage2_22[19], stage2_22[20], stage2_22[21], stage2_22[22], stage2_22[23]},
      {stage2_24[2], stage2_24[3], stage2_24[4], stage2_24[5], stage2_24[6], stage2_24[7]},
      {stage3_26[0],stage3_25[6],stage3_24[7],stage3_23[8],stage3_22[12]}
   );
   gpc606_5 gpc1243 (
      {stage2_23[30], stage2_23[31], stage2_23[32], stage2_23[33], stage2_23[34], stage2_23[35]},
      {stage2_25[0], stage2_25[1], stage2_25[2], stage2_25[3], stage2_25[4], stage2_25[5]},
      {stage3_27[0],stage3_26[1],stage3_25[7],stage3_24[8],stage3_23[9]}
   );
   gpc606_5 gpc1244 (
      {stage2_23[36], stage2_23[37], stage2_23[38], stage2_23[39], stage2_23[40], stage2_23[41]},
      {stage2_25[6], stage2_25[7], stage2_25[8], stage2_25[9], stage2_25[10], stage2_25[11]},
      {stage3_27[1],stage3_26[2],stage3_25[8],stage3_24[9],stage3_23[10]}
   );
   gpc606_5 gpc1245 (
      {stage2_24[8], stage2_24[9], stage2_24[10], stage2_24[11], stage2_24[12], stage2_24[13]},
      {stage2_26[0], stage2_26[1], stage2_26[2], stage2_26[3], stage2_26[4], stage2_26[5]},
      {stage3_28[0],stage3_27[2],stage3_26[3],stage3_25[9],stage3_24[10]}
   );
   gpc606_5 gpc1246 (
      {stage2_24[14], stage2_24[15], stage2_24[16], stage2_24[17], stage2_24[18], stage2_24[19]},
      {stage2_26[6], stage2_26[7], stage2_26[8], stage2_26[9], stage2_26[10], stage2_26[11]},
      {stage3_28[1],stage3_27[3],stage3_26[4],stage3_25[10],stage3_24[11]}
   );
   gpc606_5 gpc1247 (
      {stage2_24[20], stage2_24[21], stage2_24[22], stage2_24[23], stage2_24[24], stage2_24[25]},
      {stage2_26[12], stage2_26[13], stage2_26[14], stage2_26[15], stage2_26[16], stage2_26[17]},
      {stage3_28[2],stage3_27[4],stage3_26[5],stage3_25[11],stage3_24[12]}
   );
   gpc606_5 gpc1248 (
      {stage2_24[26], stage2_24[27], stage2_24[28], stage2_24[29], stage2_24[30], stage2_24[31]},
      {stage2_26[18], stage2_26[19], stage2_26[20], stage2_26[21], stage2_26[22], stage2_26[23]},
      {stage3_28[3],stage3_27[5],stage3_26[6],stage3_25[12],stage3_24[13]}
   );
   gpc606_5 gpc1249 (
      {stage2_25[12], stage2_25[13], stage2_25[14], stage2_25[15], stage2_25[16], stage2_25[17]},
      {stage2_27[0], stage2_27[1], stage2_27[2], stage2_27[3], stage2_27[4], stage2_27[5]},
      {stage3_29[0],stage3_28[4],stage3_27[6],stage3_26[7],stage3_25[13]}
   );
   gpc606_5 gpc1250 (
      {stage2_25[18], stage2_25[19], stage2_25[20], stage2_25[21], stage2_25[22], stage2_25[23]},
      {stage2_27[6], stage2_27[7], stage2_27[8], stage2_27[9], stage2_27[10], stage2_27[11]},
      {stage3_29[1],stage3_28[5],stage3_27[7],stage3_26[8],stage3_25[14]}
   );
   gpc606_5 gpc1251 (
      {stage2_25[24], stage2_25[25], stage2_25[26], stage2_25[27], stage2_25[28], stage2_25[29]},
      {stage2_27[12], stage2_27[13], stage2_27[14], stage2_27[15], stage2_27[16], stage2_27[17]},
      {stage3_29[2],stage3_28[6],stage3_27[8],stage3_26[9],stage3_25[15]}
   );
   gpc606_5 gpc1252 (
      {stage2_26[24], stage2_26[25], stage2_26[26], stage2_26[27], stage2_26[28], stage2_26[29]},
      {stage2_28[0], stage2_28[1], stage2_28[2], stage2_28[3], stage2_28[4], stage2_28[5]},
      {stage3_30[0],stage3_29[3],stage3_28[7],stage3_27[9],stage3_26[10]}
   );
   gpc615_5 gpc1253 (
      {stage2_27[18], stage2_27[19], stage2_27[20], stage2_27[21], stage2_27[22]},
      {stage2_28[6]},
      {stage2_29[0], stage2_29[1], stage2_29[2], stage2_29[3], stage2_29[4], stage2_29[5]},
      {stage3_31[0],stage3_30[1],stage3_29[4],stage3_28[8],stage3_27[10]}
   );
   gpc615_5 gpc1254 (
      {stage2_27[23], stage2_27[24], stage2_27[25], stage2_27[26], stage2_27[27]},
      {stage2_28[7]},
      {stage2_29[6], stage2_29[7], stage2_29[8], stage2_29[9], stage2_29[10], stage2_29[11]},
      {stage3_31[1],stage3_30[2],stage3_29[5],stage3_28[9],stage3_27[11]}
   );
   gpc615_5 gpc1255 (
      {stage2_27[28], stage2_27[29], stage2_27[30], stage2_27[31], stage2_27[32]},
      {stage2_28[8]},
      {stage2_29[12], stage2_29[13], stage2_29[14], stage2_29[15], stage2_29[16], stage2_29[17]},
      {stage3_31[2],stage3_30[3],stage3_29[6],stage3_28[10],stage3_27[12]}
   );
   gpc135_4 gpc1256 (
      {stage2_28[9], stage2_28[10], stage2_28[11], stage2_28[12], stage2_28[13]},
      {stage2_29[18], stage2_29[19], stage2_29[20]},
      {stage2_30[0]},
      {stage3_31[3],stage3_30[4],stage3_29[7],stage3_28[11]}
   );
   gpc606_5 gpc1257 (
      {stage2_28[14], stage2_28[15], stage2_28[16], stage2_28[17], stage2_28[18], stage2_28[19]},
      {stage2_30[1], stage2_30[2], stage2_30[3], stage2_30[4], stage2_30[5], stage2_30[6]},
      {stage3_32[0],stage3_31[4],stage3_30[5],stage3_29[8],stage3_28[12]}
   );
   gpc606_5 gpc1258 (
      {stage2_29[21], stage2_29[22], stage2_29[23], stage2_29[24], stage2_29[25], stage2_29[26]},
      {stage2_31[0], stage2_31[1], stage2_31[2], stage2_31[3], stage2_31[4], stage2_31[5]},
      {stage3_33[0],stage3_32[1],stage3_31[5],stage3_30[6],stage3_29[9]}
   );
   gpc606_5 gpc1259 (
      {stage2_29[27], stage2_29[28], stage2_29[29], stage2_29[30], stage2_29[31], stage2_29[32]},
      {stage2_31[6], stage2_31[7], stage2_31[8], stage2_31[9], stage2_31[10], stage2_31[11]},
      {stage3_33[1],stage3_32[2],stage3_31[6],stage3_30[7],stage3_29[10]}
   );
   gpc615_5 gpc1260 (
      {stage2_30[7], stage2_30[8], stage2_30[9], stage2_30[10], stage2_30[11]},
      {stage2_31[12]},
      {stage2_32[0], stage2_32[1], stage2_32[2], stage2_32[3], stage2_32[4], stage2_32[5]},
      {stage3_34[0],stage3_33[2],stage3_32[3],stage3_31[7],stage3_30[8]}
   );
   gpc615_5 gpc1261 (
      {stage2_30[12], stage2_30[13], stage2_30[14], stage2_30[15], stage2_30[16]},
      {stage2_31[13]},
      {stage2_32[6], stage2_32[7], stage2_32[8], stage2_32[9], stage2_32[10], stage2_32[11]},
      {stage3_34[1],stage3_33[3],stage3_32[4],stage3_31[8],stage3_30[9]}
   );
   gpc615_5 gpc1262 (
      {stage2_30[17], stage2_30[18], stage2_30[19], stage2_30[20], stage2_30[21]},
      {stage2_31[14]},
      {stage2_32[12], stage2_32[13], stage2_32[14], stage2_32[15], stage2_32[16], stage2_32[17]},
      {stage3_34[2],stage3_33[4],stage3_32[5],stage3_31[9],stage3_30[10]}
   );
   gpc615_5 gpc1263 (
      {stage2_30[22], stage2_30[23], stage2_30[24], stage2_30[25], stage2_30[26]},
      {stage2_31[15]},
      {stage2_32[18], stage2_32[19], stage2_32[20], stage2_32[21], stage2_32[22], stage2_32[23]},
      {stage3_34[3],stage3_33[5],stage3_32[6],stage3_31[10],stage3_30[11]}
   );
   gpc615_5 gpc1264 (
      {stage2_30[27], stage2_30[28], stage2_30[29], stage2_30[30], stage2_30[31]},
      {stage2_31[16]},
      {stage2_32[24], stage2_32[25], stage2_32[26], stage2_32[27], stage2_32[28], stage2_32[29]},
      {stage3_34[4],stage3_33[6],stage3_32[7],stage3_31[11],stage3_30[12]}
   );
   gpc615_5 gpc1265 (
      {stage2_30[32], stage2_30[33], stage2_30[34], stage2_30[35], stage2_30[36]},
      {stage2_31[17]},
      {stage2_32[30], stage2_32[31], stage2_32[32], stage2_32[33], stage2_32[34], stage2_32[35]},
      {stage3_34[5],stage3_33[7],stage3_32[8],stage3_31[12],stage3_30[13]}
   );
   gpc606_5 gpc1266 (
      {stage2_31[18], stage2_31[19], stage2_31[20], stage2_31[21], stage2_31[22], stage2_31[23]},
      {stage2_33[0], stage2_33[1], stage2_33[2], stage2_33[3], stage2_33[4], stage2_33[5]},
      {stage3_35[0],stage3_34[6],stage3_33[8],stage3_32[9],stage3_31[13]}
   );
   gpc606_5 gpc1267 (
      {stage2_31[24], stage2_31[25], stage2_31[26], stage2_31[27], stage2_31[28], stage2_31[29]},
      {stage2_33[6], stage2_33[7], stage2_33[8], stage2_33[9], stage2_33[10], stage2_33[11]},
      {stage3_35[1],stage3_34[7],stage3_33[9],stage3_32[10],stage3_31[14]}
   );
   gpc615_5 gpc1268 (
      {stage2_31[30], stage2_31[31], stage2_31[32], stage2_31[33], stage2_31[34]},
      {stage2_32[36]},
      {stage2_33[12], stage2_33[13], stage2_33[14], stage2_33[15], stage2_33[16], stage2_33[17]},
      {stage3_35[2],stage3_34[8],stage3_33[10],stage3_32[11],stage3_31[15]}
   );
   gpc1_1 gpc1269 (
      {stage2_0[5]},
      {stage3_0[1]}
   );
   gpc1_1 gpc1270 (
      {stage2_0[6]},
      {stage3_0[2]}
   );
   gpc1_1 gpc1271 (
      {stage2_0[7]},
      {stage3_0[3]}
   );
   gpc1_1 gpc1272 (
      {stage2_0[8]},
      {stage3_0[4]}
   );
   gpc1_1 gpc1273 (
      {stage2_0[9]},
      {stage3_0[5]}
   );
   gpc1_1 gpc1274 (
      {stage2_0[10]},
      {stage3_0[6]}
   );
   gpc1_1 gpc1275 (
      {stage2_1[9]},
      {stage3_1[2]}
   );
   gpc1_1 gpc1276 (
      {stage2_1[10]},
      {stage3_1[3]}
   );
   gpc1_1 gpc1277 (
      {stage2_1[11]},
      {stage3_1[4]}
   );
   gpc1_1 gpc1278 (
      {stage2_1[12]},
      {stage3_1[5]}
   );
   gpc1_1 gpc1279 (
      {stage2_1[13]},
      {stage3_1[6]}
   );
   gpc1_1 gpc1280 (
      {stage2_1[14]},
      {stage3_1[7]}
   );
   gpc1_1 gpc1281 (
      {stage2_1[15]},
      {stage3_1[8]}
   );
   gpc1_1 gpc1282 (
      {stage2_1[16]},
      {stage3_1[9]}
   );
   gpc1_1 gpc1283 (
      {stage2_2[11]},
      {stage3_2[4]}
   );
   gpc1_1 gpc1284 (
      {stage2_2[12]},
      {stage3_2[5]}
   );
   gpc1_1 gpc1285 (
      {stage2_2[13]},
      {stage3_2[6]}
   );
   gpc1_1 gpc1286 (
      {stage2_2[14]},
      {stage3_2[7]}
   );
   gpc1_1 gpc1287 (
      {stage2_2[15]},
      {stage3_2[8]}
   );
   gpc1_1 gpc1288 (
      {stage2_2[16]},
      {stage3_2[9]}
   );
   gpc1_1 gpc1289 (
      {stage2_3[20]},
      {stage3_3[8]}
   );
   gpc1_1 gpc1290 (
      {stage2_3[21]},
      {stage3_3[9]}
   );
   gpc1_1 gpc1291 (
      {stage2_3[22]},
      {stage3_3[10]}
   );
   gpc1_1 gpc1292 (
      {stage2_3[23]},
      {stage3_3[11]}
   );
   gpc1_1 gpc1293 (
      {stage2_3[24]},
      {stage3_3[12]}
   );
   gpc1_1 gpc1294 (
      {stage2_3[25]},
      {stage3_3[13]}
   );
   gpc1_1 gpc1295 (
      {stage2_3[26]},
      {stage3_3[14]}
   );
   gpc1_1 gpc1296 (
      {stage2_3[27]},
      {stage3_3[15]}
   );
   gpc1_1 gpc1297 (
      {stage2_3[28]},
      {stage3_3[16]}
   );
   gpc1_1 gpc1298 (
      {stage2_3[29]},
      {stage3_3[17]}
   );
   gpc1_1 gpc1299 (
      {stage2_3[30]},
      {stage3_3[18]}
   );
   gpc1_1 gpc1300 (
      {stage2_3[31]},
      {stage3_3[19]}
   );
   gpc1_1 gpc1301 (
      {stage2_3[32]},
      {stage3_3[20]}
   );
   gpc1_1 gpc1302 (
      {stage2_3[33]},
      {stage3_3[21]}
   );
   gpc1_1 gpc1303 (
      {stage2_3[34]},
      {stage3_3[22]}
   );
   gpc1_1 gpc1304 (
      {stage2_6[27]},
      {stage3_6[13]}
   );
   gpc1_1 gpc1305 (
      {stage2_6[28]},
      {stage3_6[14]}
   );
   gpc1_1 gpc1306 (
      {stage2_6[29]},
      {stage3_6[15]}
   );
   gpc1_1 gpc1307 (
      {stage2_6[30]},
      {stage3_6[16]}
   );
   gpc1_1 gpc1308 (
      {stage2_7[28]},
      {stage3_7[13]}
   );
   gpc1_1 gpc1309 (
      {stage2_7[29]},
      {stage3_7[14]}
   );
   gpc1_1 gpc1310 (
      {stage2_7[30]},
      {stage3_7[15]}
   );
   gpc1_1 gpc1311 (
      {stage2_7[31]},
      {stage3_7[16]}
   );
   gpc1_1 gpc1312 (
      {stage2_7[32]},
      {stage3_7[17]}
   );
   gpc1_1 gpc1313 (
      {stage2_7[33]},
      {stage3_7[18]}
   );
   gpc1_1 gpc1314 (
      {stage2_8[26]},
      {stage3_8[11]}
   );
   gpc1_1 gpc1315 (
      {stage2_8[27]},
      {stage3_8[12]}
   );
   gpc1_1 gpc1316 (
      {stage2_8[28]},
      {stage3_8[13]}
   );
   gpc1_1 gpc1317 (
      {stage2_8[29]},
      {stage3_8[14]}
   );
   gpc1_1 gpc1318 (
      {stage2_8[30]},
      {stage3_8[15]}
   );
   gpc1_1 gpc1319 (
      {stage2_8[31]},
      {stage3_8[16]}
   );
   gpc1_1 gpc1320 (
      {stage2_8[32]},
      {stage3_8[17]}
   );
   gpc1_1 gpc1321 (
      {stage2_9[27]},
      {stage3_9[14]}
   );
   gpc1_1 gpc1322 (
      {stage2_9[28]},
      {stage3_9[15]}
   );
   gpc1_1 gpc1323 (
      {stage2_9[29]},
      {stage3_9[16]}
   );
   gpc1_1 gpc1324 (
      {stage2_9[30]},
      {stage3_9[17]}
   );
   gpc1_1 gpc1325 (
      {stage2_9[31]},
      {stage3_9[18]}
   );
   gpc1_1 gpc1326 (
      {stage2_10[44]},
      {stage3_10[13]}
   );
   gpc1_1 gpc1327 (
      {stage2_10[45]},
      {stage3_10[14]}
   );
   gpc1_1 gpc1328 (
      {stage2_12[23]},
      {stage3_12[14]}
   );
   gpc1_1 gpc1329 (
      {stage2_13[42]},
      {stage3_13[15]}
   );
   gpc1_1 gpc1330 (
      {stage2_13[43]},
      {stage3_13[16]}
   );
   gpc1_1 gpc1331 (
      {stage2_13[44]},
      {stage3_13[17]}
   );
   gpc1_1 gpc1332 (
      {stage2_14[36]},
      {stage3_14[16]}
   );
   gpc1_1 gpc1333 (
      {stage2_17[36]},
      {stage3_17[16]}
   );
   gpc1_1 gpc1334 (
      {stage2_20[31]},
      {stage3_20[11]}
   );
   gpc1_1 gpc1335 (
      {stage2_20[32]},
      {stage3_20[12]}
   );
   gpc1_1 gpc1336 (
      {stage2_20[33]},
      {stage3_20[13]}
   );
   gpc1_1 gpc1337 (
      {stage2_20[34]},
      {stage3_20[14]}
   );
   gpc1_1 gpc1338 (
      {stage2_20[35]},
      {stage3_20[15]}
   );
   gpc1_1 gpc1339 (
      {stage2_20[36]},
      {stage3_20[16]}
   );
   gpc1_1 gpc1340 (
      {stage2_20[37]},
      {stage3_20[17]}
   );
   gpc1_1 gpc1341 (
      {stage2_22[24]},
      {stage3_22[13]}
   );
   gpc1_1 gpc1342 (
      {stage2_22[25]},
      {stage3_22[14]}
   );
   gpc1_1 gpc1343 (
      {stage2_22[26]},
      {stage3_22[15]}
   );
   gpc1_1 gpc1344 (
      {stage2_22[27]},
      {stage3_22[16]}
   );
   gpc1_1 gpc1345 (
      {stage2_22[28]},
      {stage3_22[17]}
   );
   gpc1_1 gpc1346 (
      {stage2_22[29]},
      {stage3_22[18]}
   );
   gpc1_1 gpc1347 (
      {stage2_22[30]},
      {stage3_22[19]}
   );
   gpc1_1 gpc1348 (
      {stage2_22[31]},
      {stage3_22[20]}
   );
   gpc1_1 gpc1349 (
      {stage2_22[32]},
      {stage3_22[21]}
   );
   gpc1_1 gpc1350 (
      {stage2_22[33]},
      {stage3_22[22]}
   );
   gpc1_1 gpc1351 (
      {stage2_23[42]},
      {stage3_23[11]}
   );
   gpc1_1 gpc1352 (
      {stage2_23[43]},
      {stage3_23[12]}
   );
   gpc1_1 gpc1353 (
      {stage2_24[32]},
      {stage3_24[14]}
   );
   gpc1_1 gpc1354 (
      {stage2_24[33]},
      {stage3_24[15]}
   );
   gpc1_1 gpc1355 (
      {stage2_24[34]},
      {stage3_24[16]}
   );
   gpc1_1 gpc1356 (
      {stage2_25[30]},
      {stage3_25[16]}
   );
   gpc1_1 gpc1357 (
      {stage2_26[30]},
      {stage3_26[11]}
   );
   gpc1_1 gpc1358 (
      {stage2_28[20]},
      {stage3_28[13]}
   );
   gpc1_1 gpc1359 (
      {stage2_28[21]},
      {stage3_28[14]}
   );
   gpc1_1 gpc1360 (
      {stage2_28[22]},
      {stage3_28[15]}
   );
   gpc1_1 gpc1361 (
      {stage2_28[23]},
      {stage3_28[16]}
   );
   gpc1_1 gpc1362 (
      {stage2_28[24]},
      {stage3_28[17]}
   );
   gpc1_1 gpc1363 (
      {stage2_28[25]},
      {stage3_28[18]}
   );
   gpc1_1 gpc1364 (
      {stage2_28[26]},
      {stage3_28[19]}
   );
   gpc1_1 gpc1365 (
      {stage2_28[27]},
      {stage3_28[20]}
   );
   gpc1_1 gpc1366 (
      {stage2_28[28]},
      {stage3_28[21]}
   );
   gpc1_1 gpc1367 (
      {stage2_28[29]},
      {stage3_28[22]}
   );
   gpc1_1 gpc1368 (
      {stage2_31[35]},
      {stage3_31[16]}
   );
   gpc1_1 gpc1369 (
      {stage2_32[37]},
      {stage3_32[12]}
   );
   gpc1_1 gpc1370 (
      {stage2_32[38]},
      {stage3_32[13]}
   );
   gpc1_1 gpc1371 (
      {stage2_32[39]},
      {stage3_32[14]}
   );
   gpc1_1 gpc1372 (
      {stage2_32[40]},
      {stage3_32[15]}
   );
   gpc1_1 gpc1373 (
      {stage2_33[18]},
      {stage3_33[11]}
   );
   gpc1_1 gpc1374 (
      {stage2_33[19]},
      {stage3_33[12]}
   );
   gpc1_1 gpc1375 (
      {stage2_33[20]},
      {stage3_33[13]}
   );
   gpc1_1 gpc1376 (
      {stage2_33[21]},
      {stage3_33[14]}
   );
   gpc1_1 gpc1377 (
      {stage2_33[22]},
      {stage3_33[15]}
   );
   gpc1_1 gpc1378 (
      {stage2_33[23]},
      {stage3_33[16]}
   );
   gpc1_1 gpc1379 (
      {stage2_34[0]},
      {stage3_34[9]}
   );
   gpc1_1 gpc1380 (
      {stage2_34[1]},
      {stage3_34[10]}
   );
   gpc1_1 gpc1381 (
      {stage2_34[2]},
      {stage3_34[11]}
   );
   gpc1_1 gpc1382 (
      {stage2_34[3]},
      {stage3_34[12]}
   );
   gpc1_1 gpc1383 (
      {stage2_34[4]},
      {stage3_34[13]}
   );
   gpc1_1 gpc1384 (
      {stage2_34[5]},
      {stage3_34[14]}
   );
   gpc1_1 gpc1385 (
      {stage2_34[6]},
      {stage3_34[15]}
   );
   gpc1_1 gpc1386 (
      {stage2_35[0]},
      {stage3_35[3]}
   );
   gpc1_1 gpc1387 (
      {stage2_35[1]},
      {stage3_35[4]}
   );
   gpc606_5 gpc1388 (
      {stage3_0[0], stage3_0[1], stage3_0[2], stage3_0[3], stage3_0[4], stage3_0[5]},
      {stage3_2[0], stage3_2[1], stage3_2[2], stage3_2[3], stage3_2[4], stage3_2[5]},
      {stage4_4[0],stage4_3[0],stage4_2[0],stage4_1[0],stage4_0[0]}
   );
   gpc606_5 gpc1389 (
      {stage3_1[0], stage3_1[1], stage3_1[2], stage3_1[3], stage3_1[4], stage3_1[5]},
      {stage3_3[0], stage3_3[1], stage3_3[2], stage3_3[3], stage3_3[4], stage3_3[5]},
      {stage4_5[0],stage4_4[1],stage4_3[1],stage4_2[1],stage4_1[1]}
   );
   gpc615_5 gpc1390 (
      {stage3_3[6], stage3_3[7], stage3_3[8], stage3_3[9], stage3_3[10]},
      {stage3_4[0]},
      {stage3_5[0], stage3_5[1], stage3_5[2], stage3_5[3], stage3_5[4], stage3_5[5]},
      {stage4_7[0],stage4_6[0],stage4_5[1],stage4_4[2],stage4_3[2]}
   );
   gpc615_5 gpc1391 (
      {stage3_3[11], stage3_3[12], stage3_3[13], stage3_3[14], stage3_3[15]},
      {stage3_4[1]},
      {stage3_5[6], stage3_5[7], stage3_5[8], stage3_5[9], stage3_5[10], stage3_5[11]},
      {stage4_7[1],stage4_6[1],stage4_5[2],stage4_4[3],stage4_3[3]}
   );
   gpc606_5 gpc1392 (
      {stage3_4[2], stage3_4[3], stage3_4[4], stage3_4[5], stage3_4[6], stage3_4[7]},
      {stage3_6[0], stage3_6[1], stage3_6[2], stage3_6[3], stage3_6[4], stage3_6[5]},
      {stage4_8[0],stage4_7[2],stage4_6[2],stage4_5[3],stage4_4[4]}
   );
   gpc615_5 gpc1393 (
      {stage3_6[6], stage3_6[7], stage3_6[8], stage3_6[9], stage3_6[10]},
      {stage3_7[0]},
      {stage3_8[0], stage3_8[1], stage3_8[2], stage3_8[3], stage3_8[4], stage3_8[5]},
      {stage4_10[0],stage4_9[0],stage4_8[1],stage4_7[3],stage4_6[3]}
   );
   gpc615_5 gpc1394 (
      {stage3_6[11], stage3_6[12], stage3_6[13], stage3_6[14], stage3_6[15]},
      {stage3_7[1]},
      {stage3_8[6], stage3_8[7], stage3_8[8], stage3_8[9], stage3_8[10], stage3_8[11]},
      {stage4_10[1],stage4_9[1],stage4_8[2],stage4_7[4],stage4_6[4]}
   );
   gpc1406_5 gpc1395 (
      {stage3_7[2], stage3_7[3], stage3_7[4], stage3_7[5], stage3_7[6], stage3_7[7]},
      {stage3_9[0], stage3_9[1], stage3_9[2], stage3_9[3]},
      {stage3_10[0]},
      {stage4_11[0],stage4_10[2],stage4_9[2],stage4_8[3],stage4_7[5]}
   );
   gpc606_5 gpc1396 (
      {stage3_7[8], stage3_7[9], stage3_7[10], stage3_7[11], stage3_7[12], stage3_7[13]},
      {stage3_9[4], stage3_9[5], stage3_9[6], stage3_9[7], stage3_9[8], stage3_9[9]},
      {stage4_11[1],stage4_10[3],stage4_9[3],stage4_8[4],stage4_7[6]}
   );
   gpc615_5 gpc1397 (
      {stage3_7[14], stage3_7[15], stage3_7[16], stage3_7[17], stage3_7[18]},
      {stage3_8[12]},
      {stage3_9[10], stage3_9[11], stage3_9[12], stage3_9[13], stage3_9[14], stage3_9[15]},
      {stage4_11[2],stage4_10[4],stage4_9[4],stage4_8[5],stage4_7[7]}
   );
   gpc615_5 gpc1398 (
      {stage3_8[13], stage3_8[14], stage3_8[15], stage3_8[16], stage3_8[17]},
      {stage3_9[16]},
      {stage3_10[1], stage3_10[2], stage3_10[3], stage3_10[4], stage3_10[5], stage3_10[6]},
      {stage4_12[0],stage4_11[3],stage4_10[5],stage4_9[5],stage4_8[6]}
   );
   gpc7_3 gpc1399 (
      {stage3_10[7], stage3_10[8], stage3_10[9], stage3_10[10], stage3_10[11], stage3_10[12], stage3_10[13]},
      {stage4_12[1],stage4_11[4],stage4_10[6]}
   );
   gpc606_5 gpc1400 (
      {stage3_11[0], stage3_11[1], stage3_11[2], stage3_11[3], stage3_11[4], stage3_11[5]},
      {stage3_13[0], stage3_13[1], stage3_13[2], stage3_13[3], stage3_13[4], stage3_13[5]},
      {stage4_15[0],stage4_14[0],stage4_13[0],stage4_12[2],stage4_11[5]}
   );
   gpc606_5 gpc1401 (
      {stage3_11[6], stage3_11[7], stage3_11[8], stage3_11[9], stage3_11[10], stage3_11[11]},
      {stage3_13[6], stage3_13[7], stage3_13[8], stage3_13[9], stage3_13[10], stage3_13[11]},
      {stage4_15[1],stage4_14[1],stage4_13[1],stage4_12[3],stage4_11[6]}
   );
   gpc606_5 gpc1402 (
      {stage3_12[0], stage3_12[1], stage3_12[2], stage3_12[3], stage3_12[4], stage3_12[5]},
      {stage3_14[0], stage3_14[1], stage3_14[2], stage3_14[3], stage3_14[4], stage3_14[5]},
      {stage4_16[0],stage4_15[2],stage4_14[2],stage4_13[2],stage4_12[4]}
   );
   gpc606_5 gpc1403 (
      {stage3_12[6], stage3_12[7], stage3_12[8], stage3_12[9], stage3_12[10], stage3_12[11]},
      {stage3_14[6], stage3_14[7], stage3_14[8], stage3_14[9], stage3_14[10], stage3_14[11]},
      {stage4_16[1],stage4_15[3],stage4_14[3],stage4_13[3],stage4_12[5]}
   );
   gpc606_5 gpc1404 (
      {stage3_13[12], stage3_13[13], stage3_13[14], stage3_13[15], stage3_13[16], stage3_13[17]},
      {stage3_15[0], stage3_15[1], stage3_15[2], stage3_15[3], stage3_15[4], stage3_15[5]},
      {stage4_17[0],stage4_16[2],stage4_15[4],stage4_14[4],stage4_13[4]}
   );
   gpc615_5 gpc1405 (
      {stage3_14[12], stage3_14[13], stage3_14[14], stage3_14[15], stage3_14[16]},
      {stage3_15[6]},
      {stage3_16[0], stage3_16[1], stage3_16[2], stage3_16[3], stage3_16[4], stage3_16[5]},
      {stage4_18[0],stage4_17[1],stage4_16[3],stage4_15[5],stage4_14[5]}
   );
   gpc606_5 gpc1406 (
      {stage3_15[7], stage3_15[8], stage3_15[9], stage3_15[10], stage3_15[11], stage3_15[12]},
      {stage3_17[0], stage3_17[1], stage3_17[2], stage3_17[3], stage3_17[4], stage3_17[5]},
      {stage4_19[0],stage4_18[1],stage4_17[2],stage4_16[4],stage4_15[6]}
   );
   gpc606_5 gpc1407 (
      {stage3_16[6], stage3_16[7], stage3_16[8], stage3_16[9], stage3_16[10], stage3_16[11]},
      {stage3_18[0], stage3_18[1], stage3_18[2], stage3_18[3], stage3_18[4], stage3_18[5]},
      {stage4_20[0],stage4_19[1],stage4_18[2],stage4_17[3],stage4_16[5]}
   );
   gpc1163_5 gpc1408 (
      {stage3_17[6], stage3_17[7], stage3_17[8]},
      {stage3_18[6], stage3_18[7], stage3_18[8], stage3_18[9], stage3_18[10], stage3_18[11]},
      {stage3_19[0]},
      {stage3_20[0]},
      {stage4_21[0],stage4_20[1],stage4_19[2],stage4_18[3],stage4_17[4]}
   );
   gpc1343_5 gpc1409 (
      {stage3_19[1], stage3_19[2], stage3_19[3]},
      {stage3_20[1], stage3_20[2], stage3_20[3], stage3_20[4]},
      {stage3_21[0], stage3_21[1], stage3_21[2]},
      {stage3_22[0]},
      {stage4_23[0],stage4_22[0],stage4_21[1],stage4_20[2],stage4_19[3]}
   );
   gpc606_5 gpc1410 (
      {stage3_20[5], stage3_20[6], stage3_20[7], stage3_20[8], stage3_20[9], stage3_20[10]},
      {stage3_22[1], stage3_22[2], stage3_22[3], stage3_22[4], stage3_22[5], stage3_22[6]},
      {stage4_24[0],stage4_23[1],stage4_22[1],stage4_21[2],stage4_20[3]}
   );
   gpc606_5 gpc1411 (
      {stage3_20[11], stage3_20[12], stage3_20[13], stage3_20[14], stage3_20[15], stage3_20[16]},
      {stage3_22[7], stage3_22[8], stage3_22[9], stage3_22[10], stage3_22[11], stage3_22[12]},
      {stage4_24[1],stage4_23[2],stage4_22[2],stage4_21[3],stage4_20[4]}
   );
   gpc606_5 gpc1412 (
      {stage3_21[3], stage3_21[4], stage3_21[5], stage3_21[6], stage3_21[7], stage3_21[8]},
      {stage3_23[0], stage3_23[1], stage3_23[2], stage3_23[3], stage3_23[4], stage3_23[5]},
      {stage4_25[0],stage4_24[2],stage4_23[3],stage4_22[3],stage4_21[4]}
   );
   gpc606_5 gpc1413 (
      {stage3_21[9], stage3_21[10], stage3_21[11], stage3_21[12], stage3_21[13], stage3_21[14]},
      {stage3_23[6], stage3_23[7], stage3_23[8], stage3_23[9], stage3_23[10], stage3_23[11]},
      {stage4_25[1],stage4_24[3],stage4_23[4],stage4_22[4],stage4_21[5]}
   );
   gpc207_4 gpc1414 (
      {stage3_22[13], stage3_22[14], stage3_22[15], stage3_22[16], stage3_22[17], stage3_22[18], stage3_22[19]},
      {stage3_24[0], stage3_24[1]},
      {stage4_25[2],stage4_24[4],stage4_23[5],stage4_22[5]}
   );
   gpc2135_5 gpc1415 (
      {stage3_24[2], stage3_24[3], stage3_24[4], stage3_24[5], stage3_24[6]},
      {stage3_25[0], stage3_25[1], stage3_25[2]},
      {stage3_26[0]},
      {stage3_27[0], stage3_27[1]},
      {stage4_28[0],stage4_27[0],stage4_26[0],stage4_25[3],stage4_24[5]}
   );
   gpc2135_5 gpc1416 (
      {stage3_24[7], stage3_24[8], stage3_24[9], stage3_24[10], stage3_24[11]},
      {stage3_25[3], stage3_25[4], stage3_25[5]},
      {stage3_26[1]},
      {stage3_27[2], stage3_27[3]},
      {stage4_28[1],stage4_27[1],stage4_26[1],stage4_25[4],stage4_24[6]}
   );
   gpc2135_5 gpc1417 (
      {stage3_24[12], stage3_24[13], stage3_24[14], stage3_24[15], stage3_24[16]},
      {stage3_25[6], stage3_25[7], stage3_25[8]},
      {stage3_26[2]},
      {stage3_27[4], stage3_27[5]},
      {stage4_28[2],stage4_27[2],stage4_26[2],stage4_25[5],stage4_24[7]}
   );
   gpc606_5 gpc1418 (
      {stage3_25[9], stage3_25[10], stage3_25[11], stage3_25[12], stage3_25[13], stage3_25[14]},
      {stage3_27[6], stage3_27[7], stage3_27[8], stage3_27[9], stage3_27[10], stage3_27[11]},
      {stage4_29[0],stage4_28[3],stage4_27[3],stage4_26[3],stage4_25[6]}
   );
   gpc615_5 gpc1419 (
      {stage3_26[3], stage3_26[4], stage3_26[5], stage3_26[6], stage3_26[7]},
      {stage3_27[12]},
      {stage3_28[0], stage3_28[1], stage3_28[2], stage3_28[3], stage3_28[4], stage3_28[5]},
      {stage4_30[0],stage4_29[1],stage4_28[4],stage4_27[4],stage4_26[4]}
   );
   gpc2135_5 gpc1420 (
      {stage3_28[6], stage3_28[7], stage3_28[8], stage3_28[9], stage3_28[10]},
      {stage3_29[0], stage3_29[1], stage3_29[2]},
      {stage3_30[0]},
      {stage3_31[0], stage3_31[1]},
      {stage4_32[0],stage4_31[0],stage4_30[1],stage4_29[2],stage4_28[5]}
   );
   gpc2135_5 gpc1421 (
      {stage3_28[11], stage3_28[12], stage3_28[13], stage3_28[14], stage3_28[15]},
      {stage3_29[3], stage3_29[4], stage3_29[5]},
      {stage3_30[1]},
      {stage3_31[2], stage3_31[3]},
      {stage4_32[1],stage4_31[1],stage4_30[2],stage4_29[3],stage4_28[6]}
   );
   gpc606_5 gpc1422 (
      {stage3_28[16], stage3_28[17], stage3_28[18], stage3_28[19], stage3_28[20], stage3_28[21]},
      {stage3_30[2], stage3_30[3], stage3_30[4], stage3_30[5], stage3_30[6], stage3_30[7]},
      {stage4_32[2],stage4_31[2],stage4_30[3],stage4_29[4],stage4_28[7]}
   );
   gpc615_5 gpc1423 (
      {stage3_29[6], stage3_29[7], stage3_29[8], stage3_29[9], stage3_29[10]},
      {stage3_30[8]},
      {stage3_31[4], stage3_31[5], stage3_31[6], stage3_31[7], stage3_31[8], stage3_31[9]},
      {stage4_33[0],stage4_32[3],stage4_31[3],stage4_30[4],stage4_29[5]}
   );
   gpc615_5 gpc1424 (
      {stage3_30[9], stage3_30[10], stage3_30[11], stage3_30[12], stage3_30[13]},
      {stage3_31[10]},
      {stage3_32[0], stage3_32[1], stage3_32[2], stage3_32[3], stage3_32[4], stage3_32[5]},
      {stage4_34[0],stage4_33[1],stage4_32[4],stage4_31[4],stage4_30[5]}
   );
   gpc606_5 gpc1425 (
      {stage3_31[11], stage3_31[12], stage3_31[13], stage3_31[14], stage3_31[15], stage3_31[16]},
      {stage3_33[0], stage3_33[1], stage3_33[2], stage3_33[3], stage3_33[4], stage3_33[5]},
      {stage4_35[0],stage4_34[1],stage4_33[2],stage4_32[5],stage4_31[5]}
   );
   gpc606_5 gpc1426 (
      {stage3_32[6], stage3_32[7], stage3_32[8], stage3_32[9], stage3_32[10], stage3_32[11]},
      {stage3_34[0], stage3_34[1], stage3_34[2], stage3_34[3], stage3_34[4], stage3_34[5]},
      {stage4_36[0],stage4_35[1],stage4_34[2],stage4_33[3],stage4_32[6]}
   );
   gpc1163_5 gpc1427 (
      {stage3_33[6], stage3_33[7], stage3_33[8]},
      {stage3_34[6], stage3_34[7], stage3_34[8], stage3_34[9], stage3_34[10], stage3_34[11]},
      {stage3_35[0]},
      {1'b0},
      {stage4_37[0],stage4_36[1],stage4_35[2],stage4_34[3],stage4_33[4]}
   );
   gpc606_5 gpc1428 (
      {stage3_33[9], stage3_33[10], stage3_33[11], stage3_33[12], stage3_33[13], stage3_33[14]},
      {stage3_35[1], stage3_35[2], stage3_35[3], stage3_35[4], 1'b0, 1'b0},
      {stage4_37[1],stage4_36[2],stage4_35[3],stage4_34[4],stage4_33[5]}
   );
   gpc1_1 gpc1429 (
      {stage3_0[6]},
      {stage4_0[1]}
   );
   gpc1_1 gpc1430 (
      {stage3_1[6]},
      {stage4_1[2]}
   );
   gpc1_1 gpc1431 (
      {stage3_1[7]},
      {stage4_1[3]}
   );
   gpc1_1 gpc1432 (
      {stage3_1[8]},
      {stage4_1[4]}
   );
   gpc1_1 gpc1433 (
      {stage3_1[9]},
      {stage4_1[5]}
   );
   gpc1_1 gpc1434 (
      {stage3_2[6]},
      {stage4_2[2]}
   );
   gpc1_1 gpc1435 (
      {stage3_2[7]},
      {stage4_2[3]}
   );
   gpc1_1 gpc1436 (
      {stage3_2[8]},
      {stage4_2[4]}
   );
   gpc1_1 gpc1437 (
      {stage3_2[9]},
      {stage4_2[5]}
   );
   gpc1_1 gpc1438 (
      {stage3_3[16]},
      {stage4_3[4]}
   );
   gpc1_1 gpc1439 (
      {stage3_3[17]},
      {stage4_3[5]}
   );
   gpc1_1 gpc1440 (
      {stage3_3[18]},
      {stage4_3[6]}
   );
   gpc1_1 gpc1441 (
      {stage3_3[19]},
      {stage4_3[7]}
   );
   gpc1_1 gpc1442 (
      {stage3_3[20]},
      {stage4_3[8]}
   );
   gpc1_1 gpc1443 (
      {stage3_3[21]},
      {stage4_3[9]}
   );
   gpc1_1 gpc1444 (
      {stage3_3[22]},
      {stage4_3[10]}
   );
   gpc1_1 gpc1445 (
      {stage3_4[8]},
      {stage4_4[5]}
   );
   gpc1_1 gpc1446 (
      {stage3_6[16]},
      {stage4_6[5]}
   );
   gpc1_1 gpc1447 (
      {stage3_9[17]},
      {stage4_9[6]}
   );
   gpc1_1 gpc1448 (
      {stage3_9[18]},
      {stage4_9[7]}
   );
   gpc1_1 gpc1449 (
      {stage3_10[14]},
      {stage4_10[7]}
   );
   gpc1_1 gpc1450 (
      {stage3_11[12]},
      {stage4_11[7]}
   );
   gpc1_1 gpc1451 (
      {stage3_11[13]},
      {stage4_11[8]}
   );
   gpc1_1 gpc1452 (
      {stage3_11[14]},
      {stage4_11[9]}
   );
   gpc1_1 gpc1453 (
      {stage3_12[12]},
      {stage4_12[6]}
   );
   gpc1_1 gpc1454 (
      {stage3_12[13]},
      {stage4_12[7]}
   );
   gpc1_1 gpc1455 (
      {stage3_12[14]},
      {stage4_12[8]}
   );
   gpc1_1 gpc1456 (
      {stage3_15[13]},
      {stage4_15[7]}
   );
   gpc1_1 gpc1457 (
      {stage3_15[14]},
      {stage4_15[8]}
   );
   gpc1_1 gpc1458 (
      {stage3_15[15]},
      {stage4_15[9]}
   );
   gpc1_1 gpc1459 (
      {stage3_16[12]},
      {stage4_16[6]}
   );
   gpc1_1 gpc1460 (
      {stage3_17[9]},
      {stage4_17[5]}
   );
   gpc1_1 gpc1461 (
      {stage3_17[10]},
      {stage4_17[6]}
   );
   gpc1_1 gpc1462 (
      {stage3_17[11]},
      {stage4_17[7]}
   );
   gpc1_1 gpc1463 (
      {stage3_17[12]},
      {stage4_17[8]}
   );
   gpc1_1 gpc1464 (
      {stage3_17[13]},
      {stage4_17[9]}
   );
   gpc1_1 gpc1465 (
      {stage3_17[14]},
      {stage4_17[10]}
   );
   gpc1_1 gpc1466 (
      {stage3_17[15]},
      {stage4_17[11]}
   );
   gpc1_1 gpc1467 (
      {stage3_17[16]},
      {stage4_17[12]}
   );
   gpc1_1 gpc1468 (
      {stage3_18[12]},
      {stage4_18[4]}
   );
   gpc1_1 gpc1469 (
      {stage3_18[13]},
      {stage4_18[5]}
   );
   gpc1_1 gpc1470 (
      {stage3_18[14]},
      {stage4_18[6]}
   );
   gpc1_1 gpc1471 (
      {stage3_18[15]},
      {stage4_18[7]}
   );
   gpc1_1 gpc1472 (
      {stage3_18[16]},
      {stage4_18[8]}
   );
   gpc1_1 gpc1473 (
      {stage3_19[4]},
      {stage4_19[4]}
   );
   gpc1_1 gpc1474 (
      {stage3_19[5]},
      {stage4_19[5]}
   );
   gpc1_1 gpc1475 (
      {stage3_19[6]},
      {stage4_19[6]}
   );
   gpc1_1 gpc1476 (
      {stage3_19[7]},
      {stage4_19[7]}
   );
   gpc1_1 gpc1477 (
      {stage3_19[8]},
      {stage4_19[8]}
   );
   gpc1_1 gpc1478 (
      {stage3_19[9]},
      {stage4_19[9]}
   );
   gpc1_1 gpc1479 (
      {stage3_19[10]},
      {stage4_19[10]}
   );
   gpc1_1 gpc1480 (
      {stage3_19[11]},
      {stage4_19[11]}
   );
   gpc1_1 gpc1481 (
      {stage3_20[17]},
      {stage4_20[5]}
   );
   gpc1_1 gpc1482 (
      {stage3_22[20]},
      {stage4_22[6]}
   );
   gpc1_1 gpc1483 (
      {stage3_22[21]},
      {stage4_22[7]}
   );
   gpc1_1 gpc1484 (
      {stage3_22[22]},
      {stage4_22[8]}
   );
   gpc1_1 gpc1485 (
      {stage3_23[12]},
      {stage4_23[6]}
   );
   gpc1_1 gpc1486 (
      {stage3_25[15]},
      {stage4_25[7]}
   );
   gpc1_1 gpc1487 (
      {stage3_25[16]},
      {stage4_25[8]}
   );
   gpc1_1 gpc1488 (
      {stage3_26[8]},
      {stage4_26[5]}
   );
   gpc1_1 gpc1489 (
      {stage3_26[9]},
      {stage4_26[6]}
   );
   gpc1_1 gpc1490 (
      {stage3_26[10]},
      {stage4_26[7]}
   );
   gpc1_1 gpc1491 (
      {stage3_26[11]},
      {stage4_26[8]}
   );
   gpc1_1 gpc1492 (
      {stage3_28[22]},
      {stage4_28[8]}
   );
   gpc1_1 gpc1493 (
      {stage3_32[12]},
      {stage4_32[7]}
   );
   gpc1_1 gpc1494 (
      {stage3_32[13]},
      {stage4_32[8]}
   );
   gpc1_1 gpc1495 (
      {stage3_32[14]},
      {stage4_32[9]}
   );
   gpc1_1 gpc1496 (
      {stage3_32[15]},
      {stage4_32[10]}
   );
   gpc1_1 gpc1497 (
      {stage3_33[15]},
      {stage4_33[6]}
   );
   gpc1_1 gpc1498 (
      {stage3_33[16]},
      {stage4_33[7]}
   );
   gpc1_1 gpc1499 (
      {stage3_34[12]},
      {stage4_34[5]}
   );
   gpc1_1 gpc1500 (
      {stage3_34[13]},
      {stage4_34[6]}
   );
   gpc1_1 gpc1501 (
      {stage3_34[14]},
      {stage4_34[7]}
   );
   gpc1_1 gpc1502 (
      {stage3_34[15]},
      {stage4_34[8]}
   );
   gpc623_5 gpc1503 (
      {stage4_1[0], stage4_1[1], stage4_1[2]},
      {stage4_2[0], stage4_2[1]},
      {stage4_3[0], stage4_3[1], stage4_3[2], stage4_3[3], stage4_3[4], stage4_3[5]},
      {stage5_5[0],stage5_4[0],stage5_3[0],stage5_2[0],stage5_1[0]}
   );
   gpc1163_5 gpc1504 (
      {stage4_3[6], stage4_3[7], stage4_3[8]},
      {stage4_4[0], stage4_4[1], stage4_4[2], stage4_4[3], stage4_4[4], stage4_4[5]},
      {stage4_5[0]},
      {stage4_6[0]},
      {stage5_7[0],stage5_6[0],stage5_5[1],stage5_4[1],stage5_3[1]}
   );
   gpc1415_5 gpc1505 (
      {stage4_6[1], stage4_6[2], stage4_6[3], stage4_6[4], stage4_6[5]},
      {stage4_7[0]},
      {stage4_8[0], stage4_8[1], stage4_8[2], stage4_8[3]},
      {stage4_9[0]},
      {stage5_10[0],stage5_9[0],stage5_8[0],stage5_7[1],stage5_6[1]}
   );
   gpc223_4 gpc1506 (
      {stage4_7[1], stage4_7[2], stage4_7[3]},
      {stage4_8[4], stage4_8[5]},
      {stage4_9[1], stage4_9[2]},
      {stage5_10[1],stage5_9[1],stage5_8[1],stage5_7[2]}
   );
   gpc2135_5 gpc1507 (
      {stage4_9[3], stage4_9[4], stage4_9[5], stage4_9[6], stage4_9[7]},
      {stage4_10[0], stage4_10[1], stage4_10[2]},
      {stage4_11[0]},
      {stage4_12[0], stage4_12[1]},
      {stage5_13[0],stage5_12[0],stage5_11[0],stage5_10[2],stage5_9[2]}
   );
   gpc615_5 gpc1508 (
      {stage4_10[3], stage4_10[4], stage4_10[5], stage4_10[6], stage4_10[7]},
      {stage4_11[1]},
      {stage4_12[2], stage4_12[3], stage4_12[4], stage4_12[5], stage4_12[6], stage4_12[7]},
      {stage5_14[0],stage5_13[1],stage5_12[1],stage5_11[1],stage5_10[3]}
   );
   gpc615_5 gpc1509 (
      {stage4_11[2], stage4_11[3], stage4_11[4], stage4_11[5], stage4_11[6]},
      {stage4_12[8]},
      {stage4_13[0], stage4_13[1], stage4_13[2], stage4_13[3], stage4_13[4], 1'b0},
      {stage5_15[0],stage5_14[1],stage5_13[2],stage5_12[2],stage5_11[2]}
   );
   gpc1163_5 gpc1510 (
      {stage4_14[0], stage4_14[1], stage4_14[2]},
      {stage4_15[0], stage4_15[1], stage4_15[2], stage4_15[3], stage4_15[4], stage4_15[5]},
      {stage4_16[0]},
      {stage4_17[0]},
      {stage5_18[0],stage5_17[0],stage5_16[0],stage5_15[1],stage5_14[2]}
   );
   gpc606_5 gpc1511 (
      {stage4_16[1], stage4_16[2], stage4_16[3], stage4_16[4], stage4_16[5], stage4_16[6]},
      {stage4_18[0], stage4_18[1], stage4_18[2], stage4_18[3], stage4_18[4], stage4_18[5]},
      {stage5_20[0],stage5_19[0],stage5_18[1],stage5_17[1],stage5_16[1]}
   );
   gpc615_5 gpc1512 (
      {stage4_17[1], stage4_17[2], stage4_17[3], stage4_17[4], stage4_17[5]},
      {stage4_18[6]},
      {stage4_19[0], stage4_19[1], stage4_19[2], stage4_19[3], stage4_19[4], stage4_19[5]},
      {stage5_21[0],stage5_20[1],stage5_19[1],stage5_18[2],stage5_17[2]}
   );
   gpc615_5 gpc1513 (
      {stage4_17[6], stage4_17[7], stage4_17[8], stage4_17[9], stage4_17[10]},
      {stage4_18[7]},
      {stage4_19[6], stage4_19[7], stage4_19[8], stage4_19[9], stage4_19[10], stage4_19[11]},
      {stage5_21[1],stage5_20[2],stage5_19[2],stage5_18[3],stage5_17[3]}
   );
   gpc606_5 gpc1514 (
      {stage4_20[0], stage4_20[1], stage4_20[2], stage4_20[3], stage4_20[4], stage4_20[5]},
      {stage4_22[0], stage4_22[1], stage4_22[2], stage4_22[3], stage4_22[4], stage4_22[5]},
      {stage5_24[0],stage5_23[0],stage5_22[0],stage5_21[2],stage5_20[3]}
   );
   gpc135_4 gpc1515 (
      {stage4_21[0], stage4_21[1], stage4_21[2], stage4_21[3], stage4_21[4]},
      {stage4_22[6], stage4_22[7], stage4_22[8]},
      {stage4_23[0]},
      {stage5_24[1],stage5_23[1],stage5_22[1],stage5_21[3]}
   );
   gpc615_5 gpc1516 (
      {stage4_23[1], stage4_23[2], stage4_23[3], stage4_23[4], stage4_23[5]},
      {stage4_24[0]},
      {stage4_25[0], stage4_25[1], stage4_25[2], stage4_25[3], stage4_25[4], stage4_25[5]},
      {stage5_27[0],stage5_26[0],stage5_25[0],stage5_24[2],stage5_23[2]}
   );
   gpc2135_5 gpc1517 (
      {stage4_24[1], stage4_24[2], stage4_24[3], stage4_24[4], stage4_24[5]},
      {stage4_25[6], stage4_25[7], stage4_25[8]},
      {stage4_26[0]},
      {stage4_27[0], stage4_27[1]},
      {stage5_28[0],stage5_27[1],stage5_26[1],stage5_25[1],stage5_24[3]}
   );
   gpc2223_5 gpc1518 (
      {stage4_26[1], stage4_26[2], stage4_26[3]},
      {stage4_27[2], stage4_27[3]},
      {stage4_28[0], stage4_28[1]},
      {stage4_29[0], stage4_29[1]},
      {stage5_30[0],stage5_29[0],stage5_28[1],stage5_27[2],stage5_26[2]}
   );
   gpc615_5 gpc1519 (
      {stage4_26[4], stage4_26[5], stage4_26[6], stage4_26[7], stage4_26[8]},
      {stage4_27[4]},
      {stage4_28[2], stage4_28[3], stage4_28[4], stage4_28[5], stage4_28[6], stage4_28[7]},
      {stage5_30[1],stage5_29[1],stage5_28[2],stage5_27[3],stage5_26[3]}
   );
   gpc606_5 gpc1520 (
      {stage4_30[0], stage4_30[1], stage4_30[2], stage4_30[3], stage4_30[4], stage4_30[5]},
      {stage4_32[0], stage4_32[1], stage4_32[2], stage4_32[3], stage4_32[4], stage4_32[5]},
      {stage5_34[0],stage5_33[0],stage5_32[0],stage5_31[0],stage5_30[2]}
   );
   gpc606_5 gpc1521 (
      {stage4_31[0], stage4_31[1], stage4_31[2], stage4_31[3], stage4_31[4], stage4_31[5]},
      {stage4_33[0], stage4_33[1], stage4_33[2], stage4_33[3], stage4_33[4], stage4_33[5]},
      {stage5_35[0],stage5_34[1],stage5_33[1],stage5_32[1],stage5_31[1]}
   );
   gpc606_5 gpc1522 (
      {stage4_32[6], stage4_32[7], stage4_32[8], stage4_32[9], stage4_32[10], 1'b0},
      {stage4_34[0], stage4_34[1], stage4_34[2], stage4_34[3], stage4_34[4], stage4_34[5]},
      {stage5_36[0],stage5_35[1],stage5_34[2],stage5_33[2],stage5_32[2]}
   );
   gpc2116_5 gpc1523 (
      {stage4_34[6], stage4_34[7], stage4_34[8], 1'b0, 1'b0, 1'b0},
      {stage4_35[0]},
      {stage4_36[0]},
      {stage4_37[0], stage4_37[1]},
      {stage5_38[0],stage5_37[0],stage5_36[1],stage5_35[2],stage5_34[3]}
   );
   gpc1_1 gpc1524 (
      {stage4_0[0]},
      {stage5_0[0]}
   );
   gpc1_1 gpc1525 (
      {stage4_0[1]},
      {stage5_0[1]}
   );
   gpc1_1 gpc1526 (
      {stage4_1[3]},
      {stage5_1[1]}
   );
   gpc1_1 gpc1527 (
      {stage4_1[4]},
      {stage5_1[2]}
   );
   gpc1_1 gpc1528 (
      {stage4_1[5]},
      {stage5_1[3]}
   );
   gpc1_1 gpc1529 (
      {stage4_2[2]},
      {stage5_2[1]}
   );
   gpc1_1 gpc1530 (
      {stage4_2[3]},
      {stage5_2[2]}
   );
   gpc1_1 gpc1531 (
      {stage4_2[4]},
      {stage5_2[3]}
   );
   gpc1_1 gpc1532 (
      {stage4_2[5]},
      {stage5_2[4]}
   );
   gpc1_1 gpc1533 (
      {stage4_3[9]},
      {stage5_3[2]}
   );
   gpc1_1 gpc1534 (
      {stage4_3[10]},
      {stage5_3[3]}
   );
   gpc1_1 gpc1535 (
      {stage4_5[1]},
      {stage5_5[2]}
   );
   gpc1_1 gpc1536 (
      {stage4_5[2]},
      {stage5_5[3]}
   );
   gpc1_1 gpc1537 (
      {stage4_5[3]},
      {stage5_5[4]}
   );
   gpc1_1 gpc1538 (
      {stage4_7[4]},
      {stage5_7[3]}
   );
   gpc1_1 gpc1539 (
      {stage4_7[5]},
      {stage5_7[4]}
   );
   gpc1_1 gpc1540 (
      {stage4_7[6]},
      {stage5_7[5]}
   );
   gpc1_1 gpc1541 (
      {stage4_7[7]},
      {stage5_7[6]}
   );
   gpc1_1 gpc1542 (
      {stage4_8[6]},
      {stage5_8[2]}
   );
   gpc1_1 gpc1543 (
      {stage4_11[7]},
      {stage5_11[3]}
   );
   gpc1_1 gpc1544 (
      {stage4_11[8]},
      {stage5_11[4]}
   );
   gpc1_1 gpc1545 (
      {stage4_11[9]},
      {stage5_11[5]}
   );
   gpc1_1 gpc1546 (
      {stage4_14[3]},
      {stage5_14[3]}
   );
   gpc1_1 gpc1547 (
      {stage4_14[4]},
      {stage5_14[4]}
   );
   gpc1_1 gpc1548 (
      {stage4_14[5]},
      {stage5_14[5]}
   );
   gpc1_1 gpc1549 (
      {stage4_15[6]},
      {stage5_15[2]}
   );
   gpc1_1 gpc1550 (
      {stage4_15[7]},
      {stage5_15[3]}
   );
   gpc1_1 gpc1551 (
      {stage4_15[8]},
      {stage5_15[4]}
   );
   gpc1_1 gpc1552 (
      {stage4_15[9]},
      {stage5_15[5]}
   );
   gpc1_1 gpc1553 (
      {stage4_17[11]},
      {stage5_17[4]}
   );
   gpc1_1 gpc1554 (
      {stage4_17[12]},
      {stage5_17[5]}
   );
   gpc1_1 gpc1555 (
      {stage4_18[8]},
      {stage5_18[4]}
   );
   gpc1_1 gpc1556 (
      {stage4_21[5]},
      {stage5_21[4]}
   );
   gpc1_1 gpc1557 (
      {stage4_23[6]},
      {stage5_23[3]}
   );
   gpc1_1 gpc1558 (
      {stage4_24[6]},
      {stage5_24[4]}
   );
   gpc1_1 gpc1559 (
      {stage4_24[7]},
      {stage5_24[5]}
   );
   gpc1_1 gpc1560 (
      {stage4_28[8]},
      {stage5_28[3]}
   );
   gpc1_1 gpc1561 (
      {stage4_29[2]},
      {stage5_29[2]}
   );
   gpc1_1 gpc1562 (
      {stage4_29[3]},
      {stage5_29[3]}
   );
   gpc1_1 gpc1563 (
      {stage4_29[4]},
      {stage5_29[4]}
   );
   gpc1_1 gpc1564 (
      {stage4_29[5]},
      {stage5_29[5]}
   );
   gpc1_1 gpc1565 (
      {stage4_33[6]},
      {stage5_33[3]}
   );
   gpc1_1 gpc1566 (
      {stage4_33[7]},
      {stage5_33[4]}
   );
   gpc1_1 gpc1567 (
      {stage4_35[1]},
      {stage5_35[3]}
   );
   gpc1_1 gpc1568 (
      {stage4_35[2]},
      {stage5_35[4]}
   );
   gpc1_1 gpc1569 (
      {stage4_35[3]},
      {stage5_35[5]}
   );
   gpc1_1 gpc1570 (
      {stage4_36[1]},
      {stage5_36[2]}
   );
   gpc1_1 gpc1571 (
      {stage4_36[2]},
      {stage5_36[3]}
   );
   gpc1343_5 gpc1572 (
      {stage5_1[0], stage5_1[1], stage5_1[2]},
      {stage5_2[0], stage5_2[1], stage5_2[2], stage5_2[3]},
      {stage5_3[0], stage5_3[1], stage5_3[2]},
      {stage5_4[0]},
      {stage6_5[0],stage6_4[0],stage6_3[0],stage6_2[0],stage6_1[0]}
   );
   gpc615_5 gpc1573 (
      {stage5_5[0], stage5_5[1], stage5_5[2], stage5_5[3], stage5_5[4]},
      {stage5_6[0]},
      {stage5_7[0], stage5_7[1], stage5_7[2], stage5_7[3], stage5_7[4], stage5_7[5]},
      {stage6_9[0],stage6_8[0],stage6_7[0],stage6_6[0],stage6_5[1]}
   );
   gpc1343_5 gpc1574 (
      {stage5_8[0], stage5_8[1], stage5_8[2]},
      {stage5_9[0], stage5_9[1], stage5_9[2], 1'b0},
      {stage5_10[0], stage5_10[1], stage5_10[2]},
      {stage5_11[0]},
      {stage6_12[0],stage6_11[0],stage6_10[0],stage6_9[1],stage6_8[1]}
   );
   gpc135_4 gpc1575 (
      {stage5_11[1], stage5_11[2], stage5_11[3], stage5_11[4], stage5_11[5]},
      {stage5_12[0], stage5_12[1], stage5_12[2]},
      {stage5_13[0]},
      {stage6_14[0],stage6_13[0],stage6_12[1],stage6_11[1]}
   );
   gpc1163_5 gpc1576 (
      {stage5_13[1], stage5_13[2], 1'b0},
      {stage5_14[0], stage5_14[1], stage5_14[2], stage5_14[3], stage5_14[4], stage5_14[5]},
      {stage5_15[0]},
      {stage5_16[0]},
      {stage6_17[0],stage6_16[0],stage6_15[0],stage6_14[1],stage6_13[1]}
   );
   gpc615_5 gpc1577 (
      {stage5_15[1], stage5_15[2], stage5_15[3], stage5_15[4], stage5_15[5]},
      {stage5_16[1]},
      {stage5_17[0], stage5_17[1], stage5_17[2], stage5_17[3], stage5_17[4], stage5_17[5]},
      {stage6_19[0],stage6_18[0],stage6_17[1],stage6_16[1],stage6_15[1]}
   );
   gpc135_4 gpc1578 (
      {stage5_18[0], stage5_18[1], stage5_18[2], stage5_18[3], stage5_18[4]},
      {stage5_19[0], stage5_19[1], stage5_19[2]},
      {stage5_20[0]},
      {stage6_21[0],stage6_20[0],stage6_19[1],stage6_18[1]}
   );
   gpc1163_5 gpc1579 (
      {stage5_20[1], stage5_20[2], stage5_20[3]},
      {stage5_21[0], stage5_21[1], stage5_21[2], stage5_21[3], stage5_21[4], 1'b0},
      {stage5_22[0]},
      {stage5_23[0]},
      {stage6_24[0],stage6_23[0],stage6_22[0],stage6_21[1],stage6_20[1]}
   );
   gpc1163_5 gpc1580 (
      {stage5_23[1], stage5_23[2], stage5_23[3]},
      {stage5_24[0], stage5_24[1], stage5_24[2], stage5_24[3], stage5_24[4], stage5_24[5]},
      {stage5_25[0]},
      {stage5_26[0]},
      {stage6_27[0],stage6_26[0],stage6_25[0],stage6_24[1],stage6_23[1]}
   );
   gpc1343_5 gpc1581 (
      {stage5_26[1], stage5_26[2], stage5_26[3]},
      {stage5_27[0], stage5_27[1], stage5_27[2], stage5_27[3]},
      {stage5_28[0], stage5_28[1], stage5_28[2]},
      {stage5_29[0]},
      {stage6_30[0],stage6_29[0],stage6_28[0],stage6_27[1],stage6_26[1]}
   );
   gpc2135_5 gpc1582 (
      {stage5_29[1], stage5_29[2], stage5_29[3], stage5_29[4], stage5_29[5]},
      {stage5_30[0], stage5_30[1], stage5_30[2]},
      {stage5_31[0]},
      {stage5_32[0], stage5_32[1]},
      {stage6_33[0],stage6_32[0],stage6_31[0],stage6_30[1],stage6_29[1]}
   );
   gpc606_5 gpc1583 (
      {stage5_33[0], stage5_33[1], stage5_33[2], stage5_33[3], stage5_33[4], 1'b0},
      {stage5_35[0], stage5_35[1], stage5_35[2], stage5_35[3], stage5_35[4], stage5_35[5]},
      {stage6_37[0],stage6_36[0],stage6_35[0],stage6_34[0],stage6_33[1]}
   );
   gpc1415_5 gpc1584 (
      {stage5_34[0], stage5_34[1], stage5_34[2], stage5_34[3], 1'b0},
      {1'b0},
      {stage5_36[0], stage5_36[1], stage5_36[2], stage5_36[3]},
      {stage5_37[0]},
      {stage6_38[0],stage6_37[1],stage6_36[1],stage6_35[1],stage6_34[1]}
   );
   gpc1_1 gpc1585 (
      {stage5_0[0]},
      {stage6_0[0]}
   );
   gpc1_1 gpc1586 (
      {stage5_0[1]},
      {stage6_0[1]}
   );
   gpc1_1 gpc1587 (
      {stage5_1[3]},
      {stage6_1[1]}
   );
   gpc1_1 gpc1588 (
      {stage5_2[4]},
      {stage6_2[1]}
   );
   gpc1_1 gpc1589 (
      {stage5_3[3]},
      {stage6_3[1]}
   );
   gpc1_1 gpc1590 (
      {stage5_4[1]},
      {stage6_4[1]}
   );
   gpc1_1 gpc1591 (
      {stage5_6[1]},
      {stage6_6[1]}
   );
   gpc1_1 gpc1592 (
      {stage5_7[6]},
      {stage6_7[1]}
   );
   gpc1_1 gpc1593 (
      {stage5_10[3]},
      {stage6_10[1]}
   );
   gpc1_1 gpc1594 (
      {stage5_22[1]},
      {stage6_22[1]}
   );
   gpc1_1 gpc1595 (
      {stage5_25[1]},
      {stage6_25[1]}
   );
   gpc1_1 gpc1596 (
      {stage5_28[3]},
      {stage6_28[1]}
   );
   gpc1_1 gpc1597 (
      {stage5_31[1]},
      {stage6_31[1]}
   );
   gpc1_1 gpc1598 (
      {stage5_32[2]},
      {stage6_32[1]}
   );
   gpc1_1 gpc1599 (
      {stage5_38[0]},
      {stage6_38[1]}
   );
endmodule
module rowadder2_1_39(input [38:0] src0, input [38:0] src1, output [39:0] dst0);
    wire [38:0] gene;
    wire [38:0] prop;
    wire [39:0] out;
    wire [39:0] carryout;
    LUT2 #(
        .INIT(4'h8)
    ) lut_0_gene (
        .I0(src0[0]),
        .I1(src1[0]),
        .O(gene[0])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_0_prop (
        .I0(src0[0]),
        .I1(src1[0]),
        .O(prop[0])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_1_gene (
        .I0(src0[1]),
        .I1(src1[1]),
        .O(gene[1])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_1_prop (
        .I0(src0[1]),
        .I1(src1[1]),
        .O(prop[1])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_2_gene (
        .I0(src0[2]),
        .I1(src1[2]),
        .O(gene[2])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_2_prop (
        .I0(src0[2]),
        .I1(src1[2]),
        .O(prop[2])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_3_gene (
        .I0(src0[3]),
        .I1(src1[3]),
        .O(gene[3])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_3_prop (
        .I0(src0[3]),
        .I1(src1[3]),
        .O(prop[3])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_4_gene (
        .I0(src0[4]),
        .I1(src1[4]),
        .O(gene[4])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_4_prop (
        .I0(src0[4]),
        .I1(src1[4]),
        .O(prop[4])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_5_gene (
        .I0(src0[5]),
        .I1(src1[5]),
        .O(gene[5])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_5_prop (
        .I0(src0[5]),
        .I1(src1[5]),
        .O(prop[5])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_6_gene (
        .I0(src0[6]),
        .I1(src1[6]),
        .O(gene[6])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_6_prop (
        .I0(src0[6]),
        .I1(src1[6]),
        .O(prop[6])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_7_gene (
        .I0(src0[7]),
        .I1(src1[7]),
        .O(gene[7])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_7_prop (
        .I0(src0[7]),
        .I1(src1[7]),
        .O(prop[7])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_8_gene (
        .I0(src0[8]),
        .I1(src1[8]),
        .O(gene[8])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_8_prop (
        .I0(src0[8]),
        .I1(src1[8]),
        .O(prop[8])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_9_gene (
        .I0(src0[9]),
        .I1(src1[9]),
        .O(gene[9])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_9_prop (
        .I0(src0[9]),
        .I1(src1[9]),
        .O(prop[9])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_10_gene (
        .I0(src0[10]),
        .I1(src1[10]),
        .O(gene[10])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_10_prop (
        .I0(src0[10]),
        .I1(src1[10]),
        .O(prop[10])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_11_gene (
        .I0(src0[11]),
        .I1(src1[11]),
        .O(gene[11])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_11_prop (
        .I0(src0[11]),
        .I1(src1[11]),
        .O(prop[11])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_12_gene (
        .I0(src0[12]),
        .I1(src1[12]),
        .O(gene[12])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_12_prop (
        .I0(src0[12]),
        .I1(src1[12]),
        .O(prop[12])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_13_gene (
        .I0(src0[13]),
        .I1(src1[13]),
        .O(gene[13])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_13_prop (
        .I0(src0[13]),
        .I1(src1[13]),
        .O(prop[13])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_14_gene (
        .I0(src0[14]),
        .I1(src1[14]),
        .O(gene[14])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_14_prop (
        .I0(src0[14]),
        .I1(src1[14]),
        .O(prop[14])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_15_gene (
        .I0(src0[15]),
        .I1(src1[15]),
        .O(gene[15])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_15_prop (
        .I0(src0[15]),
        .I1(src1[15]),
        .O(prop[15])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_16_gene (
        .I0(src0[16]),
        .I1(src1[16]),
        .O(gene[16])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_16_prop (
        .I0(src0[16]),
        .I1(src1[16]),
        .O(prop[16])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_17_gene (
        .I0(src0[17]),
        .I1(src1[17]),
        .O(gene[17])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_17_prop (
        .I0(src0[17]),
        .I1(src1[17]),
        .O(prop[17])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_18_gene (
        .I0(src0[18]),
        .I1(src1[18]),
        .O(gene[18])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_18_prop (
        .I0(src0[18]),
        .I1(src1[18]),
        .O(prop[18])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_19_gene (
        .I0(src0[19]),
        .I1(src1[19]),
        .O(gene[19])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_19_prop (
        .I0(src0[19]),
        .I1(src1[19]),
        .O(prop[19])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_20_gene (
        .I0(src0[20]),
        .I1(src1[20]),
        .O(gene[20])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_20_prop (
        .I0(src0[20]),
        .I1(src1[20]),
        .O(prop[20])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_21_gene (
        .I0(src0[21]),
        .I1(src1[21]),
        .O(gene[21])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_21_prop (
        .I0(src0[21]),
        .I1(src1[21]),
        .O(prop[21])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_22_gene (
        .I0(src0[22]),
        .I1(src1[22]),
        .O(gene[22])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_22_prop (
        .I0(src0[22]),
        .I1(src1[22]),
        .O(prop[22])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_23_gene (
        .I0(src0[23]),
        .I1(src1[23]),
        .O(gene[23])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_23_prop (
        .I0(src0[23]),
        .I1(src1[23]),
        .O(prop[23])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_24_gene (
        .I0(src0[24]),
        .I1(src1[24]),
        .O(gene[24])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_24_prop (
        .I0(src0[24]),
        .I1(src1[24]),
        .O(prop[24])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_25_gene (
        .I0(src0[25]),
        .I1(src1[25]),
        .O(gene[25])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_25_prop (
        .I0(src0[25]),
        .I1(src1[25]),
        .O(prop[25])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_26_gene (
        .I0(src0[26]),
        .I1(src1[26]),
        .O(gene[26])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_26_prop (
        .I0(src0[26]),
        .I1(src1[26]),
        .O(prop[26])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_27_gene (
        .I0(src0[27]),
        .I1(src1[27]),
        .O(gene[27])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_27_prop (
        .I0(src0[27]),
        .I1(src1[27]),
        .O(prop[27])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_28_gene (
        .I0(src0[28]),
        .I1(src1[28]),
        .O(gene[28])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_28_prop (
        .I0(src0[28]),
        .I1(src1[28]),
        .O(prop[28])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_29_gene (
        .I0(src0[29]),
        .I1(src1[29]),
        .O(gene[29])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_29_prop (
        .I0(src0[29]),
        .I1(src1[29]),
        .O(prop[29])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_30_gene (
        .I0(src0[30]),
        .I1(src1[30]),
        .O(gene[30])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_30_prop (
        .I0(src0[30]),
        .I1(src1[30]),
        .O(prop[30])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_31_gene (
        .I0(src0[31]),
        .I1(src1[31]),
        .O(gene[31])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_31_prop (
        .I0(src0[31]),
        .I1(src1[31]),
        .O(prop[31])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_32_gene (
        .I0(src0[32]),
        .I1(src1[32]),
        .O(gene[32])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_32_prop (
        .I0(src0[32]),
        .I1(src1[32]),
        .O(prop[32])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_33_gene (
        .I0(src0[33]),
        .I1(src1[33]),
        .O(gene[33])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_33_prop (
        .I0(src0[33]),
        .I1(src1[33]),
        .O(prop[33])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_34_gene (
        .I0(src0[34]),
        .I1(src1[34]),
        .O(gene[34])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_34_prop (
        .I0(src0[34]),
        .I1(src1[34]),
        .O(prop[34])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_35_gene (
        .I0(src0[35]),
        .I1(src1[35]),
        .O(gene[35])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_35_prop (
        .I0(src0[35]),
        .I1(src1[35]),
        .O(prop[35])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_36_gene (
        .I0(src0[36]),
        .I1(src1[36]),
        .O(gene[36])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_36_prop (
        .I0(src0[36]),
        .I1(src1[36]),
        .O(prop[36])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_37_gene (
        .I0(src0[37]),
        .I1(src1[37]),
        .O(gene[37])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_37_prop (
        .I0(src0[37]),
        .I1(src1[37]),
        .O(prop[37])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_38_gene (
        .I0(src0[38]),
        .I1(src1[38]),
        .O(gene[38])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_38_prop (
        .I0(src0[38]),
        .I1(src1[38]),
        .O(prop[38])
    );
    CARRY4 carry4_3_0 (
        .CO(carryout[3:0]),
        .O(out[3:0]),
        .CI(1'h0),
        .CYINIT(1'h0),
        .DI(gene[3:0]),
        .S(prop[3:0])
    );
    CARRY4 carry4_7_4 (
        .CO(carryout[7:4]),
        .O(out[7:4]),
        .CI(carryout[3]),
        .CYINIT(1'h0),
        .DI(gene[7:4]),
        .S(prop[7:4])
    );
    CARRY4 carry4_11_8 (
        .CO(carryout[11:8]),
        .O(out[11:8]),
        .CI(carryout[7]),
        .CYINIT(1'h0),
        .DI(gene[11:8]),
        .S(prop[11:8])
    );
    CARRY4 carry4_15_12 (
        .CO(carryout[15:12]),
        .O(out[15:12]),
        .CI(carryout[11]),
        .CYINIT(1'h0),
        .DI(gene[15:12]),
        .S(prop[15:12])
    );
    CARRY4 carry4_19_16 (
        .CO(carryout[19:16]),
        .O(out[19:16]),
        .CI(carryout[15]),
        .CYINIT(1'h0),
        .DI(gene[19:16]),
        .S(prop[19:16])
    );
    CARRY4 carry4_23_20 (
        .CO(carryout[23:20]),
        .O(out[23:20]),
        .CI(carryout[19]),
        .CYINIT(1'h0),
        .DI(gene[23:20]),
        .S(prop[23:20])
    );
    CARRY4 carry4_27_24 (
        .CO(carryout[27:24]),
        .O(out[27:24]),
        .CI(carryout[23]),
        .CYINIT(1'h0),
        .DI(gene[27:24]),
        .S(prop[27:24])
    );
    CARRY4 carry4_31_28 (
        .CO(carryout[31:28]),
        .O(out[31:28]),
        .CI(carryout[27]),
        .CYINIT(1'h0),
        .DI(gene[31:28]),
        .S(prop[31:28])
    );
    CARRY4 carry4_35_32 (
        .CO(carryout[35:32]),
        .O(out[35:32]),
        .CI(carryout[31]),
        .CYINIT(1'h0),
        .DI(gene[35:32]),
        .S(prop[35:32])
    );
    CARRY4 carry4_39_36 (
        .CO(carryout[39:36]),
        .O(out[39:36]),
        .CI(carryout[35]),
        .CYINIT(1'h0),
        .DI({1'h0, gene[38:36]}),
        .S({1'h0, prop[38:36]})
    );
    assign dst0 = {carryout[38], out[38:0]};
endmodule


module testbench();
    reg [161:0] src0;
    reg [161:0] src1;
    reg [161:0] src2;
    reg [161:0] src3;
    reg [161:0] src4;
    reg [161:0] src5;
    reg [161:0] src6;
    reg [161:0] src7;
    reg [161:0] src8;
    reg [161:0] src9;
    reg [161:0] src10;
    reg [161:0] src11;
    reg [161:0] src12;
    reg [161:0] src13;
    reg [161:0] src14;
    reg [161:0] src15;
    reg [161:0] src16;
    reg [161:0] src17;
    reg [161:0] src18;
    reg [161:0] src19;
    reg [161:0] src20;
    reg [161:0] src21;
    reg [161:0] src22;
    reg [161:0] src23;
    reg [161:0] src24;
    reg [161:0] src25;
    reg [161:0] src26;
    reg [161:0] src27;
    reg [161:0] src28;
    reg [161:0] src29;
    reg [161:0] src30;
    reg [161:0] src31;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [0:0] dst26;
    wire [0:0] dst27;
    wire [0:0] dst28;
    wire [0:0] dst29;
    wire [0:0] dst30;
    wire [0:0] dst31;
    wire [0:0] dst32;
    wire [0:0] dst33;
    wire [0:0] dst34;
    wire [0:0] dst35;
    wire [0:0] dst36;
    wire [0:0] dst37;
    wire [0:0] dst38;
    wire [0:0] dst39;
    wire [39:0] srcsum;
    wire [39:0] dstsum;
    wire test;
    compressor2_1_162_32 compressor2_1_162_32(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .src31(src31),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25),
        .dst26(dst26),
        .dst27(dst27),
        .dst28(dst28),
        .dst29(dst29),
        .dst30(dst30),
        .dst31(dst31),
        .dst32(dst32),
        .dst33(dst33),
        .dst34(dst34),
        .dst35(dst35),
        .dst36(dst36),
        .dst37(dst37),
        .dst38(dst38),
        .dst39(dst39));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13] + src0[14] + src0[15] + src0[16] + src0[17] + src0[18] + src0[19] + src0[20] + src0[21] + src0[22] + src0[23] + src0[24] + src0[25] + src0[26] + src0[27] + src0[28] + src0[29] + src0[30] + src0[31] + src0[32] + src0[33] + src0[34] + src0[35] + src0[36] + src0[37] + src0[38] + src0[39] + src0[40] + src0[41] + src0[42] + src0[43] + src0[44] + src0[45] + src0[46] + src0[47] + src0[48] + src0[49] + src0[50] + src0[51] + src0[52] + src0[53] + src0[54] + src0[55] + src0[56] + src0[57] + src0[58] + src0[59] + src0[60] + src0[61] + src0[62] + src0[63] + src0[64] + src0[65] + src0[66] + src0[67] + src0[68] + src0[69] + src0[70] + src0[71] + src0[72] + src0[73] + src0[74] + src0[75] + src0[76] + src0[77] + src0[78] + src0[79] + src0[80] + src0[81] + src0[82] + src0[83] + src0[84] + src0[85] + src0[86] + src0[87] + src0[88] + src0[89] + src0[90] + src0[91] + src0[92] + src0[93] + src0[94] + src0[95] + src0[96] + src0[97] + src0[98] + src0[99] + src0[100] + src0[101] + src0[102] + src0[103] + src0[104] + src0[105] + src0[106] + src0[107] + src0[108] + src0[109] + src0[110] + src0[111] + src0[112] + src0[113] + src0[114] + src0[115] + src0[116] + src0[117] + src0[118] + src0[119] + src0[120] + src0[121] + src0[122] + src0[123] + src0[124] + src0[125] + src0[126] + src0[127] + src0[128] + src0[129] + src0[130] + src0[131] + src0[132] + src0[133] + src0[134] + src0[135] + src0[136] + src0[137] + src0[138] + src0[139] + src0[140] + src0[141] + src0[142] + src0[143] + src0[144] + src0[145] + src0[146] + src0[147] + src0[148] + src0[149] + src0[150] + src0[151] + src0[152] + src0[153] + src0[154] + src0[155] + src0[156] + src0[157] + src0[158] + src0[159] + src0[160] + src0[161])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13] + src1[14] + src1[15] + src1[16] + src1[17] + src1[18] + src1[19] + src1[20] + src1[21] + src1[22] + src1[23] + src1[24] + src1[25] + src1[26] + src1[27] + src1[28] + src1[29] + src1[30] + src1[31] + src1[32] + src1[33] + src1[34] + src1[35] + src1[36] + src1[37] + src1[38] + src1[39] + src1[40] + src1[41] + src1[42] + src1[43] + src1[44] + src1[45] + src1[46] + src1[47] + src1[48] + src1[49] + src1[50] + src1[51] + src1[52] + src1[53] + src1[54] + src1[55] + src1[56] + src1[57] + src1[58] + src1[59] + src1[60] + src1[61] + src1[62] + src1[63] + src1[64] + src1[65] + src1[66] + src1[67] + src1[68] + src1[69] + src1[70] + src1[71] + src1[72] + src1[73] + src1[74] + src1[75] + src1[76] + src1[77] + src1[78] + src1[79] + src1[80] + src1[81] + src1[82] + src1[83] + src1[84] + src1[85] + src1[86] + src1[87] + src1[88] + src1[89] + src1[90] + src1[91] + src1[92] + src1[93] + src1[94] + src1[95] + src1[96] + src1[97] + src1[98] + src1[99] + src1[100] + src1[101] + src1[102] + src1[103] + src1[104] + src1[105] + src1[106] + src1[107] + src1[108] + src1[109] + src1[110] + src1[111] + src1[112] + src1[113] + src1[114] + src1[115] + src1[116] + src1[117] + src1[118] + src1[119] + src1[120] + src1[121] + src1[122] + src1[123] + src1[124] + src1[125] + src1[126] + src1[127] + src1[128] + src1[129] + src1[130] + src1[131] + src1[132] + src1[133] + src1[134] + src1[135] + src1[136] + src1[137] + src1[138] + src1[139] + src1[140] + src1[141] + src1[142] + src1[143] + src1[144] + src1[145] + src1[146] + src1[147] + src1[148] + src1[149] + src1[150] + src1[151] + src1[152] + src1[153] + src1[154] + src1[155] + src1[156] + src1[157] + src1[158] + src1[159] + src1[160] + src1[161])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13] + src2[14] + src2[15] + src2[16] + src2[17] + src2[18] + src2[19] + src2[20] + src2[21] + src2[22] + src2[23] + src2[24] + src2[25] + src2[26] + src2[27] + src2[28] + src2[29] + src2[30] + src2[31] + src2[32] + src2[33] + src2[34] + src2[35] + src2[36] + src2[37] + src2[38] + src2[39] + src2[40] + src2[41] + src2[42] + src2[43] + src2[44] + src2[45] + src2[46] + src2[47] + src2[48] + src2[49] + src2[50] + src2[51] + src2[52] + src2[53] + src2[54] + src2[55] + src2[56] + src2[57] + src2[58] + src2[59] + src2[60] + src2[61] + src2[62] + src2[63] + src2[64] + src2[65] + src2[66] + src2[67] + src2[68] + src2[69] + src2[70] + src2[71] + src2[72] + src2[73] + src2[74] + src2[75] + src2[76] + src2[77] + src2[78] + src2[79] + src2[80] + src2[81] + src2[82] + src2[83] + src2[84] + src2[85] + src2[86] + src2[87] + src2[88] + src2[89] + src2[90] + src2[91] + src2[92] + src2[93] + src2[94] + src2[95] + src2[96] + src2[97] + src2[98] + src2[99] + src2[100] + src2[101] + src2[102] + src2[103] + src2[104] + src2[105] + src2[106] + src2[107] + src2[108] + src2[109] + src2[110] + src2[111] + src2[112] + src2[113] + src2[114] + src2[115] + src2[116] + src2[117] + src2[118] + src2[119] + src2[120] + src2[121] + src2[122] + src2[123] + src2[124] + src2[125] + src2[126] + src2[127] + src2[128] + src2[129] + src2[130] + src2[131] + src2[132] + src2[133] + src2[134] + src2[135] + src2[136] + src2[137] + src2[138] + src2[139] + src2[140] + src2[141] + src2[142] + src2[143] + src2[144] + src2[145] + src2[146] + src2[147] + src2[148] + src2[149] + src2[150] + src2[151] + src2[152] + src2[153] + src2[154] + src2[155] + src2[156] + src2[157] + src2[158] + src2[159] + src2[160] + src2[161])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13] + src3[14] + src3[15] + src3[16] + src3[17] + src3[18] + src3[19] + src3[20] + src3[21] + src3[22] + src3[23] + src3[24] + src3[25] + src3[26] + src3[27] + src3[28] + src3[29] + src3[30] + src3[31] + src3[32] + src3[33] + src3[34] + src3[35] + src3[36] + src3[37] + src3[38] + src3[39] + src3[40] + src3[41] + src3[42] + src3[43] + src3[44] + src3[45] + src3[46] + src3[47] + src3[48] + src3[49] + src3[50] + src3[51] + src3[52] + src3[53] + src3[54] + src3[55] + src3[56] + src3[57] + src3[58] + src3[59] + src3[60] + src3[61] + src3[62] + src3[63] + src3[64] + src3[65] + src3[66] + src3[67] + src3[68] + src3[69] + src3[70] + src3[71] + src3[72] + src3[73] + src3[74] + src3[75] + src3[76] + src3[77] + src3[78] + src3[79] + src3[80] + src3[81] + src3[82] + src3[83] + src3[84] + src3[85] + src3[86] + src3[87] + src3[88] + src3[89] + src3[90] + src3[91] + src3[92] + src3[93] + src3[94] + src3[95] + src3[96] + src3[97] + src3[98] + src3[99] + src3[100] + src3[101] + src3[102] + src3[103] + src3[104] + src3[105] + src3[106] + src3[107] + src3[108] + src3[109] + src3[110] + src3[111] + src3[112] + src3[113] + src3[114] + src3[115] + src3[116] + src3[117] + src3[118] + src3[119] + src3[120] + src3[121] + src3[122] + src3[123] + src3[124] + src3[125] + src3[126] + src3[127] + src3[128] + src3[129] + src3[130] + src3[131] + src3[132] + src3[133] + src3[134] + src3[135] + src3[136] + src3[137] + src3[138] + src3[139] + src3[140] + src3[141] + src3[142] + src3[143] + src3[144] + src3[145] + src3[146] + src3[147] + src3[148] + src3[149] + src3[150] + src3[151] + src3[152] + src3[153] + src3[154] + src3[155] + src3[156] + src3[157] + src3[158] + src3[159] + src3[160] + src3[161])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13] + src4[14] + src4[15] + src4[16] + src4[17] + src4[18] + src4[19] + src4[20] + src4[21] + src4[22] + src4[23] + src4[24] + src4[25] + src4[26] + src4[27] + src4[28] + src4[29] + src4[30] + src4[31] + src4[32] + src4[33] + src4[34] + src4[35] + src4[36] + src4[37] + src4[38] + src4[39] + src4[40] + src4[41] + src4[42] + src4[43] + src4[44] + src4[45] + src4[46] + src4[47] + src4[48] + src4[49] + src4[50] + src4[51] + src4[52] + src4[53] + src4[54] + src4[55] + src4[56] + src4[57] + src4[58] + src4[59] + src4[60] + src4[61] + src4[62] + src4[63] + src4[64] + src4[65] + src4[66] + src4[67] + src4[68] + src4[69] + src4[70] + src4[71] + src4[72] + src4[73] + src4[74] + src4[75] + src4[76] + src4[77] + src4[78] + src4[79] + src4[80] + src4[81] + src4[82] + src4[83] + src4[84] + src4[85] + src4[86] + src4[87] + src4[88] + src4[89] + src4[90] + src4[91] + src4[92] + src4[93] + src4[94] + src4[95] + src4[96] + src4[97] + src4[98] + src4[99] + src4[100] + src4[101] + src4[102] + src4[103] + src4[104] + src4[105] + src4[106] + src4[107] + src4[108] + src4[109] + src4[110] + src4[111] + src4[112] + src4[113] + src4[114] + src4[115] + src4[116] + src4[117] + src4[118] + src4[119] + src4[120] + src4[121] + src4[122] + src4[123] + src4[124] + src4[125] + src4[126] + src4[127] + src4[128] + src4[129] + src4[130] + src4[131] + src4[132] + src4[133] + src4[134] + src4[135] + src4[136] + src4[137] + src4[138] + src4[139] + src4[140] + src4[141] + src4[142] + src4[143] + src4[144] + src4[145] + src4[146] + src4[147] + src4[148] + src4[149] + src4[150] + src4[151] + src4[152] + src4[153] + src4[154] + src4[155] + src4[156] + src4[157] + src4[158] + src4[159] + src4[160] + src4[161])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13] + src5[14] + src5[15] + src5[16] + src5[17] + src5[18] + src5[19] + src5[20] + src5[21] + src5[22] + src5[23] + src5[24] + src5[25] + src5[26] + src5[27] + src5[28] + src5[29] + src5[30] + src5[31] + src5[32] + src5[33] + src5[34] + src5[35] + src5[36] + src5[37] + src5[38] + src5[39] + src5[40] + src5[41] + src5[42] + src5[43] + src5[44] + src5[45] + src5[46] + src5[47] + src5[48] + src5[49] + src5[50] + src5[51] + src5[52] + src5[53] + src5[54] + src5[55] + src5[56] + src5[57] + src5[58] + src5[59] + src5[60] + src5[61] + src5[62] + src5[63] + src5[64] + src5[65] + src5[66] + src5[67] + src5[68] + src5[69] + src5[70] + src5[71] + src5[72] + src5[73] + src5[74] + src5[75] + src5[76] + src5[77] + src5[78] + src5[79] + src5[80] + src5[81] + src5[82] + src5[83] + src5[84] + src5[85] + src5[86] + src5[87] + src5[88] + src5[89] + src5[90] + src5[91] + src5[92] + src5[93] + src5[94] + src5[95] + src5[96] + src5[97] + src5[98] + src5[99] + src5[100] + src5[101] + src5[102] + src5[103] + src5[104] + src5[105] + src5[106] + src5[107] + src5[108] + src5[109] + src5[110] + src5[111] + src5[112] + src5[113] + src5[114] + src5[115] + src5[116] + src5[117] + src5[118] + src5[119] + src5[120] + src5[121] + src5[122] + src5[123] + src5[124] + src5[125] + src5[126] + src5[127] + src5[128] + src5[129] + src5[130] + src5[131] + src5[132] + src5[133] + src5[134] + src5[135] + src5[136] + src5[137] + src5[138] + src5[139] + src5[140] + src5[141] + src5[142] + src5[143] + src5[144] + src5[145] + src5[146] + src5[147] + src5[148] + src5[149] + src5[150] + src5[151] + src5[152] + src5[153] + src5[154] + src5[155] + src5[156] + src5[157] + src5[158] + src5[159] + src5[160] + src5[161])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13] + src6[14] + src6[15] + src6[16] + src6[17] + src6[18] + src6[19] + src6[20] + src6[21] + src6[22] + src6[23] + src6[24] + src6[25] + src6[26] + src6[27] + src6[28] + src6[29] + src6[30] + src6[31] + src6[32] + src6[33] + src6[34] + src6[35] + src6[36] + src6[37] + src6[38] + src6[39] + src6[40] + src6[41] + src6[42] + src6[43] + src6[44] + src6[45] + src6[46] + src6[47] + src6[48] + src6[49] + src6[50] + src6[51] + src6[52] + src6[53] + src6[54] + src6[55] + src6[56] + src6[57] + src6[58] + src6[59] + src6[60] + src6[61] + src6[62] + src6[63] + src6[64] + src6[65] + src6[66] + src6[67] + src6[68] + src6[69] + src6[70] + src6[71] + src6[72] + src6[73] + src6[74] + src6[75] + src6[76] + src6[77] + src6[78] + src6[79] + src6[80] + src6[81] + src6[82] + src6[83] + src6[84] + src6[85] + src6[86] + src6[87] + src6[88] + src6[89] + src6[90] + src6[91] + src6[92] + src6[93] + src6[94] + src6[95] + src6[96] + src6[97] + src6[98] + src6[99] + src6[100] + src6[101] + src6[102] + src6[103] + src6[104] + src6[105] + src6[106] + src6[107] + src6[108] + src6[109] + src6[110] + src6[111] + src6[112] + src6[113] + src6[114] + src6[115] + src6[116] + src6[117] + src6[118] + src6[119] + src6[120] + src6[121] + src6[122] + src6[123] + src6[124] + src6[125] + src6[126] + src6[127] + src6[128] + src6[129] + src6[130] + src6[131] + src6[132] + src6[133] + src6[134] + src6[135] + src6[136] + src6[137] + src6[138] + src6[139] + src6[140] + src6[141] + src6[142] + src6[143] + src6[144] + src6[145] + src6[146] + src6[147] + src6[148] + src6[149] + src6[150] + src6[151] + src6[152] + src6[153] + src6[154] + src6[155] + src6[156] + src6[157] + src6[158] + src6[159] + src6[160] + src6[161])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13] + src7[14] + src7[15] + src7[16] + src7[17] + src7[18] + src7[19] + src7[20] + src7[21] + src7[22] + src7[23] + src7[24] + src7[25] + src7[26] + src7[27] + src7[28] + src7[29] + src7[30] + src7[31] + src7[32] + src7[33] + src7[34] + src7[35] + src7[36] + src7[37] + src7[38] + src7[39] + src7[40] + src7[41] + src7[42] + src7[43] + src7[44] + src7[45] + src7[46] + src7[47] + src7[48] + src7[49] + src7[50] + src7[51] + src7[52] + src7[53] + src7[54] + src7[55] + src7[56] + src7[57] + src7[58] + src7[59] + src7[60] + src7[61] + src7[62] + src7[63] + src7[64] + src7[65] + src7[66] + src7[67] + src7[68] + src7[69] + src7[70] + src7[71] + src7[72] + src7[73] + src7[74] + src7[75] + src7[76] + src7[77] + src7[78] + src7[79] + src7[80] + src7[81] + src7[82] + src7[83] + src7[84] + src7[85] + src7[86] + src7[87] + src7[88] + src7[89] + src7[90] + src7[91] + src7[92] + src7[93] + src7[94] + src7[95] + src7[96] + src7[97] + src7[98] + src7[99] + src7[100] + src7[101] + src7[102] + src7[103] + src7[104] + src7[105] + src7[106] + src7[107] + src7[108] + src7[109] + src7[110] + src7[111] + src7[112] + src7[113] + src7[114] + src7[115] + src7[116] + src7[117] + src7[118] + src7[119] + src7[120] + src7[121] + src7[122] + src7[123] + src7[124] + src7[125] + src7[126] + src7[127] + src7[128] + src7[129] + src7[130] + src7[131] + src7[132] + src7[133] + src7[134] + src7[135] + src7[136] + src7[137] + src7[138] + src7[139] + src7[140] + src7[141] + src7[142] + src7[143] + src7[144] + src7[145] + src7[146] + src7[147] + src7[148] + src7[149] + src7[150] + src7[151] + src7[152] + src7[153] + src7[154] + src7[155] + src7[156] + src7[157] + src7[158] + src7[159] + src7[160] + src7[161])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13] + src8[14] + src8[15] + src8[16] + src8[17] + src8[18] + src8[19] + src8[20] + src8[21] + src8[22] + src8[23] + src8[24] + src8[25] + src8[26] + src8[27] + src8[28] + src8[29] + src8[30] + src8[31] + src8[32] + src8[33] + src8[34] + src8[35] + src8[36] + src8[37] + src8[38] + src8[39] + src8[40] + src8[41] + src8[42] + src8[43] + src8[44] + src8[45] + src8[46] + src8[47] + src8[48] + src8[49] + src8[50] + src8[51] + src8[52] + src8[53] + src8[54] + src8[55] + src8[56] + src8[57] + src8[58] + src8[59] + src8[60] + src8[61] + src8[62] + src8[63] + src8[64] + src8[65] + src8[66] + src8[67] + src8[68] + src8[69] + src8[70] + src8[71] + src8[72] + src8[73] + src8[74] + src8[75] + src8[76] + src8[77] + src8[78] + src8[79] + src8[80] + src8[81] + src8[82] + src8[83] + src8[84] + src8[85] + src8[86] + src8[87] + src8[88] + src8[89] + src8[90] + src8[91] + src8[92] + src8[93] + src8[94] + src8[95] + src8[96] + src8[97] + src8[98] + src8[99] + src8[100] + src8[101] + src8[102] + src8[103] + src8[104] + src8[105] + src8[106] + src8[107] + src8[108] + src8[109] + src8[110] + src8[111] + src8[112] + src8[113] + src8[114] + src8[115] + src8[116] + src8[117] + src8[118] + src8[119] + src8[120] + src8[121] + src8[122] + src8[123] + src8[124] + src8[125] + src8[126] + src8[127] + src8[128] + src8[129] + src8[130] + src8[131] + src8[132] + src8[133] + src8[134] + src8[135] + src8[136] + src8[137] + src8[138] + src8[139] + src8[140] + src8[141] + src8[142] + src8[143] + src8[144] + src8[145] + src8[146] + src8[147] + src8[148] + src8[149] + src8[150] + src8[151] + src8[152] + src8[153] + src8[154] + src8[155] + src8[156] + src8[157] + src8[158] + src8[159] + src8[160] + src8[161])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13] + src9[14] + src9[15] + src9[16] + src9[17] + src9[18] + src9[19] + src9[20] + src9[21] + src9[22] + src9[23] + src9[24] + src9[25] + src9[26] + src9[27] + src9[28] + src9[29] + src9[30] + src9[31] + src9[32] + src9[33] + src9[34] + src9[35] + src9[36] + src9[37] + src9[38] + src9[39] + src9[40] + src9[41] + src9[42] + src9[43] + src9[44] + src9[45] + src9[46] + src9[47] + src9[48] + src9[49] + src9[50] + src9[51] + src9[52] + src9[53] + src9[54] + src9[55] + src9[56] + src9[57] + src9[58] + src9[59] + src9[60] + src9[61] + src9[62] + src9[63] + src9[64] + src9[65] + src9[66] + src9[67] + src9[68] + src9[69] + src9[70] + src9[71] + src9[72] + src9[73] + src9[74] + src9[75] + src9[76] + src9[77] + src9[78] + src9[79] + src9[80] + src9[81] + src9[82] + src9[83] + src9[84] + src9[85] + src9[86] + src9[87] + src9[88] + src9[89] + src9[90] + src9[91] + src9[92] + src9[93] + src9[94] + src9[95] + src9[96] + src9[97] + src9[98] + src9[99] + src9[100] + src9[101] + src9[102] + src9[103] + src9[104] + src9[105] + src9[106] + src9[107] + src9[108] + src9[109] + src9[110] + src9[111] + src9[112] + src9[113] + src9[114] + src9[115] + src9[116] + src9[117] + src9[118] + src9[119] + src9[120] + src9[121] + src9[122] + src9[123] + src9[124] + src9[125] + src9[126] + src9[127] + src9[128] + src9[129] + src9[130] + src9[131] + src9[132] + src9[133] + src9[134] + src9[135] + src9[136] + src9[137] + src9[138] + src9[139] + src9[140] + src9[141] + src9[142] + src9[143] + src9[144] + src9[145] + src9[146] + src9[147] + src9[148] + src9[149] + src9[150] + src9[151] + src9[152] + src9[153] + src9[154] + src9[155] + src9[156] + src9[157] + src9[158] + src9[159] + src9[160] + src9[161])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13] + src10[14] + src10[15] + src10[16] + src10[17] + src10[18] + src10[19] + src10[20] + src10[21] + src10[22] + src10[23] + src10[24] + src10[25] + src10[26] + src10[27] + src10[28] + src10[29] + src10[30] + src10[31] + src10[32] + src10[33] + src10[34] + src10[35] + src10[36] + src10[37] + src10[38] + src10[39] + src10[40] + src10[41] + src10[42] + src10[43] + src10[44] + src10[45] + src10[46] + src10[47] + src10[48] + src10[49] + src10[50] + src10[51] + src10[52] + src10[53] + src10[54] + src10[55] + src10[56] + src10[57] + src10[58] + src10[59] + src10[60] + src10[61] + src10[62] + src10[63] + src10[64] + src10[65] + src10[66] + src10[67] + src10[68] + src10[69] + src10[70] + src10[71] + src10[72] + src10[73] + src10[74] + src10[75] + src10[76] + src10[77] + src10[78] + src10[79] + src10[80] + src10[81] + src10[82] + src10[83] + src10[84] + src10[85] + src10[86] + src10[87] + src10[88] + src10[89] + src10[90] + src10[91] + src10[92] + src10[93] + src10[94] + src10[95] + src10[96] + src10[97] + src10[98] + src10[99] + src10[100] + src10[101] + src10[102] + src10[103] + src10[104] + src10[105] + src10[106] + src10[107] + src10[108] + src10[109] + src10[110] + src10[111] + src10[112] + src10[113] + src10[114] + src10[115] + src10[116] + src10[117] + src10[118] + src10[119] + src10[120] + src10[121] + src10[122] + src10[123] + src10[124] + src10[125] + src10[126] + src10[127] + src10[128] + src10[129] + src10[130] + src10[131] + src10[132] + src10[133] + src10[134] + src10[135] + src10[136] + src10[137] + src10[138] + src10[139] + src10[140] + src10[141] + src10[142] + src10[143] + src10[144] + src10[145] + src10[146] + src10[147] + src10[148] + src10[149] + src10[150] + src10[151] + src10[152] + src10[153] + src10[154] + src10[155] + src10[156] + src10[157] + src10[158] + src10[159] + src10[160] + src10[161])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13] + src11[14] + src11[15] + src11[16] + src11[17] + src11[18] + src11[19] + src11[20] + src11[21] + src11[22] + src11[23] + src11[24] + src11[25] + src11[26] + src11[27] + src11[28] + src11[29] + src11[30] + src11[31] + src11[32] + src11[33] + src11[34] + src11[35] + src11[36] + src11[37] + src11[38] + src11[39] + src11[40] + src11[41] + src11[42] + src11[43] + src11[44] + src11[45] + src11[46] + src11[47] + src11[48] + src11[49] + src11[50] + src11[51] + src11[52] + src11[53] + src11[54] + src11[55] + src11[56] + src11[57] + src11[58] + src11[59] + src11[60] + src11[61] + src11[62] + src11[63] + src11[64] + src11[65] + src11[66] + src11[67] + src11[68] + src11[69] + src11[70] + src11[71] + src11[72] + src11[73] + src11[74] + src11[75] + src11[76] + src11[77] + src11[78] + src11[79] + src11[80] + src11[81] + src11[82] + src11[83] + src11[84] + src11[85] + src11[86] + src11[87] + src11[88] + src11[89] + src11[90] + src11[91] + src11[92] + src11[93] + src11[94] + src11[95] + src11[96] + src11[97] + src11[98] + src11[99] + src11[100] + src11[101] + src11[102] + src11[103] + src11[104] + src11[105] + src11[106] + src11[107] + src11[108] + src11[109] + src11[110] + src11[111] + src11[112] + src11[113] + src11[114] + src11[115] + src11[116] + src11[117] + src11[118] + src11[119] + src11[120] + src11[121] + src11[122] + src11[123] + src11[124] + src11[125] + src11[126] + src11[127] + src11[128] + src11[129] + src11[130] + src11[131] + src11[132] + src11[133] + src11[134] + src11[135] + src11[136] + src11[137] + src11[138] + src11[139] + src11[140] + src11[141] + src11[142] + src11[143] + src11[144] + src11[145] + src11[146] + src11[147] + src11[148] + src11[149] + src11[150] + src11[151] + src11[152] + src11[153] + src11[154] + src11[155] + src11[156] + src11[157] + src11[158] + src11[159] + src11[160] + src11[161])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12] + src12[13] + src12[14] + src12[15] + src12[16] + src12[17] + src12[18] + src12[19] + src12[20] + src12[21] + src12[22] + src12[23] + src12[24] + src12[25] + src12[26] + src12[27] + src12[28] + src12[29] + src12[30] + src12[31] + src12[32] + src12[33] + src12[34] + src12[35] + src12[36] + src12[37] + src12[38] + src12[39] + src12[40] + src12[41] + src12[42] + src12[43] + src12[44] + src12[45] + src12[46] + src12[47] + src12[48] + src12[49] + src12[50] + src12[51] + src12[52] + src12[53] + src12[54] + src12[55] + src12[56] + src12[57] + src12[58] + src12[59] + src12[60] + src12[61] + src12[62] + src12[63] + src12[64] + src12[65] + src12[66] + src12[67] + src12[68] + src12[69] + src12[70] + src12[71] + src12[72] + src12[73] + src12[74] + src12[75] + src12[76] + src12[77] + src12[78] + src12[79] + src12[80] + src12[81] + src12[82] + src12[83] + src12[84] + src12[85] + src12[86] + src12[87] + src12[88] + src12[89] + src12[90] + src12[91] + src12[92] + src12[93] + src12[94] + src12[95] + src12[96] + src12[97] + src12[98] + src12[99] + src12[100] + src12[101] + src12[102] + src12[103] + src12[104] + src12[105] + src12[106] + src12[107] + src12[108] + src12[109] + src12[110] + src12[111] + src12[112] + src12[113] + src12[114] + src12[115] + src12[116] + src12[117] + src12[118] + src12[119] + src12[120] + src12[121] + src12[122] + src12[123] + src12[124] + src12[125] + src12[126] + src12[127] + src12[128] + src12[129] + src12[130] + src12[131] + src12[132] + src12[133] + src12[134] + src12[135] + src12[136] + src12[137] + src12[138] + src12[139] + src12[140] + src12[141] + src12[142] + src12[143] + src12[144] + src12[145] + src12[146] + src12[147] + src12[148] + src12[149] + src12[150] + src12[151] + src12[152] + src12[153] + src12[154] + src12[155] + src12[156] + src12[157] + src12[158] + src12[159] + src12[160] + src12[161])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13] + src13[14] + src13[15] + src13[16] + src13[17] + src13[18] + src13[19] + src13[20] + src13[21] + src13[22] + src13[23] + src13[24] + src13[25] + src13[26] + src13[27] + src13[28] + src13[29] + src13[30] + src13[31] + src13[32] + src13[33] + src13[34] + src13[35] + src13[36] + src13[37] + src13[38] + src13[39] + src13[40] + src13[41] + src13[42] + src13[43] + src13[44] + src13[45] + src13[46] + src13[47] + src13[48] + src13[49] + src13[50] + src13[51] + src13[52] + src13[53] + src13[54] + src13[55] + src13[56] + src13[57] + src13[58] + src13[59] + src13[60] + src13[61] + src13[62] + src13[63] + src13[64] + src13[65] + src13[66] + src13[67] + src13[68] + src13[69] + src13[70] + src13[71] + src13[72] + src13[73] + src13[74] + src13[75] + src13[76] + src13[77] + src13[78] + src13[79] + src13[80] + src13[81] + src13[82] + src13[83] + src13[84] + src13[85] + src13[86] + src13[87] + src13[88] + src13[89] + src13[90] + src13[91] + src13[92] + src13[93] + src13[94] + src13[95] + src13[96] + src13[97] + src13[98] + src13[99] + src13[100] + src13[101] + src13[102] + src13[103] + src13[104] + src13[105] + src13[106] + src13[107] + src13[108] + src13[109] + src13[110] + src13[111] + src13[112] + src13[113] + src13[114] + src13[115] + src13[116] + src13[117] + src13[118] + src13[119] + src13[120] + src13[121] + src13[122] + src13[123] + src13[124] + src13[125] + src13[126] + src13[127] + src13[128] + src13[129] + src13[130] + src13[131] + src13[132] + src13[133] + src13[134] + src13[135] + src13[136] + src13[137] + src13[138] + src13[139] + src13[140] + src13[141] + src13[142] + src13[143] + src13[144] + src13[145] + src13[146] + src13[147] + src13[148] + src13[149] + src13[150] + src13[151] + src13[152] + src13[153] + src13[154] + src13[155] + src13[156] + src13[157] + src13[158] + src13[159] + src13[160] + src13[161])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14] + src14[15] + src14[16] + src14[17] + src14[18] + src14[19] + src14[20] + src14[21] + src14[22] + src14[23] + src14[24] + src14[25] + src14[26] + src14[27] + src14[28] + src14[29] + src14[30] + src14[31] + src14[32] + src14[33] + src14[34] + src14[35] + src14[36] + src14[37] + src14[38] + src14[39] + src14[40] + src14[41] + src14[42] + src14[43] + src14[44] + src14[45] + src14[46] + src14[47] + src14[48] + src14[49] + src14[50] + src14[51] + src14[52] + src14[53] + src14[54] + src14[55] + src14[56] + src14[57] + src14[58] + src14[59] + src14[60] + src14[61] + src14[62] + src14[63] + src14[64] + src14[65] + src14[66] + src14[67] + src14[68] + src14[69] + src14[70] + src14[71] + src14[72] + src14[73] + src14[74] + src14[75] + src14[76] + src14[77] + src14[78] + src14[79] + src14[80] + src14[81] + src14[82] + src14[83] + src14[84] + src14[85] + src14[86] + src14[87] + src14[88] + src14[89] + src14[90] + src14[91] + src14[92] + src14[93] + src14[94] + src14[95] + src14[96] + src14[97] + src14[98] + src14[99] + src14[100] + src14[101] + src14[102] + src14[103] + src14[104] + src14[105] + src14[106] + src14[107] + src14[108] + src14[109] + src14[110] + src14[111] + src14[112] + src14[113] + src14[114] + src14[115] + src14[116] + src14[117] + src14[118] + src14[119] + src14[120] + src14[121] + src14[122] + src14[123] + src14[124] + src14[125] + src14[126] + src14[127] + src14[128] + src14[129] + src14[130] + src14[131] + src14[132] + src14[133] + src14[134] + src14[135] + src14[136] + src14[137] + src14[138] + src14[139] + src14[140] + src14[141] + src14[142] + src14[143] + src14[144] + src14[145] + src14[146] + src14[147] + src14[148] + src14[149] + src14[150] + src14[151] + src14[152] + src14[153] + src14[154] + src14[155] + src14[156] + src14[157] + src14[158] + src14[159] + src14[160] + src14[161])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15] + src15[16] + src15[17] + src15[18] + src15[19] + src15[20] + src15[21] + src15[22] + src15[23] + src15[24] + src15[25] + src15[26] + src15[27] + src15[28] + src15[29] + src15[30] + src15[31] + src15[32] + src15[33] + src15[34] + src15[35] + src15[36] + src15[37] + src15[38] + src15[39] + src15[40] + src15[41] + src15[42] + src15[43] + src15[44] + src15[45] + src15[46] + src15[47] + src15[48] + src15[49] + src15[50] + src15[51] + src15[52] + src15[53] + src15[54] + src15[55] + src15[56] + src15[57] + src15[58] + src15[59] + src15[60] + src15[61] + src15[62] + src15[63] + src15[64] + src15[65] + src15[66] + src15[67] + src15[68] + src15[69] + src15[70] + src15[71] + src15[72] + src15[73] + src15[74] + src15[75] + src15[76] + src15[77] + src15[78] + src15[79] + src15[80] + src15[81] + src15[82] + src15[83] + src15[84] + src15[85] + src15[86] + src15[87] + src15[88] + src15[89] + src15[90] + src15[91] + src15[92] + src15[93] + src15[94] + src15[95] + src15[96] + src15[97] + src15[98] + src15[99] + src15[100] + src15[101] + src15[102] + src15[103] + src15[104] + src15[105] + src15[106] + src15[107] + src15[108] + src15[109] + src15[110] + src15[111] + src15[112] + src15[113] + src15[114] + src15[115] + src15[116] + src15[117] + src15[118] + src15[119] + src15[120] + src15[121] + src15[122] + src15[123] + src15[124] + src15[125] + src15[126] + src15[127] + src15[128] + src15[129] + src15[130] + src15[131] + src15[132] + src15[133] + src15[134] + src15[135] + src15[136] + src15[137] + src15[138] + src15[139] + src15[140] + src15[141] + src15[142] + src15[143] + src15[144] + src15[145] + src15[146] + src15[147] + src15[148] + src15[149] + src15[150] + src15[151] + src15[152] + src15[153] + src15[154] + src15[155] + src15[156] + src15[157] + src15[158] + src15[159] + src15[160] + src15[161])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16] + src16[17] + src16[18] + src16[19] + src16[20] + src16[21] + src16[22] + src16[23] + src16[24] + src16[25] + src16[26] + src16[27] + src16[28] + src16[29] + src16[30] + src16[31] + src16[32] + src16[33] + src16[34] + src16[35] + src16[36] + src16[37] + src16[38] + src16[39] + src16[40] + src16[41] + src16[42] + src16[43] + src16[44] + src16[45] + src16[46] + src16[47] + src16[48] + src16[49] + src16[50] + src16[51] + src16[52] + src16[53] + src16[54] + src16[55] + src16[56] + src16[57] + src16[58] + src16[59] + src16[60] + src16[61] + src16[62] + src16[63] + src16[64] + src16[65] + src16[66] + src16[67] + src16[68] + src16[69] + src16[70] + src16[71] + src16[72] + src16[73] + src16[74] + src16[75] + src16[76] + src16[77] + src16[78] + src16[79] + src16[80] + src16[81] + src16[82] + src16[83] + src16[84] + src16[85] + src16[86] + src16[87] + src16[88] + src16[89] + src16[90] + src16[91] + src16[92] + src16[93] + src16[94] + src16[95] + src16[96] + src16[97] + src16[98] + src16[99] + src16[100] + src16[101] + src16[102] + src16[103] + src16[104] + src16[105] + src16[106] + src16[107] + src16[108] + src16[109] + src16[110] + src16[111] + src16[112] + src16[113] + src16[114] + src16[115] + src16[116] + src16[117] + src16[118] + src16[119] + src16[120] + src16[121] + src16[122] + src16[123] + src16[124] + src16[125] + src16[126] + src16[127] + src16[128] + src16[129] + src16[130] + src16[131] + src16[132] + src16[133] + src16[134] + src16[135] + src16[136] + src16[137] + src16[138] + src16[139] + src16[140] + src16[141] + src16[142] + src16[143] + src16[144] + src16[145] + src16[146] + src16[147] + src16[148] + src16[149] + src16[150] + src16[151] + src16[152] + src16[153] + src16[154] + src16[155] + src16[156] + src16[157] + src16[158] + src16[159] + src16[160] + src16[161])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17] + src17[18] + src17[19] + src17[20] + src17[21] + src17[22] + src17[23] + src17[24] + src17[25] + src17[26] + src17[27] + src17[28] + src17[29] + src17[30] + src17[31] + src17[32] + src17[33] + src17[34] + src17[35] + src17[36] + src17[37] + src17[38] + src17[39] + src17[40] + src17[41] + src17[42] + src17[43] + src17[44] + src17[45] + src17[46] + src17[47] + src17[48] + src17[49] + src17[50] + src17[51] + src17[52] + src17[53] + src17[54] + src17[55] + src17[56] + src17[57] + src17[58] + src17[59] + src17[60] + src17[61] + src17[62] + src17[63] + src17[64] + src17[65] + src17[66] + src17[67] + src17[68] + src17[69] + src17[70] + src17[71] + src17[72] + src17[73] + src17[74] + src17[75] + src17[76] + src17[77] + src17[78] + src17[79] + src17[80] + src17[81] + src17[82] + src17[83] + src17[84] + src17[85] + src17[86] + src17[87] + src17[88] + src17[89] + src17[90] + src17[91] + src17[92] + src17[93] + src17[94] + src17[95] + src17[96] + src17[97] + src17[98] + src17[99] + src17[100] + src17[101] + src17[102] + src17[103] + src17[104] + src17[105] + src17[106] + src17[107] + src17[108] + src17[109] + src17[110] + src17[111] + src17[112] + src17[113] + src17[114] + src17[115] + src17[116] + src17[117] + src17[118] + src17[119] + src17[120] + src17[121] + src17[122] + src17[123] + src17[124] + src17[125] + src17[126] + src17[127] + src17[128] + src17[129] + src17[130] + src17[131] + src17[132] + src17[133] + src17[134] + src17[135] + src17[136] + src17[137] + src17[138] + src17[139] + src17[140] + src17[141] + src17[142] + src17[143] + src17[144] + src17[145] + src17[146] + src17[147] + src17[148] + src17[149] + src17[150] + src17[151] + src17[152] + src17[153] + src17[154] + src17[155] + src17[156] + src17[157] + src17[158] + src17[159] + src17[160] + src17[161])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15] + src18[16] + src18[17] + src18[18] + src18[19] + src18[20] + src18[21] + src18[22] + src18[23] + src18[24] + src18[25] + src18[26] + src18[27] + src18[28] + src18[29] + src18[30] + src18[31] + src18[32] + src18[33] + src18[34] + src18[35] + src18[36] + src18[37] + src18[38] + src18[39] + src18[40] + src18[41] + src18[42] + src18[43] + src18[44] + src18[45] + src18[46] + src18[47] + src18[48] + src18[49] + src18[50] + src18[51] + src18[52] + src18[53] + src18[54] + src18[55] + src18[56] + src18[57] + src18[58] + src18[59] + src18[60] + src18[61] + src18[62] + src18[63] + src18[64] + src18[65] + src18[66] + src18[67] + src18[68] + src18[69] + src18[70] + src18[71] + src18[72] + src18[73] + src18[74] + src18[75] + src18[76] + src18[77] + src18[78] + src18[79] + src18[80] + src18[81] + src18[82] + src18[83] + src18[84] + src18[85] + src18[86] + src18[87] + src18[88] + src18[89] + src18[90] + src18[91] + src18[92] + src18[93] + src18[94] + src18[95] + src18[96] + src18[97] + src18[98] + src18[99] + src18[100] + src18[101] + src18[102] + src18[103] + src18[104] + src18[105] + src18[106] + src18[107] + src18[108] + src18[109] + src18[110] + src18[111] + src18[112] + src18[113] + src18[114] + src18[115] + src18[116] + src18[117] + src18[118] + src18[119] + src18[120] + src18[121] + src18[122] + src18[123] + src18[124] + src18[125] + src18[126] + src18[127] + src18[128] + src18[129] + src18[130] + src18[131] + src18[132] + src18[133] + src18[134] + src18[135] + src18[136] + src18[137] + src18[138] + src18[139] + src18[140] + src18[141] + src18[142] + src18[143] + src18[144] + src18[145] + src18[146] + src18[147] + src18[148] + src18[149] + src18[150] + src18[151] + src18[152] + src18[153] + src18[154] + src18[155] + src18[156] + src18[157] + src18[158] + src18[159] + src18[160] + src18[161])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13] + src19[14] + src19[15] + src19[16] + src19[17] + src19[18] + src19[19] + src19[20] + src19[21] + src19[22] + src19[23] + src19[24] + src19[25] + src19[26] + src19[27] + src19[28] + src19[29] + src19[30] + src19[31] + src19[32] + src19[33] + src19[34] + src19[35] + src19[36] + src19[37] + src19[38] + src19[39] + src19[40] + src19[41] + src19[42] + src19[43] + src19[44] + src19[45] + src19[46] + src19[47] + src19[48] + src19[49] + src19[50] + src19[51] + src19[52] + src19[53] + src19[54] + src19[55] + src19[56] + src19[57] + src19[58] + src19[59] + src19[60] + src19[61] + src19[62] + src19[63] + src19[64] + src19[65] + src19[66] + src19[67] + src19[68] + src19[69] + src19[70] + src19[71] + src19[72] + src19[73] + src19[74] + src19[75] + src19[76] + src19[77] + src19[78] + src19[79] + src19[80] + src19[81] + src19[82] + src19[83] + src19[84] + src19[85] + src19[86] + src19[87] + src19[88] + src19[89] + src19[90] + src19[91] + src19[92] + src19[93] + src19[94] + src19[95] + src19[96] + src19[97] + src19[98] + src19[99] + src19[100] + src19[101] + src19[102] + src19[103] + src19[104] + src19[105] + src19[106] + src19[107] + src19[108] + src19[109] + src19[110] + src19[111] + src19[112] + src19[113] + src19[114] + src19[115] + src19[116] + src19[117] + src19[118] + src19[119] + src19[120] + src19[121] + src19[122] + src19[123] + src19[124] + src19[125] + src19[126] + src19[127] + src19[128] + src19[129] + src19[130] + src19[131] + src19[132] + src19[133] + src19[134] + src19[135] + src19[136] + src19[137] + src19[138] + src19[139] + src19[140] + src19[141] + src19[142] + src19[143] + src19[144] + src19[145] + src19[146] + src19[147] + src19[148] + src19[149] + src19[150] + src19[151] + src19[152] + src19[153] + src19[154] + src19[155] + src19[156] + src19[157] + src19[158] + src19[159] + src19[160] + src19[161])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6] + src20[7] + src20[8] + src20[9] + src20[10] + src20[11] + src20[12] + src20[13] + src20[14] + src20[15] + src20[16] + src20[17] + src20[18] + src20[19] + src20[20] + src20[21] + src20[22] + src20[23] + src20[24] + src20[25] + src20[26] + src20[27] + src20[28] + src20[29] + src20[30] + src20[31] + src20[32] + src20[33] + src20[34] + src20[35] + src20[36] + src20[37] + src20[38] + src20[39] + src20[40] + src20[41] + src20[42] + src20[43] + src20[44] + src20[45] + src20[46] + src20[47] + src20[48] + src20[49] + src20[50] + src20[51] + src20[52] + src20[53] + src20[54] + src20[55] + src20[56] + src20[57] + src20[58] + src20[59] + src20[60] + src20[61] + src20[62] + src20[63] + src20[64] + src20[65] + src20[66] + src20[67] + src20[68] + src20[69] + src20[70] + src20[71] + src20[72] + src20[73] + src20[74] + src20[75] + src20[76] + src20[77] + src20[78] + src20[79] + src20[80] + src20[81] + src20[82] + src20[83] + src20[84] + src20[85] + src20[86] + src20[87] + src20[88] + src20[89] + src20[90] + src20[91] + src20[92] + src20[93] + src20[94] + src20[95] + src20[96] + src20[97] + src20[98] + src20[99] + src20[100] + src20[101] + src20[102] + src20[103] + src20[104] + src20[105] + src20[106] + src20[107] + src20[108] + src20[109] + src20[110] + src20[111] + src20[112] + src20[113] + src20[114] + src20[115] + src20[116] + src20[117] + src20[118] + src20[119] + src20[120] + src20[121] + src20[122] + src20[123] + src20[124] + src20[125] + src20[126] + src20[127] + src20[128] + src20[129] + src20[130] + src20[131] + src20[132] + src20[133] + src20[134] + src20[135] + src20[136] + src20[137] + src20[138] + src20[139] + src20[140] + src20[141] + src20[142] + src20[143] + src20[144] + src20[145] + src20[146] + src20[147] + src20[148] + src20[149] + src20[150] + src20[151] + src20[152] + src20[153] + src20[154] + src20[155] + src20[156] + src20[157] + src20[158] + src20[159] + src20[160] + src20[161])<<20) + ((src21[0] + src21[1] + src21[2] + src21[3] + src21[4] + src21[5] + src21[6] + src21[7] + src21[8] + src21[9] + src21[10] + src21[11] + src21[12] + src21[13] + src21[14] + src21[15] + src21[16] + src21[17] + src21[18] + src21[19] + src21[20] + src21[21] + src21[22] + src21[23] + src21[24] + src21[25] + src21[26] + src21[27] + src21[28] + src21[29] + src21[30] + src21[31] + src21[32] + src21[33] + src21[34] + src21[35] + src21[36] + src21[37] + src21[38] + src21[39] + src21[40] + src21[41] + src21[42] + src21[43] + src21[44] + src21[45] + src21[46] + src21[47] + src21[48] + src21[49] + src21[50] + src21[51] + src21[52] + src21[53] + src21[54] + src21[55] + src21[56] + src21[57] + src21[58] + src21[59] + src21[60] + src21[61] + src21[62] + src21[63] + src21[64] + src21[65] + src21[66] + src21[67] + src21[68] + src21[69] + src21[70] + src21[71] + src21[72] + src21[73] + src21[74] + src21[75] + src21[76] + src21[77] + src21[78] + src21[79] + src21[80] + src21[81] + src21[82] + src21[83] + src21[84] + src21[85] + src21[86] + src21[87] + src21[88] + src21[89] + src21[90] + src21[91] + src21[92] + src21[93] + src21[94] + src21[95] + src21[96] + src21[97] + src21[98] + src21[99] + src21[100] + src21[101] + src21[102] + src21[103] + src21[104] + src21[105] + src21[106] + src21[107] + src21[108] + src21[109] + src21[110] + src21[111] + src21[112] + src21[113] + src21[114] + src21[115] + src21[116] + src21[117] + src21[118] + src21[119] + src21[120] + src21[121] + src21[122] + src21[123] + src21[124] + src21[125] + src21[126] + src21[127] + src21[128] + src21[129] + src21[130] + src21[131] + src21[132] + src21[133] + src21[134] + src21[135] + src21[136] + src21[137] + src21[138] + src21[139] + src21[140] + src21[141] + src21[142] + src21[143] + src21[144] + src21[145] + src21[146] + src21[147] + src21[148] + src21[149] + src21[150] + src21[151] + src21[152] + src21[153] + src21[154] + src21[155] + src21[156] + src21[157] + src21[158] + src21[159] + src21[160] + src21[161])<<21) + ((src22[0] + src22[1] + src22[2] + src22[3] + src22[4] + src22[5] + src22[6] + src22[7] + src22[8] + src22[9] + src22[10] + src22[11] + src22[12] + src22[13] + src22[14] + src22[15] + src22[16] + src22[17] + src22[18] + src22[19] + src22[20] + src22[21] + src22[22] + src22[23] + src22[24] + src22[25] + src22[26] + src22[27] + src22[28] + src22[29] + src22[30] + src22[31] + src22[32] + src22[33] + src22[34] + src22[35] + src22[36] + src22[37] + src22[38] + src22[39] + src22[40] + src22[41] + src22[42] + src22[43] + src22[44] + src22[45] + src22[46] + src22[47] + src22[48] + src22[49] + src22[50] + src22[51] + src22[52] + src22[53] + src22[54] + src22[55] + src22[56] + src22[57] + src22[58] + src22[59] + src22[60] + src22[61] + src22[62] + src22[63] + src22[64] + src22[65] + src22[66] + src22[67] + src22[68] + src22[69] + src22[70] + src22[71] + src22[72] + src22[73] + src22[74] + src22[75] + src22[76] + src22[77] + src22[78] + src22[79] + src22[80] + src22[81] + src22[82] + src22[83] + src22[84] + src22[85] + src22[86] + src22[87] + src22[88] + src22[89] + src22[90] + src22[91] + src22[92] + src22[93] + src22[94] + src22[95] + src22[96] + src22[97] + src22[98] + src22[99] + src22[100] + src22[101] + src22[102] + src22[103] + src22[104] + src22[105] + src22[106] + src22[107] + src22[108] + src22[109] + src22[110] + src22[111] + src22[112] + src22[113] + src22[114] + src22[115] + src22[116] + src22[117] + src22[118] + src22[119] + src22[120] + src22[121] + src22[122] + src22[123] + src22[124] + src22[125] + src22[126] + src22[127] + src22[128] + src22[129] + src22[130] + src22[131] + src22[132] + src22[133] + src22[134] + src22[135] + src22[136] + src22[137] + src22[138] + src22[139] + src22[140] + src22[141] + src22[142] + src22[143] + src22[144] + src22[145] + src22[146] + src22[147] + src22[148] + src22[149] + src22[150] + src22[151] + src22[152] + src22[153] + src22[154] + src22[155] + src22[156] + src22[157] + src22[158] + src22[159] + src22[160] + src22[161])<<22) + ((src23[0] + src23[1] + src23[2] + src23[3] + src23[4] + src23[5] + src23[6] + src23[7] + src23[8] + src23[9] + src23[10] + src23[11] + src23[12] + src23[13] + src23[14] + src23[15] + src23[16] + src23[17] + src23[18] + src23[19] + src23[20] + src23[21] + src23[22] + src23[23] + src23[24] + src23[25] + src23[26] + src23[27] + src23[28] + src23[29] + src23[30] + src23[31] + src23[32] + src23[33] + src23[34] + src23[35] + src23[36] + src23[37] + src23[38] + src23[39] + src23[40] + src23[41] + src23[42] + src23[43] + src23[44] + src23[45] + src23[46] + src23[47] + src23[48] + src23[49] + src23[50] + src23[51] + src23[52] + src23[53] + src23[54] + src23[55] + src23[56] + src23[57] + src23[58] + src23[59] + src23[60] + src23[61] + src23[62] + src23[63] + src23[64] + src23[65] + src23[66] + src23[67] + src23[68] + src23[69] + src23[70] + src23[71] + src23[72] + src23[73] + src23[74] + src23[75] + src23[76] + src23[77] + src23[78] + src23[79] + src23[80] + src23[81] + src23[82] + src23[83] + src23[84] + src23[85] + src23[86] + src23[87] + src23[88] + src23[89] + src23[90] + src23[91] + src23[92] + src23[93] + src23[94] + src23[95] + src23[96] + src23[97] + src23[98] + src23[99] + src23[100] + src23[101] + src23[102] + src23[103] + src23[104] + src23[105] + src23[106] + src23[107] + src23[108] + src23[109] + src23[110] + src23[111] + src23[112] + src23[113] + src23[114] + src23[115] + src23[116] + src23[117] + src23[118] + src23[119] + src23[120] + src23[121] + src23[122] + src23[123] + src23[124] + src23[125] + src23[126] + src23[127] + src23[128] + src23[129] + src23[130] + src23[131] + src23[132] + src23[133] + src23[134] + src23[135] + src23[136] + src23[137] + src23[138] + src23[139] + src23[140] + src23[141] + src23[142] + src23[143] + src23[144] + src23[145] + src23[146] + src23[147] + src23[148] + src23[149] + src23[150] + src23[151] + src23[152] + src23[153] + src23[154] + src23[155] + src23[156] + src23[157] + src23[158] + src23[159] + src23[160] + src23[161])<<23) + ((src24[0] + src24[1] + src24[2] + src24[3] + src24[4] + src24[5] + src24[6] + src24[7] + src24[8] + src24[9] + src24[10] + src24[11] + src24[12] + src24[13] + src24[14] + src24[15] + src24[16] + src24[17] + src24[18] + src24[19] + src24[20] + src24[21] + src24[22] + src24[23] + src24[24] + src24[25] + src24[26] + src24[27] + src24[28] + src24[29] + src24[30] + src24[31] + src24[32] + src24[33] + src24[34] + src24[35] + src24[36] + src24[37] + src24[38] + src24[39] + src24[40] + src24[41] + src24[42] + src24[43] + src24[44] + src24[45] + src24[46] + src24[47] + src24[48] + src24[49] + src24[50] + src24[51] + src24[52] + src24[53] + src24[54] + src24[55] + src24[56] + src24[57] + src24[58] + src24[59] + src24[60] + src24[61] + src24[62] + src24[63] + src24[64] + src24[65] + src24[66] + src24[67] + src24[68] + src24[69] + src24[70] + src24[71] + src24[72] + src24[73] + src24[74] + src24[75] + src24[76] + src24[77] + src24[78] + src24[79] + src24[80] + src24[81] + src24[82] + src24[83] + src24[84] + src24[85] + src24[86] + src24[87] + src24[88] + src24[89] + src24[90] + src24[91] + src24[92] + src24[93] + src24[94] + src24[95] + src24[96] + src24[97] + src24[98] + src24[99] + src24[100] + src24[101] + src24[102] + src24[103] + src24[104] + src24[105] + src24[106] + src24[107] + src24[108] + src24[109] + src24[110] + src24[111] + src24[112] + src24[113] + src24[114] + src24[115] + src24[116] + src24[117] + src24[118] + src24[119] + src24[120] + src24[121] + src24[122] + src24[123] + src24[124] + src24[125] + src24[126] + src24[127] + src24[128] + src24[129] + src24[130] + src24[131] + src24[132] + src24[133] + src24[134] + src24[135] + src24[136] + src24[137] + src24[138] + src24[139] + src24[140] + src24[141] + src24[142] + src24[143] + src24[144] + src24[145] + src24[146] + src24[147] + src24[148] + src24[149] + src24[150] + src24[151] + src24[152] + src24[153] + src24[154] + src24[155] + src24[156] + src24[157] + src24[158] + src24[159] + src24[160] + src24[161])<<24) + ((src25[0] + src25[1] + src25[2] + src25[3] + src25[4] + src25[5] + src25[6] + src25[7] + src25[8] + src25[9] + src25[10] + src25[11] + src25[12] + src25[13] + src25[14] + src25[15] + src25[16] + src25[17] + src25[18] + src25[19] + src25[20] + src25[21] + src25[22] + src25[23] + src25[24] + src25[25] + src25[26] + src25[27] + src25[28] + src25[29] + src25[30] + src25[31] + src25[32] + src25[33] + src25[34] + src25[35] + src25[36] + src25[37] + src25[38] + src25[39] + src25[40] + src25[41] + src25[42] + src25[43] + src25[44] + src25[45] + src25[46] + src25[47] + src25[48] + src25[49] + src25[50] + src25[51] + src25[52] + src25[53] + src25[54] + src25[55] + src25[56] + src25[57] + src25[58] + src25[59] + src25[60] + src25[61] + src25[62] + src25[63] + src25[64] + src25[65] + src25[66] + src25[67] + src25[68] + src25[69] + src25[70] + src25[71] + src25[72] + src25[73] + src25[74] + src25[75] + src25[76] + src25[77] + src25[78] + src25[79] + src25[80] + src25[81] + src25[82] + src25[83] + src25[84] + src25[85] + src25[86] + src25[87] + src25[88] + src25[89] + src25[90] + src25[91] + src25[92] + src25[93] + src25[94] + src25[95] + src25[96] + src25[97] + src25[98] + src25[99] + src25[100] + src25[101] + src25[102] + src25[103] + src25[104] + src25[105] + src25[106] + src25[107] + src25[108] + src25[109] + src25[110] + src25[111] + src25[112] + src25[113] + src25[114] + src25[115] + src25[116] + src25[117] + src25[118] + src25[119] + src25[120] + src25[121] + src25[122] + src25[123] + src25[124] + src25[125] + src25[126] + src25[127] + src25[128] + src25[129] + src25[130] + src25[131] + src25[132] + src25[133] + src25[134] + src25[135] + src25[136] + src25[137] + src25[138] + src25[139] + src25[140] + src25[141] + src25[142] + src25[143] + src25[144] + src25[145] + src25[146] + src25[147] + src25[148] + src25[149] + src25[150] + src25[151] + src25[152] + src25[153] + src25[154] + src25[155] + src25[156] + src25[157] + src25[158] + src25[159] + src25[160] + src25[161])<<25) + ((src26[0] + src26[1] + src26[2] + src26[3] + src26[4] + src26[5] + src26[6] + src26[7] + src26[8] + src26[9] + src26[10] + src26[11] + src26[12] + src26[13] + src26[14] + src26[15] + src26[16] + src26[17] + src26[18] + src26[19] + src26[20] + src26[21] + src26[22] + src26[23] + src26[24] + src26[25] + src26[26] + src26[27] + src26[28] + src26[29] + src26[30] + src26[31] + src26[32] + src26[33] + src26[34] + src26[35] + src26[36] + src26[37] + src26[38] + src26[39] + src26[40] + src26[41] + src26[42] + src26[43] + src26[44] + src26[45] + src26[46] + src26[47] + src26[48] + src26[49] + src26[50] + src26[51] + src26[52] + src26[53] + src26[54] + src26[55] + src26[56] + src26[57] + src26[58] + src26[59] + src26[60] + src26[61] + src26[62] + src26[63] + src26[64] + src26[65] + src26[66] + src26[67] + src26[68] + src26[69] + src26[70] + src26[71] + src26[72] + src26[73] + src26[74] + src26[75] + src26[76] + src26[77] + src26[78] + src26[79] + src26[80] + src26[81] + src26[82] + src26[83] + src26[84] + src26[85] + src26[86] + src26[87] + src26[88] + src26[89] + src26[90] + src26[91] + src26[92] + src26[93] + src26[94] + src26[95] + src26[96] + src26[97] + src26[98] + src26[99] + src26[100] + src26[101] + src26[102] + src26[103] + src26[104] + src26[105] + src26[106] + src26[107] + src26[108] + src26[109] + src26[110] + src26[111] + src26[112] + src26[113] + src26[114] + src26[115] + src26[116] + src26[117] + src26[118] + src26[119] + src26[120] + src26[121] + src26[122] + src26[123] + src26[124] + src26[125] + src26[126] + src26[127] + src26[128] + src26[129] + src26[130] + src26[131] + src26[132] + src26[133] + src26[134] + src26[135] + src26[136] + src26[137] + src26[138] + src26[139] + src26[140] + src26[141] + src26[142] + src26[143] + src26[144] + src26[145] + src26[146] + src26[147] + src26[148] + src26[149] + src26[150] + src26[151] + src26[152] + src26[153] + src26[154] + src26[155] + src26[156] + src26[157] + src26[158] + src26[159] + src26[160] + src26[161])<<26) + ((src27[0] + src27[1] + src27[2] + src27[3] + src27[4] + src27[5] + src27[6] + src27[7] + src27[8] + src27[9] + src27[10] + src27[11] + src27[12] + src27[13] + src27[14] + src27[15] + src27[16] + src27[17] + src27[18] + src27[19] + src27[20] + src27[21] + src27[22] + src27[23] + src27[24] + src27[25] + src27[26] + src27[27] + src27[28] + src27[29] + src27[30] + src27[31] + src27[32] + src27[33] + src27[34] + src27[35] + src27[36] + src27[37] + src27[38] + src27[39] + src27[40] + src27[41] + src27[42] + src27[43] + src27[44] + src27[45] + src27[46] + src27[47] + src27[48] + src27[49] + src27[50] + src27[51] + src27[52] + src27[53] + src27[54] + src27[55] + src27[56] + src27[57] + src27[58] + src27[59] + src27[60] + src27[61] + src27[62] + src27[63] + src27[64] + src27[65] + src27[66] + src27[67] + src27[68] + src27[69] + src27[70] + src27[71] + src27[72] + src27[73] + src27[74] + src27[75] + src27[76] + src27[77] + src27[78] + src27[79] + src27[80] + src27[81] + src27[82] + src27[83] + src27[84] + src27[85] + src27[86] + src27[87] + src27[88] + src27[89] + src27[90] + src27[91] + src27[92] + src27[93] + src27[94] + src27[95] + src27[96] + src27[97] + src27[98] + src27[99] + src27[100] + src27[101] + src27[102] + src27[103] + src27[104] + src27[105] + src27[106] + src27[107] + src27[108] + src27[109] + src27[110] + src27[111] + src27[112] + src27[113] + src27[114] + src27[115] + src27[116] + src27[117] + src27[118] + src27[119] + src27[120] + src27[121] + src27[122] + src27[123] + src27[124] + src27[125] + src27[126] + src27[127] + src27[128] + src27[129] + src27[130] + src27[131] + src27[132] + src27[133] + src27[134] + src27[135] + src27[136] + src27[137] + src27[138] + src27[139] + src27[140] + src27[141] + src27[142] + src27[143] + src27[144] + src27[145] + src27[146] + src27[147] + src27[148] + src27[149] + src27[150] + src27[151] + src27[152] + src27[153] + src27[154] + src27[155] + src27[156] + src27[157] + src27[158] + src27[159] + src27[160] + src27[161])<<27) + ((src28[0] + src28[1] + src28[2] + src28[3] + src28[4] + src28[5] + src28[6] + src28[7] + src28[8] + src28[9] + src28[10] + src28[11] + src28[12] + src28[13] + src28[14] + src28[15] + src28[16] + src28[17] + src28[18] + src28[19] + src28[20] + src28[21] + src28[22] + src28[23] + src28[24] + src28[25] + src28[26] + src28[27] + src28[28] + src28[29] + src28[30] + src28[31] + src28[32] + src28[33] + src28[34] + src28[35] + src28[36] + src28[37] + src28[38] + src28[39] + src28[40] + src28[41] + src28[42] + src28[43] + src28[44] + src28[45] + src28[46] + src28[47] + src28[48] + src28[49] + src28[50] + src28[51] + src28[52] + src28[53] + src28[54] + src28[55] + src28[56] + src28[57] + src28[58] + src28[59] + src28[60] + src28[61] + src28[62] + src28[63] + src28[64] + src28[65] + src28[66] + src28[67] + src28[68] + src28[69] + src28[70] + src28[71] + src28[72] + src28[73] + src28[74] + src28[75] + src28[76] + src28[77] + src28[78] + src28[79] + src28[80] + src28[81] + src28[82] + src28[83] + src28[84] + src28[85] + src28[86] + src28[87] + src28[88] + src28[89] + src28[90] + src28[91] + src28[92] + src28[93] + src28[94] + src28[95] + src28[96] + src28[97] + src28[98] + src28[99] + src28[100] + src28[101] + src28[102] + src28[103] + src28[104] + src28[105] + src28[106] + src28[107] + src28[108] + src28[109] + src28[110] + src28[111] + src28[112] + src28[113] + src28[114] + src28[115] + src28[116] + src28[117] + src28[118] + src28[119] + src28[120] + src28[121] + src28[122] + src28[123] + src28[124] + src28[125] + src28[126] + src28[127] + src28[128] + src28[129] + src28[130] + src28[131] + src28[132] + src28[133] + src28[134] + src28[135] + src28[136] + src28[137] + src28[138] + src28[139] + src28[140] + src28[141] + src28[142] + src28[143] + src28[144] + src28[145] + src28[146] + src28[147] + src28[148] + src28[149] + src28[150] + src28[151] + src28[152] + src28[153] + src28[154] + src28[155] + src28[156] + src28[157] + src28[158] + src28[159] + src28[160] + src28[161])<<28) + ((src29[0] + src29[1] + src29[2] + src29[3] + src29[4] + src29[5] + src29[6] + src29[7] + src29[8] + src29[9] + src29[10] + src29[11] + src29[12] + src29[13] + src29[14] + src29[15] + src29[16] + src29[17] + src29[18] + src29[19] + src29[20] + src29[21] + src29[22] + src29[23] + src29[24] + src29[25] + src29[26] + src29[27] + src29[28] + src29[29] + src29[30] + src29[31] + src29[32] + src29[33] + src29[34] + src29[35] + src29[36] + src29[37] + src29[38] + src29[39] + src29[40] + src29[41] + src29[42] + src29[43] + src29[44] + src29[45] + src29[46] + src29[47] + src29[48] + src29[49] + src29[50] + src29[51] + src29[52] + src29[53] + src29[54] + src29[55] + src29[56] + src29[57] + src29[58] + src29[59] + src29[60] + src29[61] + src29[62] + src29[63] + src29[64] + src29[65] + src29[66] + src29[67] + src29[68] + src29[69] + src29[70] + src29[71] + src29[72] + src29[73] + src29[74] + src29[75] + src29[76] + src29[77] + src29[78] + src29[79] + src29[80] + src29[81] + src29[82] + src29[83] + src29[84] + src29[85] + src29[86] + src29[87] + src29[88] + src29[89] + src29[90] + src29[91] + src29[92] + src29[93] + src29[94] + src29[95] + src29[96] + src29[97] + src29[98] + src29[99] + src29[100] + src29[101] + src29[102] + src29[103] + src29[104] + src29[105] + src29[106] + src29[107] + src29[108] + src29[109] + src29[110] + src29[111] + src29[112] + src29[113] + src29[114] + src29[115] + src29[116] + src29[117] + src29[118] + src29[119] + src29[120] + src29[121] + src29[122] + src29[123] + src29[124] + src29[125] + src29[126] + src29[127] + src29[128] + src29[129] + src29[130] + src29[131] + src29[132] + src29[133] + src29[134] + src29[135] + src29[136] + src29[137] + src29[138] + src29[139] + src29[140] + src29[141] + src29[142] + src29[143] + src29[144] + src29[145] + src29[146] + src29[147] + src29[148] + src29[149] + src29[150] + src29[151] + src29[152] + src29[153] + src29[154] + src29[155] + src29[156] + src29[157] + src29[158] + src29[159] + src29[160] + src29[161])<<29) + ((src30[0] + src30[1] + src30[2] + src30[3] + src30[4] + src30[5] + src30[6] + src30[7] + src30[8] + src30[9] + src30[10] + src30[11] + src30[12] + src30[13] + src30[14] + src30[15] + src30[16] + src30[17] + src30[18] + src30[19] + src30[20] + src30[21] + src30[22] + src30[23] + src30[24] + src30[25] + src30[26] + src30[27] + src30[28] + src30[29] + src30[30] + src30[31] + src30[32] + src30[33] + src30[34] + src30[35] + src30[36] + src30[37] + src30[38] + src30[39] + src30[40] + src30[41] + src30[42] + src30[43] + src30[44] + src30[45] + src30[46] + src30[47] + src30[48] + src30[49] + src30[50] + src30[51] + src30[52] + src30[53] + src30[54] + src30[55] + src30[56] + src30[57] + src30[58] + src30[59] + src30[60] + src30[61] + src30[62] + src30[63] + src30[64] + src30[65] + src30[66] + src30[67] + src30[68] + src30[69] + src30[70] + src30[71] + src30[72] + src30[73] + src30[74] + src30[75] + src30[76] + src30[77] + src30[78] + src30[79] + src30[80] + src30[81] + src30[82] + src30[83] + src30[84] + src30[85] + src30[86] + src30[87] + src30[88] + src30[89] + src30[90] + src30[91] + src30[92] + src30[93] + src30[94] + src30[95] + src30[96] + src30[97] + src30[98] + src30[99] + src30[100] + src30[101] + src30[102] + src30[103] + src30[104] + src30[105] + src30[106] + src30[107] + src30[108] + src30[109] + src30[110] + src30[111] + src30[112] + src30[113] + src30[114] + src30[115] + src30[116] + src30[117] + src30[118] + src30[119] + src30[120] + src30[121] + src30[122] + src30[123] + src30[124] + src30[125] + src30[126] + src30[127] + src30[128] + src30[129] + src30[130] + src30[131] + src30[132] + src30[133] + src30[134] + src30[135] + src30[136] + src30[137] + src30[138] + src30[139] + src30[140] + src30[141] + src30[142] + src30[143] + src30[144] + src30[145] + src30[146] + src30[147] + src30[148] + src30[149] + src30[150] + src30[151] + src30[152] + src30[153] + src30[154] + src30[155] + src30[156] + src30[157] + src30[158] + src30[159] + src30[160] + src30[161])<<30) + ((src31[0] + src31[1] + src31[2] + src31[3] + src31[4] + src31[5] + src31[6] + src31[7] + src31[8] + src31[9] + src31[10] + src31[11] + src31[12] + src31[13] + src31[14] + src31[15] + src31[16] + src31[17] + src31[18] + src31[19] + src31[20] + src31[21] + src31[22] + src31[23] + src31[24] + src31[25] + src31[26] + src31[27] + src31[28] + src31[29] + src31[30] + src31[31] + src31[32] + src31[33] + src31[34] + src31[35] + src31[36] + src31[37] + src31[38] + src31[39] + src31[40] + src31[41] + src31[42] + src31[43] + src31[44] + src31[45] + src31[46] + src31[47] + src31[48] + src31[49] + src31[50] + src31[51] + src31[52] + src31[53] + src31[54] + src31[55] + src31[56] + src31[57] + src31[58] + src31[59] + src31[60] + src31[61] + src31[62] + src31[63] + src31[64] + src31[65] + src31[66] + src31[67] + src31[68] + src31[69] + src31[70] + src31[71] + src31[72] + src31[73] + src31[74] + src31[75] + src31[76] + src31[77] + src31[78] + src31[79] + src31[80] + src31[81] + src31[82] + src31[83] + src31[84] + src31[85] + src31[86] + src31[87] + src31[88] + src31[89] + src31[90] + src31[91] + src31[92] + src31[93] + src31[94] + src31[95] + src31[96] + src31[97] + src31[98] + src31[99] + src31[100] + src31[101] + src31[102] + src31[103] + src31[104] + src31[105] + src31[106] + src31[107] + src31[108] + src31[109] + src31[110] + src31[111] + src31[112] + src31[113] + src31[114] + src31[115] + src31[116] + src31[117] + src31[118] + src31[119] + src31[120] + src31[121] + src31[122] + src31[123] + src31[124] + src31[125] + src31[126] + src31[127] + src31[128] + src31[129] + src31[130] + src31[131] + src31[132] + src31[133] + src31[134] + src31[135] + src31[136] + src31[137] + src31[138] + src31[139] + src31[140] + src31[141] + src31[142] + src31[143] + src31[144] + src31[145] + src31[146] + src31[147] + src31[148] + src31[149] + src31[150] + src31[151] + src31[152] + src31[153] + src31[154] + src31[155] + src31[156] + src31[157] + src31[158] + src31[159] + src31[160] + src31[161])<<31);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25) + ((dst26[0])<<26) + ((dst27[0])<<27) + ((dst28[0])<<28) + ((dst29[0])<<29) + ((dst30[0])<<30) + ((dst31[0])<<31) + ((dst32[0])<<32) + ((dst33[0])<<33) + ((dst34[0])<<34) + ((dst35[0])<<35) + ((dst36[0])<<36) + ((dst37[0])<<37) + ((dst38[0])<<38) + ((dst39[0])<<39);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'h0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'h781b78ad6d49ee2532823b0fb44e949e625363e2e16f2b8312f31de8218167165dd1d410536aef47384995a60daa703e634604eefb0881ff85ba69d1524fa85f285c0095b21122e1d9ce5828242e25e18b2849e2d4de8b3d6b35b1ab6602d694fcf7898c1f7bed92d519936e25d4eb9da2a323267dc98c3b68e2d108ae1660f327fe9c9ffccdbef2f387fa44ccffe499445c8b3ead8a0b336c953c91e17d8042c273824a9a67a3682d3f12fdf91bffb01549452cd0b768cdbda3fb994d1f6836d0dd8c76806eec7cb19fb6a0e81bb719a38fd48415525e2cd8bb8fa477d7cd7881b5861a01ad0c434276d624feb57574f8dd4275347a597fe40353872c57cd72f82c708ee3c6562fd2e58d8d2f6c79eac378e6da34cf8c0a6cd980fc99b86aa93d8f2341b3e32aa032ccf06e8153da9e73d62a800930db29cd68cd98a1798beb361eaf0e80956a0a4ad527e3b893b3328bdc88c8d0b2129099054a9ca888d7c737aafe0e6ccfade92f876d39aee343cd63e15a1075559c13c1b214833ab434e4124643d0ff5a4ccdfc34d215ba0c26871126680eb27379a8bb77b013c698dd06b90053124fd9f50b30f3e197214ac171c48ce8efdaf956afe8fd51237032f29d9bd75482d584f6a77bc34af017fa902921df5803bd66a50a26126d42eda14eacbd055b235bcbdae1dbce142944f65b5d4bdc80c5e14ef8d3cf4eacf55580cb2734088b8997d1ae128db8c43f6c00a12a95d4061b78293748624cd8046e1a7fb8a12e7f062ef210391b659633b788d6f93ec7ed61b4e5fdb76b49256a1a45d75a44296ac246c54e67ce2f74524586daba7423cff8e4cb6061b9074b1e0668942fe760ac71eba1d49517a6ca8ce89b4be40a04707eb67c24adc898440739d6627abe274949c81017e3;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'h371b07b4a2949d3605e701cf8c14b6f5c6569b5493afa63f6209513504b46ec53c8072009eced054ea79401ab39139dd848e545271cb571b63d39a475460d1366520e0b62457a6bc177c516ebfd7f516e211eb51b193483a44d7b1fa00f5130ba5254dbf9b2f55a40cc45ba78ff16b7c6593021615fdb26b55dcaae07f6dff67cdf617095ddc7877e2d827089d9b0f617b88fdb33748e9eff15d5e26da65c663f5d50fb3aab6d6897237999d5f7f8a1029dd8c045efc14b22812588e9c2dd34b3731ed2954651f1388f3a5262cffaf7468b750df3bfa4fe5ff43e0414115c1c8596c23553e178a431e2eff3b568468e07dedb9491522b5801a44b917ee144399828cf894a7b3f5d85be6b55686ec4f10b10837638da98bec26b5dedb814a2e5e266cbdd09c39bca376cdbab85d86f2419f7737e9d841f7bc8585e881b0c044c25d6ea8155b72fea9a2ff644b47a9f089a9f3e00a406ef1466a3affe088069588e3c3ff13c61eb148e2a745f6ecc05748bdc16a865e4c3130a59b5ef570a2f5c867c96712c22fe1c40f7f3af792e2875cf4653fd978b64daec088f8a7dc5c0fd61d42ee284ad59c5481811337f37beac2e9ca7f7830c751109c8db2de2f9686cc1b4e2336280ee0b2abdd1d1e33207c56b874c93e83e73836a5d7080ecd5b16c6cf3c6d9527b6801d2869af0d414382f6e16c64bef33dfb00438d4cc2996deafc18caa25a90128842614611de41cd4e4255bb727fbb3011d3984fb86e9c9217dcf9d2df21d9f7638983b79d18083ebeede4fd5221bdbafeeb50a815a50028e0608585b223bb34159880eb9e0c466c13c55bfcbcf2eecd605444f4834ccc69e1cdfc380af2e4547c094764cb80156e82ba8b6174fc21a2943efad5af6a7df86497adf47098c4e2ef95;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'h2e8a446d0b493ffaa4629318f921f6a192fd315d8bdb40ad52cc0e103adf7987bf76621748da04c998f98b75d0da0087038588ac9a00fbf0b1ff6808e8e196f48925608622b2271410c16212792dc2b269c158cdf771119ae9d922f9f62492472fe776c898c14a10f013a817fac13af71a05ed592c9e4bbc6af08c130d0afd2d4666daab7b3e09494dd43d45b1ecdcd6505fe81c1d962b595df6a1e0d698a00f203257eb87f752f3a45ac96f2f97261398aa474ad18f6b92bfea6844b75cdad5ff3a3dba910869a9cfa4fd8399ea55507940bd4c8b90c1e83c1a0fd3c7206af79c7dc5f13d668c10f282f8302a9e8e8160decdd50adc186d3acfaefc9a41472fbcbe163d69a88e3a090df630ac2cb41fffb81c0ebb6a93c6067f8b585f1756fd0f7bb599d9b7480d143c32db0e534210f3930ba7c58bdacb1c39e26b95d333cd0ebce202b4c4c53d65c2d7ceb84ee531693984defaa45d77dcbabd839b1c4ed6eb8607d2498cac170b5de26f2859dc7c6d31598af816ee321ca8a004f3f311f8d8dcedeb916d9bd5a26789fab6f28b2c8583de856ce2698b0cc780b9d0c67a6f48243c2e31c0aa419d1943c6b34196cc4fc80580fa203024d9a61690bfce3d1a7e37c1f42722c9b2c810a215f75606946c5f418260723fbb6fb25f061bec25675aa932d8c15a02b64dd81d14436decbdad49ba5695b03c024c2f59f8cc586f49c17535a26a3d600d0937b26fcfcfb77401356596b7d86bcc868d6e172c45f8f43f3dc089b5214a9775494789da88ed3c0759c84b9e51e9d7f36fe8f1f6ca36c0d58af57d3b5d4402d023532bd4d9f2a418145857994469757acafc1506460f59d3fdacb170773d9bf89226f216505d67bce5c774bc50d0e24081451e0c41a1c88f1bffb43678bf89;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'h665290440570aa931f8c7c3f1cfed4a97a52cd815ac0b2e10a904d0bd724bd36e876aacfd45a261a120afeb22fc945547838dee1f209334f563bf0daf2e727205e65e412e96a0085c9ed2b185db9163218418672d49e4bd19bcd88e1326c2c93eb5dc1fd263375762b71bc4d7e3082d526a487818103929f1c5696c9512456e4d017f5ef47b03c7ef344dfd7610cf4399f18444587074a61fa60369603c932dfc16112ca6ecacccbc4d39b92a00608970cdebb28dbe8d38c6af0790780fe6cf14c8f70486567f88643e09f58f860a6eb22ddbb2d9664fef96688495408bd67b1af64c2d1d00c4f711daa820ddbc79bc3cb8a6efef31d56f08b430ed54abd3d7d8d93adfb4a99f08f1e20932db96ce116ca7ef38a7f98907922a60bc0a2b016831abdf9e7f992541d1bf9849e4d5e41837b16d5a97f5e43ee1f58588204eac1178b9a0dc0ae98fb7fb39ed9e629b6a6060a5f68dc1099be150f7b81001fc1236da23e485a8ce718c0d7c9bdde655b2edadfdcca838d6d17ac5e2f17ee457a0056ed8dac43f55d60424fa29f1e1a600bfdf0bc9630c03056b944e346e54f64b4dffd49cc12f3ed3b8d5c262f1a21aa9e7c04fc52af03d8cbebfa05d8370abe288b4cf3537c1409c167b84a778f56a8b69e68d75037f6270de7afccbe1459c1ad760d244949a93d884254e0f5897cf5c7b1c15e98e73ba3a28b0fdde3bd6ede5429d58585997b9aec0adb97a5e2c803e6b6c0730c2a3391fbb3eb3c5371333f347dc87d7175a728c089a6a9ae590c8dd3c69168f4d668cc2c32229ba9d1c607042901f408ca0bbcc5dfcf68d21264a600f0f16a4f2811bbc04141b86c5332abd29bcb1ad5c81de3db7f50f5f1fa651789ac1b3e9ab82e8bed59a7d34c29de8ffd7a69342c7234bc979e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'h92eb58f680bed11baa49950c31c565f4871e33d52a51c21595400597013dff991d1515743c057c1eaa1a423aa6c775cc01753fd6469f11f20f05dee873ed4e08727c78b76c41667cafc30e18afff4e235a419a3c441523a4165374efc35309c0e0f29a07f14482e1c7c97436241892a02352e605adc64ed171e511a2dc8fa03e18308ae2256ba3cae62e397225793324dd3ab856040c9316496153e73bdd1d8b91ed79eb64c8f3a8c0a4d6f1538c873ae937c6de01b544ddd0a79d60f1d8dc72d435408d107760a5188e9ff7aa0e7fb85da81056bba95e60670df728dabf462283d1c7dd1744f5543c06c55c9dc2b48d69862c9cb2e5e108efa05595a47568b916933bd6b0060731b754c82ed536cfab31f02f5a1e2e6f4b59d90872109b12fb24a4b2b5eb0fed313f510891df3accbd16fa125ba35200b3da61112343b014f22c3082a0e0b881037217fd6aac10b1387aa949e21bc8af4175268ca64fce8423e6b2498c47a2645deff500e0573e9b704623ad3fb4feba65564a7462f1bf36c467c4fa1456fe87829c6869092b6877d136e4f23953286f66a8ec40f580010c45dedd1f1b9c01ea4eec34447d452af1be1f2457505d143592a78a66dabe3da9ee0667b15774880831ec579e2d7695dea47de6f60a9d3512a21d688e85c1f60a4facf2790a342bbd25e91100a96abb280a8453a8db54fe240648cb28a6c83c88f72975f277552be1af33c0af3f38d22556c417be84ffe870332e42a0071187d605bbf9fdbe12fea91ca7ebd539317e9f8984de14aa2928d3fbd57223210c74d3a318bd85130c8ef3edf9474d8b09b8a36776db05c0e0d7b09419d3dd4a6d58b926de8ae22e3ad823bca669c9f65fb07868da63be74a5747a7e544e79c61d66d20af7d240a402c2433e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'h2190277b55bacf984f5910f6de99643d3ab3a073e8aa2857124381f378c51a2daf6e5129aa240f6608010b4c219031b1694a99af3439fa8672d197e630712aaff563ae217e8eacffe1943b948c398539077da6e83e41491d5c99d5d52590b87e9ecbb15567394a5375153f92c84e9b3d3d929e7812d6764eb4b948f99d5665101a7ee931cf7aad29a33400b632cccae6faae4dddeec73cf44dd7e4746a2d929fa6c55a872944bea8958c59fc1a8241fe47f188e932e14223d1d073e35a0eb1da81be450fdc572ffe42f7b77e231d184f004f2c2d47e191028c97280766dd29c4ffd4572fdac41cc3b85dd855080d0d496af0bb652ca2772d54655dc46278472c301a4bd8b0dfa9d35ae168a715a12b8d9aea196d9524df49f08b8049c2a2cb564a982164b5f12c5992f5220c07ed3a79a1d5df460138c5c36b8b7cf9b00906252fc3d875f7bc706c1a4f40f9cc0652bae47f236f5e5fabb2bf14408b35e341320f874c74b715fe8881a858ddf91533ca8f4348558fed671e16b56565827fb6de7ad8a049c65877d2c7b7b9f3600e4ccf70be1df22ed87017ac493b649afc835ae07c3786fa0854bc2d35061bc1c9765c9f39b614957e2f00c509db99f5d7ed906706ff558669b41b171fa6ce444de3de02cca01a8b684a234436846eb8f695fde5c10c9294ec31ce1727e46d8ae52af68d492955f1426f87430d83a8de3d4e024c59e0ede667e524a6f9e13c955cce66284bad8269910e985ee3077bb1cc848cc30d2c4932b03c925558f7166db4599dc6ad5798fde2306e9517e4ccb1b0a41008d8e39ccac3b0c332faec779c3097f59f67ee918499311bc00235492a216fc8e98ccb4758f99d05b4880fc9cc5c2787dc8e25ae827db1cdd8adcf995797f4f501020f5295a29879;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'h5dfbcccccb774760315043f8efae1a2f3f131880a118c1d0eddae7c2d81ee297c9408378e5e4d7adf9825229cfd20c83ea06dd464f9c01282be902aa834beb5734b2fb25ebd6615e07b4c3d751b6627d80c1c8953e860561abf342cbfcd57af20d682723763173c52ad2659032ecb77619d0d73661b9605fcd5a4a591c30a82a06b16b81824801ec106e21326d3cefb0827ab69c2e631eded48f153320dc857ba4dab6306fb2f5a0d034f73d78a613eaf990e578834f122380470fdeca3979795732d50eb7a507962874f6b8fbe5a2ff7414001aedd69e5c1c250c0cca31d283f5e2119e1fa04f501e962c79e4ece232be6561d189059d45a6a8f89fcdb1b6ec75cb952e811b1a44220594240165fd4862ad0678914787d8d677f0e7f2b6d53d8a20bb62e624f0a867edf678731843544123283b4c4df356d0b1eff9da40eca990c8a93f273e851c30805836677614cdb59e85ef276490179a9590491bb83a44e7a8f5445514b956c24c167c230206417042e8123f880f25ec917fae9cf5abf76ccb57bbcc082a4b8d92f6dab0a3a5ca11cf81f2a801117b86f090eafecdb0e9bf873407326e2caf0d2be641975673427e96b75217074481b8ef62e771e423819b01441229c51d86b2a4119d41166a94a615ffdbf047a08ce2f9cdb19aaf49559ecc0543820453b85eec1d3e682addcce4f40fa5a148d0ac1fa82778d22e33413833a09de9007db3cbffa90ea4d594d40a02a6768bdd57fcb71dc8d869ec9482e0f319184a0835ab481e9bd547ef89d84ab4cda9aa5c41560c6a3c73530a9f7cf9951dc8f06f5e7ac7ddcc7fbf7f06d55cc80a8ffb94770276ced4b5ff84f1464827f8405850095d1eb3481898407875a004fbcadf0754bdc9bbb8356b99e745163fc839c6e0dbe7;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'hd2f8165f3b48c5051c066e3c1c45395d2a6e5027b354edde58c9b609055bc55bd4703fe5f5ae4f055647e3c787bf2b4c49071517903c3073a255f93d2b3a9c5d7e479a329b3b310ec16a355c999a3da40cd820fa8dbe5c37cb2071cdc2b90bd3ddbb7a7807cb35f7d466d7643de0895944d472a664af767130989f18a2e65e243bd4f933565adc1551d3a8280b8e0d969787b2b70b836410f22e399eb70c9658a7f69d051fb76eb5adf330d2352ae6c9ed0eb463b13e2c6532ca55823925b577be8975ef515fbcb0f3c1ff591e3c2482a242f41b948f7328778790a4ff188cba3d92b7810ab3b788676520f47e0a126688f94a6a920cefaa3076350240831a8a527820edae309e3a1b07995b60a7beb5722b72eb81b71dfee8528a3b1ceadbf4e303f9f172f8db68fe06b34f7b06705034bd3aba490d556f4e73c8e06adfddfa24f615ec64a5f44d03c435695fa129802c47bb73042327faf699c19114b7ba15a0fc43e3e5c2d9a024be1cd9bacad96d12bc6751d518a4eb3984b0a4216dae20233a15e1bf7e43480b39050820145db5189fedb4de1540e7cd7250a8d8aad38cff63d737329957e9e4f315167383a79c0371e9875d8156ff15bd0fce75d45385252c8ed32ba5f91d61e1cbe472e0fb8663ad7ca86c7de9351cda06bc34bbc80cb841bb0669ba748b62d9971550e17cb9259b3ff390beb6f0892efdd82c3d0ccde2d0cb8952b5a72b5b8fed133f3bb44d8353a6c8ccac7e1de1d0aee5b8e10ecbb4eca04e1b290ad69933afabbb160f16830be0b715d62fa25a29a049498882abb7b24b95e4cdcbccb0caa4f2f1c1ed9d0990398282472de6109ebcbf6e2857eaf8a5fe1b32c7929358da82e564af58ce2ea0226c4756ce9c4ce82b017c53843222a6fa9c4ebe9053;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'h4f0c65b615c0ebfaef68a89bd62c3d8aaef275b40e2d0f8081ac6b8fbbfe97912d3b78c2a9a2c5e138ed5a63c2b1d74d94c6592969708975043099ee83f94fc9bd62168a67ab4f54b67ddd633304980402b17a14ff9fda2ecccbf6208ba1716e48df880605cb82fa09669cf425426b297d930655eb87d9035a96f89b4c56a9b7eb0acae00e7f78eecc6ed5ead7c5da30886f9bcf23dbab246e093341ca3ed7c6a0135c08d72ea773e97058fbb18d06366dbab8e5d884c242c857341a7c320c4493da88fc936e6974556fb18856f00f3b18097e4cd746c0014c73fe18995467dce18db06252de77dcc7d14ea36ac0951a62b13e5b1edd5e76a75ca4ffb8f901017293b9f39e37f03011750d4f72783cdd08f590620a0c6ee7cde9369e07cfcfc6c278cbc4b3795c41d2351ee75f1c8556b42f1fdb60915843f9e01c0e73a4da48cc9328503f2d66ab5e6e63a6abd7e340ebaaa5f5d054ecc6edba8a4f49e160f0e976f8035a24594ed500bed1d1a2c4a3946d9acf0c215f67fd1ebc8e63f3cc5c81ca893c242cc0dc264853fff392424613f7ceb202fd4cdb083908dc524bbeb1f7368a273fa4d70d5e2e284c6d92f674a70c19ee96713b4a6c3a6b7af604a66357c16c25dcaaec7ce7a20ddaea90a4d8af0289c71f38ba94db6420632a307aa916e1d8fa3db2653d481201846cdda19eeec472abe51037bc802089a531b9c24f3621565176f1d79d4d3f3bb361638d6fffa04994274a1f9057bce07b5aae48a974b2b382cb41f2ade57cf261dbb81a1e29080df25b1f8cbf9ac27171dd97b33e3df5f8c30b0b5efd567970735deaf87654d5a1c9bd655e8eed8ebcefc5d3f2d362051ec196301a6c55c05f46c7aac9d22266cfd4bf67a98893c34a9181335810b40e19ce3b6dc825;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'h9897c4ae0a4bbfd33d0aed5ea90daec24a0cebba07436087df4f8e58c33706a3168d4120ad32780908f4ebbc6dfaa492ca47b94b4bd575d888ac08a63f365e7f7ad0b0fe1ec419b3681f93eff6d76bbe79ac8743ee57809fc75589ab1dd7b65a5b30c898376d0d5b77851ad70b8806c65ecd157d6d85131e188fa73db7e762c6bf3b322b1124173c9b836dc6ae6fc32ac2eb61f4e5e2b0c1925bb9673e00a3c71d9f07bf6f76e11a65893e02a1605560553a81e169178a9e6c230e6925a2ff1726864f7c07d927b2a45b28448c31f1e2568e91ce8a98b180f47eacc114ca0b856a94cb41e1b5bf5425c08aa89c2c15ac75289f0abc4bbdbc0cd632ee011eb4b240ea2c5c59bb42879e580100c2a83195d0e555e384c439708e496569038873788a9c0f61fd2102f2e167561f3e78e5499df40dbfc2d92f66844fde2dd1bec726966c1da6505623651e2a58b3f3eb3734d23b84fcbaf0a5d12678864e7d2fbc02cbceec3e8010a8c0c1f631805a443e3a0e31b348992d7134a01b0eafbaa544aea20553cdeac2b2ae44be2155efa8727f6c95c03ae5446419d97504c167caf44fedb6b12fbb8e2e21e0543d7aeba85df0a03fce7492872078b679a0dd451a399b550943b62708ac2eed4c45ee1d8bb5fec89d133236fd476e796e77501700f9f2b30a81d30366ec14c71c1b19d4042f9b3e741834f4b9795737fef73a5f47a654c32ce3e0e568fdadd4b0a2ccb25e033314525fbab2e3649737abcacc546dc541eb42a7e2e335a12ac1177b7e9cb1d5f37eecc0569c886c2cb03ac4ffe0cc31c0eb94c6aef9b599f284895112269cc8ad3fef6d637b9bf0375fa5b471cb1fea4ef0c4ad1089c9907bc564169314ad5c4e27c31af89e6518f5a6fe5b62c588c88e646c54829b35a560;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'h431215cde61a338999cefbfc3beadccc9f60e6259bf8cda3ad05429a2bc6aea331b6bbb205d8ab97a11c040ba7e5bd81633d0b75949d84fc29939681e737a80f9a1287362b16da9e85ac9dc5e844a35e1764eb70b0a1a8aeed84481760eeb0c13ce3aa16f93eb1cbf0662c924176379563bf173c1848678a11ca4af9ddf988b0db0fb455cb1b8656d22cf975aa64dda47d0825449a6791d386f4870e3a7769ff4f6268262a24629ba365bea958b943b9fe8ccde119eb48b422aa6352bec9afe3dbbecb85eb123ef56d6da60176da21e70dd7a97b43d6492c35af63ea6ce6efe8350d90a71eed616733b9417b3bdeea8b0b6af751c14634bd67c1bd0d213e637ecb6483ce2f17cd471349f771702da92a11f2f36bbd9e474ddb9102aecb0d13c61a05067018bc77dd19c161d71954394be69eb62ca114509536081f18728fb3a082d70ba8678613ab915009fb05e88f71c2ccec6d36180fbc0973e14f29993e0970367cc20b3213cba1828bd282d44fbd5c132238fbb6996d1b87f369971d3f71d8bf66451914031fb878cea1b54fbe0f626a2f7586b89a236c3c89e52cdc85e90ee984acba34498c93a0f810df03c3fdb6f4ec1e1621f621930ce1d4a399ddf0da9003f4f1f8030bd74c1ed1dcf34aadc5a669be77d901b952b206cf2891313e3e784ff252f935f6c05a80afeb6e7fe4b1a7c31444c371510cc8349d5fb73209603483e34289d5fcadb58763ed2f6a542f2fd6a432e9aa2b8f60170eee58f44dc013ec4acb12fa11b3b565a5b9fc76fe372d393d399cdb822d2827c194cf3d52038d7b6ef02a7ec3e77beb7d8f13055c2d7c870a328157b0c3c0196546a81ad6bbd209d2381601d10650538cb2420334b6448c807b8589e734b052813c610ca0248bd3c4a04d0a8f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'he4402214f1c2d3169506d4fb876bd481c0b70e67729b98231ffc05038d85b32a3f19b24602b429667b6937985bcbbfe3b8c615a2002a58df71539b8234439472ad8660f9b9041d46980a2b7d1c3c7040440eaeb8c24de75b9785da3fd3a0c6314b6b8b728bf5360c668ad89cb94fc9cdc6d4f53eb3a2585b33b27be85899357031bb7844ccff1961f834787719bac9c08c7611c50313b6c6eae84a9d4429f4b14da13fceb9c9737f9228d9a68441a1dce6d0f70517f94b775bab806be8a20a40581378763e8ea18a4e139a2224f507ec1c8042fd7d9f3739b3c79f56eda94666e9557745cba6f3792cc6e7b02145e2b8a1c967972fbe1b1fd1ee17659483bab53bcc32bddab68f50988c2f44f3de3c00460f1b41f97923c94ef4977efe061d8058ca6a160607d851b408f3f2490ee805e6bc54fdae93a8c4556456c5052b0acb2b967deb96ea1f9d3d54d31e4499803cab791346447dae4f8a6f427b3a981af81677d8a79d23a627f50493f994ce04036ef895b99ea6c28d5936ef7e469dd216cbe7c8fe3c42d163c002c0dc04545cc040ef023183c4c1f949f22dc209e77325562904ea9cca11db1b12394fe5e206edbe27210722f4b93d33cfee2b9726b97c1ccbd58766d6a8b766a9bc782747ac39bb1f6b8af7d52fb341947f50ed14d4160a1718ffd6ada03a55eaeb69cf7419206ea3d52f8799a42f3dc72a0f5e9c4307e1eb813fb79ae3f9b945470b7fa43185a637edb27e226ebf864882a2bcb5d1389535ad0ed518cd73d9c735e9df873407ca8aed5750335f645ddcf4f152f1924354d6c492a7e976ab34943b906173f4f6a1491e1e96ad96f810d13920c068cfbb4c029a075d040eb32a685a37b3a05fc5ea51b8f3366fe992439c492a77fb549f3322544806d088cc;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'h4d1be56d5cbc44de973a124d69f2a6229bf023eaea8629aa437c64b2dd453f3c0b9cb9d8d23a07859111eb71af9c817403100a0396826304730b246e8ca69425b0944611c264f0afbe95e41fbad896df4930245aeedc10c328bf62f0d042e48a14450800964201ba667781146ed9a1a6fab09e86f5a8c162eaaf39410e98ef76fbeff7faafb83a0b09e438eaac4a3c576f9b1eb3f62b83044c994be6c68e244fcb60773b63c5cdfb065bab1e5740d3267d56322f03c346fc47dd87822067321a6504db25a7f9ebec0188beea7329b2e88bb7b25e1be5df93fa37ce311b092023bd630a2f06887438ee7cce7384ce084e99506bca97e2ff1c0d32bed0e0a4cdc0f6a2f77ca8456d363082bba17c5d76a63f3215aa424f4e85bafda2c46bbeee28f7802bc1df7aa07d1e0199976a45fc6a2ec75850fe3d0453058a085d87b0a96f94b261a048cb494c3d28b483c5c75222c88172ff0d61eb56b71de336818a678d98c17ce8319beeeb952ae5b7beb6d0fdd076d99a51972c50d1acb957252192bca7fce08e907af022c032d4eea09f829256b1715e82cb9cb8978a8970288781e978a097f31a0b20238146d5e39ea671948f8b511c2481c4d755445915f29f5fb3a37388cd17da3cfc45bdee135b324c8b92140b2dbae5b18b6753c592cb5478a716236d5b3c2a39091b9bc8cdcdfd4e85e8adcaeb217d56a476bc726e1eb00b4280a87d6cfb752b39806d5e6bdab8aa1501cc697a2ce06dcd98bc6176226bca5b454950ccc9c07d3d9787d1a97aa42e748311cd029db58c98377c44b6ed2bf1d51c390ba3ba5c2f2c479b5b097a76a35541247cd286d2f51c73696d60de3342c3aa97d8df746e5890d77a9ce618409026554f0e9e63366b5677e715244f26c096e7fda6cb08ab1190;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'h647e0a88d974ad82b4184b64886a3468f8870d605161f3a50e8e6ca2dcf7599be3ec66070fc1617d4323ed7b37af6724898c403743480cbd3f285a0c11527ad7b69fec19b345ffd67de899b917f2dac84006f62c661478e8e0f9134d2ce44052ea7a6681a7050e55beec907474a37540cb9e0f7790b4509a0eb6a0a27bf1441c47a556f549749c8debfe1d1fe154ae9ee09c7179e45d3bddd92d0bb5a2716775926cc8c1aa8e550b307b15cf48d2f2626848fcdd91e4a8425800f74e54450d7a63b327d3b28cd3fd5c9b73bef1bfec477ad85c324755ff7ad712aaf34fe47494b641d30cb187adae88beda9daab52dd564ac2dc02678e5f00504ee2fbefe1cec6cbe483e79fa26f64b0cb732a58da40b8c84f4355143cd761acc5b652fdb2be88a709264abb60eb8ca4161dc87f1da2176c0f0421efdd2bae1890e5f39f969b2806dbf9e9b2150ddc60c2f8a70cbe4a0b5746b09106e323bcba992d190ca277dad2f34051db1bc55678e51eab6ed3acb5416510bab9356d817acd9c1ef3395e0eb686d1c7556bb0eaa2d8e3bbb2ac79406df34e2c8a14e12a40ba95df519ec0f94e1a0c0aacb20f3244796b6c1654d84098ec831ccf0bfc1a605dd60058cf2546a4f89ddc3a50fa2845611e37f4012331f4d64e562cb035308d2cd25b7fc9231b3007962802ee0c857d56e298bfc18ed96e62d2f7f9572e6d8f3ee8b5c7c93bf8c6e94917757c82cf107eb745be726c5b59924445ede6959244972bffd8cb7b56828b09fafff7a1ca453453ad52fab48070ec69f187c69e8712c3d6c003442551bd82d682412122f5c9fee32688446a859f2b40098cf3615059de42cf0dddbb316f5f3aef544f11d43e0c8bc89e90591fc38a845ec1b4f62606b1a3e66ff91e13b46f2489579a61c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'ha47169d450837760c33735aea3048b96cd75bdbe2f61e7cf0e9f0e3b66acfc67aa0f05002d4b882471b3b1172b1893ff1637bf412847b1074184964dbabf4898d5e3d379739c5760c51516d48676d5ca7a091a6d1c91c1de66f76abdafeb2b3ad2ecceeb992873c3c8219c6d4b0e48d5c214dda1615703fc7e741927e564aec2f81d33a289c39a0dc4227df7b49344c380ca679aef84302b7acc70ba5a6dcb7710796cf3c662045de925e168a2b22027201e0bd376c5b80e7d13df0a1aa9069f2936125e2e1fc4e7e62f954e566d349c86330aa9a212e3f021ac9fc37a0abbc6669f8cdd502fed9e2f225a258feba90fd5cc64a46268de75e9f6eee7c9fef9b55d1b750af6757a2be8294e3d84cc0cb7fc8b344cee4be0885d7cc9d760b3ef6d61e7a74eaf5968bcee6e44fa541801c78339b14d036b649ce302775513600c9b557cd2f0a000fa94d88a49afcd56fac2713629bc80a8590963e0d3e0b7eea15057ff29d2cdc20d19e5fea6531a108dd8126ba063555b86420ac8c4e62b19081b253a1448d034d85fc3e851fb66dbc847d77165651672372804b3259d853eeb454a8ec732a6c7c31a4a3f162f92178db587f2bcb617c694242a249ad71f5aaa3b6a0ccee22090cea022781d6268be8a5407e0a9059c020cbb7705c3f59f29f4ecd31be75414877df655ec2d1859752257c60ff9df9e62981d49b93afb6c505ef4314be935b0cce29c7a1d27fe679ecab98804123ee903c77e199a971e9b14daedf3c648c07672e36a8156f75662b4116a62f60dfef6c18f1851e107762789803ee5e60f60c5f2060bad8f540e5f4e5a1809c1987a8a4348a4c55ce7b2a4acec50791e632038f5d0c873367619e2ea6f4e029d74c6a87f79b9dcab4e4e6c5526a4dbe0a4a5cb6e0576;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'h5380a832e275b2b9d39dea2e8b38daf08c403ff769fff47bb25ed94a8f15c3dde009599046c79f3d2681088eb1513f36603945ee49c2aecbc699946403ce893436aa0563540728ff970ef7bce5c263485056b5c4fd3830a7c11d69649c9c04e8728438c3a4ea6aebef6d697af8406c413347413dbe1e25d18f35fdb6e145113dc754ee23f178eca560d202c29f1ea1f6dd7e2c7c4434e48ee0f579c3f5e69023683dbe70331cc2460b5fe4c99f7d00c590a986e150d3ddf754ef0d2655793e5b024af66920ad41b099ecaf38910b8809804700d0156ff066212df5fc251cd446854f8bbc8ffe21e016c30a484840c314dc4abf774fa54ae2198288d4b81f0017713e77c4834a4a1b064b890e7a7f2ebea70ee648a14bb7c1a77fef73688f3ea32bc5ce22af9862fea64d4104bfcd0713ab115e3be9c77a860147ec39beffe5660b89d4efeabf0d9a157684a713306b5c8c32f3f0f3f359cfa1566f9768358faf0448a3c9d8c3ea70a4712c7f6984b6eb2a361385d333ffebd273a4f53edf3cbe9a93ff04f8112723aa31721eb8bad482140d714b2e34c94613cdb909d2b5f8e373e07670ab56310d7cc0c6392303031249dccbb24a9cf806f7ba261fe7e1cd3718d4ef57c8ccb21c6da6d4974aac165e6f17902ac4bd44724b14522614e57b39460a157aa3537d8557e533d10b30201de4101bb9c1103fe0eaf14cc120ce05099d66686ee8bda7371bbc90dba886c9a63d57dd455660155dfc25bcd2ba430e2ba08a64e977e5599b3c5d1418e8471ab8e809a111d95fb65f867cdb5dfbaaa63ab45074558059b8ecc67da88c4073548518c308d0c8025650c577d4e508953a7519890d37574e5ad62fa79d073c9e0e6fb0c136d21b8e9e71d91c8d8ca7d12c64a25aa69650b1bd0c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'h90111b669923810087918616dabe8ff525638750b74d109c780e8fecdf9f9e1af92e86d2e3cfc9fa892279a727476de81244bdffaac89b2fba094b696beff8f6068c356dec2c8a9777f4256e91e4d4309b5cd5a64ec69168296d26f57a8b5460b9359813e7e5d0669e3e735cb31674b95d5eba7e57abc971e824356235c9e2047be42b111b3515ef078cc638eecd8020d54122c2f3652798417693125629f5497a850578024e4eae5bb3d7d7637b0ec90bdc63a1cf2f5296bf005523f7d0a8d7ad97a4f5fb6388f040e5a5d5022b5da6a375b85f3c1cf3f75f9443afcb9de0c968bfe523c7ea4d123a284cc9a38716d9d31e10f39adabaea5074b1f5aad39267e4cb1b692636e2a460345d23f32b84210e442faeaf83f92f24c5d3b67bf4353451a05dbe9e4acee732fb887482db3a9e3ccb50059c8be5c2c21e5ee80ed8c37566af733b9ec2a6f286f019c15eb2063db4c61b114712b3166873fa75b531bb0a9388efaa9e5726fe04a3631174313564b5fc3d5ba264359cff12fe666943755e7b257830160da1d4d7700c19b8f9e61e244288e8f21adc41a69e4401080a1b987a928d8d067c48e5e1e363be46b76acdfa9b950f2d90c4e3a10554da99d4ae2aa892be19a4feef787c8e5f66898c030506c849ced9d5a5d5a7f073452e73255e0d9a560aa8d2a9129ddca62b5d77016ada0aa74b6b0dc88dcfc08f8a20c01d6c325dede44a09d58606f3cb4082d48f65ed3741d0751913dab632a77bf0cef34ef6210bcbec53666fc420f3c79e8f602f6f3bac03acf75ba7b57dcb3c1ebdd4eee5d55ad9da87483bead32ddac3cecceaaf952ccb6d81e4ccfa00f235cff37e7f41dde57fc0f86ab4a2cddb9c4e6114263a74317b8e78416c58362e74fb0b7b8107aa9aef3f5b0e1;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'hda4d45bca3cc71d1ba49c1f4b5365455ad62c4588575d3e9567fd3ea9e5b88dcb5e9ecd1316aead812c297e1050e3b9b16430076d080ca2934d29ebdaf8056478d362e48ab8d88146358d2f8757b6fb21d3de9d854e69d7b19ea763969d700718631d263960901eaa7cddd371608856ec25509c9e545ba5edb379ff2f03f1a106c36745bc21e3689d1bb0a4b9f5580de6f60b9d08b7c5a7c710901d1d4f4f87f4b730be447a39eeab5088cf809b4392c772eff7f51a6c52ce7ef68682e727a431db051d0fcfec082b93314d0f73778e3660015ebd3c73e73467258ec732cb318ca3838bc42cb023ed9fbe9e22190b6ceadd0d6c09fe8d0507a953d066f5e33bd2c34f409d6c835a04406971454ece80a467f439c5e71691cd085a162357dcee0db1ddd6fc3716e3e3c91a98d119e10044905a6986802c3f0f61c99218c937bfcc190a027f27f440b4bd1e47ac6e91cbbc99dec9f96d56fc9a0ee8234cd630d478801ec1b34bd58d16119baab8840d63f933827066a28cf28ca656922c12a48e53179ad0212d89c4a8ab8593a5e56b4769080148b3b930ba4d1955cfe508e3768dc6611c2428cf5be9fd0d593d94e47d7dffcc1dfceed44c006a375a4a7052920a1d83ba32021ab1b78fa16c622d3f8ef7629c5b3da5710287d9f7243d21828c60da1b93abb895b0e90e0b8d740c7daecf13a5659b55d9eb377f4cd134327b853d5e3345fa5bf70bae1cf184fe5ada601c7e5e687b9e25f605d6174a1aed5ffa9b96d22fa0348f42e405749e286afa41da7b6e47acdb43d2c2177e61502c29ae5f2d400268858cb4e4ac99860946fb238113117a45a852a28260afc3cab2f1ad9d45178751828f7b8ef08d21b3309971de0eb20be9cc7b5cc87afb374c25d0acb46c0483ba8fcb73;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'h4478ae42d98a837cc4ae71982e8f899b4e2798e4747dca78290e37049e7a95ffe6d2ba2cbd1449e59031f2caef60238be1059166bc7dbd1dc5a60116b5dcf91ddb7e5d01ef2d2c8e123f18d5eb7e182dbc7590be4edeb13de425574b3b91ed81b20fbda68942ff3d254cb174e2db30f3fb6dacea62c0acd8f8ea47bb4aeed8874f5f2148302b76bcd414865608c5bc499babdd6fc1e80daa213b714f05b6b006ce29a14f8ed5b5af0000dda3b8b450d39a8d459820e1dfe97d3ae68bc4759e978303db7f06b79dc74bf08f259b319d657b301350c1e79ae074c533a615ecd210a733c16ac18b899c0aacf488cd379952a9673f0a465792844d7ab449892311bfc33e3d4182e59dd81b289d1356518c3127f1cfc49d776bd28e9c4f2996730f5d46374bb7cbd894baa2d13961437e539a061e5a3e781c0d96f591e9f8d76ba5193f7fa93669066c501082d9e3dea13378c337b9e26763cbe801137e31265f50cdbe296c6d3de592cae5271476b7663ccbf2ecbafcb446c7256a3a8f37b7f050f02ab3cc3ad112377cc4238a8097ff307b0e2e2d92697b1439da95df9283ac1768a2afe2faecf8ac96d6840249f1a17ab39ac2ecbbd01cf2fffacf639cd8bd9413db5f5e9fd8cb8fa60ead13a9dcbd767af65037d7a9996041d9f752810c980943f2016310edc0524dc239405ad0a31f819543d49252914e2710bc64c454484398a870b63d4db26f6d3a19d162bdbc416fe3e3bca51f53492a9068a65bb9cffc2edb7913ed45b4a48912e16c3f52931556f8b45e7e30bf3aca787a2dfef70eb91133107cd9dc4a864b0e94a8e2b2be289acbd279da65161c7eb82ce10564a68243aaba71465c49422795441c3b41324a53484c02de94b3425bc59dcb9073e67b58deb7c0c71097b9fb;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'hbf079988bc2a4b11ff8f651484c5e7dfdbb25abe767badfe193a368602fb63a71ff5c75582edb70b6bf2947ebcd22650ed726716b40c55ff3f055ea5c99c1718c8b5b2905eafc619e972d0652100aff44b20a01f7e6457a7a7bf26fad1217c40550ddb37eab8d371a27a6b8bc2eaa96734b207181b5e642ed8637b9267ab07f0b45ccf73eab1827be1c04ec9f36980272f9c0b0ff4a30d5c2206de40d0d5994db735755e4c2d601a8a94d57109cd464e92d1a2ad4eae836007d38d214948b498c02b278bd88202da89dfd8388542bb93b55b89ca80953527c3bcbefc01271334dc9132dbdc14220732256f87f375052915578473c5508078c0defa6f211291c1915044d336ebebaa0a9b0a6022715b485f0b6d6df6ad9e22dabd26d66b65d99f509a8e8c645a8666e93a9a5c8847832bf783323c8fa14f106f9b552fa53ab38d38a8c5d14eb72b47fbb01522990f2368bce4f091c2abf59267b4ee9e217704fe3e0c15fd70b7b0b46901de5c6116bba2feb9513b7701fd88ee264bac1861b9dc8cd9796dad7596c14afaf5d37bbd97ffba3c4507529a0e4dea8c0c08b0fd377245e7e23405965f754e9f0dfab52b50df26967ceb50872ee80237dc7d483777515fac18ec075e104e941340b43594d9b1ed9de5368bc47b6609b1b86e1f11d04b14de02212ec239dd9e6d02362c01fe99821afc23c97eae4e9b697dac30a68923c2577d97fcd9de0fcf6be9227fbc8201d0db56e9705ff1cfde785f37d1ebf2f21c40b5aed9dce8f32b4cbd977e88990e0a0af8042a1ed8aff12f4be3124dc98e47b6729aa79f1774a9ffe95b1245b41e4f741f7f03063f8b59afeebc6431b865c093d6388ffc694cbf53c737cb9997fe964656f6fc42aa1e1605b6339b0383307b7cac4e840af8b0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'h416656016d08f4fb3b0f99a9ac858fdbb0e960d32174e739a93e821a923cbff27f321b14ccf02e97ee9c6011e908557259dc40bd69f456bc04d79ae352590af8b9710383a1d1c41770679a3c51383828719391c26036caab40bc10d1b5d86882040cc2e0f1b43866e49e58be234af8947384951f31671eb9d869f595cfd474c50736ffac7da1d1e67cf5dbb46317935d7ff2fc8bb24d7a6c6bd4c3982cc6f927570aad70fdebffb5ac1f5b183dc504128a998f2650c667daf20d03827d4187166a71dba9a7288824cddfd8ae289e3cc0795ed418d563f55d776c66041e4d672665081ab4f54e431cf1fb91a3c0061cff7c4df86a1e9797024cb6957342e0d5e5aa02674a1ddd3ee2f16bd3f27621833a314e4178943bf999e57dcd1e755c8379c6e205a66d4d0d9229d65b57182c07e791d9a1dd517db683f6136e80fdfeec23f7583aaa793f87cc10dfdf7b22eb9ca8ab549e0b261cb1d3e84813967b078876d3c089afb4fc8ef3eeec3b16268504f8b477e7251cf7fb8cf057b6baab75f50ff21620807dad304e50670b0dbf6d6806a5f36d1e03682dd04dd5e5345899ec1f320461e323f831aff3f98cbf29e71f61238e999909f41f6c0a0c5078d6d395dfdcecc8440401fc2a8d2c795db06d16b81ea8f63915b38de8c29c72aa8ff285713210458e88162a8c911d93c9788ac5511c1b90d322e65abfc6c7af9c4ea3df196755296d6f1a3db9fcadac18c423e1f67756d116ac1b812afa4937fa83aeb318b1991f61bbcb0ca45c7176268f1b61eb9c179763489da9ac3a7fdd158e432b9e62c72236eb0f27461f16b6b9f44a4b3fdf8bb5e2c57297f18532cea69f3a21edf3dca7a6983ea87661d063d82c9f8eeb0a05e9fb3723d6e40b3feb39c494035f8fdb2a521a4aba22;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'hf52a439780030162e3d48915d2d57becc5d9667d4afb10cd699bb2fc0acd859989461e58f491db6978e08bba7f3615ec20282379afc9b58b55199669056993e5cfa24e6d6864988b79565f737116d27ac861e9de1503edf06deebc76a02e6edaaff6fc807621f22452ecfc6b59d4367d818c80518768e4e9199982df9a8ae1788241df01a0638ece08a1cc606257755c72e0df0e6be4a61fa618cc067d47205576f7fb5e1980df1dbc82c6b70ea6c612f33e004c7cad0c44745c5b15ed6ae940e879d33a34606a5a04e6e8105defaa7eb48d3dd38f3ba55c324835bf0c9e02b4130f6df7039cecfd9543e408bc65ebf062a3ae2c9e9bcf3f71cf94721117b884e42ae11928ebb63736bae276b8f7b39daf29d37292bf92426a5f3e8f8179d4b474f5cb73040bbbaf642103a39c8619b0a324cd1a06f1eba958e1a3e86db495162533fed1619a32352da5fb5aa98e70801f9f978afbde84b0d87cd2c5eb1ba4ec1bceda2859daa51cb36d2871452816b0bfc9c5cf242817cab510c6879f3627cfc29b0b63b0e25807e90b7d88cd4362cf6393727db55dcee9a0df1ba2333b48c4ab4a9554351811c6991ef0b2fa682045511204078f3466067a90bb9580d09d96a60f0663c6b7072c9dc3094f6a7fb53ad928220403027ed6ed84951eeedf4d4ef4d676d3e6b34bb1e74c043dc495f45a445f6a9a4d95617eae47964bef070ffb5f21eeea12e8f479982d0a81161362be411785ca350418a0f27b94d29e1f724d05e1e02a9cc86ed3745b6535f33996621f981b37c22ae4b1c0a057c80c8f26227d026c08eae8e513fcce2ba6962f6bc0687f8783d5f9156f0ce6b949e0f0aa50fd0ff79b8f05d07f0ae01ac52d26200a0e0a76088a6e3c5fb95d1ce9ce42421b24c47bdf66f2688c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'h27b5e36e70c20b0c941758466fb282b259640cb8d4972c44dea66500aafffbdb165ce25231ef98295473034a624d90021615c735c99758e139beca97d02dd669608f93bb23ced166491f2cd83b858731504ae926e6a5eca5e3efa747feb0bffcf17e5568430a9c87107d2318cc71e39d0d07331ca9c229579a31b31d4cd9db831f41bb062ab0541f93d7540843713b984c8baa9091218c1993ab52636f3b0906100ca906a6c0fe92aa12a12ed5181a841bdef830cd735bb0771c6ad84076ec941f0adb9fcce8bf4f72a99bb2188924501134928fdc3ec519c87abf0dd79e87b2eabafe690d7540ed08fae66ad3ae4616fd937475ec1003bd3dd97926862150fd7bf777132c01bc4dcd0489d491a5aa86154163eb55362c63c3c2992eb07130b656b7e905531bbeb08b768f4012995dee88a349346caed9da41ccfbb60904234e19937867e49b65e172f08b695a6a582f0b6096e41b014447da56c9b19c1b2afa4f2107dea9e1aded4362057b89cfa2bb35f60b32a1f36c5c7e738d19fbb8a26c3a77181bacd7fcacc282d7c1d386fe2a0727032b9c6308c9120cf56d014faeae1450d4d6276d6f2458b96e13e6de57279b475c1b53e59eebb0a84b6e86fbd2479440124949cbd590dc798424b49bfbf13bb713a91a5b6dbbabd8316e460461320f9bae2fa259a809858c6c18c499c4ddb52e1efd1dd82341fae31b4370fcabb1a3ee748a18b5ce8997e81156799bfb91f550da15419837b4da8ff4cfea260ab314be004ac7d515c78d02a6a699b0b8cc5abe07f506b3a109d50c438eab3ea085cb7b51f44e34e48062eaa50082b2a8df703056e2ad5d98f1fce5f33e1165b641334f39c2a8706e8169390d127040f6b594a6651e123f700aeb9e22be04a0b01d906e4682f93278b6;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'ha810dd8fc6ac40fabb84a62dc0ccc9bfdc43dbfd3ea0ca3561f2eeb614efb179e90bc675d8fc0ea5e1335b6544f6a018624b502683771c24d64bdd513888c4402be0efe9fb90b843173fbf83e98116bdf96a6585d03cab4d7863471eaec2595c0b49d50e08825fd0b5508c058113d843c27648e993d5da666a6b92cb5d9cc025503d799964649b9e75709919d17726ed13257005b66ca6b778c6afd75183e351c42d23c9f4f9a4f8e20f5550928435ebbe066f9bc82c3ab9fffc3342df5f2686ed24d7e4855a025bf62a4b401af3090824bbdbb36b42c1512b4effb7bfbaaa2683ca7d8097d0837bfc52227ff8f8606ac9041adef70eea1e50f996a54b3d994bb48e4631e7c3dcd707b604c3d05e5bc260ff072883c4466db90684fe7e7c60743c758c14134a6189d2bdae3077bc513638606ddae76b36c4376701723c2c5f81476a20ed478960c9d3d86dee2e929876fe3428be790daae7fd9cfc6a9911343ef18d701b91486069a01665e8f92e082f711eb511a57ab9a5977a6dde951c222dd779b5b17a0bccb3542b1d1a9f443081fbdbd9317502ea80691effc88466009cfdb209a284f52ef205a5afaed26dbbac37ba1e4edb4d96d777a9edf525db524b1e1a8de9a6c0c29c6cd9222097320ad1cf73474ccf65ec33e8fc4e7426f1b989abaf4afb330901916e6f8415959c687d4e1961547d42fa1658919e62b4b951c9581dfa5ea37fc998f26e74faa4f9a0ccc929eb7fe70250775a17f3a9c48bd877d7ed4eeb133d58121c04648e21aba50ca347ecb4d88433fc7fd69f52606a14215c65cd8e8dc0f6f0f09b6c058b86bc4bbdd76631745eee5b1cf5b52d856a145bf0f4349b43f3a4748611c35f8a2491e0eb4dff897e6b1ad25664ab9e89501ba0808f39a451f8d962;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'h54cd756423169ebf6a5a209ac11248e85817188e7ab47a97ddb682a6660d08354e05864868ffddaaa9a3dd51af686fb05ed812428d22a24ff899f253dcc070160df04c82b6c48483bafdb9442cd3a18f8a611bb2933dad53bc482f5ae39520ed6428663416cb3bf295cca4b7adde4d5309ce3560bf6efa7d47bab443eb2cecc82840fedc4fbb5907409006a3e05c8500c600aac4e7830f0a3b1e71623e963c3a4844e2930987752d7f34de8bde0f5ae88d95b5cad63f7eea638c08641b0532f1678cc07580030f61d7122ffd294529ff05a3d897dae5c6f32840034870d6539be3782013b2ffaf7a59f5bda488361a628d34aedff7283d8e02e76956590e8cbbac70ed4850ffef07e13d669dbec46b8b95507dd568fbfa039b1d1139ba23e0051662cd68a235bd60803df680a2df0a377c14162a499008d576d203c20216a60bfd92042b54050a4ef8d4e3fbd33f79462fcafff6d009673b7da85cc915ab22e81e26301fc84afd28e467894abd18c04d8ce182ff3c0b208b83718e752f4cef1f97987ec60b774bf87a80cc5ca17f329e3510a103f6d759d0b912af99d571aedbc6b1108e68ef14d9fad4d4df62d00db6ea841d0c902abb5e57b546e16c75716e5d3d2eb1e6041ba634b408278fead7aca4b5e8bcdef8832106ac40de883f2c3201589bc05a31f17efe54bc936ac7fd807d3e69275268cb6f44fd58801a04b2e1d5ed549b81acbcd2ae1ccdc2e9ff87d0c5e804e343a4182d17a1ea7ad66cc70f82a4734ce491e8114975115e74df52ac05be6c863eed993e23be9eafba864dc75b8e0bcdd1ad679bd5676ef295d378a7fa67a3985c11bf767f0d08dc8adfd8923883c70642d8bfb90d1e398b72be2080c330db92a71690ec88ffce4e82593d42039f880b4f1d0a03;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'h9f4616f98675140c42a88310ae9f0d068af8717f8b47c4f0b620175663a4c2c1dc7228693e2a662f5ccc06f3ce6e5c6aa8d56d8fb94b702416ef46fd14cd8ed4ea64f00498bff315de9fd22e7989529bfac44535788097d0527707fa3769ccf5ba50d1cf4b81566f9ffe7584d62801bdb546ffd7da88a97dfc9b52285ffdd4ff620aee0439377a654bd398926df618e0cd7d6c25e5630955cf10dcf37f9abd8755ecc75fe5216f62ebd6aa766f3b51c0585a767670a43be2d12d00947cb227cc3765ec81ce3695b2b5f417b2881661570d211ad9d285392b192ed9d25c61a5749a0225b3b0782953ea71adf7dfe2772b1c8ed87b825973a7aac304712b175e08b7bc7c8ad16e8e1aff6121ba6f5ed70ec8362005ba0bc91476c450a6a91c63462f3d10859e2437c07277444ce236d60d22ddbb089d4a07dda4c0401324ee87b625f8637c05875e70dc8bd43fbc5120e4f6164ec36e69d85b21d8ad278a1717921995713a54243d899ee4562c69d23104f55fd03df6b4da2d7232a27b76d51a22465b35ea8be558e30d4ee41b7c3fda372d43f50770cf02948a7dd7a900f4a926d50cb53ee1ce8030c7047eb8da944fa2a76597e7b4b904e54078681ce04e79a522c5d49258863a737489be8eb9f3e3ad8b5d477f74fb187320fb7562137f0e3195a61d340911694a4dfab12405912d66f258644200793405b2e5c6a8ce55cb71b089612cc4d7fb27decfd2a50cfc52cbe5ddad7a3e7cb0c5a8bb7a16d915a2cd83dfba62959d6a3e3e28a824f17081675514c430efe6e6f1c9c862c58e51779334b35f18015762336cc7e4bc38a2d93c57649878b869c9a0cda6f2f7a2503f0eeff481280f636d0a5fe478ff17902aee9415297ed40ac860b029fe6b3f876fd5f446e5cc91c52e10;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'h9722e7e4a155ce5e93024a1015a49923dddcc43ef59a39fdeb3ecc25c9fc6435b34a6cb870b6645782ecea341d5be967f99468cfaa5df031d5d627dfb517be3842b441a970d4423f4da6882ed9d1da8ae122676858ede22d88a0721ff4263ccae5d3511a44a0170b06b08d4f766fcb09c68c6476956cdce53e1276da469dc122458644958c0d488b34984e84baa9aa8d38c85a1f7252dc750fb8b4c1be7bd590f36db8c80c842d6f2c3cfc132f798c46803795e63eca99a23658c49cd155696cdb295bef5c3135a65f07a7f9c5d84373d474c699285b7de1dc1bcb243d257f8ffca146f3180209c410b3eebc46cbc5a9d67e5f71d29a4a7ebada96828723a55e7767fb757b8bb14af9e7655a645f1eb087783c9e79a6fa3353f29dca8aa7865c1fd91bd207e30479fa9e26f906a15fc5e78ba88d75e567d67a29d90780cdbea206a7032cc33d52a84c173b15ff01d5fe9861e7f8e81a9ae46f1acddacbaf708a96375e34282299a70f7f0f5ddaa1d7551dbe64fd7b9634ab396848589bc1b4f0731bba51d9f6191330bcaca6822ea974cfe8618a44018459d27c4fc9b32178e192e0e11d93e8b5dec85931da397d6081ca785ee2862bef8e2736c560e5fb97edca42cdbbaaded35225571e8d699aed17fbe4b21dde5239bbc1f5019b540a538185129fbe1c4ea01d5df7e579e97cc0f3a404f8cf85cb311b17e168661edac04f85eee46b4294fdbc67d9c533ba778344d32f36f78169b6e89d0fd9c7cd0114e3ec93a04c8d567189cbbacd4bd37fe30c0388908c05225f84eebb18995d965f551ddf2f0ffd3905dd1a08151d8efa7a950d5869d04b4456fa1deb604e84896764a2410f59efdf3c6c3240b84c382336cbcbc2455f92a776b9401f2d1fcdac2c2d06a64fb50643c2e7;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'hb4e9a234f02527f6b8174c76c014edeb2c5bba3b825a09f1406dc48a5ba32eec7858bbd95ebc0c2710ea83774e35b027c8f68acdf847471cc490f37397f9d3cf1d8507485ff426553c6069418a147da2bfe6a862efcee0b296debd952c1d3f951b2200cf994dbe9b6469c5ca62c4a57cba103238f3b22676507de433d76cfb5553b4ebe84dab500d1729d4ce5afebb1faf3649fda09f6d18837828a09a3ebea07939989162c7b6b0f0ae1fddeb4737932f2da055b51e8c6989765f117a9767d7c4ba7c748f6cc2b6f9420b9d1f0d21b71dfa6d2249ac06b5e7a2af92fb4843b2c6730378df9a0235cef1e96abb7e669314fc53d12e6bd5d8d19741f3acfd2d03bcc62f32abd43d9e8980937934cc7fc09ff72a4669ba6c1890938188bc06b73d667dd1ff34e133fcf4bfe5b7b242adb00e08445a02ad76a3b19850a9d90d6eb0f955ac9d92a1caac5b4a6eae17c991d1480d51a63e11ae8871f08e6f9a87845597b946558d321553efbc0145349ef0590372204d727cc665eb3c8c9a9040e0866e68a75939adfa13c6c4c22995c527aa9f6c531b35e3521a3996f1b54b504e0392ffa225a9c9b432b9e7bcb00011f5870464b859d95da34035a9b2204cbc38c38b8c16cffd3091bb1f0a9d391774b082cb7b5cb57a7215817d0db8ec23fa9808fa3a60ea7deff4a370073aec8437ceb8433b8988c6e1813de7e229874635a95ae43c5852de92f7fe2732cb676faf2541f65e4b610fef228603a8b18e790b7a3417d412f72aa545b626d63bc810d7d42f73c9747f73ba875043b78f3702e9457bc5c3c9e4b224a01a666c05428dd7374f71bc223a3cc28a97cf6545ff3f147a7988e7435733568460bd51b8e01e23d88aa4ff2107c5d6dcbef28bb12b0a43b6d264e80da5047a2a18;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'h7acac0f3733cd0b5e9f4cb996ac2742d2b26e4a9414e0c459e36d396703c9a554562f02a3423ce9d29d65ad12927c7a9306907cd998dc17792c899f7baef7c9de3a281f38ebc7f0895d54be47e5599f2d43819c54b75ea3993771190c2403f6c22af64d53938b33b05e7cc94db5a57d3f17f558abbc871d53bb5b379fedf0b35a48f0ef03e7e570e4ccf3bfb9aa20c9cc51bf5db5adaee6775af4a60080e26344376fdff4dcf426e68953a575a28c663a2410de3bf78dac70d021a178d63ba30c3e16ba100e627451e5ca594879664c9b1a6cb55fdabea539db4234520c18d3be7ec850d348dae381d9beeedfa3ef3743162e1d741ba2f61e7e19b93b8374a690ef5f3275172273b4a126969b14008a173bcd62058b7820ba0603ae9f1b7c5d34c0d75cf3c87bd47aae45be12e24543cdc227bf574a3f77396c611fddf707eba7e1492383b059f937a54e4091c41edef34322626ef880655a8402fd0375ccb1e477d9151bc38495e5c714570cae86a98bfcd9ced1b966f95b41118a468b139df8ed94505e2e11aba465847e7f30a123868d242ada55bd56d52c729e44a78816fd32335b5222adf1d8b7dcb038940720bf2a8687c9d154beb65d129de539995bcba3528e987c3cfb0c67b7afa56f2f150b79f51717357f765a492b8ac9035057e8fd67cf4582f789ca4df452cd732c49b1cc4cb58babbe1519c9db6b23ab35df8d816373ccbd63ce888e32aad09edd3e8df1baf604f9625c684bf1b5d298833fc4e02413e65dcc37db4622ac85ff50125517bb7dbbf31cb928a0c40c7411caefe2144fbcbf9bc300fabba35efa60fe49b6d775f13129a9bde9465364bbe3d6ac25f93fd55c38e42062e9dc20bcd3866eeeacbf2cea101eb5957b5155ec2601d9c39b9009ba4cec796;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'hef9743e4d43a5b87aad4a2f3036663f1cc012f8ec25e116088e4c44c559efc6ef567ed5f1fb69df949cbc5fe66e0bbe6a64d35fdf296ef82f883341cc4214ac8f9b067e0f8a55dd6ff0a4dbef45df5b75ac64870ee292f627de04446b4e6d5b4a4f5f6b9f1e142d18b254e7fcb0f796392d43bf583be21896cd3fd51a696093eb1fec120ac2700ef69794aa2fac286f67aeba8cf0fb9122943d5d8545c55e06328bf0543601f190c3687f5e7275b78583c093a63cf5e36fbdae129975fb9aad73c0517d37c57438c5fe7765f3a703ae2706430ae476557defa0d519336b0a727632d880394543428e9b9926386736cad3a932bcf894a6f1eb1b1683dba08e1cebfa4104a90b3296711cda19f1fdf317a48dd7616235cd83d7d21f6d441a3177878aaeb5815075d7ec734ac5ca2a31a756448ad026fae206741f31ea4243b63abcfa9d8326c870d83f1f5100e696ff49b4a130a60f62b9f9661d77dc579e28a7dbf120bb8c7c59aaac57ef39f0dfa07c40518fbb8c0332943d2e28bdfe0ce052f10e015979e7097992a84aa5b2cff8d2ae4f3edf920f8ed5f9dd2ed53244474da1d09b85366c6a91ef822b29be65d3ede98d4f6b5861026cbc07dce0f9eecda0a61274c92b6a0770fc9bb79e77db5714add3c4adee25a7a1aebc465c1c43cc51ce7834f1fcb722afe6e8afede7b51ee1bfc12bb8545291b11fdfccc85fc4e73abf3f5ea11450a011fa2cf8d9818d5911bfba42a9312d72b6a9fb45e96602b8adc13d9166f64533a54740fb667d3a6086959f46bf5c7f2d0164cbb3bde113a503c0be87165c008e775bdfaad920139ac67a799eb0aa91d7c771554e46f8227679e1c8e92e2a17672096235d599cd7307bed5fcea59172d2cdce51263c4be03864cd4d669db3e85f629;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'h985918077aebbc4a93f81f5ab9cadab0c9237217515cfd791af65a27cca91465e4af7734d0d44be302cd91215368b1c75c58b92a851e491f7f3a3b7c2604bd7edfddbbf523b79cd829c01a7db4438aca72aea295b45ff543e42ed4a72ad3b8948e4a5423aa939e174af80ab830045cb8d6d0ec7a9e755eaef0c86c7038b4a9933166bc8308a07381d2c7475c61bcc55a68fd49ba377ba197274cfe9c52deac2b382241615fb707254d404ba0553a3cbfa81fac012db46c20053ff115fb8a1e98637dbba9265b2ea099c3eae56ac83c4404e30d6021cd25a40b178fe9d6f13e221b06357b80efa685c44c9fb4beb71a7df3ce7ef1beb1ac57ffd69a5eedafe890fe2489418fd81a1aa87280c021e1cb15e978887a0b048c7214a7bebd132e493799d4d2778752f7ce45c2560d8da18dfb1e0c15b8c2f96f8f555f575f7aabc11a69f1f5ed584963f1a90f80533d6fcd911e670685f3435f39f01ed59792113bb1fc6e96c7521fb8f03f145bdfb01fc2d4af734ec79c6c8a4cb1e18d482a959f5cdf7a6cb1d1834e318afe18a3e4b3b0b5f67ddaa5b456933ffd5ca92fb87b715c779c7ad93370e67cdc945b7cb23e6f1742e3ebd2b0a2e8122f57254e75f5bd530b84a0f6306f2d92b99e64ced88e8b97b34aeb008154c25b3fb3baab158786d59a3a9cd9fa6d493655ad4ba75c40c9657a403d3b386fbc5bed4a0565f2e52707d0146fad06788ae5256ee715d2a3f9794351102f4694bfd442bd045657f8bf56d7586f29c6657c0ef2926f804da786493e722802f217e6eafc99f809c006044b2a09cf5dd9789a1037e2b315aeed3a10394d4e90d2e0d4a165f39e96d94a481f928bd07c6607461d7f419643999c25c74b7fd45c44b8641a81a1f1a5c0acb054bd8529fa6e7e3868;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'h7e9c054a8824811fdc95b818e87e21afac65b1542ce0008807a2dd0f87e1c3aef65fb97b347a2dc38f47d20f391f658b521babf9c5a8c3c34133002fe3dfacef58e2ec9873d6bcd72b714b51a4b46b32dc893c0c0da98b9c8fcb15e5de0787d690e95b3c7c3aa7c5a5fe767541ccc5c3d40a6e60674a61f57496a68718feae9dd6c8b887271a45459e855ef23985be7bb892094f8e9573e4938b8dd057be6693c064ff02ceaa16f0522327308583ec479105eb44e8ac38a83ba9dbe16cf21c39cbd2ab0ac6a7a267c08365b0bf62b1259d766803d2c99ef39a811146a2e56823135435c04852e95e410f46a1662d83d1a70844c5aef08f4c4743e9d254694ed2df84288c7ddf8143a7dd50fe65fd7b168cc7e11baf1f7b623e34c9bfd1fc0bb794d34cd76869104efe8686356006d4a398f51004992f5c60b8fc4ae2f6ab9e4d61aee6a66042681ae6c3d798c7bc49d5cc07adcbd52c4e7a888006ca1f32b956580efc6734ce341ef1d22f3a9e0eda927c8386db6b638fb252df200598e74ec78a5d9763eeeee19372cd792516b5765b63369fe6fea862d90b312dfb30fe1632e83e87fefa934bba15afd3fe1f1bb5c365742049aaf6f1611ac614c3f8703c5706753b40ed18aad2d767f892a957137ced81236e6bc3938fb112ba98d515e8efc869e8b78907721045e8a3ada4c5ff4e01cca008d5f6ba4a2be2e37bd4d9ea3b33b1c1f69e7cadb2ed99fcdf65aecce91d47a2f3612d21a5ac331d0a3ff0374d1c9a9c867c5aacea1b79cc54fa49ceb81c6a6a1309c4d80a503827ee39c3128f227e2f6b96a2d4264e4db497ed31bc903022744568783ea1b578d0eac057b3f9a2e501d3ae11f5ee68e0274002e1b034e24cb375d9799329d35726d8d5b53f1d690ae19e3a5f2b27;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'h135b718881e1b2098ce92b195b33b6e57883dd548ec81997553ab8c2ae6235f821fa5eea551957d1e39c2492c0f21a97dbc62917f650c2d43885a6cd854e03d32095d2457a3ee8cc955c7fdc8b11c08adf34ca67a64a38b1813b82c20ad608fa304d4af0c3d7c76e5cf7fd7f8657555115cea15102c6fbda2d3ed28504bfc84ac670ce896b258047b310744570b7b05f9ca4972c5d38c8f2ada39b7dd6c483f578b794128e980ca67c213cf804e558aca03b56a5d3722981b23f0cee7f8134ed3b809350233f1e8dc3f7049c76cb3b4d1ad71ae26ecd301d3a974ee0e522e961d65fcb2666bb81d11e03b0476e6e200cdf5c7cba4d99f0bc468288b7f39cd6157340d210e5a48e8f9a09d216d269eb7f412019ed07b667f767cf42d8fce9c2ba3b36089cebb44b92833d7dea6a2a060d226b692eb180af6987471963e2bdc75a91672d568a5d41353acc6a9c718ec160c3b27da7e590bdcf33da1f9dae3af6f1b69d3f6c2eb9210ccafc92fa2d5574853c4731ca4eec08e1081fa0b53d84b03696db469c6e5dbb7c4c97fde6253e41c9fe18fbb974211eddc9ac4828a6e24b91f32d7c954d795eb708190f78b97a7eb5603e50b6cb0c623e2cba05e2baa240715ad2440e3c7ddc3e908d1563ea4288e9b14c51eb212eb207210c9d8451976a58b167f823482a2b97baf55a3b6fc79e98b6cc5382d770006eaf2237c6fe7c13f7ff13b5dddfb950f6d1fd0be27fcb59e2883a8ebc82648329b39d39e43a3fa190ea2e270899b53fd17d3fa442f51ccc14b70c95e6cd0b76475d8fc2edc20a42e1b68608ded2cf5015e9e711ef8cee9614be946774f3c4ae67938edc9f8a9149b9782d68afd0f2b8bc7802d6cb2dc75fbf20f046ffa31982310ed130edcc5fd613a2a0aa775c37db6d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'h394fa6ec790542b90c7ce9391fe475c9c42b52e6d3c97f8f0115280aaf8f52ea64afdd8cfe7bfa4d2eaebe46c212933e8d0f8ac51ad5167c64f4bc3ac65d1d6b108c721d6657d2259eb4fe8569be0e40f0eba01461932045acaed99d6e06516ea90d8134c08a54c8c51587a122a95a7afd44ec0c99c944b2749307650064ad36e01fa8ec7a47f785593281b50fb49d864f2f09a730ca4b33b5ed749e30164622e2f0cb5c0a4fffcfab9677d0aa3e1075591721142058586297e0527cd3ddfb917c6f2c6e5b1e2d05e864b670496b8a7aa35e0090a6f16bd83d3bb36b645c0bafc00d12de1f9689abf38e34a980d62080b03768bfb047bed5dea5836529541432287283b06181141d8525a953ac4101a941ecdd98dc9bbd0de4cc49fc8fbbff4053af313fba609c8e5ebec9b506ea5605027be909d3d8e6f7bbf2732d4add2c2616fe0b4f21b11235b01ea9f9dc6896d029df7eabb6e2f5000eb1504dba066cd25de6c5140dd32cfbb8033007e5014918aa7e8003cdd622b7ccd89b6bb2e7fdaa08247db6df34cb4ff44008d99be5fbbaae492af3a9c266632efaf7e2acb8d76263edd962ef37cfec6d6bab80f8a8c7f22f69bc6703573c43435533f1492c9db1acc1511192d2f542717b1d29dce578f61c1f16ab525fd0056f5419ac5acf869abee0a87a5e3cff35c5a9259f367eeb023d15b357dd7db5e9574514feac8697d35d1d8b1ccbbfee7bd861c9f8c550e839ec1d649d85dc4bc849caab7f5ff02961d8ea68f7fc1517227bffab107d6011b4d23566d0a34307da411af36df206523c0a4d0d763af023f145cd67524a7173d58f95284739d0d5372019914529ee10cd193458be40228c08e47865dcd381a960b3932b0994fe5f56a92d69325297d21469a902cc3fa11a53;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'h2d7d4c30474258e7adadc5d5e90b537bc098ffe204581328f05c484ea3781793bcbd52ad013b081c3d1fed7da47fffed6b2d7e27b6060a42db3c186865bdd6914132a0f2e1de49148f6056141552f0a1357e9911178739689d0925464b3a42fc22bea2d09e3b158097b7d7eb0d7c5bece4c5d130c6c007495da16373ff5d897383e99c3541518589f836eddb12f87377237e0cfc9d8b1596c2759c6f6ef52e84d6ba122e1c28937542cf86a7721df6ef954c7d05316e25fc050e4a619a956e7c4f16f34bddd73dbd26d369c6709922002a6bf6fc44a4853f413d20df89520da42fb7cdf431cbb8f6b61ff5e875b304f9da7afcfc144069f8c781fbdf1cbf20ce60c370b446c59ccc42c4c72d48589959a9057f28442a5881b21a532967613ffcc001c00d0f02db32e723ccb04d1ce425f81954f17799c65d5994db161c708652aca92e0471ef19344cf2cbad6d1bbec582dc963bad0cbe7c31e72709309d29865180433a363688fbc9a243deb49ce97eb571ece27e425fd3f6a9354507dd99f4cdc3183d413a5f80a5381f4f93fd9c5c04e4164824e4013ee6ecdbbd33b6a8d34da082dfae8dde366ce096bcd76594ee91a59649e959bfb57a54647e1828b45b56f80b36f9e7cd1b27dd6f9e76b11ae70daddba4599256e9a398811882a4dde5398028e0b36355c3b2363f4fcc49b0f5fa3f700e193f9cf76f5854fa2542e8e58dbd446c6665994e805159919483b82a62b6e8ed38f12c6ad53a55919ffb33e40d10a1b9bcd38b8459a569702e1ece016f3f10f6911b7caed3208fe27451e2e506cd34bbccffc32e3c76591411a02c3ea852838840b4bfb0ed4e2fb4254dbad76baae27ad4c44f0561987c876fc0e3e375a29d128ab9cba8921ed3bef7eea3c7b1a1ccedc566ff4c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'h572858946da10797f87eda3aad2b734136e7d408612b99aaf513ecfab96d9b5cab0311b8b87753b385c662c5125f7e80f6f773339855e763937f3fe0909a482bb75cbe611722b3ab3423524bef418109b46a969345a696f16a39a464e35ec6b4089fa800c7168d8adfac228c86ed8cd02649af8b9b7963a5efd156f4d101864d49426f09e82e4a23786c49d923f1d78314d2f8bc19f0ad3610ff0440f45eba5eec09e0d28222a79cd2fa9d5fd252ec00e000c8d58be675e62ccbf7711f8953bde2949df5c5707ae093f0629a2498725d97218d60d09d917f260dafd3a5a6ba592776f3b8fc451d71d47767e324ca089841b93a48fc5845aad9f8eb7bbc3326564189424a1ecde53e0550b7dc141e438345f0d29ea1c1927ad0aeab0f0817af16a406a19c3a9839e086f8a086acde1f343343ab7442c4aa2a1544ffd467853ebdf996301f48a4cdc38f85399a9265d060fc0045d1adbcfbe65d49ac6042ca7c48fbeb08df5316ad83f63539d83cbec6e4beaee7dee772c4df742aa8e8b46a2ab52e97388548815bdcba555a87df9c5647910a64df1e0bfb73ef40e0bba7dd77069849237fed8b6600200781056f204f03378d1dfdfc6d671e6591290c0dc3dd46b686c60a5829e669adbdcda6876aa7d385810e66d30c4d7b033e516a9d96db8dc5374a5aca4de96482d5bcceabcb38e43a3b4d3971c8a449c22b55db52acc420027701f09045bc5960faddd3503b2b945d929ba9233e5c648391ba6881254aec35148c1ad94350d8f1c166765d55d055bf2d8658581695bf2bfb977c66759e1f8e61bb0b1f0a9054ba7b420d00a50550f754ddc28461361a6f2a622650301cb09a51d1cf71a127d6d6412c21490e3819c7660e3d45a5e0169350d53734e4032f88cc522df4bd322;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'h3823a90b339cb6a3decd7287ad148cf9727c706dec869b40e44b30091306b34158cff0c5d26fe576c127174a9d082aed403ebbc9b35bb058e0c997ba34bde060f1765403f5402d5413f1f400c1b819390ae42542fb14b842e89d965a0f898b197a325eedfea87fa5d3cd54bb2441dd3586310c278efea2b84ed2012fd13b7ba7774f1c1058aba8a07b4c9474e3d35ed155b511b857fdfc91c40e32ef0e8436c24fbc14a6bae886de94d941b823624a717d099c6ebcf0437026bf130d436ccbe66324099c6e2be5c16870268876e2a9417bad0caf61cbac102b304ef254832520e815ddb59ef6dc9a6b9341f5a4df9217146f32b641c2ab0fb177757bf29e552ac9fa21d24ff76a1bf0cce975e680d1e98963c0b65e1355ae5ba995cd6a9dd2aa84e38860afa2165662044c18bffa0ee160a0c69791e7a9905d76c624329b6c7980dc54f62972597f37b7c6b12c9a17ffc84697548e02741d49a746b0e5cc22d992810d6364be3ff08c6c24911a03bef9e1a843422acb2145e9ca32fe8413f74c961a1fd1d56e021665ab579b3b523cce078995ac95247e682c69733645a2f73b296b1f9eef4cd33c7890297018637189a96397df3744baac82dbe50f2d600bb4da3253bb200d29a3183ce0baeb3ae4bb2f80ede5feb9a51649b38edcb8f243ce43bca46f0b7db8d1e9852e0c90e70bb155b6eed3b059a4a82d8bf7c77c30811f8b430707ab5a823f520481a6f23316adc0458b937b9e8a668b9c2d397089f0f540bdb4c7934184b3a6acb2539af7514fa15bae83f067ccd4eb8dfe879a1c9c3f34d9c8099bcf8916a40e135227fd1ad3eebde25b61bfdd1be8bd73903938802dc6bef0d6014988d4ceff7d6d69614e47d9c006a0c616aa02a8d78dd31ce799406a400e8b08395c87;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'hcb81f1a024bb9d317d9afad9f538f30176c667d014fe2252261459df77325df6c89013d6dc0f0b27b9fbe10d83db8373f7561d79c23d3498b0ee864450d0d325a4d89a3dd19f76f49f193430ca8ea539cd5f359d5979459885a83979958ce1092439a0b95c27ed503e42be0682332d68f18064b5481168cfb80385d9ab4009633a13806ceddcaf8b8d47217d43513fc818cc762450b6cc4611ecb209cb649edd80e01d1ac1698a7848cd33e0eb3d04d83d343a9e626328736806e4316fed0cfff7260ad72424aeffe0fed77092be4eeb9757f32aa6cb097e8c551b779fda4b10f6a79d9a35eb65bf2f2019744a9f62aa7e1cbd584c232081443367111717635f9b1c4fe4fee08b88f9b9f929c98964a7f7ba37fdab4e867415c833baabd39eb464f431d7c0f213e7a6a040e98fde447f7fd7ff43360a68c4a7040ba2f7f29c615f634ef70f7cd3fbee3e6dea23a09c3495d419603a047597cc143f8b86ee74ffbb3016eb10bf8c2b85f61bd230bfb6466abe2624cfe6f0450c9c2abf9624d6cdaab2a36cef7f2a08567741e03ef5618ec5e03c14ca4a9aebece5183f582a4f7839da03b7fa00eb6fa8b52d70f24581b3ff56f24264928d943c3792942b31c619ab962945ba971ef25b625f13184fb61de51f6be47fc6fe3c619a2ab2e44954c214e195b8d0bbe7d0950e5250c6e1babf1d70cea72e7a41869b68f7706874211fb27444177c6871c5fa15b4020d406fc836c6160c3b7e009a0b7f80d8dd9b2bfb7d9a7ae74207c8e41ce7229a43d3c3be32ecfaeef8094d51db4a6e78f6df5aada3f4d1c84d3aefdd6f3d3eb6375c69c605ae2d474c7a175b4eed905d0f5731fbb0a7b49b798a71c89fd8d5be542e5b987fdbd4553655eb0f027ef67d2818394d9752c85eed371a44;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'h12863efe8e89f7783ab44e08f700b688c4800b1d5542b91774095886cac2ede586b673eab0cc36a3031a734c6e8b584483e7d83aba3db5dc9b7ac578901aad9e9ac756707b2587d61f13c43f25cd3c098957939761b8647fea33f849a3127f59a92c34030231d1090bbe710bcaff4b0cb44647fffa7362980a3c2fe1aadc0562f6f7532abdf839dfdfe00f0375b3f8902bd172e2f5a8a62577c9d483c34935a1fe25c2491ff8bb77cabea685324c80dff73f00995261e81e44ffab275edb706354275ddf3acc91e30226b4eefe7605908285d8436da19738949a787c2bc77b482602441d7cbce884648fb9957a66577adafdf157b8a607cf85baa945ada5c9af45c751c7ea7170beab1f42358d1060e6152280a914e40ca38d43e6e093de3c3507c8cbc3874047b71e013c1831dcb4ad3f9b39e07fb88b3df4c8cd20c51b393806e01573182aa226af31fafb35cd1c3ccbd24e27d729f007414c67a7971c441f590bdc3009b51600599d11d1e18b969daaa0261ccecdc37e583120835486a0ed6626c2ea96c884c2f4edd0721b981436162454391f0e8fe13c3f41e6bde78bd0ffb08344bea793b4d1edfda5ecf187b082e2655d88554b2ccf3b0132e1ce6b1a9c65a1d55a681fbb6fb0885bfbb6f259219ce48041b67a20f97e1794c6a25210a17130807a42f4be6e7227122ea68d2d9830fd1f6b4f258dc67ed03283dddc40ffdb4080ddf9c4e3646fc8f54f618fc6db2147f1b7e5e47e681d1c4b9289d572c2ac3e3e36480a6c84a68b4415bd020bba6d37bc3625f8fe804e7f0bf28eaae7f78364820daaad7b9dde6dcb1a5de5fbc1b7dc868bd22eaac0db7287a070ab6ca3ce10a804ea9f6e225c2e54d60a1990979186e048d409a49e67c8674ff26bcd7e4a9803fabcc720;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'h356d64786e8116d5d696d9cbfacd15e9b21685d09f5210f5c78135b36c04d32a33687be52b724c56798e45bacbb10f22097cdb75ab6ed062bf25f2380991bbb95b821cc37cac862e0074b50377e960a2cfd17b1fbdad66db040fb671219cdc5018c9fe1ca96bd05cc058b1c531695da641e5fb49488beb004dd750138d44f620b62d24f29cdec27096f1ddd3505c019b66bff0814a14d202b8289d294d4641772e845a5d8a5c5aacc07310874248e4dbfdf15c4ad33b930b4962f7475062a9d0fbf32ad26dbe2254e7c791234fabf6adcfbccdc6495a2431022d0751deab46a313c7753ff1132b5c8eeeb2b9897d8c8da22ffe0e3ded6119d473b0c9764e2d0da0066e7bd4a4393cb914f7c3ef136e2e859cc288692bf0684b94306f917ab3143ee4dac42c6fcf21c4b534bc5afb69703d4fbc9f25dfd5640895641a71c6dcfb727ca784c7cdaff9a4ae79d998935c85155f9e6035d719100c2086b714cae7d5f4cb7d719942261067e585ffa8c8e9329b75e6e182cfba264ad74280fca879abc4651fa08c52696e4237181aeafad6a7dee8059884cc27c8b22ed8d7112be3a76eaded539d33884d99793fd26ce689522257102ac1b7b834b62e99e6dced63b6d27d78ddc17bfa240c73174db96baf2f89e261f7efc3bd0e9a8285910cd3a74dca218faee2eed116d0b1421d949e5917375540a3ad31f2f4f1ecc1cf0834b543ca241ca027639a55e12614f399b7b5835c9cee423992456421370a9178606fd0499fc0110464654b437262da6f86a7d788e88e24e1cd984312148465f1c85204bdc96777a1ef755abde545555656631b5b35796cb0e51522c9529d4c687c72a22db8449c9417458413bfa33b639ef33e1ca860233438c6326b04edb4f0def1b139f19cceda55b640;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'h80cb1351f9e00b751eeb8f88401895024f285e175832f3abceced49f461503e8f1f971dab9ca06a9a5736354acc6e39285bd1ecb10c3ba15ac80a66bcc6530fde02b0ab38b9be54bd6321b00b4044f413ba0230f1e08c852c39e9e40d75d247eb0e34314f2c2a94a46084d6481b2fa39027ef8079e4d1995879842ffe71277437b7f0b29af37749a04f7a71cda44cea2e86c154e90830fc1264677dcf2b88e10e0fd0454e1a39c89e51b7b36cf179abfbdc535f49ba5f2809456e4375ba75d62eac58a3382f46dd93e330d09ab23c3ccf260733f3f0b3751221f1e2e3e6ac3bc4634dcc5e5693553bff038bebced2dde711af39dc874720f21f22faceb9aabfb025e48c3202e4f7d1a589227750c81970ee9ab6125e033219a0aeafccbf84b08b64400ba96a6888bba3e1f5f694194efff0b78350e4b9f4546606914afe432001fd1dabbc2a0e0780955edd8f5fff5cc53b07c238edae8075416b116e7de9904cd886e7803ecdd0e6b3b3850050f071bd97d8ffe9af03c04c7603997043728cb30909a139bc0c97063d55e2965feaf3406d54a9be9490244e313bd3b0dfeb0a70b7c176d25d587e4a3901df53714618e892ffdea7a5a8af50f86036e887483d374593cf1373cfd9d7dd7a0fd6fb1988f67917653c6c37f16b972a389abfd685a81c8924cbbe6cfbf9b7ebe5a86f71792506e4020c140ea4c5b33fb8030a1f9af3a534c7463d76977433ee9530ec5a2e7570910157fc8d3d11067266a4bac71731d2a47025ac3868dc3982918ffe6531a0bf1b9599fe80ae9c7fdbc3dc34e1c8ab2ed3f6e51ecd6e45ae780ea7b9fa6a26131741b4195915ffc4e3db07f98d56cd16c2d9e425fe57a3ebc4fe8d1508ac8acb3eed5820f78f2b1e040241659c98f98cb6fab70175749;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'hb5af7c2b4e24eb9a99c9c32ed7f2d70f9c0d2510dfdf01ab7a086cb7fdc018c5444b4a15ec900e3317792a93835557f35404145aced1023ecbf42c3a98883c334bb770e319fb769b6ad8cba09bc7db3ca5e7cdb5118f03a54b7953642b2ead177f790b28a362433134892985e53d6bf73e38cda37a5b01e895ce9f045f76176a2220bee69350a107842a2445eb172469367e016d1f2086798071fe3ee51c9d5b2b15d7512760491ea4c459874fe1763d4a399425087bbbd04754c390918ea9c31f343f7d86ff4370e76d20fc7adda32b7fb0aa19e653333e1794379c97925b473518361d6d3e66c54770f53bf3a5780489b8a227b549cb7bb17e39ff34ea3bb8428ffe97f7d2ed9c6b288a6a7e775640b29d37b11f67d8daf181b58eb0bddcc0aa48594e973ae5095ad329700599c21eadb0da07b455a4c5ed7d9aed676a7b54bdc759d976191dca77da9297478d6d32b98dac741950adffd1e24a87a872840a2f630e8d5c2ec0f9544e13e9d1fc76c71b06cab6bf6fa357ac9d8e99b0ca4d8d0be44caa1aef686f84c4cbaeb6e690020262dc3d64be0d0cc5f1be8bfc1e8b16fd156746d9ca4bdd238d44277f76fbb92f1f6fea53f491192d7a98eb5edf7801b2746bdf1c9fa0c548e8a278f1a84829deae61a39fde258b065005eb9e8c31560695d18307f184011eb52a6bc39ac54d948f4e760df14aebc665323d25b5a258f722ebefd539c7c656e8c2e5d24d4b1801db507c2735d9b88ca8205783424ba352771573e319e870650ba669ec4a764e7fc4eae4a33898d8edae2b88b850308aa2f9b78d7e54644d2eff44523590f9c37696d8545c2379aa1cf192af753db866c356bf4d5b69093a38020809230d295438d8f1a4a1cadd0bd79b5ec47dec61d77fa3947509f12439;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'h3cca21a6cb63edb3c4e1291910df79b6b3e4420e43e2500048a815879a06aceb66905eea16151b7becac00b1ff8b8aef88983dd7f7467f8345d9d0a980c5dcb94c5d5132388ec0ed61d6c590d196c565b81593fd44cccdc948fda4c701588d5cfb12ff621752805cef109ed0f357a9da15572c051ba02d5db8371da3dbb68d9b5d78987dde529f01510b33978a3df3ae6fbfae6b13a94a7db302f5120c5ca43625879e354d23b1181cc3106f895f190383686fedd3d45d4534f295d80a526f82edb59b3c4b15bedd55babfa2e759180d871191c2f7bc41b1d4265484b2974af20733a11e64c998f1b3179337af5a2c25e585f14ff55ba16e4a3e1f4f13a6806ec8c74e70e9bff5cbf221ba4318cc16b975d81066a66f4755f60fc599da6de3e6ff2c5e214e9a95514c6e6db71250111df1593202f545b7404905c3af38c36bfb7442535223c0472482798f4e34602724c468616c7bfa7db1c5bbbdfccc7c899636c14c902dbee45c1868330be1f4b6913705502a4d7d3662730a97446fd21f683b622be541c72aa9f9b5deb418caf984e0205429472e5f8b8cdc0a9c4c39a8bcaf38d70d6f7097d2f122c05687cfb2fb104c61b84c65767ad09eca2029b5bdb022f8d1ad58c8f81be8730995d4d7f4bbd747dcc400dd6e65622ed6fcb318a98c1f84970b0dc5d65b1aff5576fa0dcadbd58abbe8902bb33f2b489ae391ff703c185c728cf5ff6b1ff495a4192e6c22ca7733b5f3e4e05a2e3ff3d258b5358a3e55e0922c5ce3bbc306c1d75db83ff21c83034161c01e5ccbc30b39aea5d7c5532b4cdf25237cf5c81f93d1deec02101a3caf10bf8473b9ed384047e6b684d556f9f186013f6f3b7f37051b6c96ad6c1f5b3fd04644f96ca9f9a6a2c507a0986f7bd9a8bd229fca2c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'h63ce12c11e07992f276d755ddbdccfe09e27bbc986966125c74b37d85518346c9e5e115dea0c84056597edf5fb1169f0a3ddfea0f239204a4bd2f1a6ec6a37d89dda5c82a59d51382c10dad6e405560f86ea9e09d20b1eb3023d30e39a1441914fce81e0aefa9734ea1ad33413e3b3356c4640f558776790d30db51d72edf3a1f22d0b30e73da868b169a3e090988fec4a9467e96555030d3f0fef943dde6ddbcd285a3dcae9f44d4b8259ac2ed54f24435525fcb13e27e780f15ec4dd6068260250bc26ea273c88dba16e002468b4259a0d9d68cd07c49b6149fbf92e4f6b823de7e66d44fdf5d69e4dc103be78e537b9403eae70160345b08e1792d29fb938f7bdb3fe3cb8fe7b24a95c3e61969c12de8d3f9bff3db9d49ff0d2be34136cc96e38b452d4c7cd2cfc43b4594f24d48388801d0d8abfcbcd0af5b8114a243767395bd6f2846289a877396448214011ffb6aa65a9bf6f5e44a4bc8e432bb60c3fc84f954772d66d9c66f197ac5f89cd560957332e1c8feb265b3d87523489d77cf8e965c9fca6a9db47abd511be51bc7755642b85e6e06d779193284647a944b63a12f3c0958ff7f250a5fbe23b7af5c9fa4130a9aaef8275cb8e16c8f458c85e2c21363b62f5e8e0e62fd816f65b5d0cb758b1930cf229332cd23804d8ceb4363a16df231999eb65e3eb87ff2d96a0d5ca551f4b1e3364381410c72888627bc7af1d126fe89d6e9b50ae58c516cf10ab517e17cb39cba5665c2bb13cf45a1ff0d134c4a1069396698ab7be7ee9287ccde23495cf963694ba0857477949e3c0a7c1d7866dcb35812d25afad0a33c8935cdd7e8d7d47895abdf33b57e23c38586b39a94021eeee9adc43109798433058ccde240e9066f831d632590768219cde26e5075a7c35947d69;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'hd1bcbeaa29d763fbd194a03fbf6b6525958c7a951ddde622fd28a3a0be58f43903d4f5de8f98ede36fbef9544967dcc2a8b38d3f1759dcbaf40c8d1069934222398a3442cd321aba87ea5b55965c945eb2c547f3e8b23f42f2ea4dc330aed4e5742dccc8d9292a7c02660d8c032ad400f233f3da7ceb8f9b139e365f3c494bdb49ee1ed47e97eebb4bff51cbd88433552ef86e825a608be5274141d51ae4c35945868d9b4815421706c8ba87d2b1320e4a246f0e73dfc0365a78431e85a0d104fa8b3d86bbe4c39156442a5e96f612cede8ede9627e9ab7d09c89e4c26bf1f5eba85e7a2685d17d2294334af1dff06774a4930c5db27806aaea9006b5b720a5cdbdb3b72358f7dd8ce58a9d4486484f8de4149cb54b58506d2e5d34dd2cf36881c364bc87f1951573f832014dc419d74bcbd4b26f1265b1d1ebd59c250012b01a244172e79fcb86952ed25f7df952f7b02491ad2d733457c9bf218bb30f7d780c396e7eee1243c6d681933f40f06f7fef8ddd5f4eae8713c7ec5c9ff8ae7f2abc3d8dfc008063ae553fb574370a9ffefe0457a15e718c4c600720074f8ca1bfe18fcd1e6e41ecabbc53aa6bb03bed7f23b8e145ee79b08b47c444da94c8d93897fbaab8254ac924e55555c7a61f4d4453daf1ab57c68e8e103476356ccbc44df8f7f512730ca1419fda5e43ce45c3ae4c9c6610bd48504d94469171ec91abf77af952bb92c30b583a0ab71309beed965f354175897c752e267b23119bc61041e47f1718de4029763e4774dc0c0e4f01e85a337ebb5ca427471779fb6970190b23832c27e22278626724b4bceec3e17e4a1ea57fd843b77767364f9fe1e95d04f9bc459e0a52280c46ab56d9795e565eb6f78951bee51b5057e768b8a840b6168343a2e1d6e074589;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'ha179ab60cb398bc6bf6fdc8fc32aedd7b525d41a5740b7763962e266ce38d19d08b5b688e27afb271595341fd4b2e961ad1cdbb69b1710e412cff472e3ef9392afffb989cc727db1ccd4e0e693dea74aa741685b12055383f7d419c907f4427b12072f1365ac101eb66435de1d2c4484aeb31f67e4c9846344b0ec6c6588343c93347cd027187865bd6538d073be7c2dfc2d3620377dba588f97ab809ad3091d8b2c5f43273281221706613bdeb6ac81f177561c5a6ced3801bd21a6e7e968e242489fde8aea12dae68ecc8c5f04265529cd200024741f82e560b9bbc1f84f09f5a9918b92080196e12889d61ca3f40f9f26074cff4ba6dd6b1d5881536e31be4d0a2ed07faa06b83d8cc83b65011814e88831c4b4a9eeaa8da5090690f11ce7c710e0e976931e360f93254c37746db51ab5f06c2ab8bf841d10eeacfaae601661dc3ff9755b4fe7000446d968afeed898567444953652e05b204268fa76ea95cf29353b0e64dee1c37e580ad0076acd875b812144d279793a483bd84872adefe8a8c482ba7295fb55ca05100c73f255be14b714f851d6b650b71af2bf842300a062698ff8e830e98d68c56842386545ab5f34ef4018895f2bef09a5e829eaed708029a9fd761a9928eecefe8c0252b53c67656394802d40232e5baf208d1ab69f3a9f3762e4192b8c070f2669b7bde4f15c2a5fca7070005789a4da83fec7b0b887cf293739b1635ee54c471faa02096fd0101c312ec9c9d384f3b47a37e9092089e771829430ac95ad583f4549b85a0db48c89d6738e90dd766c93a7a6615d2f4a901d2927b2901cc44972b93b475bc655dbd31804527501033ea83eadbd607f3aacb5db3e0bae3d8f5811b2396f66f4a5087e3ff478fb0a5b50f722ed7b1259d5cfaf53121a4a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'ha78a9f3aa16636e004bffe34093567992623469b740c78de6b7741d7026e66f190a9fb6c2e8d4bce84895b90929a9954e3636a556ee8f5ddd5db43750cc48d8732ce6ee8e73d42651cc06dc9d205dfb0a60243478d6b11e09e5b42afb15d619e9bf355263300223e47243a514c1b8438dc09d1024c7bf602817ebcf1d1e7c685159697ecc63c1077b309a6be112c9640292ff914f831624806f3a51d7c882f7180636cca3ef0c4f944888e3f5173b1d9fa82d4f1bd0ce3bc71b40e92877a9a87111a2222a8784f6536b35b66a3cde3e62f2eb0d652ed85e3e67ff1d6743a0798eadda187fa39d0f1c2bf2c802b57dbe763a97f03f0f8de73d814243d1eb9eeeb70b93de01d8f0b5bbe98f8dee50d00eeb57532581ba6ab8ffde25ce16249a9c76cf8c9c2ae7d35c8b0fd565edaed3b0a350161ce6d74c1f47c5f12feb60b72fcab3c8dd70e9a2566b25a3807a284511dda3e152ca66676c98e133a9916f4e45653492247ff9fc6abcc50bba5c1d44e5310fb88df25e586d1a4e558a21a024f9bb55103e54f7de225e99b4def74fa59b0fcc1654f261b2cec1323db9f0a4afb35dd15a136a26aaf335ad4845204b2cca04765f5df02fa928ce7d8752e0ddc8d81560ef16a88446d8fc2277ae6a3f4a6547dfcc4543c5c1d6c5eec561283b64a5dd6eaa0a35af33049b214955aaa8cd06d08a66a2fcddf7f708e5863ab48a3f6412d1afdce6e943152e14d62511ad22e84f81f339f91b808f20249f3d52235bb9d5c516c326a8ac469e5b55938c9d02b077b1c95627f5c70de4e6f7a61e72fc07db60e5244fbd0de26461a4da70900a0ea52994749b3f1da434f2c293c107b71a5352461cec0463ee519915dddbcc66f83103726adeb004e71f1d5996f3a43a479201feecc23f21b1e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'hcc48ddb0290f27480eebbcb24b0d7598b30767e018abe28850250c75212298a70d47e8b2814949b43fcb16f01feaecc2be7af06c411524f506ac9a15f450cffb9709db89c831d623d92fa0d06f6a9e706236c8c8d7fcd5ac0b5bba2b8dc46c607b8718d4a0b44d066b829cb1c1948b147fa0215b82defb4ad424ddf95d9d2ea883fec55c55dc86a08f85d363efb378519f32142825d3c716352ee60b60db79e239f5f8f4422468b6f3ec5a22a69c5dfe174dc2c34e493acdfd1c2f61e12a9e4801a89e1515b2db03ed341febcf036066fa4aa5e54281551c3957978c1e8e6db7ce75f39650d65e883610aee6bf82883d250c881b912a3c87a157ea08bed3eeae569e85b1d59e30d729a65c16f9c89cf4fa23a30297481b8f3c732177c2c70ee005bb577236a22c77fee5f6d2de9bbe8cd80ef91fe3f3f27145e98e3d7ecd2be2a0e8265a972e61a25e4d8578d1b8bab82eb96b5630e1c4f776ec70b89cc5ec413d1f537540ed6904a7127ae90ea87f72e52c961e820bd3ca771fca5bdd475a50a4dad1d745aa2ba77a557c10e9d16b3ef6ea6d2cb55aa2c967dc7fabcb8a399d9f803e28a3912bdca943ff132c96995101ee6f425512b292362c6bb5e99fbf2bc19dd78b14f66bbf0fa0993ceec850e09613fa351499000ea08a56e42038fd9a1c5042eb4d534499baa7dc65eb74fcef27b54b2d7e506071898fd732a4822a63be456e2695ca706efdec92a171eb700d4991c91241b4ce0867848c2e60d1a8db5ca1064574d07a81cbef4ef5535675b188228d6e807a6a33d9e65d6c86421f8ef3d884a7e95c73b815dcc250d8991b1e645fe8e90cd453f6643e8f50d5416b5eb884b9f52eb626dcebf8dbc86f9c2466fc1ee9db8b705f532a836ade6573d0d003bde4031662041b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'hd1f55b7c7ff768bcf5021ed8e951f920fad31d1aeb4d1246c8e665182272e65bff92a6264ccb6dab0e3c09cd8bd599861458e34e8ecdbc3d8f0c3819d096a4d1388f8529cbfe66cd28579da064ab79cf7718ca059ec99a496b46356ca9d6e45ceca7d082f1ed0ac2cdbdd14886076e1d3a432e63fcc5765c2402dd80e4f6cf717dfaf53ce57dc0db64661c32bfb893a18d928d0e3aeaea4f96040fe280a8ba8c23133375bf0651b6a1c366894abb1b1bfd4ceff84cb9b115aed098dfb3c1808010b97a1a3c93904c84e90e334e69a614358f2476288cc266297d5e66b894aa7d9bb0e50cf96f9a968fb8b3e5928f500f1dc381cea61b1f67a23a646a09be0c5b0c3cfe344d271f736078dfaf428d738dcf161113e0fca1faaf487fb660a28209260e5e251a3f205264a9cbd2f1e149a347b6422e487652022a962fcde86c4aa97886f3f3117c757e781990c41e932bb10db5da58c994e33e8f4d7f73f7c5c428744cfb973a5ac85354a5b47945922bf980697324faca7713995d197c470beff2748ff910c05c0a1f184ecef35391fd4525f005a6f35263b8e50108e1b547021ceb342561cbaebc5650a0dafe4a5fb84097d45a08e705a4da317233949063c173ef02958f2f4588444de27f88261016e49daf08beb86856ec89ee0b8674b52241a5dadaa0dc566869203766015ab9e0c77c700a3ddb1ef8c48396ef151c0cd133289408cdaa0d6729f0445a01351d39e1cf1e66c5b7689b34871aed134b749ff5f86078295814794f1af15640e4ec0be2aa4794088aa348d99b989aa8208f30dcfb273db2f9434d249cbe665edc6093524c056b3121227af7810637c62c1b1735f63d5ec6bbda9206e4d74f01fff84edda433d5b7935090d08c6dad66fcaab3ee6764de7d5872b343;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'h4916f6f93529aac26b491b0b277dfac3973730ef9b3aaf053df3617d63251174bc030570daa058921c1a4b068ed40b0b69f784684fc74eb07a8b65e6a6668839b85a5ec0bdef4728ba14319a26e469bb8795d0c86adac45935193a75b7d825a636267b739c209092c7c7a38dfb2e5fc050a35d1092fd5e80d9de9cc86bab895a2af205e8c929b73a6f052c3bafc6325cdd2558f1674629fd563d24d0b79dac222f2ff3d9432210c8b9a5401c51937fc68c78ed0b149ba39162cf7f4c1f4efef94e0c5238bc0f3e00e6047cfda8017f3f56b9e68365e74de9dce4b7317283ee9d13efcdd8aa121a653928a5661c25f547ce14e4058e50bc1f2e38edb922a795036a3242d7209165519d38acfa48e209c31498cad5815ef371e69a4f591b558be997757a578836bc3d6a197c5f0bc0d480ab97d39a3402a9344c29ecbe60662fbd9a4659615692c37e27ca0be2f8922ef07c501cd150348335cfde42edcd34a93bbaeb01ea74f7be591403ec53121f39f2b8fc81841419b0e8f04dc9f3cc58472fff1ce8641fe912e7d7952021bc2d67247cc37899a6ce195da05c66ad27fba58736707735d19da79330ddea7c007e88661f36b3d3e3e228de6ef0694bfaa6c0dbf0fabeb64d462cc0d3290b9097e18acdbdc9c270e2ee3c4ec5721527b3385d540e3a50b1c4bd56bc4d53d82e9f43f42561b0714ae5d6289da3efc7769af47dd4f8031f8ac4438b8b1ef6aa6ab3573e179da8a62597f7e2072e52997c8da796b4290be00d73967c1d1ea078aeab8c9da326097570389816420580075d8262e063728ae4b0127363aae5c7403d98de053c98ac1c1a692593474417ec98b98b23f4fad7130ddc32d0889bba596606dbccba2254fee1487804486ee6244e6d1fa5c9f32d87d8e9a6d104;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'he3b17b902b277342a0ee8730f4288d2238b47e59f5f352a1bbf78378a5747d7e6b96c0ec93d8a0497a54c56dc21d9bc08010d3284cdfb8d60ec3797bc7e3ebb49c3bf3587e6167c5bc0ac6b10b5778f99d4eccc4a14735a0c1cbca4f32f7e9cc7e7f9d708c52d0ff6f43ecbcc35198e99b7424ab2daf433783829cd1fb145ebc8e3aaea5d9bf94817a09f995cbc5aae3f61d7f4fcae300a7fbf1098a22fcb1044afd81ef7061187946f84c7dbc24eb32660aa779f37bab66066d1278592369e9ff28514b5212cdaf3935a2f514183b9516de33f455d11757983cf1c2f8a7d4b7f3370b7435ad446b561162e0b685aa13c9c7a40545ecc6b5d313cf01a795ad23db931e6a3946516abd5affba1cca84795f71aacc76b188e1533e6672cabf635956acba40188661945b1f237fcb1b597bb3464b656fb81fc8f8bf85ef2fc28cbb1f10b1e50736b3916ea81cb1536e954d29e30f966e55c4ac8bf44f2320ebeda11c5e17e18980a406e2f4c5eba25dd7db28ca88a6dbce83857e36f8fb7f99e0256febdebb494f343f466074bc23b7ceffd237d27d02d7cd8676d5fa9604a36bb2b3e007c5874d27ea02f0ab6d6977a352a95650104aadc175468235ae8af44a8da843049269a3d7fa3efa9cc6363d55f7a253f52b2c871725f0dbad1c7e9f079e4c269ebb078c7124175682694d8b905e8d743cf25e636e80cfe01c3b6dd49ea71d75daa180d6a14eab235b75af5b8d1e99c8800babb977bb31bc9fe3a112b64e3e8283cdc7df584bf2e1bb08b5c1d0903a0e1a0c1bc183dd9eb86603a028d6b20c0e31804d8f009214e93b396705ea6dab7ed9685801681f7c759bd6e933edf8c6205ad70ab4108b6faf57b2d64c3e551bdb98101ed50da860794100e32c0ae6d5685141d70088e2;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'h6b1694282fd65a5a4166cfed7b052fe60d2c2b25b87c63378f938a55de68ef14659c2c62e3b90badf0c721bd6fb041a2b802c0056e7788577a3cc01e74a6aefda87ad63c10e514bc192915fc758a2bc52e8a6d1fbbe9a19269a4506349f579adffc000316c46ea15624fef173d99d745877bcac4da3f0961416b0169c046505684b6f6482246e32df86a54a67e3d9deadb6f819cf2ae5ca93985f1782a84ac3ad2ab260bdf29f7c303d1c8341b7e9f8ffcb8f095554b096983640a49f0af9b963a260a5e3d8e4eda9468f28bb317b583b8206536ea465d86e05e26217f7da5c74edabffcd9a5807eefa68ceb2397c3a1ec463cd05cd38174f0dcda965bc19eaa8b1113a6c169049ab230a280b9e17859990845d1d3cc47eb4fe191ab364f61fc8157771d57d20e891f05b4570806fe72447b5610136af3084c8a047873540cf731f92be733cafa316a133e10d2285f8ac639277afb53800e01a9acbf1453db91aa6c476a341e0b8d810ea475c84aedba9dd9c8d4f2777b0b879dc36897add47027dd1d2f1ccb145537c71da7fb6aa0da7e4bc63bbe0980558fc195c3fdb863702a0ada155ed48e73824fcd285d1b561cb2d2ece6d5646669e35cdf54760687683a44213b5064366866454d9613f9f7209fbbf6050ad26a7b51427044db0252726fa0cf6b27b01c35836d812f95b30811249ebd344230e6c073cfa4978a270efa73d24ba7304eab6791c1b5cf2796f5d64633ec83daf77da35b0ac2f3e76ccc023ea86bbc83db9f3cd15e46b0ee6cfd16dd4ca4f507fd3035f99d974d96b793d282a1e73634cf1c1df40a0ebc9baa69b23889d5a26bcef5f9cb8e483337f4e3ffebbed4affc81fb01f890aaabde1ba504ae14bf4ca9e0b9064bc25a79af2b0b6e8ffde2c64f189083;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'hba2debb02206afc5314458eb8c11fe51c85804121b3a1ab85ba8cba715e2e04b3ca01e7bc9a06b22d90675b3d3170685fc3b0c18093d114923140240a009263f40296b3f6a1ca9f06b303c7f4b0bdb5540b60fedc943b0c9338643e4e92d1cc2c4a47079f2a5f348dac537c37ad8501e039315cf40091b368d135294b583f6f015f65594aba29a1e0be315ee6d77fc5364e619354b8f7683220bd0501a7b85963262b4b7ed0fd0e4f07c665aaa1c83d18221883e2e11dffe85058f769b1348462cb4f64e3f4ab05c0a6c67447f67ba86327fcc46ba4547d4fba709aa97e14bb0987673a7f86dc8a5c48efd545434ed617720b8e39a8188f634cd26b24a2fabf0e3a25cfb222f88c2fb9bec76734e794ee8d73ad6095eae5666131ec199dfbc2eac2804effea8fd61e488f44f77640f527fe5a5f8b0f07b05335ca42724d51741ea3c3dd8ec607a870db826355cb5a55fefa7f02a8a97db6ed00d781e2fe1972b0951feede88951b662a0baf26d94bcb64e169bc88f23a07ca3a6aaf479ed42947013fc6d5ac96906e6b92ac519aeae39d353eee58321e570832787bf791c91050937ed1469bf32a10ccc84a76e87bc7e3e334e1db1d5a74877a2cd0205f43f39b01457ec56aa4ed0ba989aee5fd64293468f84d4f5d2ed6ac6cf5aef936dc20fd271580eda9467b2ca372f6374e6a0088766c6813a91da31c57006b1ed1ffef6516aa663be25106751d055c4b96127a95992c2ed3f6850725179f788456165fad3b0f9db3afbae2871236e094931f11fca13447df83c978b117bc6860dfdd2a01d1374ec36fa912f70ea71f4094b287835e1c5c59827608e7c3d7140727fee9ce5e53f9dd542833ce52ef3a724b613e1c342067ad0c0a63ec978209785fa25944e883c03ebee3874;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'h7565c042e35eb68c8ae7ded55b6283f6fb4c5b755ab6c85ae735f728f0beb7773cd8ba2027aa7fed4f6dbca69831c327e0b9080e456c24c9f5e27ed693bbcbc42b3fb8f1632f9174a106e3d172e4e6b2aff0c5a83d246d7bae30324ffdbdc37b6d6f9a9c3f2dad8ec7faecdf9b807c25a0d6676df56591ef510724c2a87da81051592e88843a61f73b2c19d7f45204cdc4f212eeb59d137bb4fce099dd7fe69c019bbce7b82f2639b5e1339a754fa2adaae052f721c1c6ae2587ce25fbe21746cd9b8229ef3ad8a59377ad9097ef0a4fe1855a0c5b41678a43830a13feedc762273e7ae45292de4528c42b532577ecf51aa1856e8ede4b93d7b0745a232f22fe868fae0e15a09c55d1920aebf43140ba0de22e08eec3966bad084cc3beaa902138d4ed253938240eff139d80389a5d0760e5951c3f57ec434a87c443a162720de53e172cc8c6382b4b8ed7d99d52f60bd9f9567eee25814f967a8effc1604e713f4be2349dcac1cd13d39b391677faa8aad28059c6791e5327b62d84f74b507ff3f2cf25f8cdd4a9597a235707a93138c27dcd65a1e0522fe7f8411c04185e000ddf5df820dbe235aa93c0fe75295334dbddba65964164a7e4bdb58769104b5165a4aaa666a2701ee3e90863eb6d578df7ae609e4c305f07bd63104383dc70ac217b585a7abf1bb2e3f3d83ecd33829b17277625831f9fd90a6cbc403f225201ec1e7f33c4a4e46da55fa5a50862a5287db6515dd83b4c93d6d93a92da1f8c9698deb67a8b095bf0a94a198bc20b6ee57111779e7cb3ef75933aa0e072423fe554a04d3de50827404a895987301f132720b07c327fec10a55193ef9710dc6914140387bb188b9ae125c00d1e33329c4479a0422f15a39676012123d76612ecf953ace8642d3fbf89;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'h2977ba81fa84a25a77a3c81581ad772ce62f274d85bb15935c18c3b36f9e97b6567a12c0934adde097f63975ee773df6e337bde920f2476cbe45e8a229e2d37b71895cc544dbc3beb0cc76e0bc621f0d8a557a6181552d675e97139d314909d0ec32ce25ed569f83446f2b2b3fe6128a0e9bfee379d71bb6f262bfc9c165cf96a80686ca02ea613d438779dca2425162203acb27f97ee6d4821494b9a7d82453daef77e31cf88999a8c23e13f47a6ba13f2e5647a0db5bffffc1a15b19f8572a451e1a503b8a7c06413f146880b263497153a8d0f9bdb3b414ff6df98d156b36e96d627c2ab0787d1c0bfd803e9bcbc72a11d8c76e71ebb79c7c768eba3839016d899c958ccdd3d1345278b9139146d178feb1dc6deae697ec206a535f014b839c4853d50da6b95c0d59e580560caed19bbb0c74b9946f0cf72fbaf0e9795204ddf21ee9ece5d2480db204e4f3023ff85d84123559a8aceca10acac61aabef34a47920211b249de0051a8ebcba0daef7b6225321898bb24d2d35b0faaf2332e03e8732bcf22285394b7784d8cc2228d4e221b6e5b4666e15f18637ade87064cb0430e7a242fe721292018f26eeb06fd6125e93b06a70baf19df86ca6b120748c53ab43af5918b90358e717eb57242647b19d2eeda443806bc7e21dde5c7dc3ec2f8a8058ca9f775a2d387e44778c6b4620099b861297afd36aa688d8a45ebd6d192d36099be08e0841265893627c25c294369b1deb5c19bc1e4c2cacd542dceabf0b2e2c2e7246c58aa85fa9810c84127b312ccd9f7eafe03bce40f6ee21191076a51e0d58b3fa263386ce805915d15a017a94bda5bce725dad6ac0f3d98a7aa4e02b11f23e6479f846e8030ba60ace3283599f46c74485b0325904653a3d9c520ac8edd12be23d2;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'h16f91c88e3b206a87ce02e002b83da1cecfd18a3b21c8b1fe04aab9238d4d6c3edf37fab24b4aa74a96669539099be4e3265bcb1715ddfdd81227664db8b3d0933fe82e80865ca9af9b28508a5341b8b06505707a5315ca6baf8f556b651bf62c687694bdb0bda475c8f0e5ad06abb131417412cacc8e4197bfb03edabe3d4e69840cd5332edee59d66c046c8f3c1368cd4f79db6af893f0040dc545c66e10fb09d7abc778a2ec955bcbc31da3a034c559eeeb00b70a5930a53f3ec1472d48c71b2cd902cddffe181f213b8301c1ba962beb263307a2ecf921d2117922bd0fc593e64628f56a0b0be14a63ca80efce1fe6464ad206d3d764a307868c1fc5dd05c7a249065b65db40ea783d03b2d6cbf2f9c6ed090c8c2b013e02796fb85fa5159aec5063c7dea4007a9064016e760d6e50a08a3f22d5fca48324b2f0e4b67b1aa972066b44e7a00c01edfb7ed9a5b586a91a5689727456cb029a3265a42d1cbf623120c7e87010504f9a8fdf0b4a18bbb73d066ce02f3092ebca8ba35f16112671d349d965c974b72a76c6724647f1c2ae2b5c5659a2cfdc48dae13ad69c03ef8940845773b7715ed1fb0b60176ab702c7812d82ca5e340c9ea84c0f225c05fcb8e3bca0bd93de6477eca6485792bc109549dba2460cb61ace1901bb8d8a149c8db5f53950a955d2d4a7b037c00beefa1251adc76a194ebf0772ff6ebfb14953e9efefc2ee34e609c2107a607e29b136b3ccd5da9186e3478318934f809e1a4d710092afca5966096d2eef892f977823cd001991ea3d279b8b346c4f5e3a731141a897dc36b0b58a30b2880997397e9f712e20e9caedaadd95bf31c3e76994663b5f54c0bc9955f432130ce9873ccfc42b219404d74ea7a76559484f9176d5d0981672381de97e1b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'h9df61c0c49a1197d1987f1250c39395ee668fc81a111f1b8857a85f0621c3403aaa0647cc25b51dd1292b61a844638d92c23d4ea834bf13a0e6fb62b5861f7403c14956934a6e75808a4228974c8ba1f80a603cf23f2d0898ac14b46540552639d5f4b336a3192cf3b27efbea2df1ece56b84a599f7c8e6c68de02d9942a194aed2897996f7f3af695e31ee3678c14ae39ce8ccba7caa331020ddb1c91ced51757f982647604ca3e9b290615adf22e13548640a81f6f214bcffce5773c68edd5cd02df817ea26d13451641a6b91866e83a740d17c7d313212880c6b8f0924450a3acf7029dc1fa1e9592b4d94bee1348cb8cb7bc20cbdfcf77574c118a86a3f4adaadcbd04f2386d3b4ae4eaf0dd2eb175d5d52e67d690f5f129f1a8a9c188d66e5e7ca3c36ad797624ca514774d516adcea1d6c59367398e53abedbd9fb04171252a7e05262e0d9ff476d27257499df337afa0aaaae2c182f96a674f9cfcee42822d9e2a925872a5dbe1cca1c911a4e4f4cdf41fdf4222e1c6a0cce195eb12a1fe90c30f97d06b631d4056b900205cf0a1d1a5ded58d44d8014c587ca7df8ce369c7dd4cb144cb760ac751d882ef072c5a988c8b45552872b019c7a126900c5d831ad987f52338f6cb48e569687ccf1491175ef6f1fb75d4bd1bd9f57a233706abf58265310047278615415a3601d7800fa7dacf1b218e2f88cf88dbedda4d224e7c349615e06ad0b93a03ee7c6998aa3bfd9fc7297534189b68dba66b8781f55ff5f7445b68793178063a6e81e4fa80644bdcaef869fc0d73385645f7bf92fa8b671d070831cae8ac3c72ee5dad5abf1ecd972d99c141484b91b5ce161048b90a1d4fe73b657d80b47332af1daca59fa7831ecc3e306fab92ecfd49464fccf703704d99eff7390;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'h274c53122c0aff4767a9dfecf3f5a9de4dc3856a5cf32d1dfc369ee6cf1e2df7cba586d691d1a33cd4b0b530b97141292016ae6af94e088051d8141beec0ab35c270277c9abdb788478317991a54e8248db5edec2aea71f44588294fde3b6a737ff90593f6571f20e8229a1fc9cc94aef555b36f74da4805fe658e859863a5d67f9dfcdf3fd354a8fe3bdf161e21309ad0ec8c0b24d8715410bf2c048e29f0a7859b39485af971be8b27008d05e2a96595eb63709e8ad49f8994b3e92345ba9febbf6007fe0013779826aa51274ec2addc72c82207cab983425cd09747db0149ecaa8938090c2008ffa0d2e0be0026313e0768306022974dc65d3b816ab5381161483eabee7203a1b4119b12c1b0c4588c380a91cfb30308f4dbdf484aacc00a049a1481b5618c82f80a3a03b87e8e17ed2cfe600c6768d214bf4129c3fd85582c1b6b2e493b84676dfb587ec44f93385f4768c4b66334b8c7782c356b6c213f9add3ab5fa5537fedf56705895ef5cccda344c34d2abf9467ec40037cc94387e7b8e1afc55cc7fc48fcbc1b2ff365817df7ecb6846c2c3e5ee68d1829e4a2b26b9ca3a325a020932f892885632c3cc70c5ba1ea1db0ffa62f2183b6fec84112edc4bb42610e44cd9bc93d110e8893851465c5c92b5039a7eef868a570137a321d08e8465324f03692c7d3608076ba67a15ce675309954d3c57a1cf60914cbe7787e06ac23bde5f5b472acc9689bc6ee0217996dd2d45977b608c62f221b6d0eece43c244194b1d4adae5a43635a3772c07d0f3cbe602bcba08e37e76f1591b8ebf951faf49a6e9ec04c625fb84daae96e433fddf82239fc7b2297c37c0391fc44cca030a4d61a965937593f08717383fd45beff5356c9fe8634395743624a3ce8dc1369269b4a461;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'h13330da4b99cdfcef9e5df2c4402a9270c2ff0b90cc7cde9c370bb3a63e34db3538233ff5b54ab3344d41aa0dd2efe142102c5d3462897d5bbce95427f85be13865fc8964e4099fe4d4b685eab8dbd33672f54957945a353213f2ee30258bc5545fa3b70307c76a84d81cdf24d3430a1d235e36747dedc64faa0a89690c8ad7f0a484e54eb4a7f2144a12ddeb888b5b701d91130abd641b9ceac8904fa7d89236e171e64afdc3bc9f0a71c551c5411c31909cfd8a4537da278e5bec10238b81aa43248d2e26b2040a081a287c566ee838049afd738f1867f04e1a18a7b24f6aed1c9c3b001e1d4cee53790adbfa939dcfeb35cbd9a2eec1ad2e10ee1907e01d8d92df685dc6f818e1f009b68f52f16ddea18bcfd748fc436171191c8e33660585e0d8cabcf551d2d96396e2c87450de00dadf179eaf1ff2597de4c449ac329b58b3f98ebec8a1f02dc5fba246dd550a84e4199ee84d5a8ea9ec3bfc8ed2cde41bfe0c12d62e1e0ca3c44f57f37e49447c2ef6b127f760336273b17c04a7714e824ff6206a7b5169dbfeb0e0239bc7619c2c741f578f3d75603485783832757881abbfe7f9119ef66d758f5aeb69c298d48d84cece749575ce0b7e2827254f3712fd5a5113b39f44dddad974597dd3bb64b01a174f4c197acba6fc40c6ac6b66ccb42a9a318e3364d811d28ff38a038ad423429899fe5b1318c1b6279ffbdce62501d85dd344aa7a9d335b6d988d62cc21495555da6eabbe1319b142446d6738a6cf10e32c0aa5bf9957524b45d6ba6af8812ee3856c2dab8e19328f9465b468504d4dbf2eca1bc953c47aad33b313533f3afa32a87c953809aa1e46314c47d002f4160dd069db487994465fbce4a0710dfa1ab3c41548e886f111db7502c6fc885215453ca0ef908;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'h11ca38ddb0f12361c8ac23690b0ce0d93fb49458835280aa1f9cc73431db5afe9caf13a452cddda74fb3d0eb3392c91e4f36c33a739923e6af13b4deb9298f28971e3afd7eecdcfe9521792e2fc5653bbfca175af8a847886b3c77060c4976c81745919fbd80b1f196d42daab6823f517add68bc3984a63ba4f4d7f9b1058096db720184b1ed15464164a05ff2d03f1529f24c7aa684f2a101ad975fef2ced1c09b55311eec267e1a97d7ad3183fb4fdfd4b106d8af7cd4c6e4a884597a9271728889e10b60c6a3afd641b441d4d0520da5b7e137ef51a13420d0ef57c2febe40eb13fa3605f8f1020ed189afdabe951b73ccfa282a02180873c986419aa2eea8cc0c50caa31ed6b8f1af473101877b7815484d6ea4a0784accc156e1a2fe11b81d14e0dcc5132431776b37c6e9de116bfe0562a8b465eb0d13e114fad284ce8dc3be01e55e3f3802394fc44e97f43ec62ee73094392806bf8324bf0298877cd97cdd7ae71b14b6a8a2302d54a48fff2cfc04f87b55c9da16261a34a473f13107c3ec2d74515df6ad2c6389e0c1aa20a4dd903648a60b4a38f6aafce9c9d8e13e996bdb7045037a0ec0490c9c77225306cec2c1a530f3223fb435462291de58ce91fe0a539e232c57e5370191d30d6bab3aafc960f4ad96c2f8d8e5097abaf1bf6027019818c546e1bc21347166870f78ef2e0e6e4568ca33912e27e6d80927ebb6d4f7e38272e96fc8d45c2ab5be6eb69afca1e2c26bfc75c64e129949105a9cc89e22497bd4bbfb04fd5aaac62b639d85115db5a7a7b8e1f6dbfe6ea872f52a0d038e78e0d163b04cde05877e2d9bafb84d0373f909acd86245d74ba24d0c239a50c1adff46ea0e039ecf409ac8a83dd6bdef95924d50e83285436aea5d70ad1dc843f861e1645;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'h6941ddac020a9599fb1eaacda6650287ea55569f1d528b544f1f08fd93dd89dd42417b26ad5a57b859a4008790c5dbcbad2594efe1a26920a459d4733449bbefc3752d0c2fdf4541676bf4d8201998b5bb77966cf9cd30590992fc55f2a1088993dc286bc59dc038a543e920dde1749a414e10343ec882641a5a236fe292d8f834bc72a6888ff6c8dbba5ad884c9880b1047c2529f58937b8035eaf471e8f0402eb693cc683d93052dd87a5e728f3139a71a82ac1a0f53936bf304547dd79a8bfc239ef245b51f99cff53057b1efc8db0e97f52ed43a8e8f679cd50753d83e852c7ed5e12a48b502456b42b4efe00652ab1259f965a411438e6c370fe18eb078983998a20877729ae9bb643e6ede6b5fa305ad2b92b7c0bde597e99c1483a58f6a506f952407119db8381620e02659a721053660240ff1674b95742a13a5967f1c802fcc0ecb0415ec016f5a2b6b7bd1a71397c48721e9687e6d97ca07511c522d1494e76d4bbd977d93fd7c3ecd07d04e93931054330c3ed011a4efb8c80c1aeb31fd9e82f293381317edf6d03404931fd2974d0941a01639e61233cc2d37b074c756a4fb196a3cd42a85648e04a71d6b74e1618f4190514094ef670bf8fba4fcff40b54275a4af153e602dcf898cd6a75212011067f194d36a8a36c6a2cb390b454ec87d8cdd9a478e32d6267c989b79681580ce041f95b9ad351c6df7f8fe243e56b88dc8c6d73f04dae6f14a01985d4facb3ba5bdd096677e1513f745922ae3f90a3a40500c0edffb79a2e3355d950c530c852b86d01b09bf3c96668f75360d42433035732a6f754135e96b3a460c459a17ac92ff14fc928c3a412bfa56893d417663d0943a9c4e80ab13c133582db6ca67f0291c05954e742d959069bb72314309a0717f41d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'h7bcb4a672db2adce601ca9b7c6373367665961f6e89bad348f4559a22e84dc1b0a48ae67c5cf0d14d989913e337d5f13ab3f006f7d49e86d6655b731a2c0b4dab4c32ea8f4ad1c2b40ed4dbcb16ea739aefbf47c058be1bad1eb1d95bae2a64423e9546d4b929e273db3e73161379216e7e10a26d5eb2b0c698c37f020ef846d30ae1cd642ffbb325d2100ff2772718f04fce3231b1359947337e86c698cee32f2eb149ffef3acb4817ff4797ea8524157c3d2a43cd98ed7fa57cb9de23f9ac39068d75030d6c8f2ce5a40153e8971a21679b740c0d8b1f0a746c79a828c08233a12e1806e799bfea5cb9e02c0f3fc454d614a9fc08f66234ddc62f37c4b7f432901efbd4c88fdfa6ffebf5f3ee7a94278c0aad9952981a347900f258ed7c5c5e30ab64abe4504da935d20db82d640684972dcd3d696392f25ec63b5210a4df1e29eba673067d620aa3461236e150d068f9f8d8aa23e70d22ed5e02cb4e626b707e5b2ee233ad1dab462b49be9622dcceae008ee1c6c96868042fe14a6bdb8028918454fa94f0d33e7e597044c4f1b70bddd01ae68640432cd9f028441ac1e2567d789479bb7d563e4e66d2b082ba885a18571ac7ca8f42f9806064d4624ffd93d261242c55991609c8a8cc3bda3649674107dec64f680864d841af9a1c2af026ceac7ebd29a912ff5071f1282aea99960ca92302949f9a2b76e1b232d0329b4bef990bda48c8428a30b5e8a29d9209e8085a9ad51e7780dfa0d0688683e04aac5aa65a0ebe67e4058ed77f0428a334e1b6dd1d54f6187964b5d7cb72210e5fd80ab75425e3c4c2cf6757e90682edbb0fac212af95759c81c8a626dd68766b11c7a95e76c005755ba02b4b8db3ae2fe8c488e7d5df3b5da86b43cee296e419281b495c0bcb6956b4;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'he7ce05af95245735bec1aba0d692ea11fd71d5373a124240ee233ebeb094260ed63df0317a23be93ba0d1387297471807aa713d1b0d89f5f2eca9eaf7d8338a7c9012eb3a35907bf2352ba846efcefa96c40060d3e5f55e79d1f09d01867faf00e984dca62ff307a791b74d1ba076be0408521f211c10b139c2402091fdadcdee1658f5fd53fa4aaf8eed6c6b49931118959929aceb42094f746de8ccf98da16266ccf1db17e69822fa7275fc3bbc8da403b5ab475342ce067996638de6b6fcb7d66c6cb966c55b53126283da2cc3015bbc7290016b06a1063b0495281408e5378721bbcafecb781fda3fb1996b83769823ecfa324ba5013f9f1fa31e196f443783ccc99a54f57b99d39d759da42300d760fee920a0e1a8713e66dbeab5591ad0513a7c322169440a67ea6dc4d5642a48d5b4b277e33f2f635b0d976e39a3cca81dcaf4fd3af94cddb75bd1953ea8b31feefef14a01a166c480be877312aad3166bcd52fd496f1e86f24a19273a530a071b1aa56c934ae7d8a169a7d4738433e7a8e440e1a2c0dd97ac55aab8c444fe27a7eb44d889415d101122fe14a6ceea548a6d1e249010aa238028c619e752cc46b78b6071e1e11ed616094d40537a67639cfcace5ff39218983f405de33e7d21d09ba05197f7f406a4336d629ca545c767979916547ca4ff85a3256398f29b401091608965afebbe1324b74406288fc710dc9f7d8e1c2a3747bb55fda1af678306c1e364fbd0616798d83ab63ddea718b36d2d1981166b1d326081961414119dd5a632b98ca6d2f3fcb430102d0e783e32b6cb4818f1c6780bb09805677350471735b66513e9ce3618ecf0a845506ce6aa55d17fc01f947841f73fea553388be7e54f413d054a79922b43204c41b396e36a01340fcc0969f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'hc3c4f2974b38163fa6b48aa62d94efdfd848ffd918065253db97fabadec08d01ea231f6f82f118473c4526c7b8f379d9824c84de8a5e1b15cee5e08746d7579d45269f558b5ced134007de8d31b44c3ab98026cd441521429305583f9607a91f9f6fa1c927aeae346f98acb5dbbbb7ba3e6ceb9340dd26a5dfec2d2f1c63f06743ff081687db4b6f1b8d0048c474433966aa982df069562972ebd8fc5f5548edf4a1457bfad478772c473b793a919a6e8ac0e6da4878189061aa0d74389856b79215553571321742cb6915f8c434f4f793c5fb5232bbb615a757bee42cfe585fbb3b7beac507215d420ec28a087b55c7d504492fd53bdea333f4281fcab06ecb66ceb191db155295c154ffd14d68ea0f9b06e225156e3076542703b8e13dfd3f93a8135e73a7d2c7deebf1d0f0153a9399324e11089ebcac967223169da922125c17a15d7ae9af98a7a768fc6091cea013fa2838b189a505dd9cccecc070e3b07eb609d9a5ba136586f01dcc91e76bacce4ba6035f6ebc98578c3be22e291970fa18f8abcefa9466ef211ba115e06ccaf4a80a0847f2bef8129b2a3446a32db66588e6917cac20209c2f3c7042da8b605d55403d148b906b65310b05df5d83b35965337e14b774225041af25b39f4d0e59593467fc7c40e763361e3bc7f7537ec41767e7d05ab5b10230992883cf141c7af409fe1770da4e5fc1ea8eb47d0f5f01fc11c7f328c5c763a75957263c3a48e15c7775721fb13f2b9b13ab9bc7f4d5558639cbdb9d3a310cae0f2c598eb5636d9c243fcd1edb6a430dd5660261636100818ad07eabd2ab6fbf49f00d4e8d3053ba64675c6801024ad9f4cf0911a6311bb38255e42988268b856056129dcb106304a391287c5cda0ecca6d5765d4b3db30326eea375e5d6;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'hd69a2141c73e86c454f6151552b816ae7b9fef6f7b0d9651037f6920a37be340f614a5011289c070e12e0c9583e696378601891bda5da4014b53f2d8cc934afb1d6e5330ded42a58685489cefecf1f1a6d1ec7823111312bf785b0d180a98a7c33742979e6e619ba556a9006cb9503ce12b2ccb4e53b9ae3a7f24f1f4377acf4458f8cfbaf9aaa4e26fbdb7d847af3f57ed4f51a25515a66af5f3b287892fab4376c4e4376f91eb7c4481815bdf23a3ca3f67f5d0aa63647ed7e16211199b69e84bb9982a40b6b7ca839955edd511bcd79f8c022568cd9b6ed8a80a5ef7386a1bb9d992bc46aebfef39838edb33f4d1288ad149d022953b7f412461ea0cd31bfe6a71fc25dbbee8f34431145ff7e8ff610b92f662fc06d301d3d81f50556db1a249bbaba8abef3df47b9853b19b98dd0952be98197674cef49950074ff0e429edbc2655eecd6e12d6dc5b2be05b7bbe3b018082cd89883f31fe102af0a6ed4485bbb31a780ec62aec5a4503cb053caa8c62e3cd657739c8d95b322e92d38495aa0849e074a0758a3f9949f6c664174cfc500d487abbb09fb1137d3d02c717d910ea1cc7fa2d40f18e310ca6e61181c55dbf965d82217629bf80e6846721bff940c0db0ec4f66832e016a7819a3941d08e77d099e90b4a80eed87f8abab3b3b8af05e26516786f484dfb317b5c429777c3c6af0245036c56b5f112d433855dd6f71d0fca336751d78345121977c9aea75ac49cbd3aaf65788f09bdf880b8211d24eea95dd98561bba4a363de7ccbb2a94260281863c458ad4c25f7b87adf506aeec6de04987e839f45218960a08b96339ac17e1e1a166fc336dccc74733823f5b70ea8cafeea6a4c5e2d2bccc5d7089fc022ebb35f7578c365ffa18790430785474b7b9299899c283;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'hf4bf8cc0e2940d2207c9ce77ee1eb0a6aa5511663d6e4fb7ef1936c12d0a8c351764abff21eaaf2704d1a2713a3fb0126bc1127d276a8af5dbb79259b45a9943e11d7936cee8a4758e35b99ccbac707e92bfcc2ced36be8ea0a99db6e81bcb4cf0b605660a728616dd76731951bc4e43aa7715c70b578eac712531517ec224748b70e9df2aeff73b4c1002bbf7196ae4c1dc57d8c9462bc924b901f86e0f3c0106d20f2cafd47c5d01411db28228a7d57da9aef34945ba5466e2b54e9cbf285966625489681616883f0fd84aa2293f6483f627eb39ccc9287b074b6174dd523fcca13d89efa0c60837908f2afab796565e1571c87f54ffe2cb013687cab502e426d365fbe510ea04437253d68d2113e14f6f0270c1665b56d982439b2ece185897657de26e6ae6b5e58d3fc86e40a50807e495a5e81c28c61a5739691d56f9049d8e5687cee99b676125cf11a9648e9ad5df8e4ee932ba37b679acf90b5e370a294cef1d2bb5f8c22aa022009684a01af5568624ed197ef93899a10b2b1dbc7a4450417e5de22633187d074ce8d9604c239af701cdfb7cd96a433582a1f02acfde81d9e7ecdb1e43be4ca634f117c6c2b3fbb2855bdc77bc5eecfd36e8af661e5af6808db411a922a7d9e8f74b7c03fd1abe5b7143ecff3287d59c082a72fe853f93fae2d929a9d6278707dc4880c274a00b435ed074fd23a291f4e321f32b324fbd6dedf331c6c080e7953ef74354832b38aa1a8238f8fe8e366527ed58fdf85dbd926263b99b34bcfab0b0a8215114ade1a7fee73aa668ecbb1828ff735fdce2bd5fc9dfe80c6757998f423ea94ac69bda98e1a9c005ae1df123fcbc0796a5afa65abfad39100d672c17e1c6a4793dc6a264cb0843d42ef3a1e018db53025732bb80d50511c054;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'h36db40015527db4156a84f3807ef68683eb37511bc0a9b2d817e8a20febbf44720f6372afc8789607a06e21b6c36c758ed08ed7cf7cb4c559fe1aba0bbde6cc29b5455c15418f70b4eb14eb0fca726344e27a6e42bbf91241c8a37bf26f8e70bdb29eeaac21f67ec131e0d021a9298dbe61fd8a8ef57276c3c5d1f914fc8d9cd206d2c9a7c9067730419285d899f45ba99c2bd959b505818c463ee4a2340139f3689be2ee2bcf8eb696e3139b9511d70de964c9afdcaa6890ef88cfa26d8e3352436f2203abdaddf30d00601a7854be9a34ab068ce940f406e1198f2e5a1ddcdd01f8c0b64c811584c6cae467434bbd9290b772828993402ef3615f68ee24fd3ff4c65ae551daebc25771a12c5f08bbdef5f06bbd5b5b905c9973ffdf34b368725c6a3c70d52971ad097cc5fcbfe7930fdaf1cb3d0514c177fac137efd551a5020d67351500346ecd2afe6ebf277aed47c8cd1cf5ebc5ef3fb14677f10f54f7ef476264fe21d9aede12100658d6ddceaf40bb9fd69d51d969489f5a3f16f525511b10ae5b941c722a9e17ed958dcb2cbe9533570355ce8b456dfb4b052441d38d358832ea296138e750d20281fd81822fdb85c15c613beabe0029fa07727c433bee870f0c7e1ff40d1384b77dbfb6304af953fa904428790903df5aa7f57f1838730c4cd09f06af69579e98be100d95080e3239fe6db5c34b53b59bcf2395b1a8422a422e35d6f6d2ef601c8d3299955c564ac4fddb53a86810538e33a3193d1bd858389e026571044b4a619d4d72632f9b4630d1e4868e7b561ad791cdacd33b8f533cb56a4cebea582933c1bd1359e9a5ccf0751074a3b94bf1a83a4801e5f5ab3545be6759d7109ae7b1d5347eeaee14fba64e58b2e4384a7832d1624ae8551739906b35bd9d7;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'h3948109dc12ce4a62f01164b34d3d3e7495907fec8debf9ed2f25ff9005e6f08717e1cde61c5d428f589ed167901acefdc37c79b8e8713bec6c323c77b563ad837dff56dcf1d97fc6ba9a31a7df737540f0715b04aa66dbb2a3394127cdac2610a4b9bf5a268550c3326c0eff0eb7a75f1507edd22725e2c283a914317007f01ec6553f0405728fcb9c1b98d7004cb1c8d7124eac27f09bdf095e16dbdf233cd3c7d362181a2ca4b14e71965c35d7dda750a10a2f61a044042e7a180205bd24e4631504962008d44d324788e8db38444900a6fe1baa07a950697099c686efceed5bdbf88cd196c3774df1915c67675805c74b29df56dd92bbe87524aa4689c8a97fa71af0eac0fe28d1511af2e01271ec3d82583f412143aebabb291a645bb63372bcf68d130f31bca914bfbeb4c33d87474be6cc801ebdeb7398fa6353784098b5f298f94ec61f00e00efe93a2cc100151d779e2ce4cd9756ef1101334dad2217c9b8af4940ebaf7a0ecb7b4e5b12bc82e513388ac5a8703e756fbd8736a5935e4d0814c6466a99f6b6af200ef1d708ca8fa5273f554ee40fb83a8a067693c42c4eb56a0ab3c9497133eb94b9a4807473140286d215654a27f48eda1436e8956461f7656b1e11f27f1d3d42d1bd438372bc5e0b20f64605ee3d1cab0b981efa07d0103974dfae4d179930cf56cb4f722ec81881829f71072e1ebe111c25ddb20c9fa0fba5ff8e1135c18f762bcc034d79bca34df89ed73ace00cd4a35897dec558c70d3411656d4b1ae8a0a0a60ebd7f42899bdbc8123fb47aa8d9d0bef45cf55eafa2d1996a52fe8e1a09eca25bf43b08f8d3e334616d2678d9d53227aa18677e611a4552f34ed0fa6f7de7e62bb35cbd8dcf8ecddaa4d8019e067f13cb811ae73b18a0ff70818;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'hb43cbf69ed8501eced0fa7012c7d929169d0ba4b2142220f82afaa068eca3226b4edb509fe3ed4bd7f9d176750212086137bda705c05e6eba2c50b5b6d3151c4c74344f707bdebb34ef0ff97fcf5d6c6f94af58065521c43c01e20b38d020c9a9a6ec3c6937b4b220980b9c85afe32b02de844092a2c8310ece39bf1afbff6d8cf8dd4c396b12cd0a257b7b23a1fa568aa7f7a079076a77326252b9ffbe41e42edb7327450d60333655aef9d71b7d41d8969fb29f28d4ce48c1907283817b2f1040092db3f87903dcc819afa4326d8f9cf73b164b215cbce35374e63aa2aec99184833fce5f36012055bcdaa8a5fa11175c1af3d7880e2f7e583eba3496f7aeaaac68d172743084e72524bad979b02313efc3851b42559e3198697f713ee850755dffc3da30421ba71de59936900e7d6a544e2121cd6747c75008fd3e25a3e788671659dedf7ab523f64a70d8c7c590ad33f241ff7e95737199effb9327267bdcef4e9e18547a31d4802902531adb004455c062dafc9040a8a4919f94ff9f501f8ff6001d7a5c76455fcfd844f441a0b9cf63b53892a2897a1a2375f3a0797c95e723b7c2d270069323c54b68ce4510135e491e37cdbe513ab661e182fc7de625e5cb0196aa8d5346b9e96353436e0fa14b249a39bc432b1e3439d9ac16713d0f7398347b414d9588030fc604ac4e5b505c81354f55de61da154a308e58e114bf03e339b5f0068c4783cb55ad5295305ac0d7bb83947a653895faa5dd3b94cb4175fe270b286d511fa7884b8db425381ba7ecfbc679b894c9a01d16d5027996bf743c836a73dd597315854132c13b8b6469db9be409efa71a48f06d3ba2e6fb638ee8bf9b77ebadfe2f4a0881af846545c75792c7ce832ec005b39f4d005db5b0815d9dcb48aad89;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'hcb84daa24a795f8e492fcee3b0ac2cf4990caf946be1be3c3ddfc17a6d57dd4d3bfd944e3bf93c56405b82d0c12bccf9aaf0d0654096d509bf65ddcd13b4fa8b583c691f8464a1bae59f7794618d4e6c319e9e2539c6eae3b609a2db86ef0bee2847dd74f5bce88ccedc7919dcfd57e28f10c665a46d60d9a1c892d5aca595a87104c6384b341be09e16bad4de7c71a504af039680e088d29c0f519545d41b44681a234a056a08252dc0f351f5319f4dd585f742ba3eb010f4259bbdaf3c5c8d5b765bb04460c5d693c2e7a6f2a4a69e894f4c2df43f39375d7d0e51f09dca002836887fa826374261a9a6a57dfc7145de0103b3dc4271a33190e64ace437a2f97166edddd75569a375ba878dd0323655f89786f5a01449ef763118ad9684bc7ebfa020e3709077f7e50e690871977fc7d4e9ea774a439a1d7fc477fdc68cc142bba0a607630d685833be5d85c0bab7c8058be704775dfa4d126dcc51b78325530cb52649160337d3a9158a3c1e2b06bdbe96674a1a17e78c87024a4b17d11bb5cba3d124d840d2b94fe82fd6145383e439e3a7db4b389631ad9277e7671966bac5c2719feb8e224b0608623c37062221a9fbb11f9c5be208ce27d722cee5ba92a530ad7202f4e59abd847f10162a891a5c103dd03137741bc67f87b80692b867f1ba9f577ddde32f70ca33cc196a082fe5194a8b40138b588898144d3b5a01664caf7ee982871e9ca9c5a75e1821225857f7edd3602b2b6d5c236bbc13e922696392f494c29950a62717890ac1703ab7cc29555917c22350d0cf49231f1f4bf3106f0471ccaa2249b3e9f98e2a690dc89b81695896696a576a0c2fa0502e4371461fab5a599a2cfd1e4decb728f12cf58c8be0fc320b7343441622ce58f1ffdf6a70ffe82665b07;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'h7498e92c35361c0e10f6b23a203da9f391ddaea2d2890859e59dc1744f5a3d64933c74f5f0be3b16da3754d14b54e425e13c759dcce503805f452251a94304c3c516d34625a7483757643a46238e8daf21d0f748feb1079902961bf7510f1ef9416e3a2784bd27edeefc551ce2b91e3d217c3944b42637c0848810ee7667c74dd9d9c73c6395dc8bf772588d51ca0b8d1b6f7624eecdf40b24a0c38b06b32a41f123fd1f9df2f1bcbb842b5cedaf57c131778d6d766e929a7d18b620240c3345169dfda630b8541f044b690d71d295e698bbb8dd6dcccfdc7aa81b26e04dfed8bc233551a01a8c8edb988764ffce01566b85a1431b8d35e6b4abaa91d491345b47bbe6fc77bc4adc318a3abd0e0a6d16da40b1c23922ba7b2a68dfc79227359b672db118757050b6e5f9a66733d52bb773dcddc1b96b6fffb1452aaff19154f2be3ae5ad463c2e86bd11bb1b258235841e0848736c5dcb43a9a481c2040ac6b01eb7000ef05063a1bcd7b40d7e42f96b589562122232cd60e0b3ea6c1f8e0cd904c7ffa6d7c01fd3d1ea7e30fcb4380777e4b9251c6a98c8f96f6e44eea64e2741facd7be1f8a5f83a90b4821e926db97ae6f882c142ce52a04a6aa40a981a0eba3cc638865e188a7fcfc0feea829524e09754d7ad2336753be6e651c79bc070a3d6e81a49fc4c651435bfebc2546597e4a6a62e0c48e9e1b30ebfa6b4d195dfc725dc5a31477e68cca5d0e6a80399ce4226a5fac70f63ac5daebe769cf98afe43ca81a17eb186c55bd9692065191ab67b51b09c4016e0ffebd7debfd2b4c8b44720626f6bb29dfc40592f154b7b2cec242b29a455c3dc7ab01cf42668685cea379ef593c299bc1c624214f3ddadf618e108c697f839c56397342207505567aa564bfbbd3f7a8c11;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'h28b04c7d58c23c1408f784724c9fae8885882ffe5bfce3e95f3130f42adac713b435a842378acdb9b2a77c4cc11d53960ab1f06eebeaafbb594321eae367af95f69b7fee9c0ef691b051377ab1c36b2634e54b8da6586f34e8d2cbc22573e48330c18ca6c3ed28040f20a8d02ffea1090f11b68cd392b5e9e49909ee7893d34ac0fcdb07dd96d9246403b028db6722fcb964b8c085927fae2fa3eaa3865aacfbd226ce5c649eed8de862aba8f68a7efc59d043b5e9d56ab61bafd9858c3e55576024af30137964623ce886fed9b02a04c9e02ba954a19ae7ea60e0014b013ac8a70a994a606c7c9182f69b7319f307edd261a1d62becb174b187d2d2136c86d810d8137121bdf648741847759776dd918a4d6bf16916d0c5df5b32fd7dac33b2cffd86a5fd84ba90ab96caf5b88906c11d97c20cfcb9456b92a69b04cf372eb67c0d0c7fecc2169f7cc2ae2f908ed716bd9b0852cc3ca7bc8fdd85b3f6606086863ee266195ae97ce600cf33a18140cd32de1b7d3eb34004b6601e386229d06246c48985401ab006e2d397b6e9404927a97b958cd754137d1c9c0b00ea640e124c869c7d6f14607490b5cffbb0cc8f8d353782c2db5c4c45c6d59766b809326b9c62a636cdb58ce89e0c73745d96ce49a8ec700e0fe1e072cc528f263cc16b21a375e9e78914e939f5629eddcf93dd63834add64db3f46beae3b94e769aff32bee7470d33cf582384861b1aec6930f3952985c6a7b277e942f7d356d720ae226e264a2cfca4845f002859f640f65ed06e6c8b946511b56118540153fccc6091af20c6dc0bb8b9dfb4b1dc6460d13182fa9233cb31e4b155f4db001437f1f5769fc84c840872134ce19ea67887a5152b034fe07deaf759fe4f957aca37d680d2c4bac8af1c434ff50;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'haba2682d799f9f76092bf26819124ee5d93e077d9ece7350ca69e2dedd1995db57c0afebde029f8541029769ec331acce581a1f09e96fe1052206c94da50cff70469182881997d02e4fa23d10e027f9c46c0d0e917d34a6a0bf4eb6e28ecb073309c3589d2204451acd3b9901c75de9a94aec19a868c0cd6e456dbed687512ce3f40ce1ca3e582c7b0b471881c70b33c9482139362ca48d037025e814a87088b9f928148dd9ccf1af0de7d72a8b379c5a675f347ee510ab31fffbe9050765e3dc60c178e9dcf6ab963264efbefbac03c9d200b94926e380e8d12d14ee822632fb6c2f4b29b4ec54ddb26bcd7c00d0dc315e516d2b1a4f1926770fd7afa5683b7096eb5bee405d2830c2d59be98f71296a27c9b3c626c4783c72e70b47f30d83f1027cc1daf80a7fa6abb16c1d8d0c2cda4a6c968420d66b2b5586681c0461a59430b6102d82f23dcd5ca72a558472c83940d3adb533e7421726d75706c8703d50d2e826a681a53eab0fb0405cc9d382a87bf54c13590d730b1a4db0ab29af07175b64da32a468e81e6a334b133b6536a3713a4adb5ead2102138e9ca4a496730920f4ac157bd2418707cb949d920e306d50bd8a2ede08e6dfad1423a34d825446b4c823ee415ab41d19a05f6c379fc08abeaea7a9f5decf9746d3ca36a6388cc32783b6ae67ca1bea9af5c529aed2122980fd419760857ed7f627330d8cb78eb44c46f3c31c287065855382c987d5303db6c121dd290e89ca9b446311ff47af64527e2bb3175921ba8c5f103120ff4e57182364df616506b2ed444b5b2b44d3b63df53c223d5b1056a589ddfce179ee65ddfa7fc088956d85bbbf94bf0d33673240618ac97f0889961c0f9e7e2f2c6e0f001333b9f062163ddf6e3b0fc6c558e5f801e81ada092db;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'h5d4491a3f2ea2be55cd79bc5f5e9aefb2a8bf11f7fde21c0d4c2c62a193401696d1909b1401dac35c4d6733cf8d080e8b5c553bca37a516daf722be7ffb4b20f704c988a623ae03d029d75a1e47433d771aff495eedab9800e98981ad908370ba3c6afaba409bc1f73a03a11415f65d03da6dad6f6c464f3e91a8375270267c18a22ec944ad7e3627c0d3ad64fb327b496a37492680f03b7c4f09e5c6b60f9da00b2cb5204896161776a045a9c8a123644cb777c5525bc8049e836fd1e2ed385df53b12edc4ee83941abf7c7611f94eda430a50048dc282ce6f71c719879484969ae4070c0d49c860a784262c2e0bb3d3b184ae070e975ce0d4aca52f282dd1e4fb9415b8888dc6b883874279f5976dc2df499f6784734748e6ea531d80a32e29b05d5c1e5ff57e4f8683e531c495d738435a7484c7c9df16dbf9b19fae314fedb4622e451d06df9d99fe00ec1e9b6cada9243cd0daf5d10093021d11a17352ca8fce9a8c1b19bbd67bf117c4899a11b98462af43045a30ca06317fbd3c013efd989b25fb0c519a8fcf609655b3484715404848506cf1d96757da48a36b676d0cf341b76e6d338d0b8a9ca4071f052369ad23a50bfdc807e23f668b08e3b00e59ece8bc888df4ce9dd4f675d56ee4351fc780855c41c6ee05151fc3af0d6b0643b9e58486648a98e8e34ecf9e7de71100beeca2326764b65250258b3689dcb61e9661c55db992f8f709db3101324c4f00c824028f7da4f1f74073fa3e3eb8e6f3047ced869d2d3b61dc7ddc99528c234ee2cf915900fbd7ae94d4cb02ae81fea6832e452b5a3940a47880e07eeab0aaae502e5c128bfe6e0c1ad3590361c8f76a8bb97f59baca27b9581ec8fa6b0223816407726875f7431622ad1497e6967568ebbaef1b001156;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'hc61f65b02dbe401d20ec99d622dd880415b2fbe5e68e834949437ca16028ed25cc3fcce34570c6f132ad6209c9e12bc5359725bc5cf62a4d3044c335930af9b9ae2b7088c2a8cf44e168da560392780e9c3902c3dfc07ba65e7c0e30cadf50036602cfa2e6905b258957a0c11aa773550f21a818852886557f7310126ac14854d14f00f93327b377278653c547e951ef15129e04f538ac726ee1f01d75b93b7a1bc41d09438e314ddb74182b1a7cd6ff6564ec4ac42b59d1566f9b06b845cda0d402ff7c3c27e2367e96c077dcdb25c4a80c0687289fb560a726eabfefc5585a2416e5874f3dc03afe1a07aa95f43edc839004833e4e7cca604e5eef32241cfb33334d9c62af24167bfa31096ff19cf085a70be4149664e4b23c500b40ae7a660be2508694b0a2862a3b80f17527a59e5ad8391440bfe48d5676b12fbcda4f15f12afb1519471a1ef0c49f957492acecfceaa768f43f82ba0e8d9b5066495b50feea5cda1f81279958a6252b5d8da7324a61a01144bc39d62b985198f040dcc7cc2777c8fbd1a3d071a72e766611d9dd68ea8876f5f665f1f06726e58b260e85b61641137020a610230e22a07102d944e5a8e38de7ff54765c77f3dba7dbfd78907ddf046bc7f51e6c1a93667b4806aecadf04468d993daf42e109e24b269dd2dfb86f0b3def75d790f82149a911b809164d1e207997eca42c056b18d615ba12eedbdd6847aa1a8d6e7f0e4a18a8ea401be9bbb64682b9157a48f0ecfeaec8da3569cfe6774885d4887b23e4bd97615c2d6a9de72dd3fbda14eb56490ca204cd87364df343ebd2f2fb3f4b980df7d3cefec7e3206d13e7c46d8a4eb12c8f75f69340f5b41894b9f43ec081a2c1162ad978dee7d0b7597ad609281ac9981af851dfba8bb60e1bb4f5;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'hac96c776197d265146903fbfd881b20b7a6a838b357f0a6eb70d545fdeeb374534cb5d386cd46ba43d34039ca77f601102cd79f826cc7b16c66cd4f7514b100565d5a6ea40b2dd3340c2a0904e5ee952b3baf5345a43cc0b46fcebd310cedae2b6c18f5feeb270592c907d35eef1ce81b216d0f3bdc98923f8fe501e5600aa81f0f63a4d5e3fe5cfaa92a68e1ac5a96f517b5ea3eadd4dbec778a035f1018b6da7f0ab8c2be8a9ae6b5091a8c1cd0aea726d001624f5e9b6e1ca69fe05fa902ebbe1813515cccc122ec61b473f0cfc44476bc243429e10506f9d5702556dedcecf6e960caf3bac416a7082e0fe42f7f7a04095f88f80a0d11a9aeb41616e2ce70c10bf263846a2d83f3eaeaa2cf6db0ab65f00a672e7c3a2eaa0e370fcccfbb3d1f8e91d2b7b4ebc9b634a32879e8f748f6c0b599deaeb3f7d0ee2a27c5162ddb1c9a9c3488578d14f8b7cce7223da0e3b98255c62576b29883650bc19db7297b54bcebd4a19e9fefbb8751a8e792289366b4e4ed6033aed09338f4e05be573b279882f1b1ec99ce3d53354876c363b4fa88ea3865c72e0906499c5062832760dc0ac98df511157a133cb829947eff770212e7bcb95ea590b0f7efa7a02eefdf7a1a029f93d257f0de633b16a3b62930d3a9f11f04fdd2434a9656b124572901de9b1a857edef33ad7dd535dbbeed2437b2dec32f638e0a914ead221fe3a5d068630a0e2a7ae53a7de4ececf77035308f9bf337d0f46d3d555cc896f3f0bd508c1609280c5853d013f25d3ad7df05ee308e8cfa99bb98257e7a469196008e31f347dbd8f8d843b548960162e41dcbd865a71f2d56d5ec70a94c4485ac35bde7507e8ea88f7b8a171eebffca9ded64b97aba93b2c1470aa377dbd8151663701993231d9f681549d1;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'hbce220562433e4b53b5aad7e409f806f15792106f71d75030e2a47cf4fa31e019b4b1f403069a9376c624ad0f0843b2c4944b333f17872e3c62d2062a15e4ca1def95375f6867f73d924e1fd36ad6a9b01e61073ac689821cd0e71aa9fec779d94c0bfb75439d258fa4aed115fb199838c8a34fda56f6dda9bb0d449dce5db12a70a4b1b70ee785a679950ec14389213020ecb17445fd31cba9e55ed98160c5a7b297fb6cd67f4030e460fa63e47b9e1439a8921ca840bbadd6d449622a4d5faa2b3c1d0d6168efc27d23cf4c09e3026a42028cc8cb193659b550c42b0b5a3467df028908596ffad67b5577fab2726edab2c4f30a0f5e288a17793afebb10a1d712147936139469386d10ca40aaae3dd8d120b41614d31e545b86d516dfb2d75b5bd85a6e5d0563d16ba89b1b3867f3f3cd808a1a85c254b3d46383ae7c04da3790fd41ecdc3d9d6bc8a025b528bef230edda4d7908cf175ea719931f957ec86e4a783060c379584ba1a417289b27acdeed582331575dbb6111201c1757292c99f79fa266e0bef87287f9b0639e286522170050c628c7ffc5fd85b1b5d89afde0a072d8636c10518f1fce56302ef96da78909547a3d2c4ce3c41bc93abf460c549e95ebf140f41639213f49d561164f752415ba59812630e7a70454da032400d2fac1b14fd51dbd99fca8ba456b6e4e7a18577f8f7c16e312273299a14f5b719b334786d3cd59b1b5b77de8eaee7fd6116d51fe0a902c4c2890dbbae7a329421199fb61eb4c3c1111d62e5480d74086a38d089fe3d178a1502b365cb62925507af29219deb6f2c369206c8684fb458160904439283277eb9944d42af01f627171e862fa967d44a687aa0adf306b9dd7264c77ec22c11bac31e265dbfe48f44c2f157e5d44b99c83;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'h176fac2bbbd2f2180c49215b20cb11e61783ed1d2d0bc0adaba62db112aa4c615fa5fd56dbc5708a25966d77512e71d7b9bcebbd24779ea18008ce8cf0a152694797f8589fdf0906d8dde5fc7320eb084c639a89c72a2af476570aad19e28b59af326883fdf744c39c5edc08148b43ed1306543ce0d148a8b592921e229216471a2c821fecab25b137edd210076b487406beda719ccf8a12792db09cf349680f3f72525e8b8586f35bcad99205892df75286b9a7b18131f5c5f7848510b24ebae27d9a779f2635aa9621e1c011313a023610d169569d61c0bc6fd26a750d51bf05ffb7df5fd9a71644e21f038bc9f1e5f2a29d388476a8c9be77c2a07d06de265c0969421b1ad01294e2d8ca6de5688bc5fb908aa15db8b3c448273cd7d1823bd738e78ad23937c2eb0aa89427453028e8780ec9f6c433cd819c44a78177cee66a1df446b94848121294f5a7013263d5f97c4a28e2bee695d3cfb8c4039debc485d7064aaf5a8701f46a0a53fc911d3da4d0b3711a5da82f67014e0f0160708161b9bca1df81409af8fc260aaba7f5f085d8f797525486f6fdd18995709f34c32f3daaad7c109a5c2161f3fee26fc57cb2e4931886bba1b7a7544b7972f81f4a3aadf556b6f39fa18bafe351fdea75e35ab1530cd63a6dd01d5ef16d27f43167ecb271833632a36e49b5b5e0a3cda73651e70f0cbbb7818531de1146b6aa15585a12949b887e2dcfaffb5baeaa9ac85ec7e93ed1c7bcfb6126f9e1dd673af789531a586a004497e4f549cf5bb2b4e8181ca15cce0a5b7a469d90604dedff2efd2385d2632389aaaf9b19583426e05ff743710f6e8c0b5c0be586e166680bac6ba4459e475bff0575c0fd61335fabd7c139a7a6c38122e45852814d66ab30b230e6cb49c99ade9573;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'hbdeed3e8869e41d7d99442c67ce8c66fb225f52d60cd1e64e674c1a3f1a90a060fe0e314ec94b35b36763d5c5a370892b1742e1fac04eea0297876632d8aa1c5ea05e90f53b0b8dfb43a77d97b54d294ae9ca3f2fd4025de78f126dc3b82e209c4ad020c9e8e5a2aef4fdfb8c05d5c42f69b76046f2f5072afad8c8a1140c9474f862be45e85ddacab2fcddd7264e6caea4987a10106c2984dd216364c99f2405ac71422c67706619e499aafcd1a419e76fe3bdc077067833c2c544acd0c16a17349e08a9fdcd79cd2d7ed423b71b181e0d4f22ee8de7295453bef3cde3f2a11d9b56ad632fe4e269bb41d200c8f1ab94ce2ab6cd470449798a78339ef4efaa161de85efffc942024b602ade600dc32bf5195d6404ceebe05bf243ba46fd5ff74a5a1abfba6886b922c8a9f50bdec4523b2cc8c9ee34a922505410f767fad0c3c3837139c7cfa6c272bbb74c1ee61801c9c6e9bdd7e1df47419818c7d291ae3fa99aaeeccabb2cbd523527156ba3ce4ab1c4c547609c5e9f60f931d6bf6c253ae4680139b52b1879567b584d21a8fed52d2ef64e4dfbb2e6f4f8217dfd08c6d6dfa38a9b5b30d351e82a6b458de1ebe6e877c1effafd02a43217edcd63c36a73f4047ef2cf0ad21d667ebb62b436d4a5443c35d2726ca200b7f1b38a14d8ba0cc0317e503a664e1220a68a685ad3de358b4c85e1bef0ce2d06fa1da659a193a33e0b0a29a7e26c3e3b08556d002d4cd145f97e1ab29d90255025d75c281bb19ff2b0aca57de1ae564fc22225398b086e6baefaf77b293def7a0a096ed53fa21c4bbc4e3ade5a9128817917f945d515d3c3ad28137ae32a7a83a8fd08534686bbf7fa4b86303c72597eeafae73cd0dea64c3b465348a33a4470894ccb1baeaf5bceb3be64d526c3db;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'h8a80be108905fc70df7926942e18d3aee843e6d6ed8f54a9180ec3eb647b0d759d8555c7a9d905b00430ab6c1bfae6b70669ea10ca5d362b62a37b4f513783040c85a5650e97cbfa53bdb363b8a3762d13d1ccc8a712fbd517d3a461507de07db8e2859adddf696b925b881a4fd7885513eae8dbf2e2d4ad08bf3fa106467a14944835c66abc10dd249234f06e69cb92a4f9900bfbdd46502d74582023ee40a978af6fa3785eed7c1971535f210937495edbd21d63e2de1acf8966e061a02fb9ca1d832854f54a1a880a6e58407d0d15b0c3284c4a83e200dc2e4d97fef314054a96978fc8ed3c6d16fe7622bc210c5d92b53a070c9682463955461c80c7961dd589c1833e71a76732037a1801769361b0037e03b3760c9e11eff849a00a3986792d7d9cab2c0073dc31fc54e5d4e6cd3582e64fb3db6b77529f6fdb6527dcc62f600e68b2e9d9f38e0c92efcda23844087a48df9ee4b6da4d4cde95b3f01858607fd877b3f496db2f8e2632c198c4a809beb73627444484878dd63e483a48b620b8c1e52824afd91f343e53c5ebf7df47e177181fffa7007446bb17fb010d26901df21b5a4c14806543109da6c82c1f2e83eafa7b7f16d1e65d6f7ca51ba58526e28b9d324784aaef10626f4c3f87007545c99e724e24418a249862865eb6b5f186ccbc062196831ce8d6ee6f6d22ee9b02e80e998ded17cfa5e2ebebd8a54612337c00e072f381c07607f223f8bacd6b9d1d8dfc2ce61a511e142262fb56a66e672bdce0e5356fe02be8dea89002b49e089bc3e93c960a93c4545fcc2d71215d533125f33642ee36bc728d411410083011034498179bd3996b88b91ef4361bac6b42730b4381f1e139aa231ed56f94a8fdde7d43f8847b8219a7bff0f46b1ff3e3a413024b3fe5;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'hd23e493e3c9639b20e70b6952c81f68213cbd1ef95e594430b85e888ce0ad137b1f8afb5ed21cefa2e80327dfef8799c0ef9d3e56bd0a2daebe17af594039e8163603a55a67faa2055006862d7d7b21292c6adce095b21388c4b6c8ccb66994724348bd6e982d6af4a8b075a184ef42f42fbd0fadad97c829fcf9f7584b912a1abc95194d837a24452ced67404589660fc8efb586f45d931dc99de0e63e7abd4662cbbb9aaaffd3b71fd7a7b96a89fea3e6a6b91e9e5b0a24c70e97f0bdbb6c04ee5e94baf4df17efdbfd0ac55f3d03b27cb6af01a1efe60dc7815972f32aafad2492e9336a4926d0dba6eaa3b6500f73ab85f46b0b36f7e9a7c0abc1dac5f7c2236f590224adf767eca6b14e1ef7601864a3a2eb46b248a0b873e546b30d862da4ce1f07402d1cd1d9d48a0fdb2f821a126282579c72b2d2606871d4720fc340de2fd40b76d1980c857462bebe9861330ac391d845bc1164e11ba7a63b3e81f240d85059e3ac3a5f38025dd54a346c0b5734b1b87457f97c9946e66fb6c939708b780761312abfcac01473dc4fc72ea03627cd7716b3dbf26090032d9d638c2161025ce20b5523467776def3603d9b353a7491c4b171fcaff741879780f7840693d037b87dc8a17cf5a5996870f3f6778aa8ced7425e8841358ec4e9df1b989bcf1464a3ccedf14960c2a1762040cc37c4d5fb214c1536434e34a8d9ebb8e463a7903484933400e4bd122bc01358d28879e5cc94e14a9729c8d4eec0376fd7538e7bd1618294758d80fb770f1766014bdcaaa9d23b98e9667f0686ded3a6e6d7796e07042b6ac592755749fd50907ad04a63aae741769c6710914ba796e7a7632d555b0c59b299f8a88e9c6969749b60643d4665468f9895441abbef1faf6df81e0453a49155dcb;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'hb9bf3f4993a15000da60eb5cafd2b6a54645020efb1d071f45b943bb1d95a2a98fc7e545024c65cb67a8f9551cebd7a67ebdbd9b2fcbda81299b8613fffc7968049d30aed56e7053c0775d9edcf0220571960c6cbfa486f065808f7678d1708cb8aad8b9fd876d1286b3ec24dece53697bc9ba87d9219f784e9dc5173893d8da7ac0436bbc99cce447b22305df66a8d949098aa3bb5df59377310084520a2bad406b0c876f6c16c62f9b5e77a13e10a8fe1d8ea327c900fa2e6108c623df964cfa7dbfc19db44b2dc7d9cd71308994055f996cbdaf4a1a2f69b9a754f7842ae3e90011e9b030ff51de4d8c9d79077eb4fc9b35a6edbf58aa4f37fd3adf95d025e5b16944955b0b9547af3a291b4585a1f8177bd1c50f3b6eeb4b7df7b22dbd337160c172611c739247f16ebdc38da09846c52b719a5ea74f2801ffcd9560aaadc5c14296ef7e4a42eeca22f90e63513a1ee7e49379a1bf23e9eff9f3ad3552dc9d6e764225d8842777e85b1078cd442d03eef6961296e27f5c43888d98ca8b70181be5b6cb4fa3465c7731b043e691cf32365e305ea5f634b0ca06569665b856fd93e8fe3b8a63c9d261e627a36199e8fd5b1d5eb81aa8280177b41f6cc9a3ee41759de7a33a2eee7855b0bbf920cd9a9c0fd7a3b79208e31f5ad72c5e39c527f9c6a2eb4ab0ad7a49149f95e3cf571d83fae7fa7574c612576d87a367741fd460f0d07ba1804ba931e7b2a8c608a7e3363b862174745f66f3df2328e2dda58671916542a740b28519ae10bedfcb28bc5e09e4ae449491329c9ac28ba646ec97006a873586707e55fb2504aff149e21b73b19b22f368c679fa8d1e2150194d54f829645be7ef073d669c05c02732f07d9d2799dfee29bd3486759b5bdef714f85a8b42329d5a6269;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'h3fc1ca94f6faf97932f8b7ab4eff2509527ec6a997baa13560a3c8fc56d59df9b81401a779a86d7b1f54a432bb93b8d1ae057920e23ea938ea1b457b79f9963df7a4ccbf09350ca5e9851d959005a773e28e8f0ae54e5b2cbb580b84ec26b915225f40fb56a8e1a96b875cd6c9e44ca2b225afc18ae0a71435838d9dede9cb36c6dab35e6ef1d945fcb564b37bcd36ba5e6cc907c0380ddfd8c038e915429fbf5773be93b1a5aacaf01fe4520cf78fe537e71ea09955c1bce97a1ba67b836de2122cf2d25d675e1e29fb2f0b5fff5e1a2894b8008fbb500a9814f4221ecf88776866bf44426186847fdbdc2572d3047305fbf0b94d3368250205919d23ae0b1ae2155af709d7a321279ac35276c71d2cd21bb63b83efa69b43e65dfb3bb5fbde71a54d0bde036ec57052c03e4f5a4d8177c8915aca59280fc4d3be08ba9082a144074f06753e129b7b5bfced4453ef402c71298b9dbf1e34c60a662d9ea89acb801c6bfcae3bb7cfa8d4c522db9b0a0d7d65fb58575e4b0a9384080e0726a3b7a84472f73b149abfc51ba4781ea761026df5fa12c3ba011a5c8145ab16c651f3cf4f6cb3c5159e6c34d166c5d33ade97493f3f9607f9ed63b579d418ecad338bfe092da6308253921183f23f7765aa83be950ec922a4b9f1b1d8fc8a52e4a629133c0f8b9949a7148ddbed07219c96b024ad23018ae096abefc33010351b939504eb458058108ddc86d79537055ae6885d5f8557139416fc24a4ee353ca903e703642004c5b4d35600e1ddd9fea5b80f2644f970da40c9e155236c6c39307f7f1a1a462c458b89a407c8883e926d6d4257bcfe44a2b2f8699217c26c00648fdd2b6a2ec9a60b56cb0d050978fb8dd7547a071ff2f3b58df66d687079fcec94fc721fd707c6d08a64;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'hb01d945af610eb411896eccba2c7c58f45698dcd90c17c7753dbe962241d4cb692714e685246bb9ec19ec61a32582d65f48ee071c44821a6bec5c7a31876df8918a63da698f3048818417d438dc0a68e9564303d5f2fcb411046a975807ea6e87be26ca974d16197b9a29a7e36fb7e0a474797766860e314102a366e7f2e87715746db66155c1ee30f12d7aec84799ce8065bd6c4e91e63c3aca1f29cb36fa684efcb2070d0570851d523932a7cb42ed022b659a81f709affe149f9581e88b8200bc5d713a81bd24de70dcbd3f30af908e6ee7f12ef2ef49fb555cc7308a9d07ad31815f881a872ba3a84e811c3fb1529b90d4c9b85f7e3737ff29327d322475c435b6c5c22c20e76a7d776dedb3b56fd01516d3abe665792ce0b6a5b1d947f03385b4555541e5ae3b5d029b27681ec481d3d24791e3cfb9559688579faa24b1d802e5c9c2218c06728b25940de68eedacc8dd82a01b80ca775ec5dca11ae060e19b92e2eae0c04cab80d5f010760632e696311d9f098d1746c4686099689e4e09367270dbdd38b0839b84babc2e4380ae332bc77061c1abeb02e69bb944a6d7e32c69888ffa55632f256b13e60293b69457dec28d2ebb07e24c0020e4acb294d6dc906612e49bb477a6f2b9ab6e75d71831241567f95137f77b7185dc8f18931303f0b8bf1f10c73d55c0d8f306ef3d4244d7a8ad9a45d98c8d8f753447f9d021142d243b0a9889522aa85fc3808ad532369d29c31ad1ab9caae0ed1d2b84d210ebb3adc0390fb32d90e995274de4ffa93351c35b7c7fed29a2abd221d861f3ae4dc9cdf94f035d559a71b3659a9c9beb1207c07ac0c124ff55cd1772e7b92b80ecf78527a30e455bf28d391073d3cc0bbf9ad44f813c11a02201007215fa6edbcc6f24d469c9cc;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'h946a397540f3c5619abff6bfa8a413658c827263131411bcd839f23718c3bd91419557d308552d2a7a0ce56acab12305ee72632114b8dcd675eea7f444affe0ffae1d201f6732a54946ce7f0a0302541f40ce25a63f323e74ebf01fa0f93537558b3e4b01661a3561519fbe1f54929d1422c43b7fd06c4817258299592e9f0d1625e6ee2d3e733336cb0bd1d9a6b5639f81d4e427a5c2ee2c219e387a99d435099adddabb8bbdf6e634eccc13c056a8e6def339cff3e4eeb4207b06aae6a5dd6b23e8ccafcf0122a627ed99b01a2f6cb0b0150fef2d25452ece66f2cbc058090de914cd51b5d13fc19027439d535488dfe1a143389f91cee5cb7116a7f0dd330fb6444a25ce386b6cd8450298f12f039981914830e113461e1b3646af19db59d308a692a113ee1c9ac908d139378bea664eb38d74e10ddf007eb3c2dc8884d3b50cf963266aedfafbeb8f9e9faf39c62343921c71327c8f94c3eae6ff8c86ed6a30255470db6cf8b601684bd002b7f2ffeeb319af90912771bdefdf06d797490631a211917b504e590b1605b12e39b306b1a3bbb01c5116e0cd6bc4ff4229b44300bdf222829dd9583eb78828b323ea37c244cbee054773421b31b89c8fbd85aae51f9e3c22ce3307ad612fa4b538d4672db964160f2aa163e42f76e864aecd0e2321d480b79a31e796d0b6b5c3835eb6aa182ab26c55b8d0889e5c4616ba1225a4eb5429cc40012443f69a41580c1618a711dd450a8ba57e369659ad82b09084feb307ced5d599f0c2e542581e5d62238ec990066f8eb6013713c15ec39e7e6ebab6aab754efc754fb670b378bda282ad6eb2106add8a3fa704aa092fc0610d200192c68c082650c5912a4255e0afac5bef8f9323e7f8ac605a9f79010c9b922e1e0cf1b223a43c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'h5fe05fa05d75f656d1ab1c602db6df47cec56c0cf484b552254e7c1b7675ec7e671095d8bae9bebe41548784161440fa8e9b2561c750e01ee77e8ec3ba788e04bc2d64ebf0094c4fca8be2ba9a8b4eeaf64b0df9239a5b3e4c174eb850b95a3be50ec50936ec2ae83787e872c7c75076ccfab01fb64f6f5dc0ed6dd6b1adae264d909c6005e8b1a042a8027090a8b3811953f20fa3b546a3b0911bdf265e72a1d1e8d449ba1b580947314caf201f239fa1355a52aafb48b4ba1b82173793dc338b376d830de3c3574ab4121d98242afb0265ce60b846210db7e15a8e58db80e617be0b86fe430ff4db0c08251b7cf90427f3ad900c3028441c72c88fbe565ea24a25c0759a6a9ebe2d92ec2eb3c6fbdcc81b59f97175c30e2cfb9defba83c8c8fc913b878e3abcaa4c033ad316ec9f1c3bfd60c5875d492cab9612060e59308438e7a3ca12aa4097145d73f21b492fe5360df763a85b9d70ad8eb3ecd2663e04d68332c500bb79161782db3270cf2b69359cc9b7c3b96d02e98bedeed14ee7d8694f4d620cab4780baa69dcd44c8a464776e13096bf304e01520116b6b6838051bac552e37152830de1192ec5fab132a0bcfcf6d2af132106a531466f6bbd30be628d9afa76abb5921cdee3a3a0a923905389c44b5541e64080d524085e367e860e1ef41d3382a2680dd5fb76e6d01f818ad76abb8238a2790039bd0874d93db25bcd93c2438ae95de33f58030c63a281829fee3841e9a07dd7f582a45298e165f3c454adf094f991e2e019c051b3068dded31ac29297efb46d703a0e7f82a4d42010a2c29b74ca5091b73548e51b5e7b64632d95e4049e7d199618bb5344f70c16688fb4d68576d6650ce294a4cc8bfab1af45c97ed297a3bc5f6f0a3e416b75fe405044f86f7d6;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'h7efeb1631beacd9ae7e44033d4561b2cf1781efb89ea6a4b6a494f11fe7aea9e9113ffe3de9e6f00917e5a411cfc8e43d096aa68757dc5d7cac3a4022c03386e4bb1a9c31f38c6c47f3b284c6870ba860f39f94752d6062890e70bffdf6146337a87a7536709140b7bb2e233210b6d5b70025dc17be1e8bf2500e35f39a724083b171a10bc630828c9f18fbf02aaa5765e7a99b2c6bbc24b098896bf58d1e7ef33d138c71b5287c180a01aee3748519de6aeb8a223fa49ac3a1414df3b8deceecae06212fb667747c20f3c8a6ae821db039d64a2d11d32a9d379ca3640b943f5c35b7ba5ff9a2fed9967a7c865052d03bbf230eee067f92e74ea549a637b0694731431909498f7fb7424bacf3e89f965794f37df4a3b8398c2a4aa87743a4e7e37171c8d11c40b589cb2d61035f4fc1b7ef335bc3bd9dc8acdd79c75d7a434681d85048954f3e2d4578b4963e34d41878788fe96001e5b3536385010c3304513efa8fe4476017087c7098a052e40d2f58af32f44a2b0bd1560324c795e82cac439c7391e7c951789543c08b278ba3ed606ce92300a3db53aa84680ec5d67669e433aab514ebeeb275fb972eee001dcfc382881c440d3102ac716b64b5f61e38e821b1858de204f9fb506563f2052724f636ce455535e0dc44133e57be54e4d4bc4a3cb285abfdd920d96d3c21eb224f24a9381fb14bbf4e744dfe783b199b4a49fd55a295f2511449d8d7ee781c11b9eada5af755a8d7a47a811f49150e943784712bc8868ff0498bb99811ae71dfa0d64090642da982f3fab30c0c4372eadea4ef6ed7e8a9f22ab7249619083749c7331d25a3ce39634647db6690d26dd365bd672e3717e8e994494601d1b0a894e8e9f3854614fc42b215b2623a3a0df0b7316f05d19d75da12b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'h45b3238a66b484971a8b896683435efa8d12f94a637758dc5fa8ce26ac92ce4c81e19d7a38cb914bed896e08d310838fc0a2e62122852d24697eeafb8954e4665a78e6c068fb24c1017dfd46c3bc4660fd2213eb220b37a6e57b2f0d8eecd064c6f7fd1ab0b04f8c58496ca2aaf9794960693a5388c15537e9eef1e0046130747009b3827a8b9b26893d9c47391d35aae32d3ed8f50d91e46fa49e023de48e43d74a4ed9eb38e35879e36b84d33d8cb41853e20121bdf26d179f798db790754eba1061bc5f00743b02b657d776070ef9201958808c1533118f5234041a065143c4f894f64fbcbc4c919ff9201fc65eee488f53896019efb5c5dc34a6b56a1f89728f04a70cb5598bf5be4191aa724dfb47244c8e7259fd9240fc660a1c2deb89316952111ae395ac3b9fd08990d62f4ac83ad221baa1831aae0792821f3f532546f79cef9c428383625cbd2f7482aec46b490a5b3fd8c28f424084a50347ef081aca1ebf00bb0b1aa5357f4f13942f63547749424baffe8f5686898cf6057f61bae442a247701d22298f88e289db6107dbdcc4c2a7d3d773e682fd84d65e81c680717de06b90b9c1eea95151dfe2cb948484bd23a16e7a2561083f9e6b65d1cdf2ca48f48ce77d1791cdf908fc5c115af4e63950a84af650710781737cafc92ba64f07fa9aa36ad23152606fdf433dce7f44a439e69694f03ccd8c4c87f9a19a0dfccd703415181c2a7978ad605ef704d2e8f9bd2daf5135df7c6205cb3f62b9843155d422089bb40922293976030787acfd0d98214d5c9a0ff5d2a957c3e6439936e9afd8355c1e724c6acafae47555c29112fd30af920c63262b20077804f736143bee5d351d5efa3f56c31da37bf1c9deb3f9aceab9ddd5c35470659668e4e7286077b73fe828;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'h5d68e50343ebe566add2f84679eeb0c686cb3650686658b2ee19de32f01027c65abd33f6f8f8499758b93632cbd9aeb64f9f766a91e4f140e30bce2c42ccc9586619cfad8adb802615d796dddb5814fb0f9d375e9d2afc4612f41338e1c6e68ac5a76e1a7e8b1e253cf1d28f83ff8811dd3c3a0afca7fce4206d092d22523cf1ca9534101a46a121c6ccb679e5b8e3f75b846138e461a0205dddf8f2fa319d5638c555fc476b701b3082e4c011cbad05563969b52ae0380cc8a95a453fd95dc46a061f3b7bff021302e694305ee7d824fae86c4edebede55b8f9ce92fa5f6bae8191d5a06e53b2d15a151f10e3c6e1db112de770ce87f7318528e15629be477b99e577bf531fad947fa577d1785e6f8cae68a8f157bc3894719c43422e3e438ea025a3e877dcb2e2cd3a82fbc6d14f2a61a01f6d162ddd32ab9629170993754f4fc039fbb66f5bf1f83102b561e117daae9dd8758caf71cfd47b205b55638e5e51131e336bf39473a0714a4ad49c605d70086d5acae8dafc09b009b7b228d61a545c1ccb9dd386395deaf717b37792d4a75221d911b360a971dae4bc7f8264fc26b0b2bed2855d954c89dba8400e774e170f3fafa0b1320795d42ba4292314f82fc159ec4ea5976dd154c839e25c1cb96d752eeb62cab06086877fba988362f1fab3f769c409743b994be99b7bea1e4f3a6ca0045a080ee550d89d027f0b8e77c6e39d0f6bf20e8c4187b461a7f374e5dcaabd95e5e438e717ac9bbf12ef2de8c9d4ba68afa8d805039484f06b4c0f6f72f4729c52835f6830b642346a92be59fcbac7bfc2238aa273a95754781b00818006bf363b987433062ffafe26a9521c1949d65ca0b3e4579bfc4265b7415bcce7650dbaeba6eaa8963c5d07579cf3f43bb34b133f3081bd;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'h147222f6bef95394abf2d528b179dbc4a509b6326779d651df499da27acc552d2f2c28fbb1e1326cf12b86b589438b4ada1cc303efd66ba01e2f0f7fcf2da9c8a6e89791c1ec0f5545f8c69cb97e2355a5d9d1c7b6c5fa903eb443becd25c42f9ff09d34859a9c9e0e04a9bdd687730afb7dabd1b884e830f9c6ed83d49692fe6ddd03be785e09276f5400c829bfaaa1dbc8aea140e5683842715ec643f3aebc6ce9a4cd98271df3ef35fa830fd9546f0031a78bf75710b1b6a1ab227037b1da535194b2b451b7926852f3a0f914f44df2d08d7b9b7ec74b10ec91a1e30af19a4da01898154a9a172fbbae088621bf4437318ade1078104e31e1650484a4f8caae0d1f010639a32ecac4addde0f164b9a0f92360838e9fd13975a7ce71b9ae5d8f91b1eeb5831422de67312702ee5383b8cc21823632682890cc676e7ca035acaca5adbf0a0aaf757b7d09cdd8740ecc7ec2840697237abbbc8c753f3e8b7771c9878de617368bacfb25417d0c755c852f3e4a64f79587d5f984c51c06e95140721e1954b0435bef83a9a3933413e907c7b712b087bbb8703ea5f8d73e683b86e745d64c2d726276d416949e674480c9c31800d38124927c31a313e814a55e7865a339eaad1080e7cd91253ad504843078e61f0576b6760a42152f7b8a5fbdafec9b94690b975bc66e3dff0faf5f13f2343e40b1d0522e23d2a772f15e73dbd912c61a8400ae55472e68c17ceb6d577ce6ddf06f064480ec40de273550311f218b23dcc6636a6c9758c4541dc3e3d89254e6d472b7a93be0926b2b7a0d2e3844fd4afec9ec4a6909660635128af470571010f3e87ec4f10575ffbd161018996623d8618398de3626abab5c39658a50d98b1187fae11fa25ce347da7ec85d44f528d108a4b5a03f7e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'hd5638eb9c50fa6c387860a8ad07c48addc918e795615cd69b0924fae34526ac3844cb0559547532d95338eb391827784e77ffe31254b373c72307d8a98ccf1d41f1501a93c3962a2083f29d390c3c61c2f5886adfb090af69a66de74ae6fde614fbbb02ddb033a218b09a2495ad33254aab4f5adb19668e7462629d27573aebd1cc0821353e3527bd1e8a593fb27df71ac535d540c8f779122781e0f0b76d2d75db33e189b7fb2f10c7d7be143328e8b4155a29f48dc96d5c98d0ae9d5ef226601b557cfee9f52d5b862611a0cb10adedc14b3acfadd97691b2e917774172e478c61880e851873d0112f1eef3877280c21718d74f55954ef519c6846fb83c6d0726b0ca860982ae5132c9f04f735d0d4725b935f514fdb02dc2aac025278837c6d6fe3099a43377a8925936b01c35c6ad020a2cfa32781df7a27af8d10c535184390acfbb57b41dded2898c7140c9e0491d71694f6e02b946928e076095dd4596a596537f198a79d242eb05e1fe10843068f75b4b8199610fe7f188370506a1193a73bee1398d837ee5799e439d00331d0d2da1f32eb382dec8edab2a14b7d16993dad9d236061a821075d3e91654bda6115fad1c2228001a96bb113ec88e9a91774985dded093f2bab69b3ce304517e126a280063c58dd7bdc647655ad2345048c4b11180c46b1921692b4ecb88569cc8e5912dd02d62b6dce1a179c2bfeee73dd60f0a43f3a3bd2da565b8d01c80f64cf03588b80068e47cbf6ce1653d485cbe7f8aef2cab67c040e28278c8e794a96a9ee1a7d6fdefbcb5b07499c8612a00c2a3d764e4d33662996ae3f7575dd528b88b8a1bdbde0be0a5cea48d7347bf1c45d057a133c43dcc61091e36408d93283a8c67432e6164a9668142457f38f5d67aaf9900ee36a3ca;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'hcfbb92f95548197eaa7ec0a2c99bfd32363688ffc64cdfa03512cafedf0331da9de2055380f106034468c12dd4926cc01ebbd865fb9f582dc3123bc66715d3e706f26481e53b1f5cdc96c52894a55f99957efaa8165241c4e931295c91dabf85dce09ece4d7540648eec007751972a9005c93f759581d01aa40791d33eda89e320df4d2efe0d1023f60b632f1a4e414597a0b6a28536267f915d631b0012c04ee1fb6d8c6e1681738fd1705719be7e52ff21e96958d9b023e49a572702f373e327c1ac26c13a02147e0f53ddb7c8db86795741727fd059ab3062a50ff3fcbc0232779703c4490dd873a38f5ad26c48b7cd55b3332042d0b77c5eb68e8f81cecdf78381da4e0dcf6e69b3f421c0e1324b3c2359981f51bd96932562eefefe22dc7bfac7bc5ff1e9cb1fa7a1f378f835590fb1883cad954a727d632492b10dab16da4f73d1c18a2b4ed5f3f8acd6282c2365287baf0380635c99c3db2596f592b311c166b0fba947c33b591ba3932cc2ce645bc6359dfa912c29f8f9f2276b8e9706e32f57007aa12c2385b2b15abf7797fb6446b37b75a9f0c8372214bf19a52c26e189b1711f01bc4e536d5ff984b56136771595b0067672aa3bf56882b5927c86c34bfd54ba45fa7c44c029304c49dad8be850260a67730c84cf99ecd23ba1b24d7a82935ac2dd4eb2aa80f5fd9295a5388f052338a0279e9d7dd389021f870801acc1a846b02e71cf603c43b6d8fbe459fab906bf5cda0c275bc80ffce63656cfcf49130ea131f57f90e6be82d96d4db00ae624757a9dc4b05637329a8cadbe0afdb91af665a08ba1336f3c5dc3adcf6ac1105420f99dc968bf43fc4e73752dab10f6bc09df732815ddcfcd6e337d2de4a2d4d41056e3c97c3784d5a5243861d900cb1b3ecd851;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'hb7ca3969ac031b1fb3b3e9a28da4acf117c3822e02f3d8ff4c7a7daae04d550e5c536c4a4dce98fe8703f28d602c44959be7f4d833491b051e2cde6135ce4cdcf53f2f08cd25f2dbeb184d477013310a5e43f5df4895cf1ffa9bfd471e7c90399d878be057dbae91d5f7a56cfd608d2a6c11ff0e2017e34c4080cfbbc66215f07c3772072e0514f75699256ea5e663ef924b48cc283a51649f381f8e54470309abbc0feb4804165e4dfea90c6a222f32c60c2722c0199571ee3b3d7465b08aba64554ba3608dbcb0e89299682d7b90c73f0978a6f56fdf74e10532a101fef1ba663ae5e45df895be7a4be87c04531c7d45b47e7ddda6fc21d46169d6580d192320196ebe45724414ad04f7e054407b60729bdb3646607667b4bc779848a2ed2900c008ab7f217af5dd5d57e7343768e68bd08511d8de07036b5140361c3160ebfeea3cec20b3c0dcfcface6326409c3e06c23bc390692721180e0643326255d0abcba7a38714a1c67e9bd24d71abd9b0141ae3f66453568fa475964c7f317e40920f6d603c381fcc7350a1e2fd470e4fdb771a616ed6380d8a0ff4bf59f83dd31d3859a88f52aff6502c9c8a398978a7279a1b9bfff8dc4b5cc790a7eed6fe3e978b4b00e533c75cd3422d8b713c843547174a37b8019747518c11a342cb1d9f1fd95d23da5e4d929aa9b9081305adc9d365f31d4e07666444d41cb615be53dd29f7f88fdfdebe828fd00cee89f0c15ac4a3d4cf3abee28ca22d1348436f979c47b21e524053bf5b712a7d138a989894584a550cdb6f00f08eeb93df94a46d27abf07d5856f3e36a29c4d074f5bc7ac675bbaca8eab9d09786c11395bbd676db4c7b355a8d9ac12e329579ca85b80ddc1c4439f096c841136caa14b039b507b1e98f1dd70ca9ef16;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'hb912ed0fd7036c4fd96ed67e5225ceb8af2be4e0e9f14f96d2f4a0a37416a1937b96860cac9db07eb2868a443fcc7382468e1eb143bd35ed470a43d556e5425ea154fff433daaa44ba47d4e9c08e12512f898589674f6cd3965af8bcf9e423852d1c56a652ee0b7a63262b4316ecc66ff600420374194875322905a7d3f079598edef12c69f97fdfd9d72e97e54109fb2b2f8e0ca9263eb6cd2974f5a76c57de7b8fb76b3ef76930e439bd064d84e9505ba05c94ed0a480db2072b235f23c651de8efa5a2b4980e5c33b0cb636a8c8438750d7f62229524bf3700895a7e6adb94649531432134fc6b5ccd94f7bd4bac53d1699b576ee8509f2c0868fe01600b19f3a7f00f15f375fda321d9d94b4172c86412f652e7ffa03f1a650ad6a209e3a133031f68aa013095d6000d71393796ba360acbd27ea1799cf071ae4c17b318dcca88e63af91760a1e4264ff880672b1fbc8c2bded6f832c87083dfb520a314b93047c67d2623da2cdd747e22c6ed3c645149734396171461e35114b0da45e4974101eb3a70b195f8f426bc593866fe0d339a7e9a7bcd08093a4ace3d2fc64ec314b6d2bb4bcf273f35d51c83a874dd382eac894ff63cbfd9cf5ea7c7007898110e88230e881cbf8a7b4e1d5e2ee745f86a9af76f3d0ca15f3cdc529bbf23b4960b5421c55cb848bb8f2237a7072a85b3bd70774d4652bbffd26446b4762e9b373d40b20f868c53443e9864462270c86a9d3c8f7d4d9e5ba5e185a642798ca1dce45b832938990a6928223419162972fd852ff63748bf67ef045c1885b1023f99c9825bc124ae7f72a65ca83f7684beae9e22e827acbfd39edc8bd7496150ac3ae27aab9785a9fe772423b91b27852123141a9e55c6e47b2df5c3349f9fc9a1afd214df258fe5f03;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'hc0d17092af1192afcd1c7209baf16f93f1cfa3231cc2727c42c1cd329d471036c2fce4f7ef36faa2fcb96a732c2fb86f8b363fa3bd0c5ab43f9c5ae82e01d30f93d129ef37a975931461311c1d7336c8e85cd06634c58f9f4d000849bfc9e562d1af0f803187f4b5f83a610a8a92d42e9087def9d3f8ce596e79eccc80c88a5a46f22688b6ab9910b10987a5848151800bd5e321d80a3f1980d27506d6164eb014280aefd94b4b06946d1dbc134d5992885e5f9a3093365363e4f9db3d939fdcce3aa27df329affd5a2c89c76ea976ebc28e5497580a57a59aa7c356b9d21bd6ae22a57eab5feca77348935a910d501c8983d94d969c277b745fc2a8a63b6eeaa050d10b25069e01be077c84e4e0fd27af9e108d616c042f378ec44fcb8b055056560aceb1c369aab561628f714272d675db316cdb11a60d13a1c7d406d50d1583d2872e5841dbf8c267240d88db56c7d7053e368a0fe1999c619d326feffb67c4fd5faaa5e737dba0b5bbdef9a35b0775b24917f434a43eb5bf8df7867b922dc5a26f6dfbcc6a9d5c0ef18866a1e2208f2402c08b3346aca57e607d8fbe5604a27bc6d4f9a8feba5a2437550456b9687fcea84093374e118e495daf4373743390159505e00d8b05b82b34d07fe8c7a3fd9638723e0d7c895c05963d040581654182a966e6e82956ad3e682e3906c0c0a27e6bb0fde1bf93bc69005f1d7d9917218fea1f5aa57fdd5597f32c1dd495ead26c20890418d382a534cc35055b7c0dab59b3648f68a321bb91030ab3bdc6844de74cbf85b229c36518614cee63fbd1f6e2dc93d46c7230173ed862dee4650a2e25d52dce724be25c8fa5a8a4c8df0a5cac2f456b22cd2f50347e5abe5ac8b54a7743c2e3045c6078628ec0c8a203c17c80ae739e8ba1f8;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'ha2212701deda954a97ada895ba608f9f7f17850d2931329ff732d0e5db0e9df508c12f2f58cbd87bd25870dc75c5bcc4d900c09a986e400b14ebf01ab4e4ea288e90a7bd06b1b2e877ddd2bb2763da80341acf7321ddce4ca0f557045c76ae2dfa06c6088fe72178795316499218d1a772f8b25696aa675d50fcdc21a6532900306671d09ff0c5fdac0ac42161a42cf22c922caac5c5bd3ea01a65a2cd010b04d10ad1c7b5f32cfc57723f62e00a940aab47213c5ae611cf7508327f1ec718deba489ddc4acd6152918849ec2e356a6455f9303ad2db44f57a8ceea5bb4242fcd7c91c044998f00f0c9fc5a2438f2026e850a64600bfa388fbbb16d9599ef502db04013f135fce0c01cf464629dd4181165c4bc0facfbfb535f40aa309cdcb98db2b0c6cff46bc3a077f5603e1cbb8ad79fda89b20fd844b881a8c85fb83fe0f02d968113df1aae561601d22f45cd2d4a1d40a3a910aefc07863ddf3ce240746dc802cf30d71727a7dca95c83496a0a87ce454bfc2b31e188fdc1cc2e0adba9b93bebe84bdddfbac7c27b4d2dda401f0c8f874719f60c7702e2fdb2ddaa165da9512ba9bcb8a7907db630a9d2dcbd323c0f44157cba1156fa61b8d8f1b5e042bf1c43a24e92a9ced6985a0db66d3de350471db0aa883b7f9bce3b8c24689f4b5ccc1051420444f0af93bc0bf718f3f23bac835fcfc4c25e1ee1715f934cf61ab8ce07e0da8b24d168c2f13729f6c135ea92e137c9828281b7102627aefac2e65f5db83abade68df1581a81d0b639224d03d391356a16117c9834f27df440da48226dfe20bb62f803e05844ecf3ef56ab842091a097e0a1aa09934e06f95e6f24781e050b63c3be5be1545fa780492495c7b7a03f76fb2c7b50135c8704b8c4d322f87d5672400d9c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'hd18d0caa0d874110350f4b432b3740908d795ab3624f96d0a615b7b6feeff870338729932010b0e228407992e02d40bdcf663b35954f67ad1f00813941e2f4b60d84d6b0f98c65eafb84421fd89e901111f43aea9430cb1d623fed2d34a31f9783c58b6a78665cd81c535b1cbf1c64c15f6c6a31225e8c4488a0b922b921716b63b39c660c5239d8900c4c7bc1274caed68542b9e22fb5566b22bc978231903a1f4ebb15aad1439e0f24da767b7d6596b44de8084e74b2b717a7f2fcf17b6a94aefa846fe161b7114b8cd43cf0197e520ebdbe5fd9167d7770703ceb00fa093367e17f04d385e4787ac664a016a42900a17373c3462f70f7fee0bf27e76df502d4aaa787c6c9912f85e497f2e7bc113d006097c66a10e71a8281a97fb0bf1ae4e1d7bc0334402507a698ddb5f09b6d0ed7993abc52e0e5faf12d54d779f8bf4ab9df12c42e7adb2940aa274298777549d06f2edf74955510725b24922cfac41d8c7e8e8c60800b237a22f94cc9bab770011ddf1144e98d472442189de131d5e489e96a915809ade6838065b11a590e7d4501082cf179e73d4318e15188592790f09c2eba38b39877e9be73e1c5d1e1b92a0dc5aa503e7ea1ca66445b75e0a3d5a1569f5417f36a722c33f8afcd0a9507dc1cc6e77e34d5127e9c84e23193a4d32c7db40af1dce97f6c91581b90fab31dc7b880b6b33668cb5e387fa1084978f9ebe33dcfa186956586ee24580249ec977dcae19a13232717ba52f5e846ec3033e55248226d942b56ba11c592c9c5945d44ff6f3636f9b1cc4bd1e759973493758dadee26ea43e7c38da08a7e8a7fccf58f06c2f3b3dcc02157c335ecf44b4f753c1314a403cd34752b941553ab17a36bd45c46c222c745d7d5c831a048f968b3cdeaee53891d2eb8;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'h4c626761bbf1306f7d8663c4bddf74e1282f76f7b4f9d2c81377c0eb028dba9d76f1eff253cbce001565d39ece61c854cd4cebbd6b894a8814bac8afd2f316685c53405fff11bb0aa7b98749dcc16ab815a950d7cc4f2dec92cb75960db1d0a4df1aeb9d49c13ecd187ea32f7d0c069279d29e19f2e0291697b090143dee93f4b3d0ad481e4027dc94e7de87b2e47f5afa73c58322a87ca470fd2196379f02c68122b267aa743eb8d64d1b2694c96bf1c5c1c697d11f69ed05bcf7d1db4ec635c7527b1f9f6cd464f4082676c998f9e7a861cff95b96cc0626d05b9b068212dc58632781381112605a3621213b2de38897fed9931055c3c0262642321f1924571f1445ebd3690c340a3d6721da6369cde84e94219e8b8f8635683d8c86b995b53e697545d4087ab7a18f638ee9d87102773d52d36928b201ecafbf94a99e573089f329d1d091d66d8554e150a7f968abbb1fbda4fd12a969774717bc116a84b0984f67153fafafbbc270ce0d20e72388bfd8a691201f8967aceb34485ee470bffcffa5d9478f8d60ce420a89272e6d92c869e7eca8cd4f33833576748472c6d09f564122ec8662404f2077e022fa240a3c83554544e5910c24facaae34a2254247840cb55e658295765a1c388e99095e835543686d9e208f74fc49954b7bd6689f0d39702ddb41fad050d5df0f8f1efaf5d0677003f3c49076563f78150f04270a5914798276da09c91e5cd8318299665790e0078528e4b1a31399cfd86faaf5c6c674627de335157b9da5e03d90ec60891319d0a4f14ee09d1338ccbf732c1f5b67df178b08b8420253377ff58f29b7c25d10f1abecae288b13c18477fdeb4b3ca75357596771dc57c1591f18917ca5287e263af000b653eca7b076931de6d1a1f105f8e8725a36;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'he667fdb67479ce57f55dfbeef9db5b93d5f397d9e06e6ba73260cd6cb89a4defc71b7557e0163cd07e0823e5ae9c376df5b2bdb03ad15667d6eee3dbacaedace5791139bd8c26a8aa5249fe424115c48db8899abb62c5eab443b382c9ce6d6d70b5089967a4d3dba56a9548341868bf6b28d1902bbb2bd41041b720a44c23840d9b69dc823966902312b68b3e21d420ab19e34c36c6d581d5b65424d18990606f62e13afffddfc32b014aa6cb8a06545c1dd6ddafe0e0cb341835b52e47fa7d3871e5476e45a2529e0d0f647cf7a1fb317c876d7e198aac3c83032ef9fda974716bedc85ea22ca3911f8d90ea28e54356044e75f687ab0d6b1865fcc7ee0018de2e730dbd759684c08104e358024fadd4c8cbeab0734f7b4595a479d81be511702fec621c3ebc621d5bc051a2d03929a413c08e57223a63af5d21605dddc63f3ea451beb6d6a97312bf6b5f7d5b85839d1672b2919e0be9944606e65b223383e88c1f76cf02101246e5fcf6bee9bf8fccf8fc27d95681c3ff8d644c750775851b5ef0dcd958c82eb55fe1486e50a77e47433e348c761c30b80cba613b4638a1be1f0b6d9ddf24b3df4be21de92d7830fd60874d37457d304af4610a2b80dad9b1d3b62919fb381f2aeadca2434fab4934cf74313563de5118ce8a156535896d5c9671e8756b171044c4dbbf682ab2ca2e5bb43be5e763e60c53151ae2c262287d4a0aef7a395a1086d911c130df2936c9f56e8209cd5802bf7c6e8ed163808bd81fba082d19727461f8865573d64949229cb5f2668dbf5e3932105129fd11332331adb2594e83aa4672300e7df5f2f7bc4dffc7c8b7aa35a027f05868d21a8c946519b06515f68878835cfb0effa02756edb8c2ae12ed4c97f214c7cdd6f1df13a2fa1bcc6a8c06e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 5184'hd5e67dcaadf58ab3d728f866b73b4ca1cffddea2e60d5155979bcc36bbaf473d89a93293f91634c9dc577fffb75124414b47108d3295496ece540de87eb068a817b2d98af043e6b47b64635c63efb52e2cc0879d7886527ffe59dc5452b4c85a02e1379d79d86acb68c01af5637512ccfe337aa38ddde5c2435560a3589491fd000ad9b93589384fc77a982ac8523ec175562ab0c81f1c45f2f8476ebd8fc3052a7abd067fd95d9395461d89e5aee31bf3411dad21934354cb4066e9f04e87de40e424848b346980f430779cb51338eea514f8ee9ee41ca8262cbf06a3f0131e9f62b119982da54986455ba3a76c697a73d4717f66bd29ab44dd244c5b6abd23c00f908e8fd7097941102103a48a65161cfe63e215f43b099fac5358a72c2be8e8cab001fec6ac9cf78fefa878eaec113fb81fc4a223d19e3c133e576d5619218c5c8dc6e789e51261bc6c0213bbd252be1de22090c45461aa4128ff31b7a3caeeeb12cc60d7ca93a032b0f2053cfead1088a325c5dc9e877719d560a807e795fc42167ebe025cd2be2de98c9f5ac1eb9479293d9c4555b6a2ac556e1715e2da78ea592a9318c3356fc8515b6c1287549a68fbe6d771a07701cb571a249aa48658c1692cee8b4880914535f9a4276b643c2e2a97d81d085bd70f18d915dc59c137361603288b266e7d7795084407d8b8698c8067c707219435887794aa8228638a0d627b36d029602ad392043c13824e457f1ebcd427c20539ca3eb7d8a1f6fdc8da474f33517c86b66c94e183cc86a2f6e53c7d432713c2531da24c845d1b204d4baaf570a7eba4a1b425818bfeee3e6b7d811b44b55c1b533f7249374a1606ba3957db36b7560ee45464bd069d5cb3a08350ed2e4944803f119ffb90584aed51e3d9ae0d73370;
        #1
        $finish();
    end
endmodule
